module layer_10_featuremap_214(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b2cdf),
	.w1(32'hb7583992),
	.w2(32'hb79a295f),
	.w3(32'hb88e608b),
	.w4(32'hb76a63b0),
	.w5(32'hb76ff9fe),
	.w6(32'hb8ad3374),
	.w7(32'hb7c1dc8a),
	.w8(32'hb816b745),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba70ba2),
	.w1(32'h3ac7c910),
	.w2(32'h3b840fb5),
	.w3(32'h3b30ddfc),
	.w4(32'hba91942c),
	.w5(32'h3ab86b02),
	.w6(32'h3b027b20),
	.w7(32'hba8b195e),
	.w8(32'h3b115a83),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f6220a),
	.w1(32'hb629f44e),
	.w2(32'hb7ad1346),
	.w3(32'hb7b27436),
	.w4(32'h36ead680),
	.w5(32'hb73c48d6),
	.w6(32'hb7e932ad),
	.w7(32'hb6a714bb),
	.w8(32'hb7d59949),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c777),
	.w1(32'hba77a174),
	.w2(32'hba6dd503),
	.w3(32'h39538f68),
	.w4(32'h397310c8),
	.w5(32'h389edab2),
	.w6(32'h389061b9),
	.w7(32'h389c0e40),
	.w8(32'h37e99175),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e6e1e),
	.w1(32'hb896dab8),
	.w2(32'hb75902fb),
	.w3(32'hb9a26ca1),
	.w4(32'hb8faebca),
	.w5(32'hb8eec697),
	.w6(32'hb9b7aaa9),
	.w7(32'hb97d50f3),
	.w8(32'hb99e8ef4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a14ad),
	.w1(32'hb636576e),
	.w2(32'hb82289ee),
	.w3(32'hb85702f4),
	.w4(32'h34d4be12),
	.w5(32'hb817cd09),
	.w6(32'hb88ab28b),
	.w7(32'hb587db6e),
	.w8(32'hb820bb83),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba072561),
	.w1(32'h3b36beb5),
	.w2(32'h3b84970f),
	.w3(32'h3a350714),
	.w4(32'h3b7076a9),
	.w5(32'h3ba03275),
	.w6(32'hb9b4fc7d),
	.w7(32'h3b274065),
	.w8(32'h3b9011cf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef6d9e),
	.w1(32'h3b800184),
	.w2(32'h3b31ca92),
	.w3(32'h3c082d51),
	.w4(32'h3c113cce),
	.w5(32'h3bb07d6a),
	.w6(32'h3c0ddf08),
	.w7(32'h3b584982),
	.w8(32'h3b6a4db8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e40c3e),
	.w1(32'hba22cf99),
	.w2(32'h39be41a6),
	.w3(32'hb9a132b3),
	.w4(32'hba7c331e),
	.w5(32'h396823c7),
	.w6(32'h392b45d9),
	.w7(32'h37b13496),
	.w8(32'h3a7cd35f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beebcb0),
	.w1(32'h3a615a2b),
	.w2(32'h3c2779c0),
	.w3(32'h3ba896be),
	.w4(32'hba71399d),
	.w5(32'h3bb0dfc6),
	.w6(32'h3bd33ded),
	.w7(32'h3abdc176),
	.w8(32'h3c15f875),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba93aa),
	.w1(32'h3a10aa04),
	.w2(32'h39cf62ae),
	.w3(32'h39773772),
	.w4(32'hb6073771),
	.w5(32'h39406655),
	.w6(32'hb80cb15e),
	.w7(32'hb91f59ab),
	.w8(32'hb740e8de),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ca996),
	.w1(32'hbb20c43d),
	.w2(32'h393df56e),
	.w3(32'h3b8886b1),
	.w4(32'hb984ef8c),
	.w5(32'h3b270d89),
	.w6(32'h3b714bc2),
	.w7(32'hbaa89ec6),
	.w8(32'h3b6bdc31),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be14770),
	.w1(32'h3b36112f),
	.w2(32'h3c267797),
	.w3(32'h3bded279),
	.w4(32'h3b13cbed),
	.w5(32'h3c0212b8),
	.w6(32'h3bb74a26),
	.w7(32'h3b9bf64d),
	.w8(32'h3c15d895),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e7e93),
	.w1(32'h3b180bbc),
	.w2(32'h3b7385a0),
	.w3(32'hba73abed),
	.w4(32'h3aa02e5f),
	.w5(32'h3b05a44c),
	.w6(32'h386543d5),
	.w7(32'h3a844c2b),
	.w8(32'h3aabaa55),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501005),
	.w1(32'hba885aeb),
	.w2(32'h3b21b782),
	.w3(32'h39267203),
	.w4(32'hbb960b9b),
	.w5(32'hbaa30c02),
	.w6(32'h3b0559c4),
	.w7(32'hbb2ba16a),
	.w8(32'h3abf4c14),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be68ce5),
	.w1(32'h3b5cfe9f),
	.w2(32'h3c25d641),
	.w3(32'h3b947772),
	.w4(32'hb9fbef9b),
	.w5(32'h3b7ad41b),
	.w6(32'h3bc7a730),
	.w7(32'h3b6d15da),
	.w8(32'h3bf50776),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb858482e),
	.w1(32'h398463a2),
	.w2(32'h392816b9),
	.w3(32'hb8f67bc5),
	.w4(32'hb6068aa7),
	.w5(32'hb925d4d3),
	.w6(32'hb8e4e2d8),
	.w7(32'hb8df6df1),
	.w8(32'hb9a2e3a1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7e5cd),
	.w1(32'h3b5774f5),
	.w2(32'h3bbf082e),
	.w3(32'h3bc8fd88),
	.w4(32'h3b284f6d),
	.w5(32'h3c027235),
	.w6(32'h3bf64a97),
	.w7(32'h3b5cd274),
	.w8(32'h3bd46d53),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b365c0b),
	.w1(32'h3b001115),
	.w2(32'h3bbb48cf),
	.w3(32'h3b0ef3b1),
	.w4(32'h3b32ca66),
	.w5(32'h3bbdd246),
	.w6(32'h3b5d7117),
	.w7(32'h3b532142),
	.w8(32'h3bc08064),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c685bd),
	.w1(32'hb9168ec2),
	.w2(32'hb891e503),
	.w3(32'hb89f12b8),
	.w4(32'hb9605980),
	.w5(32'hb9073116),
	.w6(32'hb8818669),
	.w7(32'hb93c4129),
	.w8(32'hb86767a5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92faa38),
	.w1(32'hb8102ec9),
	.w2(32'hb8b8c436),
	.w3(32'hb9158b17),
	.w4(32'h36996cd5),
	.w5(32'hb8a3bfb4),
	.w6(32'hb943798f),
	.w7(32'hb871e499),
	.w8(32'hb9439ab6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3abfcc),
	.w1(32'hbac152f1),
	.w2(32'h3acfb455),
	.w3(32'h3963d7f1),
	.w4(32'hbb204edc),
	.w5(32'h3a578eb5),
	.w6(32'h3aa29f56),
	.w7(32'hbaac3731),
	.w8(32'h3aa510e4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c434869),
	.w1(32'hbaa90d11),
	.w2(32'h3bc03bf8),
	.w3(32'h3bd5681e),
	.w4(32'hbba1f5ae),
	.w5(32'h3b7f91ef),
	.w6(32'h3beaba30),
	.w7(32'hba5fa02d),
	.w8(32'h3c3387d5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca5449),
	.w1(32'hba5f628e),
	.w2(32'h3bff38e6),
	.w3(32'h3b0b4d52),
	.w4(32'hbb95e1dd),
	.w5(32'h3b54c967),
	.w6(32'h3bb2c689),
	.w7(32'hbadc89a8),
	.w8(32'h3bd7bcb3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3baf4f),
	.w1(32'hb9facd54),
	.w2(32'h3be0ca4b),
	.w3(32'h3c11f07d),
	.w4(32'hbb76ff3a),
	.w5(32'h3b2884ea),
	.w6(32'h3c5450be),
	.w7(32'hba1d8e55),
	.w8(32'h3bb8b2dd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4435c),
	.w1(32'hb8c418c7),
	.w2(32'h37e1c57a),
	.w3(32'hba14e4c0),
	.w4(32'hb98e43e1),
	.w5(32'h389aa013),
	.w6(32'hb9b39fca),
	.w7(32'hb96a8d23),
	.w8(32'h39804df8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0529d),
	.w1(32'hb9553700),
	.w2(32'hb9b75aa0),
	.w3(32'hb97a30b9),
	.w4(32'hb915e26a),
	.w5(32'hb993d4cc),
	.w6(32'hb9a1b3ed),
	.w7(32'hb987cdee),
	.w8(32'hb9d5d067),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b8f7e),
	.w1(32'hbb83fdca),
	.w2(32'h3a23be0b),
	.w3(32'hb9447e99),
	.w4(32'hbb626c73),
	.w5(32'hbb7926e9),
	.w6(32'h39301d05),
	.w7(32'hb8b0d503),
	.w8(32'h3a9b4d63),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b452a),
	.w1(32'hba88dd27),
	.w2(32'hba083155),
	.w3(32'h3b27d08d),
	.w4(32'hba92a0c8),
	.w5(32'hb84a8916),
	.w6(32'h3b8def17),
	.w7(32'hba2f909e),
	.w8(32'hb96bccbd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fcaea6),
	.w1(32'hbb8c2881),
	.w2(32'h3b77f16c),
	.w3(32'h3a5e832c),
	.w4(32'hbba66eaf),
	.w5(32'h3a57595e),
	.w6(32'h3b56fcb3),
	.w7(32'hbaec2937),
	.w8(32'h3b8ea746),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8891917),
	.w1(32'hb8278ad3),
	.w2(32'hb87ebb12),
	.w3(32'hb8987b59),
	.w4(32'hb83ac3b4),
	.w5(32'hb877e84b),
	.w6(32'hb8bc829a),
	.w7(32'hb88c8896),
	.w8(32'hb8a1f995),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ac3e09),
	.w1(32'hb7f99e87),
	.w2(32'hb85581d6),
	.w3(32'hb899d5f4),
	.w4(32'hb7da4d4d),
	.w5(32'hb8a7fbe4),
	.w6(32'hb876d21b),
	.w7(32'hb816d4d8),
	.w8(32'hb90d98ca),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1b6c),
	.w1(32'hba509762),
	.w2(32'h3b4dc947),
	.w3(32'hb976c8b0),
	.w4(32'hbafe2258),
	.w5(32'h3ac9afc9),
	.w6(32'h3aa1fd3f),
	.w7(32'hba6605bd),
	.w8(32'h3b1da52c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5736cb),
	.w1(32'hb9b5ff94),
	.w2(32'h3a80fef2),
	.w3(32'h3b1df67c),
	.w4(32'hbae5e6bd),
	.w5(32'hb9961fa6),
	.w6(32'h3b6f94a5),
	.w7(32'hb9fb4873),
	.w8(32'h3a48209a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a4006),
	.w1(32'h398f1d08),
	.w2(32'hb88d73ed),
	.w3(32'h3a8daa80),
	.w4(32'h3a76d3a7),
	.w5(32'hb8271ea3),
	.w6(32'h3a30cf52),
	.w7(32'h3a4b051c),
	.w8(32'h3a2e7d12),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30c80f),
	.w1(32'h3b00f999),
	.w2(32'h3b23028e),
	.w3(32'h3a53bf73),
	.w4(32'h3b18e305),
	.w5(32'h3b43e645),
	.w6(32'h39b949eb),
	.w7(32'h3ab992a5),
	.w8(32'h3aca9ba2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96b4c8),
	.w1(32'hbafb8cc6),
	.w2(32'h3bccf380),
	.w3(32'h3b4e2a72),
	.w4(32'hbb8a2a08),
	.w5(32'h3b835f55),
	.w6(32'h3af89cea),
	.w7(32'hbbf37356),
	.w8(32'h3bb337a0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f8e31),
	.w1(32'hbbc79628),
	.w2(32'h3ab87309),
	.w3(32'h3c3b4ce9),
	.w4(32'hbc29928a),
	.w5(32'hbb416597),
	.w6(32'h3c8bf54e),
	.w7(32'hbb7b2191),
	.w8(32'h3b6eb339),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc65d42),
	.w1(32'hbc250b25),
	.w2(32'hbb5d3a51),
	.w3(32'h3c1732ed),
	.w4(32'hbc1147c4),
	.w5(32'hbb9561d5),
	.w6(32'h3c5cdff2),
	.w7(32'hbb387356),
	.w8(32'h3ae50aa0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27de72),
	.w1(32'hb9b1774f),
	.w2(32'h3a0d893e),
	.w3(32'h3ad77aed),
	.w4(32'hba9c2cd1),
	.w5(32'hba099988),
	.w6(32'h3b288b1e),
	.w7(32'h36cd2678),
	.w8(32'h3a7d53c7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925a0b4),
	.w1(32'h3832f85f),
	.w2(32'hb8814e23),
	.w3(32'hb8ebb07f),
	.w4(32'h38927ae8),
	.w5(32'hb7e1c27f),
	.w6(32'hb96844c0),
	.w7(32'hb82a1929),
	.w8(32'hb92242f8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a7052),
	.w1(32'hb8a4b7db),
	.w2(32'hb99ba565),
	.w3(32'hb95f29b9),
	.w4(32'hb8600d5b),
	.w5(32'hb998993e),
	.w6(32'hb9b69005),
	.w7(32'hb95b1588),
	.w8(32'hb9d95f00),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ca084),
	.w1(32'hba0aa8dc),
	.w2(32'h3a0a01c2),
	.w3(32'h3b0b95c8),
	.w4(32'hba66a64c),
	.w5(32'h3ac44429),
	.w6(32'h3adbf58d),
	.w7(32'hb9f58aeb),
	.w8(32'h3b261892),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ee027),
	.w1(32'h3b2c8fcd),
	.w2(32'h3c206602),
	.w3(32'h3bf4e5f2),
	.w4(32'h3b20efd9),
	.w5(32'h3be18393),
	.w6(32'h3c1cadc8),
	.w7(32'h3c007cdd),
	.w8(32'h3c3308e3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25d9d),
	.w1(32'hbadec1c4),
	.w2(32'h3bdccc46),
	.w3(32'h3b1e25f7),
	.w4(32'hbbb7160a),
	.w5(32'h3b051db8),
	.w6(32'h3bb20e00),
	.w7(32'hbb3a94ea),
	.w8(32'h3ba61c03),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b3789),
	.w1(32'hb9fbefb8),
	.w2(32'h3c02813e),
	.w3(32'h3b91060d),
	.w4(32'hbb8093d1),
	.w5(32'h3b728adf),
	.w6(32'h3c0b3043),
	.w7(32'hbab4a5fd),
	.w8(32'h3bdf4d68),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd6df4),
	.w1(32'hba05fa17),
	.w2(32'h3b94c415),
	.w3(32'h3ba514b5),
	.w4(32'hbb38c61c),
	.w5(32'h3a993d3f),
	.w6(32'h3bb6efbe),
	.w7(32'hba4badd1),
	.w8(32'h3b8ebf2e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12839),
	.w1(32'h3b6d0ba1),
	.w2(32'h3bfaed33),
	.w3(32'h3b79c71b),
	.w4(32'h3bbe1a1a),
	.w5(32'h3c0b1ad8),
	.w6(32'h3b9012b4),
	.w7(32'h3baeb87b),
	.w8(32'h3c0276c3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39305c8f),
	.w1(32'h391b39cd),
	.w2(32'h3945e398),
	.w3(32'h393e5292),
	.w4(32'h395a8e61),
	.w5(32'h398c4bf4),
	.w6(32'h394d3ac7),
	.w7(32'h3971fa49),
	.w8(32'h39297cf4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e46281),
	.w1(32'h384862e0),
	.w2(32'h3893ad09),
	.w3(32'h397158e4),
	.w4(32'hb9125c49),
	.w5(32'h396f67ac),
	.w6(32'h3a031a0c),
	.w7(32'h39c56a9d),
	.w8(32'h3a32cd72),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d9c26c),
	.w1(32'h37b36350),
	.w2(32'hb7d66886),
	.w3(32'hb8339e69),
	.w4(32'h3860304c),
	.w5(32'h38e291c8),
	.w6(32'hb93bbb1f),
	.w7(32'h371cbd1b),
	.w8(32'h38cc5910),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4a7fe),
	.w1(32'h3a1ba70b),
	.w2(32'h3b83e580),
	.w3(32'h3b43294f),
	.w4(32'hba7a4a4f),
	.w5(32'h3b01af65),
	.w6(32'h3b382d29),
	.w7(32'hb98d2bb5),
	.w8(32'h3b08823b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954703),
	.w1(32'h3951979b),
	.w2(32'h3aa94825),
	.w3(32'h3a3a0c26),
	.w4(32'hb8f85d42),
	.w5(32'h3aadf3ae),
	.w6(32'h3a59d659),
	.w7(32'hb982b334),
	.w8(32'h3a6e8a6d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beea5e2),
	.w1(32'h3b46f3e9),
	.w2(32'h3bfaafb5),
	.w3(32'h3b94e0da),
	.w4(32'h3b175f2d),
	.w5(32'h3bafdc09),
	.w6(32'h3bb0165a),
	.w7(32'h3b0283c7),
	.w8(32'h3bbee6c1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a623c3a),
	.w1(32'hba3ee923),
	.w2(32'hb9e6064c),
	.w3(32'h3a921f46),
	.w4(32'h3974f8e8),
	.w5(32'h3a3fb3f3),
	.w6(32'h3abae9c6),
	.w7(32'h38f1b4bb),
	.w8(32'h39e24adc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38120673),
	.w1(32'hb80e99fb),
	.w2(32'h381c360a),
	.w3(32'hb8f2a6b7),
	.w4(32'hb9411a4f),
	.w5(32'hb962bfd9),
	.w6(32'h389b0f23),
	.w7(32'hb90a7229),
	.w8(32'hb9224920),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb838c3be),
	.w1(32'hb80c1219),
	.w2(32'hb785ab75),
	.w3(32'hb89b9165),
	.w4(32'hb87534a9),
	.w5(32'hb80fc665),
	.w6(32'hb88bf9c1),
	.w7(32'hb89706de),
	.w8(32'hb8490ad1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbcc77),
	.w1(32'hba0044ce),
	.w2(32'hb538be16),
	.w3(32'hb9941454),
	.w4(32'hb9910959),
	.w5(32'h379a8766),
	.w6(32'hb8a247d7),
	.w7(32'hb846b690),
	.w8(32'h394fa0de),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6c9b3),
	.w1(32'hbaa12d14),
	.w2(32'hba0c30d8),
	.w3(32'hb909d4eb),
	.w4(32'hbab59e84),
	.w5(32'hb9e2f4a7),
	.w6(32'h3a50e6ca),
	.w7(32'hba063d3c),
	.w8(32'h38f04085),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3973606f),
	.w1(32'h38dfbae4),
	.w2(32'h39b4c628),
	.w3(32'hb68a35c8),
	.w4(32'h38c162e9),
	.w5(32'h39dc1c65),
	.w6(32'h39030bea),
	.w7(32'h399d8cec),
	.w8(32'h3a21e53a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd49dbb),
	.w1(32'h3b3b0c75),
	.w2(32'h3b594a89),
	.w3(32'h3bb0b6bd),
	.w4(32'h3b41c9a2),
	.w5(32'h3b454961),
	.w6(32'h3ba121ce),
	.w7(32'h3b5cf4ec),
	.w8(32'h3b0c435a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba737d),
	.w1(32'h3aa2e33f),
	.w2(32'h3ac40af4),
	.w3(32'h3b6a0a60),
	.w4(32'h3ab52411),
	.w5(32'h3a03f7f5),
	.w6(32'h3b6a421d),
	.w7(32'h3b3ae4c9),
	.w8(32'h3b0b2372),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880dd50),
	.w1(32'h378a4cfb),
	.w2(32'hb84e8720),
	.w3(32'hb87971b2),
	.w4(32'h37b372fc),
	.w5(32'hb862f8c1),
	.w6(32'hb8c6dc30),
	.w7(32'hb757ca75),
	.w8(32'hb8d0aad6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bcbe44),
	.w1(32'hb78a0603),
	.w2(32'hb857b879),
	.w3(32'hb899af04),
	.w4(32'h36a1edc6),
	.w5(32'hb80900d3),
	.w6(32'hb8f0cc74),
	.w7(32'hb82c4716),
	.w8(32'hb8a78cd3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a491dc),
	.w1(32'hb639aed0),
	.w2(32'hb6fe4977),
	.w3(32'hb8c8fbe9),
	.w4(32'hb794134c),
	.w5(32'hb87011c0),
	.w6(32'hb91168b4),
	.w7(32'hb87259dc),
	.w8(32'hb8b6f8de),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c573c),
	.w1(32'hb89470a3),
	.w2(32'hb91845f9),
	.w3(32'hb9330cd0),
	.w4(32'hb8638b44),
	.w5(32'hb8fef16c),
	.w6(32'hb95f0cd6),
	.w7(32'hb8fb5d0a),
	.w8(32'hb94d32fb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4c571),
	.w1(32'h3ba00612),
	.w2(32'h3bf2a0dc),
	.w3(32'h3c06f22c),
	.w4(32'h3bcbb456),
	.w5(32'h3afabb9c),
	.w6(32'h3bbb8940),
	.w7(32'h3bb4a8a4),
	.w8(32'h3bbec849),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042625),
	.w1(32'h38e0191d),
	.w2(32'h3bd4c274),
	.w3(32'h3bab9219),
	.w4(32'hba37e89a),
	.w5(32'h3c0758b3),
	.w6(32'h3beabe31),
	.w7(32'hba6767cd),
	.w8(32'h3be8edf7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e0d8),
	.w1(32'hbb18c68c),
	.w2(32'h3b0d8a75),
	.w3(32'h3bd36ece),
	.w4(32'hbb886955),
	.w5(32'h3af3f0fb),
	.w6(32'h3c1c53a0),
	.w7(32'hba72d392),
	.w8(32'h3b603014),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36f9e3),
	.w1(32'hbb95b82f),
	.w2(32'h3c21fce0),
	.w3(32'h3bcb891d),
	.w4(32'hbc315b91),
	.w5(32'h3b2f7ee2),
	.w6(32'h3c559cd1),
	.w7(32'hbba60dee),
	.w8(32'h3c0a6462),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e2cf2),
	.w1(32'h36d668bf),
	.w2(32'hb8b3d435),
	.w3(32'hb92ce373),
	.w4(32'h3813b400),
	.w5(32'hb822b0a6),
	.w6(32'hb96e768a),
	.w7(32'hb83ee7c6),
	.w8(32'hb90d1808),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b0d09),
	.w1(32'hb84a72df),
	.w2(32'hb95fd727),
	.w3(32'hb987b135),
	.w4(32'hb73921a1),
	.w5(32'hb9395c76),
	.w6(32'hb9c1e633),
	.w7(32'hb916af9d),
	.w8(32'hb9a43de3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950d35d),
	.w1(32'h38fab8ad),
	.w2(32'hb80a49c3),
	.w3(32'hb9507a41),
	.w4(32'h3921f69e),
	.w5(32'hb6f7aa25),
	.w6(32'hb9b73964),
	.w7(32'h37a605c5),
	.w8(32'hb925d848),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04a14f),
	.w1(32'hb8e98c0c),
	.w2(32'h39c4f9c6),
	.w3(32'h3ae22a64),
	.w4(32'h393779e8),
	.w5(32'h3a3a9e5e),
	.w6(32'h3b2108c6),
	.w7(32'h39f2ff88),
	.w8(32'h3a05904f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94b68cb),
	.w1(32'hb86b8810),
	.w2(32'hb91c5d85),
	.w3(32'hb92c788c),
	.w4(32'hb764eb78),
	.w5(32'hb8ebac8f),
	.w6(32'hb9887d99),
	.w7(32'hb8c8b278),
	.w8(32'hb93de4c3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad395b),
	.w1(32'h39f5620f),
	.w2(32'h39bf36c0),
	.w3(32'h3b141edf),
	.w4(32'h3b208be6),
	.w5(32'h3ac65e32),
	.w6(32'h3ad4e9c4),
	.w7(32'h3a90a2b0),
	.w8(32'h3a3c1fbf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d498c),
	.w1(32'h3b94d94c),
	.w2(32'h3bb861b2),
	.w3(32'h3bca8d08),
	.w4(32'h3b6b9251),
	.w5(32'h3bd14dd8),
	.w6(32'h3bd4948d),
	.w7(32'h3b4e86a0),
	.w8(32'h3ba7098f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8f368),
	.w1(32'h3b24ee57),
	.w2(32'h3bff7f28),
	.w3(32'h3be8c163),
	.w4(32'h3a8d5fb7),
	.w5(32'h3b9e8e87),
	.w6(32'h3bee791b),
	.w7(32'h3b21f4ea),
	.w8(32'h3bb6336f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a3b1),
	.w1(32'hba01978c),
	.w2(32'h3b37e725),
	.w3(32'h3ace375b),
	.w4(32'hbacb1176),
	.w5(32'h3a6198d1),
	.w6(32'h3b4bda11),
	.w7(32'hba042255),
	.w8(32'h3ad0e046),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de4721),
	.w1(32'hb8bcab9c),
	.w2(32'h3b4b01b0),
	.w3(32'h3aaaf5e2),
	.w4(32'h3ab00089),
	.w5(32'h3b0f93fd),
	.w6(32'hb9dc8a9e),
	.w7(32'hba02ef39),
	.w8(32'h3b5720bf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44e58c),
	.w1(32'hba2d8fe4),
	.w2(32'h3b031c00),
	.w3(32'h3ad1f8db),
	.w4(32'hbb001bf9),
	.w5(32'hb8d0ba7a),
	.w6(32'h3b372312),
	.w7(32'hba1be4ae),
	.w8(32'h3ab0d24b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa204b8),
	.w1(32'h39e7a488),
	.w2(32'h3b433d01),
	.w3(32'h3aa9e4b8),
	.w4(32'h3ac82519),
	.w5(32'h3b75dd22),
	.w6(32'h3af63fdd),
	.w7(32'h3a882b4c),
	.w8(32'h3b43f317),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a5fb65),
	.w1(32'hb64a2d8f),
	.w2(32'hb7de6281),
	.w3(32'hb7843309),
	.w4(32'h36a279ab),
	.w5(32'hb7b2ce25),
	.w6(32'hb80367a4),
	.w7(32'hb68b2b54),
	.w8(32'hb817925d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76ff71a),
	.w1(32'hb6910500),
	.w2(32'hb6e1b533),
	.w3(32'hb81e5d81),
	.w4(32'hb824eced),
	.w5(32'hb8334215),
	.w6(32'hb7bcf16c),
	.w7(32'hb7b261fd),
	.w8(32'hb7d477ba),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ebb436),
	.w1(32'hb838dbe0),
	.w2(32'hb88594f8),
	.w3(32'h38f1663a),
	.w4(32'h3880c468),
	.w5(32'h36207cff),
	.w6(32'hb7ad7720),
	.w7(32'hb7be4d81),
	.w8(32'h3882d298),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2e344),
	.w1(32'hba1cf5d7),
	.w2(32'hb9ec281b),
	.w3(32'hb9758ecf),
	.w4(32'hba027dea),
	.w5(32'hb9d24db5),
	.w6(32'hb7c103f4),
	.w7(32'hb9ac2278),
	.w8(32'hb965ac92),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be233b2),
	.w1(32'hbaffadba),
	.w2(32'hb9b402e4),
	.w3(32'h3bbb521d),
	.w4(32'hbb53d213),
	.w5(32'hbb2871a7),
	.w6(32'h3bd7634c),
	.w7(32'hbb566116),
	.w8(32'hbabd73c2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7678045),
	.w1(32'hba1f3a41),
	.w2(32'hb997f5b2),
	.w3(32'hb9204097),
	.w4(32'hba734e26),
	.w5(32'hb9ec7f13),
	.w6(32'h3a24ab22),
	.w7(32'hba11293c),
	.w8(32'hb800c968),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b884dbe),
	.w1(32'h3aab9766),
	.w2(32'h3b88b3d1),
	.w3(32'h3a92e8ed),
	.w4(32'hbab4cf6e),
	.w5(32'h3b1e90ea),
	.w6(32'h3b3d1f91),
	.w7(32'hba0c79e0),
	.w8(32'h3b5cb243),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9e65),
	.w1(32'h3a9773e8),
	.w2(32'h3b2574e5),
	.w3(32'h3bee2b0b),
	.w4(32'h3a51d47d),
	.w5(32'h3b1ae4fa),
	.w6(32'h3c157ad8),
	.w7(32'h3b2866ea),
	.w8(32'h3b3c3eef),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc6835),
	.w1(32'hbb9e4978),
	.w2(32'hba440361),
	.w3(32'h3b5c71be),
	.w4(32'hbb8734ed),
	.w5(32'hba24522c),
	.w6(32'h3b86643a),
	.w7(32'hbb57145e),
	.w8(32'h3a5cfee4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab8c84),
	.w1(32'h3b91d585),
	.w2(32'h3bea614f),
	.w3(32'h3baf1b7c),
	.w4(32'h3a79c7ce),
	.w5(32'h3b27d719),
	.w6(32'h3b1c7361),
	.w7(32'h3a9ecc76),
	.w8(32'h3bd32ef2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba498434),
	.w1(32'hbb80967f),
	.w2(32'h3a07af33),
	.w3(32'hb9227450),
	.w4(32'hbb39d115),
	.w5(32'h3a3da7ca),
	.w6(32'h3abb5054),
	.w7(32'hbb238b3c),
	.w8(32'h3782179a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01e2cb),
	.w1(32'h3b136d5d),
	.w2(32'h3bd96500),
	.w3(32'h3ba15c63),
	.w4(32'hbacd51f5),
	.w5(32'h3ac8bf81),
	.w6(32'h3bc3e8f3),
	.w7(32'hba9b4738),
	.w8(32'h3b846b39),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d4d5f),
	.w1(32'hba3807a8),
	.w2(32'h3b353e99),
	.w3(32'h3acecc03),
	.w4(32'hbb4ce477),
	.w5(32'hbab041f1),
	.w6(32'h3a33d34d),
	.w7(32'hbb0e3859),
	.w8(32'h3a895fed),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3976b),
	.w1(32'hbb1544aa),
	.w2(32'h3b7cab15),
	.w3(32'h3b6cd2c9),
	.w4(32'hbb8a3129),
	.w5(32'h3aa6b499),
	.w6(32'h3bcb9d4a),
	.w7(32'hbb1cf340),
	.w8(32'h3b27cdaa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df22c4),
	.w1(32'h3a138991),
	.w2(32'h3a4bd6f6),
	.w3(32'h3a08df2a),
	.w4(32'h3a496f61),
	.w5(32'h3a3368d1),
	.w6(32'h3a0edaa8),
	.w7(32'h3a284e12),
	.w8(32'h39e98dc4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbb0e4),
	.w1(32'hb4236c30),
	.w2(32'h3bd98a5a),
	.w3(32'h3b6310e6),
	.w4(32'hba9603c0),
	.w5(32'h3b9c7d48),
	.w6(32'h3bd0d34e),
	.w7(32'h3b10ca46),
	.w8(32'h3c078a53),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e65b4),
	.w1(32'hbb05abca),
	.w2(32'h3b3623f6),
	.w3(32'h3ba38cd2),
	.w4(32'hbb2005d2),
	.w5(32'h3a225d82),
	.w6(32'h3b5965a2),
	.w7(32'hbaa23d84),
	.w8(32'h3b886f21),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10213a),
	.w1(32'h3a81db1d),
	.w2(32'h3bdf02d9),
	.w3(32'h3b95d545),
	.w4(32'hbb0e8a82),
	.w5(32'h3b967207),
	.w6(32'h3bc08527),
	.w7(32'hbb30a26f),
	.w8(32'h3b9ee8c4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d71fa),
	.w1(32'hbc20931d),
	.w2(32'hbb84bff0),
	.w3(32'h3b9dd8ac),
	.w4(32'hbc9ec771),
	.w5(32'hbc5d6e1c),
	.w6(32'h3be8d0ca),
	.w7(32'hbc458b7d),
	.w8(32'hbb8dd0a8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9be6bd),
	.w1(32'h39104239),
	.w2(32'h3c1a0db7),
	.w3(32'h3b06c4a8),
	.w4(32'hbb1f1fc1),
	.w5(32'h3bba6cea),
	.w6(32'h3bcb53a9),
	.w7(32'h397afe50),
	.w8(32'h3c050c17),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0841),
	.w1(32'h3b3397be),
	.w2(32'h3bcb9f2a),
	.w3(32'h3ae62ef0),
	.w4(32'h3a6ac1c3),
	.w5(32'h3b253095),
	.w6(32'hba819290),
	.w7(32'hbb346921),
	.w8(32'h3ba6fb6e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bff9d),
	.w1(32'hb8ba55e9),
	.w2(32'hb91a9dc6),
	.w3(32'h38989dd2),
	.w4(32'hb9b252d2),
	.w5(32'hba04edf5),
	.w6(32'h391b9e4a),
	.w7(32'hb98c68c6),
	.w8(32'hba115f7f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d6d38),
	.w1(32'h3b9cf381),
	.w2(32'h3c0f9a78),
	.w3(32'h3bf9dcb7),
	.w4(32'h3ad13846),
	.w5(32'h3b9d858b),
	.w6(32'h3b43cab7),
	.w7(32'hbb606a59),
	.w8(32'h3aad850c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adac69a),
	.w1(32'hb8bb5910),
	.w2(32'h3b80662a),
	.w3(32'h3ba2be24),
	.w4(32'h3b048ce4),
	.w5(32'h3ba70f82),
	.w6(32'h3aff55a1),
	.w7(32'h3aa01989),
	.w8(32'h3ba59723),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a69f5f),
	.w1(32'hb92397e5),
	.w2(32'h3938b1a9),
	.w3(32'hb88c04fd),
	.w4(32'hb9a5964b),
	.w5(32'h3811f9c1),
	.w6(32'hb86e0b12),
	.w7(32'hb99e8c32),
	.w8(32'hb7444c62),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22ce95),
	.w1(32'h3ab74454),
	.w2(32'h3ad39700),
	.w3(32'h3a9c4a93),
	.w4(32'h39d855e7),
	.w5(32'h398a4287),
	.w6(32'h3af53b54),
	.w7(32'h3a1e8097),
	.w8(32'h3a21b82f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25555f),
	.w1(32'h3af7658a),
	.w2(32'h3bdd56d1),
	.w3(32'h3b34e448),
	.w4(32'h3b2048f9),
	.w5(32'h3bcbf54c),
	.w6(32'h3b8333bc),
	.w7(32'h3ba262b9),
	.w8(32'h3c0c42c3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b4122),
	.w1(32'hb9ef6ca9),
	.w2(32'h3baca417),
	.w3(32'h3b049b97),
	.w4(32'hbaa55b1c),
	.w5(32'h3b390de8),
	.w6(32'h3b88e2f5),
	.w7(32'h390c69d5),
	.w8(32'h3b8721b2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2982cb),
	.w1(32'hbae2b941),
	.w2(32'h3ad826d7),
	.w3(32'h3b090304),
	.w4(32'hbb57bfb7),
	.w5(32'hb9b08538),
	.w6(32'h3b2ca036),
	.w7(32'hba9150a0),
	.w8(32'h3b228471),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819ae5),
	.w1(32'hba55a85b),
	.w2(32'h3b3d5456),
	.w3(32'h3add8ce6),
	.w4(32'hbb2df80f),
	.w5(32'h3a64019f),
	.w6(32'h3b096f94),
	.w7(32'hbb0e669c),
	.w8(32'h3b2ec103),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b072),
	.w1(32'hba9efa24),
	.w2(32'h3a02bf13),
	.w3(32'h3b350b35),
	.w4(32'hbab96b20),
	.w5(32'h3abf4680),
	.w6(32'h3ba6d1ec),
	.w7(32'hb92d23c6),
	.w8(32'h3b131695),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96e928),
	.w1(32'h3b0470c7),
	.w2(32'h3bbe4778),
	.w3(32'h3b092f94),
	.w4(32'hbacc54ae),
	.w5(32'h3a382f9d),
	.w6(32'h3b233d44),
	.w7(32'hb911521a),
	.w8(32'h3b494a2f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d71e0),
	.w1(32'hba20ac20),
	.w2(32'h3b175871),
	.w3(32'h3ad84724),
	.w4(32'hbaaeba3f),
	.w5(32'h3aa46f5e),
	.w6(32'h3b56434d),
	.w7(32'hb797a56f),
	.w8(32'h3b3b25c9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5c385),
	.w1(32'h38b72341),
	.w2(32'h38a965f9),
	.w3(32'h389401cc),
	.w4(32'h37ad416b),
	.w5(32'hb82c8163),
	.w6(32'h37fb42f6),
	.w7(32'h382f6ed7),
	.w8(32'hb842254e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a282275),
	.w1(32'h39cfa6a3),
	.w2(32'h3997ef6b),
	.w3(32'h3997d747),
	.w4(32'h387b7943),
	.w5(32'h3691f879),
	.w6(32'h39d906a9),
	.w7(32'h3841b0bb),
	.w8(32'h3902d141),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6f917),
	.w1(32'hb9922866),
	.w2(32'hb96864b2),
	.w3(32'h391192d6),
	.w4(32'hb94a7258),
	.w5(32'hb95a14de),
	.w6(32'h38aa08ed),
	.w7(32'hb94445e8),
	.w8(32'hb935aca0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fd07b),
	.w1(32'hb97a4fee),
	.w2(32'hb98b8ed6),
	.w3(32'hb783d7b5),
	.w4(32'hb8bde6e3),
	.w5(32'hb92bc158),
	.w6(32'hb8c7b1e0),
	.w7(32'hb962e21e),
	.w8(32'hb9daae7a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c47d2),
	.w1(32'hbaaefd4c),
	.w2(32'h3b3a72a7),
	.w3(32'h3ab10c9c),
	.w4(32'hbb50b131),
	.w5(32'h3ab2f51e),
	.w6(32'h3b56f257),
	.w7(32'hba9bdc56),
	.w8(32'h3b61c728),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d376f),
	.w1(32'h3a6c8490),
	.w2(32'h3a956e60),
	.w3(32'h39eacfd4),
	.w4(32'h392f3c13),
	.w5(32'h3a39d6e5),
	.w6(32'h39eeb878),
	.w7(32'hb81fe47c),
	.w8(32'h39d2da10),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ebb70d),
	.w1(32'h3a692ca9),
	.w2(32'h3b6dc6d8),
	.w3(32'h3aa465a3),
	.w4(32'h3acabaae),
	.w5(32'h3b3c1908),
	.w6(32'h39948c77),
	.w7(32'h3a922ced),
	.w8(32'h3b2723ba),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08cb44),
	.w1(32'hb994e290),
	.w2(32'h3b8e0ec0),
	.w3(32'h3bb5f487),
	.w4(32'hbb39ed1b),
	.w5(32'h3b02f162),
	.w6(32'h3bcf7456),
	.w7(32'hba84b171),
	.w8(32'h3b9d0dde),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a26d7),
	.w1(32'hb8c1a55b),
	.w2(32'hb784ecbb),
	.w3(32'hb9785f5c),
	.w4(32'hb933e981),
	.w5(32'hb9302fc4),
	.w6(32'hb9a1d63c),
	.w7(32'hb9886c49),
	.w8(32'hb95fe0e8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a14c82),
	.w1(32'hb72e83fe),
	.w2(32'h39895412),
	.w3(32'hb9cf88cb),
	.w4(32'hb9c17ec4),
	.w5(32'hb885344d),
	.w6(32'hb8bc27e2),
	.w7(32'hb81111b2),
	.w8(32'h39958cfe),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893c20b),
	.w1(32'hb82fae0b),
	.w2(32'hb85b6a73),
	.w3(32'hb8ae8ff1),
	.w4(32'hb8508aa7),
	.w5(32'hb865ec73),
	.w6(32'hb8d054e2),
	.w7(32'hb885b6d3),
	.w8(32'hb8a0d376),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39831e94),
	.w1(32'hba56edb1),
	.w2(32'h397e7b1b),
	.w3(32'h3a49c493),
	.w4(32'hba924c64),
	.w5(32'hb8a400e1),
	.w6(32'h38a759c5),
	.w7(32'h3a36fe7f),
	.w8(32'h39dc8950),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2943f3),
	.w1(32'h3b9119f0),
	.w2(32'h3b6bab30),
	.w3(32'hb91fe002),
	.w4(32'h3b99d41a),
	.w5(32'h3bdc487a),
	.w6(32'h3b27bbcf),
	.w7(32'h3b442548),
	.w8(32'h3b61e90b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b756835),
	.w1(32'h3b390bcf),
	.w2(32'h3bfb1eea),
	.w3(32'h3b045a21),
	.w4(32'h3ae21702),
	.w5(32'h3bc493c8),
	.w6(32'h3b844864),
	.w7(32'h3b75758d),
	.w8(32'h3c13a11d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b959d),
	.w1(32'h39eae664),
	.w2(32'hb985ebb1),
	.w3(32'h3b47c91a),
	.w4(32'hb93c9d5c),
	.w5(32'hba8422f5),
	.w6(32'hb79c6c9b),
	.w7(32'hb9be359b),
	.w8(32'hb9232797),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fffed),
	.w1(32'h3a795856),
	.w2(32'h3a8d869f),
	.w3(32'h3a9b75f2),
	.w4(32'h3a8892d9),
	.w5(32'h3aec27de),
	.w6(32'h3b48b5e2),
	.w7(32'h3a46ae9b),
	.w8(32'h3aa89693),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba977e),
	.w1(32'hbacb1d52),
	.w2(32'hba731e05),
	.w3(32'h3af38f04),
	.w4(32'hbb54b04a),
	.w5(32'hbb17f41c),
	.w6(32'h39deea24),
	.w7(32'hbb3aa175),
	.w8(32'hba28d21c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12d595),
	.w1(32'h3aea7bfc),
	.w2(32'h3b504206),
	.w3(32'hbaadcfe8),
	.w4(32'h3a8331c5),
	.w5(32'h3ade15c2),
	.w6(32'h3b8750bd),
	.w7(32'h3adc8a93),
	.w8(32'h3ab906e5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0e3f),
	.w1(32'h3b82fc8e),
	.w2(32'h3bbfd841),
	.w3(32'h3b85d41e),
	.w4(32'h384a24b9),
	.w5(32'h3a969d93),
	.w6(32'h3baf2e7f),
	.w7(32'h3a9ff1ac),
	.w8(32'h3b5b2592),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ca9e9),
	.w1(32'h3b254a9b),
	.w2(32'h3b9309b3),
	.w3(32'h3bc204f3),
	.w4(32'h3b2f7731),
	.w5(32'h3baba95b),
	.w6(32'h3ba7c336),
	.w7(32'h3b354925),
	.w8(32'h3bf7b982),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3f72),
	.w1(32'hba5d0643),
	.w2(32'h3b45d537),
	.w3(32'h3b342e84),
	.w4(32'hbb05deb7),
	.w5(32'h3acc2110),
	.w6(32'h3b3f29b8),
	.w7(32'hbab74eee),
	.w8(32'h3b41b54e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881668),
	.w1(32'hb9339bae),
	.w2(32'h3b652f40),
	.w3(32'h3b33314d),
	.w4(32'hbad7ab27),
	.w5(32'h3a52b2e4),
	.w6(32'h3ac5994f),
	.w7(32'hb92865bf),
	.w8(32'h3b40763c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d2773),
	.w1(32'h3b37d38f),
	.w2(32'h3b4e41d8),
	.w3(32'h3b42fa76),
	.w4(32'h3a9065aa),
	.w5(32'h3b775216),
	.w6(32'h3b9bf89e),
	.w7(32'h3a54c54c),
	.w8(32'h3b8bf189),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27058),
	.w1(32'h39b9aadf),
	.w2(32'h39f21fbc),
	.w3(32'h3b877cf7),
	.w4(32'hba49c596),
	.w5(32'h38c949a8),
	.w6(32'h3b556705),
	.w7(32'hbb2f063a),
	.w8(32'hba9befe7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cab25),
	.w1(32'h3b0c57ce),
	.w2(32'h3bd22606),
	.w3(32'h38ec785a),
	.w4(32'hb8b2fcda),
	.w5(32'h3b4ca7a2),
	.w6(32'h3a81efdf),
	.w7(32'h3a23ec52),
	.w8(32'h3ba3140f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a13ca),
	.w1(32'hba42788d),
	.w2(32'h3a3b3a95),
	.w3(32'h3a8ba159),
	.w4(32'hbac3e87f),
	.w5(32'h37c19bca),
	.w6(32'h3a3b3b4b),
	.w7(32'hba054d11),
	.w8(32'h38c5999d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432a4a),
	.w1(32'hbb8f7f1b),
	.w2(32'h3b9d773e),
	.w3(32'h3b851b77),
	.w4(32'hbb672fb3),
	.w5(32'h3b8b83e9),
	.w6(32'h3bb89075),
	.w7(32'hbb459b5a),
	.w8(32'h3ba327f5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad572),
	.w1(32'h3b2f699b),
	.w2(32'h3aba462a),
	.w3(32'h3b443e8d),
	.w4(32'hba214b86),
	.w5(32'hba8b1cc4),
	.w6(32'h3b8d2528),
	.w7(32'hba8236ce),
	.w8(32'hba675392),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35baa6),
	.w1(32'h399fddb5),
	.w2(32'h3a115144),
	.w3(32'h3a2eb97f),
	.w4(32'h3a0728cc),
	.w5(32'h3a2a7640),
	.w6(32'h39b45f6b),
	.w7(32'h39e48bae),
	.w8(32'h3a380fb3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a539d5f),
	.w1(32'hba8cb98f),
	.w2(32'hba1c4648),
	.w3(32'h3a68d5f0),
	.w4(32'hba0f9f18),
	.w5(32'hb98283de),
	.w6(32'hbaa8f50c),
	.w7(32'hba56374b),
	.w8(32'hba530e03),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae15450),
	.w1(32'h39e5fc1e),
	.w2(32'h3a23bc8c),
	.w3(32'h3b0e00c6),
	.w4(32'hb89bd431),
	.w5(32'hba70fe42),
	.w6(32'h3b135436),
	.w7(32'h39a5c3a8),
	.w8(32'h3a8df2e0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fdbdd),
	.w1(32'h3919e0b8),
	.w2(32'h3b46620a),
	.w3(32'h3adacdd8),
	.w4(32'hbb36b147),
	.w5(32'h3a5b0bb3),
	.w6(32'h3b9894fe),
	.w7(32'hbb03b9b9),
	.w8(32'h3b7aba6c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e56fc),
	.w1(32'h3a91e952),
	.w2(32'h3bdc4512),
	.w3(32'h3c230554),
	.w4(32'h3adbbd43),
	.w5(32'h3b913941),
	.w6(32'h3c04e120),
	.w7(32'h3b6bb176),
	.w8(32'h3baf08b9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd10d5),
	.w1(32'hbab28f0f),
	.w2(32'hba754bd2),
	.w3(32'hb95dedef),
	.w4(32'hbaa1308c),
	.w5(32'hba75ba6c),
	.w6(32'hbaf318bd),
	.w7(32'hbace6208),
	.w8(32'hbb2c2117),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dcd8b),
	.w1(32'h3b2323ac),
	.w2(32'h3c231340),
	.w3(32'h3aa10f79),
	.w4(32'h3aa1dadc),
	.w5(32'h3bc58be8),
	.w6(32'h3bc511c0),
	.w7(32'h3b3caf54),
	.w8(32'h3be8bfdc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad288),
	.w1(32'hb9e59201),
	.w2(32'h3b689a61),
	.w3(32'h3b484f37),
	.w4(32'hbad77ef6),
	.w5(32'h3a830fd3),
	.w6(32'h3adaebf1),
	.w7(32'hb906f06c),
	.w8(32'h3b54bca0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81f62b),
	.w1(32'h3bab7284),
	.w2(32'h3c1490ad),
	.w3(32'h3b0b6f47),
	.w4(32'h3b4433c2),
	.w5(32'h3babe819),
	.w6(32'h39be20ad),
	.w7(32'h3aeba375),
	.w8(32'h3b8d1dea),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73537c),
	.w1(32'hbaf1071f),
	.w2(32'h3ba95f63),
	.w3(32'h3afd57c0),
	.w4(32'hbb8c3935),
	.w5(32'h3aedbf50),
	.w6(32'h3b9cabe4),
	.w7(32'hbb094abb),
	.w8(32'h3b9751b2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8606d6),
	.w1(32'hba3a92ee),
	.w2(32'h3a0326e2),
	.w3(32'h3b5a7365),
	.w4(32'hba45d4a9),
	.w5(32'hb870ee77),
	.w6(32'h3af9740b),
	.w7(32'hbab5b129),
	.w8(32'h39577d09),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000438),
	.w1(32'hba72a377),
	.w2(32'hba96bc03),
	.w3(32'h3913d8ce),
	.w4(32'hba8da4f5),
	.w5(32'hbab1ce1f),
	.w6(32'hba457d57),
	.w7(32'hba5bbc3c),
	.w8(32'hbacd80d1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5dd26),
	.w1(32'hbb0c0685),
	.w2(32'hb8a1c95e),
	.w3(32'hba1ef00f),
	.w4(32'hbb76ad8a),
	.w5(32'hbab86fa6),
	.w6(32'h3b87906f),
	.w7(32'hbaca2874),
	.w8(32'h3ac2fec5),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd238fa),
	.w1(32'hbb61c92e),
	.w2(32'h38b21ce7),
	.w3(32'h3b91a906),
	.w4(32'hbbdb830f),
	.w5(32'hbb0ec5ed),
	.w6(32'h3b585d0d),
	.w7(32'hbb8519f3),
	.w8(32'hba303002),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae760d4),
	.w1(32'hbb946204),
	.w2(32'hba1332ee),
	.w3(32'h3aed9b0c),
	.w4(32'hbbac9d5e),
	.w5(32'hbaf6ee3b),
	.w6(32'h3b2375a6),
	.w7(32'hbb34a1e3),
	.w8(32'hb9cc1179),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b44f08),
	.w1(32'hba20e0f7),
	.w2(32'hba30559e),
	.w3(32'h38c8946b),
	.w4(32'hb86a8bf8),
	.w5(32'hb9ec95e9),
	.w6(32'hba6dad35),
	.w7(32'hbaa6a8fa),
	.w8(32'hbac9ca2c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf08d3),
	.w1(32'hba2a8ffb),
	.w2(32'hb9e41bb3),
	.w3(32'hbae746bc),
	.w4(32'hba6af9df),
	.w5(32'hba33d344),
	.w6(32'hba58795a),
	.w7(32'hba53c03c),
	.w8(32'hbaa36d3c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca53b),
	.w1(32'h3aeb77aa),
	.w2(32'h3ba3d4de),
	.w3(32'h3abcef18),
	.w4(32'h397d932d),
	.w5(32'h3b571fc9),
	.w6(32'h3b1d4f7f),
	.w7(32'h3aaa18bb),
	.w8(32'h3b6fd673),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71cd5d),
	.w1(32'hba28be93),
	.w2(32'h3a04da4d),
	.w3(32'hb9c73b3e),
	.w4(32'hba3175f4),
	.w5(32'h39f3e16c),
	.w6(32'hbabde260),
	.w7(32'h37fc4ca7),
	.w8(32'hb91a4f39),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7af4b4),
	.w1(32'h3a0250e3),
	.w2(32'h3aeb23d0),
	.w3(32'h39141e4c),
	.w4(32'hb9c9ecab),
	.w5(32'h3a839355),
	.w6(32'h3b8937b5),
	.w7(32'h39d09c5b),
	.w8(32'h3b3ad401),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5a4a8),
	.w1(32'hba2c75c6),
	.w2(32'hb9d4d31c),
	.w3(32'h3aaf106a),
	.w4(32'hb958b323),
	.w5(32'h373dcce1),
	.w6(32'hbaa71da5),
	.w7(32'hbaa9b273),
	.w8(32'hbaaf19c6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a86a),
	.w1(32'h3a8f437a),
	.w2(32'h3abf5384),
	.w3(32'h3b9b589b),
	.w4(32'h3b2631dc),
	.w5(32'h3b7efb6f),
	.w6(32'h3b9cda28),
	.w7(32'h3b21f2ba),
	.w8(32'h3b89a308),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d00edd),
	.w1(32'h3a0a33d0),
	.w2(32'hb9821760),
	.w3(32'hba6852fb),
	.w4(32'h38c9efac),
	.w5(32'hb9dcc9fe),
	.w6(32'h3a256236),
	.w7(32'h396a6c4f),
	.w8(32'h392abe86),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7a438),
	.w1(32'h3a3b3291),
	.w2(32'h3a01c02e),
	.w3(32'h397f1ca5),
	.w4(32'h3a5bc95f),
	.w5(32'h3a3130d7),
	.w6(32'h3a320eb2),
	.w7(32'h39a7ce67),
	.w8(32'h392319c9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bdbcb),
	.w1(32'hb971219b),
	.w2(32'h3b1174af),
	.w3(32'hba27f32f),
	.w4(32'hbb2c647c),
	.w5(32'h38722c01),
	.w6(32'h3ae48bcc),
	.w7(32'hbaa080dd),
	.w8(32'h3b2c8700),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be17701),
	.w1(32'h3887bd9b),
	.w2(32'h3bfc8b2b),
	.w3(32'h3b8ced12),
	.w4(32'hbaae7def),
	.w5(32'h3c1652dc),
	.w6(32'h3b8cd242),
	.w7(32'hb9f78a1b),
	.w8(32'h3bfddd3f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241608),
	.w1(32'hbae934df),
	.w2(32'hb9df1665),
	.w3(32'h3b2e40a0),
	.w4(32'hba03b1ab),
	.w5(32'h3a4022fb),
	.w6(32'h3b5cc6b7),
	.w7(32'hba8fc89e),
	.w8(32'h3a843e09),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f9636),
	.w1(32'hba5cf27e),
	.w2(32'h3ba8cbbe),
	.w3(32'h3a95ceed),
	.w4(32'hbb421579),
	.w5(32'h3b4b1f8d),
	.w6(32'h3acd4c90),
	.w7(32'hbab18d5c),
	.w8(32'h3b84faf0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c4836),
	.w1(32'h3ab3d17a),
	.w2(32'h3b018d8c),
	.w3(32'h3941c1a3),
	.w4(32'h3ab4a45e),
	.w5(32'h3aa470ae),
	.w6(32'h3b3820ad),
	.w7(32'h3aebcdf8),
	.w8(32'h3b585a2c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46984c),
	.w1(32'hbb39d1a4),
	.w2(32'h3bb8f9dc),
	.w3(32'h3c2882e9),
	.w4(32'hbb9edda4),
	.w5(32'h3b1869bb),
	.w6(32'h3bb8670f),
	.w7(32'h391b54d8),
	.w8(32'h3b6f4595),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2630f4),
	.w1(32'h3a0ffcf3),
	.w2(32'h3b89811d),
	.w3(32'h3aca6617),
	.w4(32'hbaf258d5),
	.w5(32'h3af8e19f),
	.w6(32'h3bb00b10),
	.w7(32'hbab793cb),
	.w8(32'h3b2db3c4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b70c),
	.w1(32'h3aabcb5e),
	.w2(32'h3bcda8ac),
	.w3(32'h3a8d8e90),
	.w4(32'hbb2289da),
	.w5(32'h3add396f),
	.w6(32'h3b6d5e18),
	.w7(32'h3aac268b),
	.w8(32'h3bafb116),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a572412),
	.w1(32'hbaf151cf),
	.w2(32'hba26795e),
	.w3(32'hbaaec610),
	.w4(32'hbafd1b0e),
	.w5(32'hba5dff24),
	.w6(32'hbb1771aa),
	.w7(32'hba8b53a7),
	.w8(32'hba689cb1),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908dce),
	.w1(32'hb98beefc),
	.w2(32'h3b1f48f7),
	.w3(32'hb9c9ef25),
	.w4(32'hbb0db51e),
	.w5(32'h3816d7fc),
	.w6(32'hba8d5d42),
	.w7(32'hbb170047),
	.w8(32'hba16e7d4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86eac7),
	.w1(32'hba04c4a3),
	.w2(32'hba092dff),
	.w3(32'hba8a6c03),
	.w4(32'hb9a05f58),
	.w5(32'hb992597c),
	.w6(32'hba6543cc),
	.w7(32'hba377068),
	.w8(32'hba9b7cc6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1b6a3),
	.w1(32'hbb63c2de),
	.w2(32'hbb104380),
	.w3(32'h38efb224),
	.w4(32'hbb69c63a),
	.w5(32'hbb27c6e9),
	.w6(32'hbb5a5984),
	.w7(32'hbb7d5cb2),
	.w8(32'hbb50aa0a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299726),
	.w1(32'h3acf1208),
	.w2(32'h3b2464c1),
	.w3(32'hbb0301bc),
	.w4(32'h3abe389f),
	.w5(32'h3ac58a65),
	.w6(32'h3af58378),
	.w7(32'h3ad443e5),
	.w8(32'h3b309dfb),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be078ea),
	.w1(32'h3ac09263),
	.w2(32'h3bb4c173),
	.w3(32'h3bee1f3c),
	.w4(32'h3a0462fe),
	.w5(32'h3b2c4da3),
	.w6(32'h3bdc5132),
	.w7(32'h3b15847d),
	.w8(32'h3bad7346),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d033f),
	.w1(32'h3b81c20b),
	.w2(32'h3b65bd1f),
	.w3(32'h3a6267f1),
	.w4(32'h3b794a16),
	.w5(32'h3b6cdfe4),
	.w6(32'h3b8a6c30),
	.w7(32'h3b85713c),
	.w8(32'h3b5bb1c8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ff359),
	.w1(32'h3aa42cf2),
	.w2(32'h3ad74067),
	.w3(32'h3b656c86),
	.w4(32'h3a8cd1b2),
	.w5(32'h3ab06497),
	.w6(32'h3adb04af),
	.w7(32'h3b0e38a9),
	.w8(32'h3aef2182),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83301b),
	.w1(32'h3a210b18),
	.w2(32'h3aaf7b00),
	.w3(32'h3b2219c5),
	.w4(32'hb9155d95),
	.w5(32'h39bbb7b9),
	.w6(32'h3b21f422),
	.w7(32'h394ef380),
	.w8(32'h39f9041a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8734ee),
	.w1(32'hbb683f68),
	.w2(32'hb9994277),
	.w3(32'h3b8af7cc),
	.w4(32'hbb6f47ab),
	.w5(32'hba842b4c),
	.w6(32'h3a9d2c09),
	.w7(32'hbb1fd4bb),
	.w8(32'h38cd58c0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0525ea),
	.w1(32'h3a457c44),
	.w2(32'h3ad624e1),
	.w3(32'hb9953aeb),
	.w4(32'h3a8ec1ba),
	.w5(32'h3b54e4c1),
	.w6(32'h3a36d94d),
	.w7(32'hbaa2f6e9),
	.w8(32'h3aedbdbc),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6b058),
	.w1(32'h3ae086ba),
	.w2(32'h3ab9d5f2),
	.w3(32'h3b134a88),
	.w4(32'h3aba31bd),
	.w5(32'h3aa2f39e),
	.w6(32'h3b408d69),
	.w7(32'h3ac5325f),
	.w8(32'h3b13fff1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d8943),
	.w1(32'h3c04d798),
	.w2(32'h3c8a0b39),
	.w3(32'h3c5a5ac8),
	.w4(32'h3bfd1fd6),
	.w5(32'h3c668751),
	.w6(32'h3c12cb91),
	.w7(32'h3c0ef353),
	.w8(32'h3c2b895b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31336a),
	.w1(32'h3b0cdd72),
	.w2(32'h3c14bc68),
	.w3(32'h3c053d6e),
	.w4(32'hbb6075d7),
	.w5(32'h381f24c0),
	.w6(32'h3c11116c),
	.w7(32'hbb54c290),
	.w8(32'h3b928bb2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f547f),
	.w1(32'hb90f12c5),
	.w2(32'h39d84eff),
	.w3(32'h3b3aac99),
	.w4(32'h3a51c28c),
	.w5(32'h3a3df94f),
	.w6(32'hba4c0a3e),
	.w7(32'hb979d9d4),
	.w8(32'h39dc7f88),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c949e),
	.w1(32'hbb016796),
	.w2(32'hbab3af6d),
	.w3(32'hba593905),
	.w4(32'hbb271442),
	.w5(32'hbae0691c),
	.w6(32'hbabe2357),
	.w7(32'hbac56e56),
	.w8(32'hbb248953),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb088aab),
	.w1(32'h3ab5c119),
	.w2(32'h3a27d2fd),
	.w3(32'hbaeb25ad),
	.w4(32'h3aa8f553),
	.w5(32'h3a5377b0),
	.w6(32'h3b0b5506),
	.w7(32'h3ad8e4df),
	.w8(32'h3b1514ee),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa39f70),
	.w1(32'h3a8dfbef),
	.w2(32'h3a331de2),
	.w3(32'h3ab98ce2),
	.w4(32'h3a797baa),
	.w5(32'h3a5461d3),
	.w6(32'h3a963d33),
	.w7(32'h3a8853fa),
	.w8(32'h3a5a621f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c53814),
	.w1(32'h3aa37d48),
	.w2(32'h3b4f700e),
	.w3(32'h3a85c32a),
	.w4(32'h3b0c913b),
	.w5(32'h3b8ec337),
	.w6(32'h387de189),
	.w7(32'h3b0e69cb),
	.w8(32'h3b826289),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde629d),
	.w1(32'hbaf277a8),
	.w2(32'hba0655bf),
	.w3(32'h3b91694e),
	.w4(32'hbb8471c5),
	.w5(32'hbaf7355a),
	.w6(32'h3acb6967),
	.w7(32'hbb0b9982),
	.w8(32'h3ae8d760),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd28d35),
	.w1(32'h3b03a6e6),
	.w2(32'h3c0621d4),
	.w3(32'h3b7ec06b),
	.w4(32'hbad20dd3),
	.w5(32'h3b6143d8),
	.w6(32'h3bddf3e6),
	.w7(32'h3a272362),
	.w8(32'h3b65280f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad877c6),
	.w1(32'h39847e90),
	.w2(32'h3a8f4468),
	.w3(32'h3a79f07b),
	.w4(32'h39435088),
	.w5(32'h3a01fb77),
	.w6(32'h3ae2d81a),
	.w7(32'h397925de),
	.w8(32'h3aa0fbbe),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2e92a),
	.w1(32'h3aad2b2e),
	.w2(32'h3baeac82),
	.w3(32'h3b7b8adf),
	.w4(32'hb9ed4836),
	.w5(32'h3b92263c),
	.w6(32'h3b4737a0),
	.w7(32'h3ac16dde),
	.w8(32'h3b9ba3aa),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62979),
	.w1(32'h39ee2e35),
	.w2(32'h3a56ca98),
	.w3(32'hb92d9eff),
	.w4(32'h3a850ea0),
	.w5(32'h3acfbfbe),
	.w6(32'h3b47da03),
	.w7(32'h3b0d480b),
	.w8(32'h3ad7ad3c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba426a72),
	.w1(32'h39810c54),
	.w2(32'h383481e2),
	.w3(32'hba06a21a),
	.w4(32'h3a2452c9),
	.w5(32'h39c92b84),
	.w6(32'h389c37f5),
	.w7(32'h38161fa3),
	.w8(32'hba00a5e2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65dd7c),
	.w1(32'h3ac86579),
	.w2(32'h3a866721),
	.w3(32'h3a3f53c5),
	.w4(32'h3a63545e),
	.w5(32'h39d22eff),
	.w6(32'h3a89d2f1),
	.w7(32'h392028ec),
	.w8(32'hb97d1bb0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9083dbe),
	.w1(32'hba99d0c4),
	.w2(32'hba99eb9c),
	.w3(32'h3954c2b7),
	.w4(32'hba616703),
	.w5(32'hba55b755),
	.w6(32'hbb0f98fe),
	.w7(32'hbaf0d96a),
	.w8(32'hbb2451b6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73565a),
	.w1(32'h3b0c4b98),
	.w2(32'h3b9f4035),
	.w3(32'h3ae9960e),
	.w4(32'h3aa8ce37),
	.w5(32'h3b674291),
	.w6(32'h3bd14765),
	.w7(32'h3b3a897c),
	.w8(32'h3bae70c0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20f5b3),
	.w1(32'hbb1aa3c1),
	.w2(32'h3b16ae5a),
	.w3(32'h3bd3f0e5),
	.w4(32'hbbcdde18),
	.w5(32'hbadbe443),
	.w6(32'h3bafad8e),
	.w7(32'hbb85826c),
	.w8(32'hb88a1fb1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bade4be),
	.w1(32'hb90ff6cf),
	.w2(32'h3b8f780e),
	.w3(32'h3b0e3995),
	.w4(32'hbafba882),
	.w5(32'h3b185395),
	.w6(32'h3b896b97),
	.w7(32'hb91865fc),
	.w8(32'h3b8a34b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf7f84),
	.w1(32'hbabc0e75),
	.w2(32'hba5b7055),
	.w3(32'h3a578e86),
	.w4(32'hbad39df9),
	.w5(32'hba88e1cf),
	.w6(32'h3ab749e9),
	.w7(32'hb9915f0b),
	.w8(32'hb88853c0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa1b1f),
	.w1(32'hba4250d1),
	.w2(32'h3bba124a),
	.w3(32'h3b2d68d5),
	.w4(32'hbb622af6),
	.w5(32'h3b30ed73),
	.w6(32'h3b876b22),
	.w7(32'hb9a8e453),
	.w8(32'h3bb1159b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a1d6),
	.w1(32'hba554843),
	.w2(32'h3afc5ddd),
	.w3(32'h3b269ca6),
	.w4(32'hbad6736f),
	.w5(32'h39837701),
	.w6(32'h3a4f49a5),
	.w7(32'hba1d4b48),
	.w8(32'h39e0b401),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bbe5c),
	.w1(32'hb92ff7c6),
	.w2(32'h3bcb8849),
	.w3(32'h3c2c3749),
	.w4(32'hb9c1e0d9),
	.w5(32'h3bb30073),
	.w6(32'h3c0de876),
	.w7(32'h3abdb658),
	.w8(32'h3bb0e705),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba851160),
	.w1(32'h3b11139c),
	.w2(32'h3acb5816),
	.w3(32'hba532963),
	.w4(32'h3b03e6f0),
	.w5(32'h3aa3cfae),
	.w6(32'h3b119c01),
	.w7(32'h3ad75efb),
	.w8(32'h3abc91a0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f9b72),
	.w1(32'h392f3251),
	.w2(32'h3a3ddd27),
	.w3(32'h3ab69905),
	.w4(32'h39c671c1),
	.w5(32'h3a8457c3),
	.w6(32'h3898e275),
	.w7(32'h3992d02c),
	.w8(32'h3961bc23),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd805f),
	.w1(32'h3ad6ddd8),
	.w2(32'h3ba09229),
	.w3(32'h3bb0546c),
	.w4(32'h3a8c3dbd),
	.w5(32'h3bc5cdd0),
	.w6(32'h3c0dda56),
	.w7(32'h3aef2260),
	.w8(32'h3bd7e5b7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43a19),
	.w1(32'hbb37d198),
	.w2(32'h3ba52d6a),
	.w3(32'h3b98546a),
	.w4(32'hbb78cf54),
	.w5(32'h3ba23bba),
	.w6(32'h3b989955),
	.w7(32'hbaed8839),
	.w8(32'h3bae5afd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36c58),
	.w1(32'hbb02693e),
	.w2(32'h3b12f8ea),
	.w3(32'h3b7c82d9),
	.w4(32'hbbae07ba),
	.w5(32'hbaa36e94),
	.w6(32'h3b587193),
	.w7(32'hbb6d3ac0),
	.w8(32'h3a963b97),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839ce3),
	.w1(32'hbb1e75f4),
	.w2(32'hbb0874ec),
	.w3(32'h3a46d4ea),
	.w4(32'h38cad0f4),
	.w5(32'hbaca52f2),
	.w6(32'hbbc05ed4),
	.w7(32'hbb3c1d78),
	.w8(32'hba0bc0c7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514b55),
	.w1(32'hba5782a9),
	.w2(32'hba340a59),
	.w3(32'hbb3dd61e),
	.w4(32'hba210404),
	.w5(32'hba2f1031),
	.w6(32'hbaa67b7a),
	.w7(32'hba90cca1),
	.w8(32'hbae63440),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba002990),
	.w1(32'h3b490346),
	.w2(32'h3b34a1e5),
	.w3(32'hba321b0d),
	.w4(32'h3b2ebda2),
	.w5(32'h3b267fcf),
	.w6(32'h3b5c0ebf),
	.w7(32'h3b61366f),
	.w8(32'h3b3ab660),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b053d2c),
	.w1(32'h3a8b1646),
	.w2(32'h3b92b76a),
	.w3(32'h3ba71bf6),
	.w4(32'h3b9bb7e6),
	.w5(32'h3c0866d2),
	.w6(32'h3a34cef8),
	.w7(32'h3a9420b6),
	.w8(32'h3b90be86),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10c78a),
	.w1(32'h3bae4e54),
	.w2(32'h3bcd7725),
	.w3(32'h3bec8190),
	.w4(32'h3b9b2b0e),
	.w5(32'h3be73fc6),
	.w6(32'h3bef1a23),
	.w7(32'h3bbf80a0),
	.w8(32'h3ba67d93),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa16e1b),
	.w1(32'h3ac56a61),
	.w2(32'h3b33dffb),
	.w3(32'h3a6e5c22),
	.w4(32'h3b04880c),
	.w5(32'h3b55829c),
	.w6(32'h3af0625e),
	.w7(32'h3ab0f2b1),
	.w8(32'h3b7cb428),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada4e06),
	.w1(32'hbba9b361),
	.w2(32'hbb052df6),
	.w3(32'h3b1517c0),
	.w4(32'hbbb1a223),
	.w5(32'hbaf247d0),
	.w6(32'h3bb46cbf),
	.w7(32'hbb2c45e0),
	.w8(32'h3abfe199),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73ca5),
	.w1(32'hba2f2555),
	.w2(32'h3b9f84d5),
	.w3(32'h3b7c97e1),
	.w4(32'hbb8fd608),
	.w5(32'h3a390605),
	.w6(32'h3baac0aa),
	.w7(32'hbb3573c3),
	.w8(32'h3ab9992d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380e2352),
	.w1(32'h3a5b0383),
	.w2(32'h3a251915),
	.w3(32'h38a56aa2),
	.w4(32'h3a3ffce0),
	.w5(32'h3a2bf29a),
	.w6(32'h3a486d14),
	.w7(32'h3a195ed5),
	.w8(32'h3a3bb8c4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2209ee),
	.w1(32'h3b341c3b),
	.w2(32'h3b231f1d),
	.w3(32'h3a23c5a3),
	.w4(32'h3b54035b),
	.w5(32'h3b3c8ed0),
	.w6(32'h3b58c145),
	.w7(32'h3b432861),
	.w8(32'h3b57da15),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc1fd8),
	.w1(32'hba4a7b9c),
	.w2(32'hba8d6ac5),
	.w3(32'h3b15fb37),
	.w4(32'hb87d2145),
	.w5(32'hb95a9a3c),
	.w6(32'hb9e66cb5),
	.w7(32'h394a16fc),
	.w8(32'hb9961c34),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60ec4c),
	.w1(32'hbb30d83f),
	.w2(32'hbb60bd7c),
	.w3(32'hba2a4a15),
	.w4(32'hbb3d7d87),
	.w5(32'hbb5d74af),
	.w6(32'hbb1f308d),
	.w7(32'hbb22e5f9),
	.w8(32'hbb203845),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323589),
	.w1(32'h3b823545),
	.w2(32'h3b6daf44),
	.w3(32'hbb0db417),
	.w4(32'h3b7cee8b),
	.w5(32'h3b88be4a),
	.w6(32'h3b6d8608),
	.w7(32'h3b64c78a),
	.w8(32'h3b836b23),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea9096),
	.w1(32'h38e0d939),
	.w2(32'h3b785e02),
	.w3(32'h3b630deb),
	.w4(32'hbb43631e),
	.w5(32'h3b04c62b),
	.w6(32'h3ada4a52),
	.w7(32'hba5713aa),
	.w8(32'h3b88ea4c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f27f4),
	.w1(32'hb7be7b1e),
	.w2(32'h3b4f8131),
	.w3(32'h3b517188),
	.w4(32'hba3a231e),
	.w5(32'h3b44702a),
	.w6(32'h3b23c0b8),
	.w7(32'h3ac30bcb),
	.w8(32'h3b5ae524),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb886ba59),
	.w1(32'h3a80cb24),
	.w2(32'hb7cdb337),
	.w3(32'hb9c28d86),
	.w4(32'h3b06821e),
	.w5(32'h3aa4d216),
	.w6(32'h3afc5eee),
	.w7(32'h3a953bc7),
	.w8(32'h39bea9c6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ada4d),
	.w1(32'h3b201cd4),
	.w2(32'h3baff99b),
	.w3(32'h3b363578),
	.w4(32'h3b62531f),
	.w5(32'h3c054b67),
	.w6(32'h3b528daa),
	.w7(32'h3a6b8308),
	.w8(32'h3be80578),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade62b7),
	.w1(32'h3a855b8c),
	.w2(32'h3ae42999),
	.w3(32'h3ab36603),
	.w4(32'h3a63a06b),
	.w5(32'h3ad6afc1),
	.w6(32'h3b03663a),
	.w7(32'h3a98e670),
	.w8(32'h3ac9bf8d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb856748e),
	.w1(32'h39a6a26b),
	.w2(32'hb888b585),
	.w3(32'h3959e608),
	.w4(32'h3a0edbca),
	.w5(32'h39697fb6),
	.w6(32'h39193055),
	.w7(32'h397923a2),
	.w8(32'hb92de8c5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f1fa),
	.w1(32'h392de1df),
	.w2(32'h3ab665cd),
	.w3(32'h3aca9dab),
	.w4(32'h3a1ee009),
	.w5(32'h3acdeab2),
	.w6(32'h3a5f66fc),
	.w7(32'h3a6e8bf8),
	.w8(32'h3ac73d37),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27834b),
	.w1(32'h3a7d94ad),
	.w2(32'h3a5236ae),
	.w3(32'hb9fef3a4),
	.w4(32'h3a16ab47),
	.w5(32'h3a43d381),
	.w6(32'h3a84fb54),
	.w7(32'h3a458b6c),
	.w8(32'h3a218e70),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dc49d),
	.w1(32'hbab1374d),
	.w2(32'hbaad3b33),
	.w3(32'h3a883f48),
	.w4(32'hbab5db3e),
	.w5(32'hbaaa2fdf),
	.w6(32'hbab4912d),
	.w7(32'hbaddcbbc),
	.w8(32'hbb0b9ce2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18e2c0),
	.w1(32'hb8417320),
	.w2(32'hb8cb11a9),
	.w3(32'hbb14f0a0),
	.w4(32'h397f944d),
	.w5(32'h3976539b),
	.w6(32'h388d6cda),
	.w7(32'h38ad43a1),
	.w8(32'hb9d12520),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdfd0f),
	.w1(32'hbb21718f),
	.w2(32'hbb29ad2e),
	.w3(32'hb8ab231b),
	.w4(32'hbb271df8),
	.w5(32'hbb0e80a5),
	.w6(32'hbb3b053e),
	.w7(32'hbb46e097),
	.w8(32'hbb5a0297),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9fb92),
	.w1(32'hb9a9b72f),
	.w2(32'hb8be96d2),
	.w3(32'h38ae65c4),
	.w4(32'h388f06aa),
	.w5(32'h3a11d4c8),
	.w6(32'h3b7b8e96),
	.w7(32'h39c7402f),
	.w8(32'h3a8b0705),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b464ed0),
	.w1(32'hbac1814f),
	.w2(32'h3bdec006),
	.w3(32'h3b40ef01),
	.w4(32'hbb46e5b2),
	.w5(32'h3b28359b),
	.w6(32'h3a92accb),
	.w7(32'h38ad7d68),
	.w8(32'h3b949c86),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29e384),
	.w1(32'h3af81379),
	.w2(32'h3b848fe8),
	.w3(32'h3a1b356a),
	.w4(32'h39ae48a0),
	.w5(32'h3b2e3f4c),
	.w6(32'h3aa6a010),
	.w7(32'hba022da9),
	.w8(32'h3b2ba74e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7dead),
	.w1(32'h3b4c4ddc),
	.w2(32'h3bd927bc),
	.w3(32'h3bb9c9d0),
	.w4(32'h3b4f1e73),
	.w5(32'h3bb74bf0),
	.w6(32'h3b528da6),
	.w7(32'h3b87d1b7),
	.w8(32'h3be0cd59),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999d402),
	.w1(32'hbb6f4084),
	.w2(32'hbb51e622),
	.w3(32'h3a25e1c4),
	.w4(32'hbb70a8b3),
	.w5(32'hbb540e38),
	.w6(32'hbb64dce4),
	.w7(32'hbb72f35f),
	.w8(32'hbb89aa74),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f0268),
	.w1(32'h39ecf5e1),
	.w2(32'h390bfda1),
	.w3(32'hbb6e202e),
	.w4(32'h3a363c42),
	.w5(32'h39e3fe77),
	.w6(32'h395db41c),
	.w7(32'h39b17b25),
	.w8(32'hb9c0d264),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6eb60),
	.w1(32'hb93b7386),
	.w2(32'hb9b28425),
	.w3(32'hb4869133),
	.w4(32'h39b72d3c),
	.w5(32'h3920060a),
	.w6(32'hb8d4590a),
	.w7(32'hb923f06f),
	.w8(32'hb9de163f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011a12),
	.w1(32'hb8f5a631),
	.w2(32'hb9b1d541),
	.w3(32'hb9287dae),
	.w4(32'h39d1366f),
	.w5(32'h3947d03b),
	.w6(32'h3871dae8),
	.w7(32'hb7f3ad89),
	.w8(32'hb9141685),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38d89),
	.w1(32'h3b3f0352),
	.w2(32'h3bc127fc),
	.w3(32'h3b18e83d),
	.w4(32'h39245f6d),
	.w5(32'h3b452250),
	.w6(32'h3b91737b),
	.w7(32'h3ab66312),
	.w8(32'h3b8205c8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a951efb),
	.w1(32'h3a3c00b5),
	.w2(32'h387ebf7b),
	.w3(32'h39edb185),
	.w4(32'h39b5d557),
	.w5(32'h39be6c5f),
	.w6(32'h3a167f0a),
	.w7(32'h39ee1b85),
	.w8(32'h39ac5a0b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35eff6),
	.w1(32'hba98e76e),
	.w2(32'h392556fe),
	.w3(32'h3a984589),
	.w4(32'hb9e3dca1),
	.w5(32'h39854ae8),
	.w6(32'h3b1ed751),
	.w7(32'hb9f90d61),
	.w8(32'h3a4a0f2f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1399c7),
	.w1(32'h392c363c),
	.w2(32'h3a1b12dc),
	.w3(32'h3b160afa),
	.w4(32'h39931ddb),
	.w5(32'h39ace074),
	.w6(32'h3aebd788),
	.w7(32'hb98c157f),
	.w8(32'hb8957223),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d0c847),
	.w1(32'h393b4112),
	.w2(32'h38928cb7),
	.w3(32'h3a2e33ef),
	.w4(32'h3a028b26),
	.w5(32'h39d3e452),
	.w6(32'h38c73a8f),
	.w7(32'h37ed2f56),
	.w8(32'hb9ac02bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3f390),
	.w1(32'h3a997ed2),
	.w2(32'h3b385cc4),
	.w3(32'h3abcb5e9),
	.w4(32'h39c6ddff),
	.w5(32'h3ad504c5),
	.w6(32'h3ac4569d),
	.w7(32'h3ad83c12),
	.w8(32'h3b2c4507),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9ce1),
	.w1(32'h393ea9fd),
	.w2(32'hb8974060),
	.w3(32'h3a02934e),
	.w4(32'h3a0f0574),
	.w5(32'h39dcda98),
	.w6(32'h39d9a40e),
	.w7(32'h39a79ba2),
	.w8(32'h3a8a112a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a7694),
	.w1(32'h3b68ca6b),
	.w2(32'h3c02b3fc),
	.w3(32'h3bbe1e25),
	.w4(32'hba0a5085),
	.w5(32'hb9f00c69),
	.w6(32'h3b7099c5),
	.w7(32'h3a6667b6),
	.w8(32'h3aa63821),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeec25d),
	.w1(32'hb8128560),
	.w2(32'hb8a63952),
	.w3(32'hbae5da1e),
	.w4(32'hb8a1ba3a),
	.w5(32'hb8e97b2b),
	.w6(32'hb93b1075),
	.w7(32'hb792b5fc),
	.w8(32'hb83c578c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b3e06),
	.w1(32'hbb72058e),
	.w2(32'hbb688f5a),
	.w3(32'h3ad18655),
	.w4(32'hbb9282c4),
	.w5(32'hbb88e87e),
	.w6(32'h3bec89ed),
	.w7(32'hb9120a9c),
	.w8(32'hbb7de31f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule