module layer_10_featuremap_468(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09364e),
	.w1(32'hb942e9f4),
	.w2(32'hba257d95),
	.w3(32'hba4b1c31),
	.w4(32'h392343f7),
	.w5(32'h39c10f05),
	.w6(32'hba181a99),
	.w7(32'h3aa97794),
	.w8(32'h3a1829ce),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b0b9c),
	.w1(32'hba4d276d),
	.w2(32'hbac4a642),
	.w3(32'h3a652648),
	.w4(32'hba90e04f),
	.w5(32'hbaf2ba15),
	.w6(32'h3a853ff1),
	.w7(32'hba9f143c),
	.w8(32'hbac88102),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4a7c4),
	.w1(32'hb9335300),
	.w2(32'h3a11fdc7),
	.w3(32'hbaa4499e),
	.w4(32'hba2a1c1a),
	.w5(32'hba29253b),
	.w6(32'hbb087b3a),
	.w7(32'h399c9f63),
	.w8(32'h3998c9e7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a427972),
	.w1(32'hba9b2bcd),
	.w2(32'hbae4bf42),
	.w3(32'h389137e4),
	.w4(32'hbadd08ec),
	.w5(32'hba689301),
	.w6(32'hba8b21ef),
	.w7(32'hbab389e3),
	.w8(32'hbab84740),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0883f6),
	.w1(32'hb861b95d),
	.w2(32'hb9f831b2),
	.w3(32'hbaf80b4c),
	.w4(32'h38f67da7),
	.w5(32'hb8c5e2f4),
	.w6(32'hbaa2e7e9),
	.w7(32'h399aad95),
	.w8(32'hba2127c4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41ca24),
	.w1(32'h3b005c70),
	.w2(32'h3ac28ace),
	.w3(32'h3968808b),
	.w4(32'h3a0108c7),
	.w5(32'h39571592),
	.w6(32'hb8d42cf7),
	.w7(32'h3a6d9679),
	.w8(32'h3a419b83),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1f871),
	.w1(32'hba42f75b),
	.w2(32'hba5ecc3e),
	.w3(32'hba13e38b),
	.w4(32'hb9f2392f),
	.w5(32'hbaf6d761),
	.w6(32'hba11659a),
	.w7(32'hba7e231e),
	.w8(32'hba8c4c7f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59e84e),
	.w1(32'hb9d716ff),
	.w2(32'hbb0be895),
	.w3(32'hbaf4421d),
	.w4(32'hbaad1da1),
	.w5(32'hbab93045),
	.w6(32'hba4894b3),
	.w7(32'hb9888002),
	.w8(32'hb9e77ed3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852b1f),
	.w1(32'h39813342),
	.w2(32'h39ee40b9),
	.w3(32'hba3b8d99),
	.w4(32'hb9e7c527),
	.w5(32'hb9724638),
	.w6(32'hb9b19bbb),
	.w7(32'hb89183e1),
	.w8(32'hbacdc576),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a5a90),
	.w1(32'hba4aa9f9),
	.w2(32'hba5a6269),
	.w3(32'hba81c6b1),
	.w4(32'hba88af42),
	.w5(32'h3a2060ca),
	.w6(32'hbb1d91f8),
	.w7(32'hba41c77e),
	.w8(32'h39cee920),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a4484),
	.w1(32'hba91634c),
	.w2(32'hb8bffab6),
	.w3(32'h3a3ed41f),
	.w4(32'hba125d2c),
	.w5(32'hb927cf69),
	.w6(32'h39cbba96),
	.w7(32'h3a0fda28),
	.w8(32'hb82489ff),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996e702),
	.w1(32'h3a2edd4c),
	.w2(32'h384b0935),
	.w3(32'h3a4fd87f),
	.w4(32'h3841d257),
	.w5(32'hb8947217),
	.w6(32'h3a61d04f),
	.w7(32'h39aed216),
	.w8(32'h39beb771),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9071795),
	.w1(32'hbae00ad2),
	.w2(32'hbb219621),
	.w3(32'h3994563b),
	.w4(32'hbb18e91b),
	.w5(32'hba580944),
	.w6(32'h3ad1d584),
	.w7(32'hbb2eda1c),
	.w8(32'hba91e037),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e2699),
	.w1(32'hba9d5874),
	.w2(32'h3880066a),
	.w3(32'hbafc39c6),
	.w4(32'hbaaef670),
	.w5(32'hba3d061a),
	.w6(32'hba773fd1),
	.w7(32'hb891cfeb),
	.w8(32'hba455d68),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aef050),
	.w1(32'hb874e59f),
	.w2(32'h3995ff2c),
	.w3(32'hb96ff10d),
	.w4(32'h3a2e2996),
	.w5(32'hb9b3d1f1),
	.w6(32'hb9f78e20),
	.w7(32'h3a92a958),
	.w8(32'h3a85080f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67fa70f),
	.w1(32'hb8f6232d),
	.w2(32'hba588609),
	.w3(32'hb9d974a1),
	.w4(32'h39102775),
	.w5(32'hba4541a7),
	.w6(32'h39faa408),
	.w7(32'h3a2bdc5e),
	.w8(32'hb9037ed5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8b430),
	.w1(32'hba916917),
	.w2(32'hba9b283d),
	.w3(32'hba96bb48),
	.w4(32'hb8217c95),
	.w5(32'hb9c97484),
	.w6(32'hb8100d18),
	.w7(32'hb7531587),
	.w8(32'h3a4666ff),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad043a),
	.w1(32'hb9a1eced),
	.w2(32'hbaafff1d),
	.w3(32'hba3b8101),
	.w4(32'hbab2a240),
	.w5(32'hba88d6d8),
	.w6(32'hb97c0e7e),
	.w7(32'hba7c5a14),
	.w8(32'hbaa9264e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba828f82),
	.w1(32'hbab5b30e),
	.w2(32'hba807b0d),
	.w3(32'hba1e38b8),
	.w4(32'hbaaf1aa5),
	.w5(32'hb8fe30af),
	.w6(32'hb927749d),
	.w7(32'hba4a86cd),
	.w8(32'h376d10d5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38915e47),
	.w1(32'h3b0aefea),
	.w2(32'h3aa86d6c),
	.w3(32'hb81c1691),
	.w4(32'h3abb81cc),
	.w5(32'h3b086342),
	.w6(32'h38b0287e),
	.w7(32'hb8b81c16),
	.w8(32'h3a2c6e3d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ed6f),
	.w1(32'h3819c589),
	.w2(32'hb98b61b0),
	.w3(32'h3a95819f),
	.w4(32'hba4810c5),
	.w5(32'hba384766),
	.w6(32'h3aa5264f),
	.w7(32'hba7e3e64),
	.w8(32'hbac2c262),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75757a),
	.w1(32'h3aa32e32),
	.w2(32'h3b210262),
	.w3(32'hbb065513),
	.w4(32'h39976082),
	.w5(32'h3ae74d7b),
	.w6(32'hbac5b413),
	.w7(32'h39874dcc),
	.w8(32'h3a885acc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294a46),
	.w1(32'h3a17e177),
	.w2(32'h3ad2731a),
	.w3(32'h3ae1904f),
	.w4(32'hb9c3d97e),
	.w5(32'h3ab13b6c),
	.w6(32'h3ada5522),
	.w7(32'hba5fbdea),
	.w8(32'h39866a7b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8198679),
	.w1(32'h399d5143),
	.w2(32'hbb12cbe7),
	.w3(32'h3a9e4e3a),
	.w4(32'hbb313cd1),
	.w5(32'hbb644949),
	.w6(32'hb9d436dd),
	.w7(32'hbb0f47e0),
	.w8(32'hbb4da906),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8feab2b),
	.w1(32'h38fd6437),
	.w2(32'h3aa9e5df),
	.w3(32'hbb1e5693),
	.w4(32'hb8e17c3a),
	.w5(32'hba68a133),
	.w6(32'hbaadc98b),
	.w7(32'hb9516df0),
	.w8(32'hba37d634),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26ae71),
	.w1(32'h3b17065b),
	.w2(32'h3aef91a9),
	.w3(32'h39b0538e),
	.w4(32'h3a51ae88),
	.w5(32'h3a7dcef7),
	.w6(32'hb9a9e24a),
	.w7(32'hba26d98f),
	.w8(32'h3906216f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00fb59),
	.w1(32'hbabe1981),
	.w2(32'hb6c590ad),
	.w3(32'h3afac984),
	.w4(32'h3a89a182),
	.w5(32'hba001bf2),
	.w6(32'h3a9a3a6c),
	.w7(32'h3a15eff3),
	.w8(32'hba542128),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de9273),
	.w1(32'hb983c78a),
	.w2(32'hbab9e162),
	.w3(32'hba8342ba),
	.w4(32'hb9dc2bcf),
	.w5(32'hbaa80a02),
	.w6(32'hba9abc1f),
	.w7(32'hba0b95af),
	.w8(32'hba512b5d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e3f10),
	.w1(32'hb89c457d),
	.w2(32'h3a4b044f),
	.w3(32'hb9c399ed),
	.w4(32'h3a985933),
	.w5(32'h3aafcd54),
	.w6(32'hba0161c1),
	.w7(32'h3a8025e1),
	.w8(32'h3a40b6e6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e8152),
	.w1(32'hb7e459ff),
	.w2(32'h391f5a5a),
	.w3(32'h3ac39448),
	.w4(32'hba2278dc),
	.w5(32'hb9a305bd),
	.w6(32'h399129af),
	.w7(32'hba01f137),
	.w8(32'hb9af8e75),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9803ddb),
	.w1(32'h3a921965),
	.w2(32'h38947c67),
	.w3(32'hba85052f),
	.w4(32'h3b2a0f21),
	.w5(32'h3afc8250),
	.w6(32'hba59d916),
	.w7(32'h3adb8880),
	.w8(32'h3accc243),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395aebd8),
	.w1(32'h3a484d80),
	.w2(32'h3a89b692),
	.w3(32'h397e50ed),
	.w4(32'h39744247),
	.w5(32'h3a7ea497),
	.w6(32'h3a89fbf7),
	.w7(32'h359c6798),
	.w8(32'h39ac65de),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f0e30),
	.w1(32'hb8d1153a),
	.w2(32'h3a436724),
	.w3(32'h3a1c1d91),
	.w4(32'h37301d34),
	.w5(32'h39ec9d5b),
	.w6(32'hba947183),
	.w7(32'hba4a3458),
	.w8(32'hb96fb61d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c07a0),
	.w1(32'hb9e7f2a7),
	.w2(32'hba2a5ae7),
	.w3(32'h390d4299),
	.w4(32'hb84cedc0),
	.w5(32'h39debf56),
	.w6(32'hb9d3ec0a),
	.w7(32'hb9dda0bd),
	.w8(32'h3aafb794),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f154e3),
	.w1(32'h3aabe810),
	.w2(32'hba2fa74c),
	.w3(32'h39df5f85),
	.w4(32'hba8501d9),
	.w5(32'hbae98122),
	.w6(32'h3a3cf857),
	.w7(32'hba4299e1),
	.w8(32'hbb0beed9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256dde),
	.w1(32'h3a7942e8),
	.w2(32'h3a57919b),
	.w3(32'hba51dc85),
	.w4(32'h39a0b224),
	.w5(32'hb95fc168),
	.w6(32'hba08395e),
	.w7(32'hb86ee696),
	.w8(32'hba172183),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb814ce36),
	.w1(32'hbb329e03),
	.w2(32'hb96cb228),
	.w3(32'hb9d46496),
	.w4(32'hb986b5ec),
	.w5(32'hba6135b7),
	.w6(32'hba0d0813),
	.w7(32'h3a74d5ff),
	.w8(32'h397257ad),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c2f8d),
	.w1(32'h3a2284c5),
	.w2(32'hba5c1336),
	.w3(32'h3aa9d84a),
	.w4(32'h3a1fa87a),
	.w5(32'hba97844c),
	.w6(32'h39fe9683),
	.w7(32'h385d08da),
	.w8(32'hba3adc07),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf20e99),
	.w1(32'hbb1be6b8),
	.w2(32'hbadc36b4),
	.w3(32'hbb1f904d),
	.w4(32'hbb26697f),
	.w5(32'hbb64d391),
	.w6(32'hbb3f9cf7),
	.w7(32'hb96869b6),
	.w8(32'hba985ce4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb759337c),
	.w1(32'h39d2907d),
	.w2(32'hb8e04e61),
	.w3(32'hba35fe91),
	.w4(32'hb8e7fdd5),
	.w5(32'h3a25dd28),
	.w6(32'hba088963),
	.w7(32'hba3f6a15),
	.w8(32'hba0f1183),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4f907),
	.w1(32'hbaecd7e9),
	.w2(32'hbb0c33c2),
	.w3(32'h3a6bc34b),
	.w4(32'hbaa4c5a3),
	.w5(32'hbb0d2536),
	.w6(32'hb9b5fc9d),
	.w7(32'hbb04df33),
	.w8(32'hbb066009),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43f88b),
	.w1(32'hb9078951),
	.w2(32'hb8c013e1),
	.w3(32'hba87ab0d),
	.w4(32'hb92d83ba),
	.w5(32'hba280fc6),
	.w6(32'hba075f5b),
	.w7(32'h379cb615),
	.w8(32'h39435a3a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265e1a),
	.w1(32'h376d268f),
	.w2(32'hb994c5a2),
	.w3(32'h393347b9),
	.w4(32'hba88e541),
	.w5(32'h374d7a2c),
	.w6(32'h39d185c9),
	.w7(32'hbacb328d),
	.w8(32'hbaa17a5c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3580f),
	.w1(32'h3a10c828),
	.w2(32'hb9bf3976),
	.w3(32'hbb025072),
	.w4(32'h38868bac),
	.w5(32'hbac7e596),
	.w6(32'hbae64f74),
	.w7(32'h3997e8ab),
	.w8(32'hba95ca7f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9577f7),
	.w1(32'h398b6387),
	.w2(32'hb69f27e8),
	.w3(32'h3a31df8e),
	.w4(32'h394c32e6),
	.w5(32'h3a586d83),
	.w6(32'h3a1bf72f),
	.w7(32'h385d3ed1),
	.w8(32'hb8c6fe0a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3864fbb2),
	.w1(32'hba6ccdde),
	.w2(32'hbb1cefeb),
	.w3(32'h38181a34),
	.w4(32'hba327f86),
	.w5(32'hbb1b62bf),
	.w6(32'hb96eb02d),
	.w7(32'h3876ca14),
	.w8(32'hba6da99d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba888d1d),
	.w1(32'h3a703344),
	.w2(32'hb8d2d246),
	.w3(32'hbb0aa486),
	.w4(32'hba0fe094),
	.w5(32'hbab537b6),
	.w6(32'hba7fffd4),
	.w7(32'hba4885f6),
	.w8(32'hbad2e94d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111765),
	.w1(32'hbb60cce3),
	.w2(32'hbb2e52d6),
	.w3(32'hba9b1317),
	.w4(32'hbb430636),
	.w5(32'hbb164de6),
	.w6(32'hbaa32822),
	.w7(32'hbabb55c9),
	.w8(32'hbaa9b24f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba936c39),
	.w1(32'h3a98f45c),
	.w2(32'h3aaaf895),
	.w3(32'hb9ba0769),
	.w4(32'hbaa14638),
	.w5(32'hba70c7a7),
	.w6(32'hb995e832),
	.w7(32'hb9cb4184),
	.w8(32'hba26e91b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d11b6),
	.w1(32'h3b5289c7),
	.w2(32'h3aee7b03),
	.w3(32'hba6fb12b),
	.w4(32'h3b06ccf5),
	.w5(32'h3a4b2d03),
	.w6(32'h39c43710),
	.w7(32'h3ac39afc),
	.w8(32'h3aa52b8e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcb050),
	.w1(32'hb9d9be55),
	.w2(32'hbaf31a89),
	.w3(32'h39d84931),
	.w4(32'hbaccac8a),
	.w5(32'hba4c6411),
	.w6(32'h3b0ad0e8),
	.w7(32'hbadfb329),
	.w8(32'hbaae0228),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6d935),
	.w1(32'hba7651e8),
	.w2(32'hba52c299),
	.w3(32'hbacca5bb),
	.w4(32'h39a1f225),
	.w5(32'hbad1c993),
	.w6(32'hb9afa380),
	.w7(32'hb9eb39e0),
	.w8(32'hbac0347f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c73b10),
	.w1(32'h3a22e742),
	.w2(32'hb9c5242c),
	.w3(32'hba5f79dc),
	.w4(32'hba7e956a),
	.w5(32'hba1a384b),
	.w6(32'hbac66cf1),
	.w7(32'hba35c1bf),
	.w8(32'hba777926),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e78e0),
	.w1(32'h3a793025),
	.w2(32'h39b9c8dc),
	.w3(32'hb86fb918),
	.w4(32'h3a5f4ada),
	.w5(32'h3a9400a2),
	.w6(32'hb829c753),
	.w7(32'hba4f5473),
	.w8(32'hba3943c8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bfb6b),
	.w1(32'hbac61d0b),
	.w2(32'hbb03a317),
	.w3(32'h3a9c9530),
	.w4(32'hbaef1ab0),
	.w5(32'hbab9e371),
	.w6(32'hb9dfe4b2),
	.w7(32'hbaff70cc),
	.w8(32'hbaaf16d0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd0af2),
	.w1(32'h39809181),
	.w2(32'hb9e5eb31),
	.w3(32'hbaf8ff1b),
	.w4(32'h39b99642),
	.w5(32'h3a10b322),
	.w6(32'hbb4bcb49),
	.w7(32'h39bd08c4),
	.w8(32'h3980a544),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fb90f),
	.w1(32'hba9c3bcb),
	.w2(32'hbb400e99),
	.w3(32'hb9a4bb70),
	.w4(32'h3a1d3b4c),
	.w5(32'hba44ecea),
	.w6(32'hba055f3d),
	.w7(32'h3a5ea5fb),
	.w8(32'h3934ec1e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2f33),
	.w1(32'h37edec70),
	.w2(32'h3985b4df),
	.w3(32'hbac7792f),
	.w4(32'hb9413319),
	.w5(32'hba66e5b4),
	.w6(32'hb95a2cee),
	.w7(32'hba8655c9),
	.w8(32'hba96e54b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a3580),
	.w1(32'hb9060d0b),
	.w2(32'hbab9ca09),
	.w3(32'hb953a601),
	.w4(32'h3a0b7ee7),
	.w5(32'hba86dd5a),
	.w6(32'hbac6142a),
	.w7(32'h3a4d6ed5),
	.w8(32'hb9b2992e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9e1fe),
	.w1(32'hb79aa421),
	.w2(32'h3a6bce79),
	.w3(32'hbaa20fde),
	.w4(32'h3a5fed67),
	.w5(32'hbab46de2),
	.w6(32'hbad46ceb),
	.w7(32'hba78a9ac),
	.w8(32'hbaa90974),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37637a60),
	.w1(32'hba497a8b),
	.w2(32'hba1c18a7),
	.w3(32'h39eae8c1),
	.w4(32'h393dc453),
	.w5(32'h3aa63681),
	.w6(32'hb907cb91),
	.w7(32'h397300c5),
	.w8(32'hb9594569),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d6c70),
	.w1(32'hb7f81282),
	.w2(32'h392149e3),
	.w3(32'h39b855cd),
	.w4(32'hb9b1aa2d),
	.w5(32'hba2c0acc),
	.w6(32'h38fd678c),
	.w7(32'hb93afd66),
	.w8(32'hb9ca518d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9f8ec),
	.w1(32'hba6bf674),
	.w2(32'hbb0e9c7b),
	.w3(32'h39a4d413),
	.w4(32'hbaf7735d),
	.w5(32'hbb3b16f6),
	.w6(32'hb97d7137),
	.w7(32'hbb13e9f5),
	.w8(32'hbb732aab),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe30ab),
	.w1(32'hba9ce32d),
	.w2(32'hbae86672),
	.w3(32'hbb0e1b21),
	.w4(32'hba020417),
	.w5(32'hb97f87f9),
	.w6(32'hbb0d3aa4),
	.w7(32'hb95daee7),
	.w8(32'hb969134f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1da0),
	.w1(32'h3b629968),
	.w2(32'h3b00b4e3),
	.w3(32'hba8909c3),
	.w4(32'h3b189dbd),
	.w5(32'h3b0ffcfd),
	.w6(32'h398b2ff7),
	.w7(32'h3b208986),
	.w8(32'h3ab59a94),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05810a),
	.w1(32'h3a0926d3),
	.w2(32'h38832f0f),
	.w3(32'h3acf10c5),
	.w4(32'h35d44f4d),
	.w5(32'hba743bde),
	.w6(32'h3b18e08d),
	.w7(32'h39cc3a1a),
	.w8(32'h3a061ad2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16fb38),
	.w1(32'hba6f8820),
	.w2(32'hbac3215b),
	.w3(32'h398a9a3d),
	.w4(32'hbadc0554),
	.w5(32'hb890510e),
	.w6(32'h3a1c37cf),
	.w7(32'hbabc98a0),
	.w8(32'hb90b5e1d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4efa8),
	.w1(32'hba46008c),
	.w2(32'hbb2d9bb7),
	.w3(32'hb9fab416),
	.w4(32'hbaf84a86),
	.w5(32'hbb43d71f),
	.w6(32'hb91005bb),
	.w7(32'hba98f8f6),
	.w8(32'hbae72c2e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28005c),
	.w1(32'hbab0e72e),
	.w2(32'h39c69d15),
	.w3(32'hbb4864d6),
	.w4(32'hbab4a185),
	.w5(32'hb8032fa6),
	.w6(32'hba9244df),
	.w7(32'h38b18fc9),
	.w8(32'h3a426349),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adeb6bc),
	.w1(32'hbb3b6871),
	.w2(32'hbac8eccb),
	.w3(32'h3b2d2d8a),
	.w4(32'h38a2c70b),
	.w5(32'hbb353aa7),
	.w6(32'h3b2d5679),
	.w7(32'h3a669a6d),
	.w8(32'h3b0e9b79),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104f0a),
	.w1(32'hbc08e6df),
	.w2(32'hbba9ae63),
	.w3(32'hbc0c498a),
	.w4(32'hbc451c9d),
	.w5(32'h3b65c9c6),
	.w6(32'hbb1680d2),
	.w7(32'hbb9877f7),
	.w8(32'h3ba76948),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11ca97),
	.w1(32'h3a5b3b1b),
	.w2(32'h3ba992c7),
	.w3(32'h3aad4089),
	.w4(32'h3ae18a78),
	.w5(32'h3c196b1c),
	.w6(32'h3ac5ebf5),
	.w7(32'hb98512bf),
	.w8(32'hba356f7e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b006e7e),
	.w1(32'hbba0dc8f),
	.w2(32'h3b10c336),
	.w3(32'hb70d925e),
	.w4(32'h39d7d292),
	.w5(32'h3c7e0d78),
	.w6(32'hbb1f2772),
	.w7(32'h3b56f3fc),
	.w8(32'h3b6f85a0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68e0f2),
	.w1(32'h38d3ca4d),
	.w2(32'h3b2bce74),
	.w3(32'h3bc44792),
	.w4(32'h3b4f6bda),
	.w5(32'h3bce5b43),
	.w6(32'h3bb82384),
	.w7(32'h3b11c866),
	.w8(32'h3b0feb2d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06941c),
	.w1(32'hbb8bb54c),
	.w2(32'hbb5421db),
	.w3(32'hbaa69bb2),
	.w4(32'h3b2f762a),
	.w5(32'hbbf1cb59),
	.w6(32'h3aa334d7),
	.w7(32'h39113e51),
	.w8(32'hbaa4c269),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7d726),
	.w1(32'h3b83c597),
	.w2(32'h3bd33813),
	.w3(32'h3b8e7420),
	.w4(32'h3b452005),
	.w5(32'h3bed20a8),
	.w6(32'h3b0e1b89),
	.w7(32'hb9fa1d8a),
	.w8(32'hba9f5878),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b9a3),
	.w1(32'hbc22161f),
	.w2(32'hbbf8d004),
	.w3(32'h3b600fe9),
	.w4(32'hbba48565),
	.w5(32'h3c2ea671),
	.w6(32'hb9909b8c),
	.w7(32'hbc1d53ac),
	.w8(32'hbbb2d311),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2861b5),
	.w1(32'hbaf0db51),
	.w2(32'hba74f56d),
	.w3(32'hbc0cb5ed),
	.w4(32'hbbb7423a),
	.w5(32'h3a8a9417),
	.w6(32'hbbf30a5c),
	.w7(32'hbc01bfe8),
	.w8(32'hbb994454),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b496b0a),
	.w1(32'h3b07aefa),
	.w2(32'h3b56e7d3),
	.w3(32'hbb407005),
	.w4(32'h3bf3b209),
	.w5(32'h3bec592d),
	.w6(32'hbb6e88a5),
	.w7(32'h3b17d97b),
	.w8(32'h3af683cc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c837d),
	.w1(32'hbb5e66ee),
	.w2(32'hbbcccd97),
	.w3(32'h3b593433),
	.w4(32'hbc234af5),
	.w5(32'hbaacffd7),
	.w6(32'h3a0ee89f),
	.w7(32'hbbb20629),
	.w8(32'hbb1db6fa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d05a3),
	.w1(32'h39f7902f),
	.w2(32'h3b59c814),
	.w3(32'hbbf8776b),
	.w4(32'h3bfb0efc),
	.w5(32'h3bbdf92e),
	.w6(32'h3983c5df),
	.w7(32'hbb1f9125),
	.w8(32'h3a1031c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6939e),
	.w1(32'hbaae164d),
	.w2(32'hbb17c1ec),
	.w3(32'hbbb0cf56),
	.w4(32'hbb8daa3b),
	.w5(32'h3a013c91),
	.w6(32'hbbd6cc2d),
	.w7(32'hbb127718),
	.w8(32'hb9b26f38),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bfc68),
	.w1(32'hbafe3225),
	.w2(32'hbb290529),
	.w3(32'h3ba76112),
	.w4(32'hbb33f025),
	.w5(32'hbbe8943f),
	.w6(32'hba555f45),
	.w7(32'hbac1403d),
	.w8(32'h39ff9772),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1c6d3),
	.w1(32'h3a7cc51f),
	.w2(32'h39bfd252),
	.w3(32'h3a95eca9),
	.w4(32'hbab65a7f),
	.w5(32'h3c0484e9),
	.w6(32'hba838d7e),
	.w7(32'h3bec6771),
	.w8(32'h3bfd7199),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed2db8),
	.w1(32'h3b10e424),
	.w2(32'h3bb01fda),
	.w3(32'h3ac3137a),
	.w4(32'hb9712aee),
	.w5(32'h3c7bf2eb),
	.w6(32'h3ab854a7),
	.w7(32'hba82d68f),
	.w8(32'h3b456e98),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc77865),
	.w1(32'h3c202e11),
	.w2(32'h3b8764ae),
	.w3(32'h3bdf211a),
	.w4(32'h3c5f70a7),
	.w5(32'h3bf72bdb),
	.w6(32'h39976ee7),
	.w7(32'h3cae2a5f),
	.w8(32'h3c50b4f2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc265bd),
	.w1(32'hbb413468),
	.w2(32'h3b89b061),
	.w3(32'h3c4df5bd),
	.w4(32'h3bb0a76b),
	.w5(32'hb88846f4),
	.w6(32'h3be5c879),
	.w7(32'h3b90821e),
	.w8(32'h3bd7be8c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257d91),
	.w1(32'hbb9a35da),
	.w2(32'h3adb8bd3),
	.w3(32'hbaa04e15),
	.w4(32'hbafed93f),
	.w5(32'hbb846cf3),
	.w6(32'h3b1dc2ad),
	.w7(32'hba563f3b),
	.w8(32'h3be98210),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1296d),
	.w1(32'hbbb4b5c2),
	.w2(32'hbbe9dd71),
	.w3(32'hbb8badd0),
	.w4(32'hbb88d1be),
	.w5(32'hba5bd3d6),
	.w6(32'h3ba842e0),
	.w7(32'hbb71927f),
	.w8(32'hbbc31005),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb214431),
	.w1(32'h3c3358f0),
	.w2(32'h3b78ebd6),
	.w3(32'hbc0045f7),
	.w4(32'h3c114979),
	.w5(32'hbb6ce9bf),
	.w6(32'hbbab1bd5),
	.w7(32'h3bb5068c),
	.w8(32'h3b4d815c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba214f0),
	.w1(32'h3b807ecd),
	.w2(32'h3ba17d6d),
	.w3(32'h3c00a307),
	.w4(32'hbb3e5290),
	.w5(32'h3bbdf0fa),
	.w6(32'h3ae34c3b),
	.w7(32'h3aef8aa6),
	.w8(32'h3ba852de),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f6709),
	.w1(32'h3a71c441),
	.w2(32'h3a7c47f2),
	.w3(32'hbb5365d8),
	.w4(32'h3b8eab9a),
	.w5(32'hbb63a591),
	.w6(32'hbabeac26),
	.w7(32'h3befcb1d),
	.w8(32'h3b588b8b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df310),
	.w1(32'h3b12a6ff),
	.w2(32'h3a2b7ae2),
	.w3(32'h3b7a70a4),
	.w4(32'h3bb6d401),
	.w5(32'hbb55b052),
	.w6(32'h3ae85544),
	.w7(32'h3c06094e),
	.w8(32'h3ba05fe4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1c3b5),
	.w1(32'h3ae16397),
	.w2(32'h3bb2751b),
	.w3(32'hbb7cfd24),
	.w4(32'h3b0f35b9),
	.w5(32'h3b6419ba),
	.w6(32'hbb0dab52),
	.w7(32'h3b535301),
	.w8(32'h3b4ac551),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37f424),
	.w1(32'hbb70f009),
	.w2(32'hbb65d325),
	.w3(32'hba997437),
	.w4(32'hbbf815f5),
	.w5(32'hbbb3bb0c),
	.w6(32'h3b4efea6),
	.w7(32'h3b1bb87f),
	.w8(32'h3b96bd89),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27af56),
	.w1(32'hbbd3191a),
	.w2(32'hbbab406c),
	.w3(32'hbbbe12c9),
	.w4(32'hbbb4ae42),
	.w5(32'h3ba222ed),
	.w6(32'h396aa8b7),
	.w7(32'hbafc9d1b),
	.w8(32'hbbaa1a57),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9645a5),
	.w1(32'hbb1a7113),
	.w2(32'hbb94c575),
	.w3(32'hbc3501fb),
	.w4(32'hbab7d87e),
	.w5(32'h3b9548f7),
	.w6(32'hbbb9bede),
	.w7(32'h3ae12dcb),
	.w8(32'h3bc161d5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b2ffe),
	.w1(32'h3c21c406),
	.w2(32'h3bb70860),
	.w3(32'hb7d3cbdb),
	.w4(32'h3c24983f),
	.w5(32'hbaa23a21),
	.w6(32'hbb8181e5),
	.w7(32'h3c1208bc),
	.w8(32'h3bcd8b5a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096836),
	.w1(32'h3ad78418),
	.w2(32'h3a401a1f),
	.w3(32'h3c118260),
	.w4(32'hbaa8cc1f),
	.w5(32'h3b9cc3b1),
	.w6(32'h3c40b850),
	.w7(32'h3b481c0e),
	.w8(32'hb9cc7711),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eec86),
	.w1(32'h3b32ec8f),
	.w2(32'hb7edcfc6),
	.w3(32'h3ba2b408),
	.w4(32'h3c12fb4f),
	.w5(32'h3a044521),
	.w6(32'h3bd0b482),
	.w7(32'h3b514413),
	.w8(32'hbac35f94),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba190937),
	.w1(32'h39f62d9e),
	.w2(32'hbab353dd),
	.w3(32'h3bb00133),
	.w4(32'h3aa27b0e),
	.w5(32'h3b0fe265),
	.w6(32'h3a14c3a8),
	.w7(32'h3bf8d6b5),
	.w8(32'h3c29190b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01edb5),
	.w1(32'h39755084),
	.w2(32'hb9d93f62),
	.w3(32'hba3cc2c0),
	.w4(32'hba99eeec),
	.w5(32'h3b1bfeb2),
	.w6(32'h3bcc7a72),
	.w7(32'h3a67f2ea),
	.w8(32'h3b2cb612),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29744e),
	.w1(32'hbbb45c51),
	.w2(32'hbb42cb48),
	.w3(32'h3b99b1e4),
	.w4(32'hbb89033a),
	.w5(32'hb91e3307),
	.w6(32'h3a578318),
	.w7(32'hbb97f279),
	.w8(32'hba6ab171),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb15aa5),
	.w1(32'hbb41fbef),
	.w2(32'hbb4b6671),
	.w3(32'hbb949891),
	.w4(32'hbb639370),
	.w5(32'h3a9c6db4),
	.w6(32'hbbeeee38),
	.w7(32'hbbe33e1f),
	.w8(32'h3bb47f35),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e32d5),
	.w1(32'hbc3c19b0),
	.w2(32'hbc094c92),
	.w3(32'h3b08c709),
	.w4(32'hbb866071),
	.w5(32'hbbfd3214),
	.w6(32'hb7b4d36d),
	.w7(32'hbbef160c),
	.w8(32'hbc2f3d76),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf888b4),
	.w1(32'h3b4ac02e),
	.w2(32'hb9e909ce),
	.w3(32'hbbbbe540),
	.w4(32'h3b74ed9b),
	.w5(32'h3b92b970),
	.w6(32'hbba7eba1),
	.w7(32'h3b831feb),
	.w8(32'hb87e5b3b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a576cd1),
	.w1(32'h3b8c9ed6),
	.w2(32'hb9dfe86e),
	.w3(32'h3b808a01),
	.w4(32'hbbd504e6),
	.w5(32'hbb61aa3c),
	.w6(32'h3af510af),
	.w7(32'hbba5ca78),
	.w8(32'h3aa1536a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ce2d),
	.w1(32'h3a989f78),
	.w2(32'hbc009dce),
	.w3(32'h3bd9b3a2),
	.w4(32'hbad8ba6e),
	.w5(32'hbbd5b239),
	.w6(32'h3b7132c2),
	.w7(32'hba54bcff),
	.w8(32'hbadaf061),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab8c0d),
	.w1(32'h3bb5b021),
	.w2(32'hba47a609),
	.w3(32'hbc512be7),
	.w4(32'h3c3ab738),
	.w5(32'h3bbda52b),
	.w6(32'hbb533dc5),
	.w7(32'h3bbdb7b2),
	.w8(32'h3b0afa7b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c1de),
	.w1(32'hbba43717),
	.w2(32'hbba5ff86),
	.w3(32'h3c1ae0a6),
	.w4(32'hbb8458f0),
	.w5(32'hb8c10b4e),
	.w6(32'h3a92a593),
	.w7(32'hbb6faca2),
	.w8(32'h3a4996d8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d93e9),
	.w1(32'h3b8fe2d2),
	.w2(32'hbb137243),
	.w3(32'hbba9cb7b),
	.w4(32'h3a7d6a94),
	.w5(32'hbb053887),
	.w6(32'hbb343606),
	.w7(32'h3937c243),
	.w8(32'h3af67156),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43029),
	.w1(32'h3b299ac8),
	.w2(32'h3a05e2ee),
	.w3(32'hbb0d9ca6),
	.w4(32'h3b00165d),
	.w5(32'h3aff26ff),
	.w6(32'h3b709ff6),
	.w7(32'h3abbeba3),
	.w8(32'hba7a8dba),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb352d),
	.w1(32'h3bf73409),
	.w2(32'h3b91e4ce),
	.w3(32'hbb2b6d1e),
	.w4(32'h3c1fc2e5),
	.w5(32'hba5d3d18),
	.w6(32'hbb657633),
	.w7(32'h3bb843d0),
	.w8(32'h3a1153fd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88268f),
	.w1(32'hbb18c543),
	.w2(32'h3a494b59),
	.w3(32'h3ab5f198),
	.w4(32'hbb997d9f),
	.w5(32'h3bcb2b51),
	.w6(32'h3bf7273e),
	.w7(32'hbb1b65ed),
	.w8(32'h3b840ef4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c29a),
	.w1(32'h3c51b505),
	.w2(32'h3c23cb34),
	.w3(32'h3ab4d7a1),
	.w4(32'h3c902aac),
	.w5(32'hbc66e6da),
	.w6(32'h3b3c9cad),
	.w7(32'h3c7635ee),
	.w8(32'h3baad879),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48d5af),
	.w1(32'hbba731a2),
	.w2(32'hbab51c16),
	.w3(32'h3b5e90f2),
	.w4(32'hbb088b01),
	.w5(32'h3bdc3047),
	.w6(32'h3c576864),
	.w7(32'hbba27afe),
	.w8(32'hb97101c8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8189),
	.w1(32'h3bd830e7),
	.w2(32'h3c3f39f0),
	.w3(32'h3acf95bf),
	.w4(32'h3b9e02ee),
	.w5(32'h3b7adf4b),
	.w6(32'h3b534c51),
	.w7(32'h3c0b067d),
	.w8(32'h3bd89a3c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fe358),
	.w1(32'h3aadc7b6),
	.w2(32'h3b1ba914),
	.w3(32'h3c109afa),
	.w4(32'hbb71f7c0),
	.w5(32'hbb76a785),
	.w6(32'h3c1c9936),
	.w7(32'hbaca6971),
	.w8(32'hbb3cc496),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba28784),
	.w1(32'hbb837fea),
	.w2(32'h3af99820),
	.w3(32'hb9c76278),
	.w4(32'h3a955cb9),
	.w5(32'h3b22521e),
	.w6(32'h3a6c9525),
	.w7(32'hba543b8a),
	.w8(32'hbbc0a3db),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a1f7),
	.w1(32'hbb8503bd),
	.w2(32'hba227244),
	.w3(32'hbb919a6f),
	.w4(32'h39c3410f),
	.w5(32'h3b1d2983),
	.w6(32'hbbc72ad1),
	.w7(32'h3b1d3638),
	.w8(32'hba99a044),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad85f38),
	.w1(32'hbc1045ea),
	.w2(32'hb8cd95a6),
	.w3(32'hbba9e248),
	.w4(32'hbbc8e24e),
	.w5(32'h3c366421),
	.w6(32'h3ae71991),
	.w7(32'hbc2a2197),
	.w8(32'hba52e475),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda126a),
	.w1(32'h3b44306b),
	.w2(32'h3b12b7d1),
	.w3(32'hbb9011e2),
	.w4(32'h3c036ed6),
	.w5(32'hbace28dc),
	.w6(32'hbba52f86),
	.w7(32'h3c022408),
	.w8(32'hbb244fd7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b690),
	.w1(32'hbbaa72b6),
	.w2(32'hbb8a4505),
	.w3(32'h3b03c2e1),
	.w4(32'hbbe42b01),
	.w5(32'hbb65bf99),
	.w6(32'h3adf3fa2),
	.w7(32'hbba5744f),
	.w8(32'h3b236568),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd85d26),
	.w1(32'h3a50d210),
	.w2(32'h3a90b109),
	.w3(32'hbb8448c9),
	.w4(32'h3b811d2e),
	.w5(32'hbc33da30),
	.w6(32'hba7c2cfc),
	.w7(32'h3b50d0da),
	.w8(32'hbb8cd829),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad6ee4),
	.w1(32'h3b8d6592),
	.w2(32'h3a0097e2),
	.w3(32'hbc14e23a),
	.w4(32'hbad4da3b),
	.w5(32'hbae1e3f9),
	.w6(32'hbbb3b0b7),
	.w7(32'hbb51290b),
	.w8(32'hbbb55bc4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bf4da),
	.w1(32'hbb6cb585),
	.w2(32'h3b6d033f),
	.w3(32'hbadf70e6),
	.w4(32'h3b195543),
	.w5(32'hbb1bd5c7),
	.w6(32'hbbc1091a),
	.w7(32'hbb078f7a),
	.w8(32'h3a50284d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00b6c0),
	.w1(32'h3b9918f9),
	.w2(32'hbb81e59b),
	.w3(32'h3a501095),
	.w4(32'hbc08bc53),
	.w5(32'hbc42284d),
	.w6(32'h3a56abc4),
	.w7(32'h3b1e02af),
	.w8(32'hbb8fbaf4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af22f04),
	.w1(32'hbbedb0d1),
	.w2(32'hbbb15751),
	.w3(32'hbbc470c6),
	.w4(32'hbaa73ee0),
	.w5(32'hbb1b3364),
	.w6(32'hbab5d149),
	.w7(32'hbb15ae5a),
	.w8(32'hbbd50cf7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32e917),
	.w1(32'hbbf1f8a5),
	.w2(32'hbb8e96ac),
	.w3(32'h3b5ee739),
	.w4(32'hbb565f57),
	.w5(32'h3ac8b045),
	.w6(32'h3ada4e36),
	.w7(32'hbbac59b2),
	.w8(32'hbb97f3c7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc070801),
	.w1(32'h3b8fd830),
	.w2(32'h3bb9f19e),
	.w3(32'hbbaea588),
	.w4(32'h3b14fe9e),
	.w5(32'h3a9f9a77),
	.w6(32'hbbc2e98e),
	.w7(32'h3b8baad0),
	.w8(32'h3b8bfd83),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b34ab),
	.w1(32'hbb276526),
	.w2(32'hbb744e9a),
	.w3(32'h3b84074f),
	.w4(32'h3a09d3ac),
	.w5(32'hba160895),
	.w6(32'h3bff5122),
	.w7(32'hbada6915),
	.w8(32'h393ca10b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9580da),
	.w1(32'h3bc4250b),
	.w2(32'hba973cab),
	.w3(32'hbae4cbc9),
	.w4(32'h3b5831d1),
	.w5(32'h39b39c7a),
	.w6(32'h3b311b67),
	.w7(32'hba1b2d02),
	.w8(32'hb90baea1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8db193),
	.w1(32'hbb562072),
	.w2(32'hbaf99b34),
	.w3(32'h3b07250b),
	.w4(32'hba40729f),
	.w5(32'hbbfa2d90),
	.w6(32'h3ae32b28),
	.w7(32'hbb541b04),
	.w8(32'h3982990c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b2b81),
	.w1(32'h3c266a8a),
	.w2(32'h3bc55f7a),
	.w3(32'hba9515c5),
	.w4(32'h3c34b5b9),
	.w5(32'hbc7e1285),
	.w6(32'hbb0eb2ed),
	.w7(32'h3c5a3aba),
	.w8(32'h3be7929f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc1a37),
	.w1(32'hbbedd96e),
	.w2(32'hbbe9f227),
	.w3(32'h38bd1b1a),
	.w4(32'hbbb4be1f),
	.w5(32'h3b41ff03),
	.w6(32'h3beb980f),
	.w7(32'hbba2dd24),
	.w8(32'hbbeafb32),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2ffa9),
	.w1(32'h3b11d69f),
	.w2(32'hb91eb4a8),
	.w3(32'hbc060884),
	.w4(32'h38ee5633),
	.w5(32'hbb8edc01),
	.w6(32'hbc0f68bf),
	.w7(32'h3ac90e60),
	.w8(32'hbb180805),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920d60b),
	.w1(32'hbbb15c75),
	.w2(32'hbba232df),
	.w3(32'hbc223b98),
	.w4(32'h391a7223),
	.w5(32'h3ac89c92),
	.w6(32'hbbebc5da),
	.w7(32'h3abe90ab),
	.w8(32'hb9ee224b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba22d06),
	.w1(32'hbb1dcf8f),
	.w2(32'hbbdafa95),
	.w3(32'hbbc5ccfc),
	.w4(32'hba9f1dd5),
	.w5(32'hbb8ced0f),
	.w6(32'hbb3d9118),
	.w7(32'h3971185f),
	.w8(32'h3afd4d42),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12899a),
	.w1(32'h3ac1e823),
	.w2(32'h399b7598),
	.w3(32'h3adaf92d),
	.w4(32'h3baf0c9b),
	.w5(32'h3b5db292),
	.w6(32'h37e1090e),
	.w7(32'h3b11d824),
	.w8(32'h3b28a870),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9163f5),
	.w1(32'hbbb80e79),
	.w2(32'hbb1ef88f),
	.w3(32'h3b595556),
	.w4(32'hbadbca8a),
	.w5(32'h3c9ff8f3),
	.w6(32'h3b259f5b),
	.w7(32'hbbd395ca),
	.w8(32'hb7c54389),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c5ab3),
	.w1(32'hbbcd2406),
	.w2(32'hbb893059),
	.w3(32'h3b296d99),
	.w4(32'hbbd362a6),
	.w5(32'hbaa5f7d3),
	.w6(32'hbb8d248d),
	.w7(32'hbbd66dfd),
	.w8(32'hbb4271a8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36c0b7),
	.w1(32'hba0cbb85),
	.w2(32'h3a085797),
	.w3(32'hbb114954),
	.w4(32'h3a6c774f),
	.w5(32'h3af963f0),
	.w6(32'hbba33a53),
	.w7(32'hbb8cec62),
	.w8(32'h3b9cb8ac),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1046a),
	.w1(32'hbbfaa03d),
	.w2(32'hba2ff4d1),
	.w3(32'h3ae4c641),
	.w4(32'hbbe7d01d),
	.w5(32'h3c021786),
	.w6(32'h3af2fd14),
	.w7(32'hbc01df54),
	.w8(32'hbbd6fa5b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55872),
	.w1(32'hbb752806),
	.w2(32'h3b28bb1a),
	.w3(32'h3bc94bab),
	.w4(32'h3a09014a),
	.w5(32'h3d0207c3),
	.w6(32'hbbb5f2dd),
	.w7(32'hbb4930b2),
	.w8(32'h3bcb04c2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407383),
	.w1(32'hbb8d1f23),
	.w2(32'hbb4792be),
	.w3(32'h3bbf6e46),
	.w4(32'hbb9d3735),
	.w5(32'h3a97c887),
	.w6(32'hbaefc5c7),
	.w7(32'hbbfb636d),
	.w8(32'hbb61b246),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44dc3c),
	.w1(32'hbbd18560),
	.w2(32'hbb9c854d),
	.w3(32'hb99558a1),
	.w4(32'hbbbb2cb0),
	.w5(32'hba853cc4),
	.w6(32'hbb566c18),
	.w7(32'hbbf0311c),
	.w8(32'hbb0d3b35),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42d41),
	.w1(32'hb861f043),
	.w2(32'h3a187b44),
	.w3(32'hbbda2c96),
	.w4(32'hbb789b24),
	.w5(32'h3bcea7ae),
	.w6(32'hbbc259a5),
	.w7(32'hba8e54a9),
	.w8(32'h3b460944),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0742c),
	.w1(32'hbb2455af),
	.w2(32'h3b863ff0),
	.w3(32'hbae69295),
	.w4(32'hba76e3a5),
	.w5(32'h3c0c6e32),
	.w6(32'hbb288827),
	.w7(32'hbbdf40e2),
	.w8(32'hbbb23109),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c6896),
	.w1(32'h3bc468f4),
	.w2(32'h3b13c285),
	.w3(32'hbb1b321e),
	.w4(32'hbb16a44b),
	.w5(32'hbc6292cf),
	.w6(32'hbb7b34b0),
	.w7(32'h3b4bc6b4),
	.w8(32'hbaec56c7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba389f24),
	.w1(32'h3b249765),
	.w2(32'h3b3d0a72),
	.w3(32'h3a57a2f3),
	.w4(32'hbb842247),
	.w5(32'hbc06db6b),
	.w6(32'h3983f304),
	.w7(32'hba17162a),
	.w8(32'h3778806a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5febfb),
	.w1(32'h3af3fa7f),
	.w2(32'hbb4b3299),
	.w3(32'hba23f84b),
	.w4(32'h3bdac8f5),
	.w5(32'h3bb28c86),
	.w6(32'h3b2e3aad),
	.w7(32'h3b5c07b7),
	.w8(32'h3a2413f1),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9571a),
	.w1(32'h3712646b),
	.w2(32'h3ac91d99),
	.w3(32'h3ad906a4),
	.w4(32'h3a63ac16),
	.w5(32'hbb6a5a2e),
	.w6(32'h3b942e91),
	.w7(32'h3b7407bf),
	.w8(32'h3b47abd7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ee9e4),
	.w1(32'h3c3cd255),
	.w2(32'h3c6f4925),
	.w3(32'hbab24a5a),
	.w4(32'hba8fa713),
	.w5(32'h3c108495),
	.w6(32'h3aeff0d8),
	.w7(32'h3c289426),
	.w8(32'h3c962451),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04492d),
	.w1(32'h3cd78886),
	.w2(32'h3c5e0193),
	.w3(32'h3b7fb946),
	.w4(32'h3c4e5112),
	.w5(32'hbc86ac15),
	.w6(32'h3c1d38f8),
	.w7(32'h3cd7f4b8),
	.w8(32'h3c7e0af6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf8e2d),
	.w1(32'h3ad33e7b),
	.w2(32'hbafe9923),
	.w3(32'h3bf84e1c),
	.w4(32'h3ae2f3e7),
	.w5(32'hbba79140),
	.w6(32'h3c9cd7ed),
	.w7(32'hbbcff41f),
	.w8(32'hbbd57ab5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969061),
	.w1(32'h3a83c351),
	.w2(32'h3b74028c),
	.w3(32'h3aa9142d),
	.w4(32'h3b100c5f),
	.w5(32'h3ba7b144),
	.w6(32'hbbb14ecc),
	.w7(32'h3c1668c2),
	.w8(32'h3bc34b10),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2252db),
	.w1(32'hbb18f877),
	.w2(32'hbb2d607f),
	.w3(32'h3bc23e16),
	.w4(32'hbbe22c85),
	.w5(32'h3bd5434b),
	.w6(32'h3bbc623c),
	.w7(32'hbb553c44),
	.w8(32'hbbfaea7f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932b2b7),
	.w1(32'h3b60ca1e),
	.w2(32'h3a8a62f6),
	.w3(32'hbaf6372f),
	.w4(32'hbc041b77),
	.w5(32'hbbdbeace),
	.w6(32'hbc1eed1d),
	.w7(32'hbb9eb054),
	.w8(32'hb95be259),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b811428),
	.w1(32'hbc08dc42),
	.w2(32'hbb7075a0),
	.w3(32'h3bb3951e),
	.w4(32'hbb9ab9e0),
	.w5(32'h3bd375b8),
	.w6(32'h3b8daa1b),
	.w7(32'hbc07ceba),
	.w8(32'hbbbe7936),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139079),
	.w1(32'hba83fe93),
	.w2(32'hbb6db665),
	.w3(32'hbb6469ee),
	.w4(32'hbb072f79),
	.w5(32'h3abe14e5),
	.w6(32'hbc01cf49),
	.w7(32'hba63f1af),
	.w8(32'hb9e64c4f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb764506),
	.w1(32'hbb82c893),
	.w2(32'hbb07a52d),
	.w3(32'hbb8ac73b),
	.w4(32'h3a8d58aa),
	.w5(32'h3b527a2c),
	.w6(32'hb7fe8a02),
	.w7(32'hbbad1c3e),
	.w8(32'h3af18df9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb846f2f),
	.w1(32'hbacf85a9),
	.w2(32'hba978d70),
	.w3(32'hb9ebfb53),
	.w4(32'h3a6095df),
	.w5(32'h3c101db6),
	.w6(32'hba272838),
	.w7(32'h3bce916b),
	.w8(32'h3b934274),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae24be),
	.w1(32'h3b97d87b),
	.w2(32'h3bb440fe),
	.w3(32'h3bf7a3e5),
	.w4(32'hbb5b0228),
	.w5(32'h3b94c18f),
	.w6(32'h3c20079d),
	.w7(32'hb9ddb605),
	.w8(32'h3b626ada),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22cb1d),
	.w1(32'h3ac0fa6c),
	.w2(32'hbabc72ca),
	.w3(32'hbb3f5a22),
	.w4(32'h3b81c1f1),
	.w5(32'h3b9ee936),
	.w6(32'hbb064048),
	.w7(32'hbaf19b48),
	.w8(32'hbaad9b8a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc6a0),
	.w1(32'hbac04d27),
	.w2(32'hbaa7e427),
	.w3(32'hbbb4387f),
	.w4(32'h3ab25cca),
	.w5(32'hbaa9ade6),
	.w6(32'hbb500ded),
	.w7(32'hbb2b7055),
	.w8(32'hba9c8ed4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86e181),
	.w1(32'hba968760),
	.w2(32'hbb47b5b4),
	.w3(32'h3929944e),
	.w4(32'hba82b09b),
	.w5(32'hbb8ec23c),
	.w6(32'hbb65deb8),
	.w7(32'hbba1b14e),
	.w8(32'hbb3fe2e3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb131f6),
	.w1(32'h3ac8686f),
	.w2(32'hbba952c5),
	.w3(32'hbbf3048e),
	.w4(32'h3a521683),
	.w5(32'h3b483b38),
	.w6(32'hbb243c1a),
	.w7(32'h3a98ef8b),
	.w8(32'hbb8d8607),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe9759),
	.w1(32'h3aa07762),
	.w2(32'h3ab301fb),
	.w3(32'hbc54fec4),
	.w4(32'h3b25f561),
	.w5(32'hbc1f6613),
	.w6(32'hbc015d2e),
	.w7(32'h3bba611f),
	.w8(32'h391e8944),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa31f2),
	.w1(32'h3b2be384),
	.w2(32'h3b0e1a5a),
	.w3(32'h3b0ff01a),
	.w4(32'h3bcca806),
	.w5(32'h3be1a54d),
	.w6(32'h3b653f03),
	.w7(32'hbae29b01),
	.w8(32'h3c1a0260),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfba0e8),
	.w1(32'hbc033b0e),
	.w2(32'hbbb4f01f),
	.w3(32'h3c17765f),
	.w4(32'hbbbaf3a5),
	.w5(32'hbbc67bb2),
	.w6(32'h3b09211f),
	.w7(32'hbbab4895),
	.w8(32'hbbb7f7c4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1de052),
	.w1(32'h3b369be2),
	.w2(32'h3bd8e1c9),
	.w3(32'hbc0c5bd8),
	.w4(32'h3baf20dd),
	.w5(32'h3bde06e8),
	.w6(32'hbc396743),
	.w7(32'h3bc07afb),
	.w8(32'h3b990ebf),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aada37b),
	.w1(32'h3ad897cc),
	.w2(32'hbb9f16de),
	.w3(32'hbb1126f2),
	.w4(32'h3b13b2ef),
	.w5(32'hbbc7ec83),
	.w6(32'hb9d268be),
	.w7(32'hba479118),
	.w8(32'h39f7cdb0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb921c33),
	.w1(32'hbb2150fa),
	.w2(32'h3b61a085),
	.w3(32'hbb3f0b09),
	.w4(32'hbb2c9738),
	.w5(32'h3c4a931c),
	.w6(32'hbb31eab9),
	.w7(32'h3a3c6528),
	.w8(32'h3c322ab5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad67e0b),
	.w1(32'hbb878573),
	.w2(32'h3ae97504),
	.w3(32'h3bc2ad45),
	.w4(32'h3a58334c),
	.w5(32'h3d26b867),
	.w6(32'h3c5f0867),
	.w7(32'h397bd8e7),
	.w8(32'h3c10eb59),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7d518),
	.w1(32'hbb71610e),
	.w2(32'hbb085d6b),
	.w3(32'h3c1dfd8b),
	.w4(32'h3ba37726),
	.w5(32'hbb10bec5),
	.w6(32'h3b58ab4d),
	.w7(32'h3bb76e74),
	.w8(32'h3af13b05),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10ae4b),
	.w1(32'h3ba8130e),
	.w2(32'h3baf1aaa),
	.w3(32'h3b88f221),
	.w4(32'h3be72128),
	.w5(32'h3c807f9e),
	.w6(32'h3a43ae4f),
	.w7(32'h3ba8cfa4),
	.w8(32'h3ae0833c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d8d6),
	.w1(32'h3be3f1ac),
	.w2(32'h3c056015),
	.w3(32'h3b362c89),
	.w4(32'h3c15e885),
	.w5(32'h3c0d2bbd),
	.w6(32'h3804c391),
	.w7(32'h3bdde786),
	.w8(32'h3bd0c0a0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8345),
	.w1(32'h3bce3bf0),
	.w2(32'h3bb23d36),
	.w3(32'hbb6f1f62),
	.w4(32'h3c0102a6),
	.w5(32'h3c16eb64),
	.w6(32'hba69e90b),
	.w7(32'h3bfe0e1c),
	.w8(32'h3b94d99b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548aaf),
	.w1(32'hbb37388e),
	.w2(32'hb9982919),
	.w3(32'h3a803995),
	.w4(32'hbabbf6c5),
	.w5(32'hbaaf7c4b),
	.w6(32'h3b18e896),
	.w7(32'hbba4c27c),
	.w8(32'hbabfa985),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75c257),
	.w1(32'hbb632c2f),
	.w2(32'hbb80f83a),
	.w3(32'h3a7281b1),
	.w4(32'hba294072),
	.w5(32'h3b8f9fb4),
	.w6(32'h3a6c82f8),
	.w7(32'h3b9c8bdf),
	.w8(32'h3ad60610),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69726d),
	.w1(32'h396e4b29),
	.w2(32'h3b4d9438),
	.w3(32'h3b5ef0a5),
	.w4(32'h3bb4b979),
	.w5(32'h3a6457f6),
	.w6(32'h3b40d637),
	.w7(32'h3ba23186),
	.w8(32'hbb01b674),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cdef0e),
	.w1(32'h3ba5bd06),
	.w2(32'h3b229b09),
	.w3(32'hbb2d6ec1),
	.w4(32'h3b2e0948),
	.w5(32'hbbd33ba6),
	.w6(32'h3a578a69),
	.w7(32'h3b4b1980),
	.w8(32'h3b94f66e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e4e72),
	.w1(32'hbbfb95cf),
	.w2(32'hbb1b26e2),
	.w3(32'hbb698cc3),
	.w4(32'hbb925932),
	.w5(32'h3b6dc9a0),
	.w6(32'h390effc9),
	.w7(32'hbb3ab7f1),
	.w8(32'hbb45910f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83482),
	.w1(32'hbbd81191),
	.w2(32'hba599c72),
	.w3(32'h388549c4),
	.w4(32'hbb193edb),
	.w5(32'hbb95a1cc),
	.w6(32'hbb76d265),
	.w7(32'hbb938251),
	.w8(32'h3a8971ec),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7af0b),
	.w1(32'h3a86ebf3),
	.w2(32'hbb05c4f7),
	.w3(32'hbb98cbe4),
	.w4(32'hb55751d1),
	.w5(32'hbc44910b),
	.w6(32'hbb1f8ea7),
	.w7(32'h3a156456),
	.w8(32'hbba574be),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01a9b8),
	.w1(32'h3babf808),
	.w2(32'hbb040ee7),
	.w3(32'h3a1d1a7f),
	.w4(32'hbb9a8863),
	.w5(32'hbba1b3ca),
	.w6(32'hbb68e20a),
	.w7(32'hbb560938),
	.w8(32'hba299aa5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02628c),
	.w1(32'hbbb111d1),
	.w2(32'hbb35e4df),
	.w3(32'hbb2437fd),
	.w4(32'hbb06fe27),
	.w5(32'hbc0cdf3a),
	.w6(32'hbb980beb),
	.w7(32'hbb0b7d52),
	.w8(32'hbba2dcf6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad299ae),
	.w1(32'hbaef6687),
	.w2(32'h3bad5b4f),
	.w3(32'hbbc31a11),
	.w4(32'h3ba5f41d),
	.w5(32'hbba91e67),
	.w6(32'hbb0a733d),
	.w7(32'h3b806d38),
	.w8(32'h3be4c104),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62d497),
	.w1(32'h3bfd0120),
	.w2(32'h3b338811),
	.w3(32'hbb158dd0),
	.w4(32'h3bd3c0df),
	.w5(32'hbbab6859),
	.w6(32'h3bb801c2),
	.w7(32'hbbad7ed7),
	.w8(32'hbb21fca2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c041313),
	.w1(32'h3a1f10e5),
	.w2(32'h3b0d93be),
	.w3(32'h3c3240ee),
	.w4(32'h3af4ba54),
	.w5(32'h3aab98e8),
	.w6(32'h3b8d4db5),
	.w7(32'hbabff665),
	.w8(32'hbb75f80f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b8005),
	.w1(32'h3b6ab407),
	.w2(32'h3b2c1c2b),
	.w3(32'hba7b1da8),
	.w4(32'h3ace2e0f),
	.w5(32'hbbab542b),
	.w6(32'hbb4916a1),
	.w7(32'hba8306f4),
	.w8(32'h3b083e9a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5453bc),
	.w1(32'hbbb01e10),
	.w2(32'hbab1526b),
	.w3(32'hbbe004ec),
	.w4(32'hbb67d58a),
	.w5(32'h3c067262),
	.w6(32'hbb0cf379),
	.w7(32'hbbc97495),
	.w8(32'hba2b3528),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5a10f),
	.w1(32'h3bb4b0e0),
	.w2(32'h3b64e14b),
	.w3(32'hb959b22d),
	.w4(32'h3b0879e8),
	.w5(32'hbbd3ff1d),
	.w6(32'h39319b97),
	.w7(32'hbb1e7f08),
	.w8(32'h3a007ce4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6023),
	.w1(32'h3a8139c6),
	.w2(32'h3a239290),
	.w3(32'hbb093f7c),
	.w4(32'h3bbaabb4),
	.w5(32'h3c2f3a89),
	.w6(32'hbb5114d6),
	.w7(32'h3ba92298),
	.w8(32'h3ae37545),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02f872),
	.w1(32'h3b503572),
	.w2(32'h3a0c1b3c),
	.w3(32'hbc285829),
	.w4(32'h396eb3a5),
	.w5(32'hbb9879f5),
	.w6(32'hbbcf552f),
	.w7(32'h3b292f6c),
	.w8(32'h3b10d2ec),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29e50),
	.w1(32'h3c649d65),
	.w2(32'h3bfb2796),
	.w3(32'hbbc22385),
	.w4(32'h3c20ee97),
	.w5(32'h3bf5e51f),
	.w6(32'hbb8fe6ac),
	.w7(32'h3c105dc7),
	.w8(32'h3bd00c9b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0c82c),
	.w1(32'hbbfc0368),
	.w2(32'hbbd48134),
	.w3(32'h3c0b8418),
	.w4(32'hbba420a7),
	.w5(32'h3af0818b),
	.w6(32'h3bc86ef0),
	.w7(32'hbc1497f1),
	.w8(32'hbbefa2a6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab8a4),
	.w1(32'h38b739f4),
	.w2(32'h3bd559ef),
	.w3(32'hbbc4aaca),
	.w4(32'h3a7d0841),
	.w5(32'h3c0ba36b),
	.w6(32'hbb966dd7),
	.w7(32'h3b196997),
	.w8(32'h3c1ad880),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f32386),
	.w1(32'h39d8fa7c),
	.w2(32'h3a304835),
	.w3(32'h3bc5710f),
	.w4(32'h3ba5f794),
	.w5(32'h3b9a9abd),
	.w6(32'h3b566790),
	.w7(32'h3c02bc4c),
	.w8(32'h3b99b3dc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bbcefe),
	.w1(32'h3b169663),
	.w2(32'h3af5e211),
	.w3(32'hba855810),
	.w4(32'h3b991929),
	.w5(32'h3b5ff20e),
	.w6(32'hbace412b),
	.w7(32'hb9cd5447),
	.w8(32'hbab418d4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43103),
	.w1(32'hbb3360b7),
	.w2(32'hbb299f8b),
	.w3(32'h3b850375),
	.w4(32'hbaa671af),
	.w5(32'hbb6a8dfc),
	.w6(32'h3aaba370),
	.w7(32'hbb107337),
	.w8(32'hbb1efb44),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6366),
	.w1(32'hba3e33bd),
	.w2(32'h3a60dac8),
	.w3(32'h3ad79ce5),
	.w4(32'hbb019ede),
	.w5(32'hba7816e1),
	.w6(32'hbac568fb),
	.w7(32'hb938fbba),
	.w8(32'h3a090e8f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0bd0),
	.w1(32'h3a116da7),
	.w2(32'hb918aaee),
	.w3(32'h39e2934f),
	.w4(32'hbacc953d),
	.w5(32'hbb0bc3ab),
	.w6(32'h3b09e695),
	.w7(32'hbb318923),
	.w8(32'h3a92810e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b86cf),
	.w1(32'h3b308502),
	.w2(32'h3b78ef1a),
	.w3(32'hbaf8eb41),
	.w4(32'h3b10c8f1),
	.w5(32'h3ada36fb),
	.w6(32'hbaf6c21e),
	.w7(32'h3b542159),
	.w8(32'h3a4ff2d1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2345b9),
	.w1(32'h399cdfcd),
	.w2(32'hba66fcbc),
	.w3(32'h3a2cf204),
	.w4(32'hbadd4634),
	.w5(32'h3a280697),
	.w6(32'h3a7d514d),
	.w7(32'h381615dd),
	.w8(32'h3a95a148),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10307c),
	.w1(32'hba8be28e),
	.w2(32'hbb572885),
	.w3(32'hba98eae6),
	.w4(32'h3b09a0a3),
	.w5(32'hbb95d2a7),
	.w6(32'h3ab4a146),
	.w7(32'h3a12a16e),
	.w8(32'h3aaefbc0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fcb2f),
	.w1(32'h3b3dd91c),
	.w2(32'h3b18feb1),
	.w3(32'hbb371fd2),
	.w4(32'h3b38a099),
	.w5(32'h3b38c4f9),
	.w6(32'hb915a4aa),
	.w7(32'h3b91975a),
	.w8(32'h3b8dd65e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152638),
	.w1(32'hbaf82540),
	.w2(32'h3aeeeb29),
	.w3(32'h3b069c7e),
	.w4(32'hbace2e5a),
	.w5(32'h3bc6b095),
	.w6(32'h3b294136),
	.w7(32'h3a711f25),
	.w8(32'h3a4f00be),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9932159),
	.w1(32'hbb1cd92c),
	.w2(32'hbb11bcc6),
	.w3(32'hb9dbc91c),
	.w4(32'hbc07424c),
	.w5(32'hbbf0c9bd),
	.w6(32'h3a1e4416),
	.w7(32'hbb8a30b5),
	.w8(32'hbb44f01a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33739d),
	.w1(32'h3a908678),
	.w2(32'h3915852a),
	.w3(32'hb9c0891b),
	.w4(32'h3a9b4be5),
	.w5(32'h3b718808),
	.w6(32'h3a96eecf),
	.w7(32'h39ae9a51),
	.w8(32'h3ad7252a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4725e),
	.w1(32'h3b135dbc),
	.w2(32'h381c72a9),
	.w3(32'hba67418e),
	.w4(32'h3b3c8dbf),
	.w5(32'h3a98bbaf),
	.w6(32'hba986fef),
	.w7(32'h3a1f2ce2),
	.w8(32'h38dbac7b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17df40),
	.w1(32'h3aa97a38),
	.w2(32'hbb9983fa),
	.w3(32'h3b2615c2),
	.w4(32'hba93b28a),
	.w5(32'hbb4946e6),
	.w6(32'h3aa90b70),
	.w7(32'hbb266efc),
	.w8(32'h3a349aaf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb580e),
	.w1(32'h3b0460b3),
	.w2(32'h3ade75dd),
	.w3(32'hba07c160),
	.w4(32'h3b0baf66),
	.w5(32'h3bc60ab1),
	.w6(32'h397288e8),
	.w7(32'h3ae58688),
	.w8(32'h3a76cc07),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b2830),
	.w1(32'h3be515f4),
	.w2(32'hba48114f),
	.w3(32'h3af5714b),
	.w4(32'h3bccc23f),
	.w5(32'hbb23728f),
	.w6(32'h383a8628),
	.w7(32'h3b1bad1f),
	.w8(32'hbbb98336),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d835e6),
	.w1(32'h3a33f64e),
	.w2(32'hbb076560),
	.w3(32'hbac9f023),
	.w4(32'hba4f5b34),
	.w5(32'hbace6b1b),
	.w6(32'hbb4dd7eb),
	.w7(32'hb9f8e312),
	.w8(32'hb91dd806),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7765d6),
	.w1(32'h3a2a6af3),
	.w2(32'h3aa8fba7),
	.w3(32'hbb42daa7),
	.w4(32'hba30ab62),
	.w5(32'h37c1798b),
	.w6(32'h3a8d4470),
	.w7(32'hbb3ad4f0),
	.w8(32'h3b6f90f7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901afe3),
	.w1(32'h3b0e2609),
	.w2(32'hba8f2ac0),
	.w3(32'h3a7d6406),
	.w4(32'h3b12e838),
	.w5(32'hba455fe0),
	.w6(32'h3afb5012),
	.w7(32'h3a27c163),
	.w8(32'h3b965ca1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b1e3),
	.w1(32'h3b98ca0d),
	.w2(32'h3a9ccf21),
	.w3(32'hb8a7cc10),
	.w4(32'h3bb77f39),
	.w5(32'h3b1c5041),
	.w6(32'h3b433f44),
	.w7(32'h3baecee1),
	.w8(32'h3b22056a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b3c9),
	.w1(32'hba46ff1c),
	.w2(32'h3b829487),
	.w3(32'hba7c503f),
	.w4(32'hb9ed9f7f),
	.w5(32'h3be68768),
	.w6(32'h39dfc189),
	.w7(32'h399319c2),
	.w8(32'h3be16983),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb791ee),
	.w1(32'hbaa2ffaf),
	.w2(32'hbb00e4bc),
	.w3(32'h3bd8d662),
	.w4(32'hbba122c0),
	.w5(32'hbafe010f),
	.w6(32'h3bf35ab4),
	.w7(32'hbaa23195),
	.w8(32'h3ae139f1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad81389),
	.w1(32'h3b8fb0ca),
	.w2(32'h3b1abd86),
	.w3(32'hbb2c309b),
	.w4(32'h3b7b568f),
	.w5(32'h3bfc410d),
	.w6(32'hbb0ead30),
	.w7(32'h3b3abf57),
	.w8(32'h3b26721c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374933),
	.w1(32'h3b4dd3da),
	.w2(32'hba696038),
	.w3(32'h3b7428a8),
	.w4(32'h3ad8cb3a),
	.w5(32'h3abc9265),
	.w6(32'h3ac4ea79),
	.w7(32'h3aed7797),
	.w8(32'h39190b8e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06deab),
	.w1(32'hbb1b012d),
	.w2(32'hbb633840),
	.w3(32'hb93fc056),
	.w4(32'hbab66091),
	.w5(32'hbb787aeb),
	.w6(32'hbaa8bf1d),
	.w7(32'h3b836bff),
	.w8(32'h3b7792ac),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251f32),
	.w1(32'hbb0c2597),
	.w2(32'h3b1606a0),
	.w3(32'h39d28982),
	.w4(32'hbb655bfc),
	.w5(32'h39617829),
	.w6(32'h3ac0fe68),
	.w7(32'hbb3d908f),
	.w8(32'h3a334f89),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e3c86),
	.w1(32'h3bcfd267),
	.w2(32'h3b46bdaf),
	.w3(32'h3a7e7570),
	.w4(32'h3bd78e2d),
	.w5(32'h3b776fd5),
	.w6(32'h3b5daa24),
	.w7(32'h3b799a95),
	.w8(32'h3b1eb0cb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25296d),
	.w1(32'h3be0e611),
	.w2(32'h3b3f6d34),
	.w3(32'h3a8a7961),
	.w4(32'h3b3fe201),
	.w5(32'h3b0aae58),
	.w6(32'hbaa1aee3),
	.w7(32'h3bdb4508),
	.w8(32'h3adf04cf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5ebd5),
	.w1(32'h3a82cdee),
	.w2(32'h3b0cf1a6),
	.w3(32'h3ad2007c),
	.w4(32'h39816ff5),
	.w5(32'h3a67203c),
	.w6(32'hb908d5d3),
	.w7(32'hb98f5b8e),
	.w8(32'h3b0b475b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba307420),
	.w1(32'hbb2c5095),
	.w2(32'h39440fde),
	.w3(32'hb9e1086b),
	.w4(32'hb73d4cd0),
	.w5(32'hbb4306c1),
	.w6(32'h3b501f73),
	.w7(32'h3b010807),
	.w8(32'hbaa7d7c1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8312f73),
	.w1(32'h3b5d3fcb),
	.w2(32'h3a71db3a),
	.w3(32'hbb22e9ad),
	.w4(32'h3a985a5e),
	.w5(32'hbae58eba),
	.w6(32'hba98bdec),
	.w7(32'h3b6ddc00),
	.w8(32'h3b34b506),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaac51),
	.w1(32'hbaadba0d),
	.w2(32'h392d2bd2),
	.w3(32'hb9e67c56),
	.w4(32'h3aea9234),
	.w5(32'h3b97b3a4),
	.w6(32'h3aee52b1),
	.w7(32'h39ffaaa0),
	.w8(32'h3ad30d3a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d47f),
	.w1(32'h3ad555ed),
	.w2(32'hb91bf299),
	.w3(32'h39308750),
	.w4(32'h39f4011e),
	.w5(32'hbaed514e),
	.w6(32'hb87bdd33),
	.w7(32'hba92f760),
	.w8(32'hb9c1b942),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9612b),
	.w1(32'hb9439cf9),
	.w2(32'h3a585030),
	.w3(32'h3b10e442),
	.w4(32'h38b794b3),
	.w5(32'h3ba5c596),
	.w6(32'h39640caa),
	.w7(32'hb9cc3891),
	.w8(32'h3b1c63c0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79253),
	.w1(32'hbb359baa),
	.w2(32'hbb94687a),
	.w3(32'h3a12ea64),
	.w4(32'hbb943050),
	.w5(32'hbb7c9645),
	.w6(32'h3a9077fe),
	.w7(32'h39807f1f),
	.w8(32'h3a97fa17),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ecae8),
	.w1(32'h3a36fa26),
	.w2(32'h3a9abab7),
	.w3(32'h3b0ffb74),
	.w4(32'h38922c55),
	.w5(32'h3b7f8912),
	.w6(32'h3b8851a8),
	.w7(32'h3a2663a9),
	.w8(32'h39ce8302),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d7581),
	.w1(32'h3afed7c9),
	.w2(32'hba9326d5),
	.w3(32'h3b2d4453),
	.w4(32'h3b54d87a),
	.w5(32'h39b71d00),
	.w6(32'h3a0e91b7),
	.w7(32'h3b1a96dd),
	.w8(32'hbaef10f8),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfa852),
	.w1(32'h3a67a872),
	.w2(32'h3bb27f1a),
	.w3(32'hba84dd62),
	.w4(32'hba466282),
	.w5(32'h39fb51e3),
	.w6(32'hbade453e),
	.w7(32'h382077e6),
	.w8(32'h3b24f0b4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bdea7),
	.w1(32'hb92310b9),
	.w2(32'hbac7543b),
	.w3(32'h3c31c9a0),
	.w4(32'hba3cf0d0),
	.w5(32'hb8eff9b7),
	.w6(32'h3bd59405),
	.w7(32'h3b344ef9),
	.w8(32'h3abef9a2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa1846),
	.w1(32'hbaa2161c),
	.w2(32'hbbaa0199),
	.w3(32'h3ae7cf05),
	.w4(32'hbb0bbd8d),
	.w5(32'hbb0c2047),
	.w6(32'h3b2007a6),
	.w7(32'h3ab0b869),
	.w8(32'hb98d2209),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39065b76),
	.w1(32'h3c4f3272),
	.w2(32'h3bdfba03),
	.w3(32'h3ad635f3),
	.w4(32'h395d600c),
	.w5(32'hbb128791),
	.w6(32'h3b2463db),
	.w7(32'hb9af1739),
	.w8(32'hbb3adff9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459a8a),
	.w1(32'hb9c7a0c6),
	.w2(32'hbb739953),
	.w3(32'hbac84d70),
	.w4(32'h3ae53c9f),
	.w5(32'hbb91c4b3),
	.w6(32'hbacd8da7),
	.w7(32'h3b53ef50),
	.w8(32'hbb32b63a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1df8f),
	.w1(32'hbb91ba62),
	.w2(32'h3b1d3263),
	.w3(32'hbb08470a),
	.w4(32'hbb47ffa4),
	.w5(32'h3ab705a1),
	.w6(32'hbab565a3),
	.w7(32'hbb55de01),
	.w8(32'hbb204ac1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade052c),
	.w1(32'h3b9d9f54),
	.w2(32'h3b20cfea),
	.w3(32'h3955a966),
	.w4(32'h3b4f5887),
	.w5(32'hbacd0f36),
	.w6(32'hba68dca2),
	.w7(32'h3c0972f9),
	.w8(32'hbb5fdc18),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e4a6),
	.w1(32'hba181c5f),
	.w2(32'h38fe53bd),
	.w3(32'hbb835232),
	.w4(32'h3abea085),
	.w5(32'h3b81b19c),
	.w6(32'hba3c42fb),
	.w7(32'hba564649),
	.w8(32'hbaf0caa7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945238b),
	.w1(32'hb90fb7f8),
	.w2(32'h3b0150bc),
	.w3(32'hbb1c3ccd),
	.w4(32'h3a8e4f66),
	.w5(32'h3bf5122c),
	.w6(32'hbb09f42d),
	.w7(32'h3b47fb72),
	.w8(32'h3b7bcaea),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5b96),
	.w1(32'hb93b3f61),
	.w2(32'h3ae17742),
	.w3(32'hbaff119a),
	.w4(32'h3a10b3a1),
	.w5(32'h3c079659),
	.w6(32'hbb318625),
	.w7(32'h3ae9a8dc),
	.w8(32'h3b09787d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3445e0),
	.w1(32'h3b9812d4),
	.w2(32'h3b09fe1d),
	.w3(32'h3ac70108),
	.w4(32'h3b58631d),
	.w5(32'h3b4a1278),
	.w6(32'hb74ae172),
	.w7(32'h3b122cae),
	.w8(32'hba70a234),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c457f),
	.w1(32'h3aeac53a),
	.w2(32'h3b3fb520),
	.w3(32'h3ae00e01),
	.w4(32'h3b39c40e),
	.w5(32'hba379ddb),
	.w6(32'h3a2e86a2),
	.w7(32'h3a5f7465),
	.w8(32'h3b268c4a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7daf7c),
	.w1(32'hbad1d365),
	.w2(32'h3ab6c387),
	.w3(32'hba668246),
	.w4(32'h3aa20ab8),
	.w5(32'h3b4fda74),
	.w6(32'h3b09a4bc),
	.w7(32'h3b097c8d),
	.w8(32'h3ab9b103),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbd45),
	.w1(32'h3b0bc938),
	.w2(32'h39dcd2df),
	.w3(32'h3b6f5aee),
	.w4(32'h3a9bd2cb),
	.w5(32'h3623c41b),
	.w6(32'h3b0d9796),
	.w7(32'h3b0bb244),
	.w8(32'h3afbf945),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4fd58),
	.w1(32'hbb23b4a5),
	.w2(32'hbb631bf6),
	.w3(32'hba07caed),
	.w4(32'hbb170c91),
	.w5(32'hbae54ba3),
	.w6(32'h3a882b3b),
	.w7(32'hb7f0d553),
	.w8(32'h3bb27047),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1d11),
	.w1(32'h3ab678b3),
	.w2(32'hba4aca85),
	.w3(32'h3a1eb134),
	.w4(32'h3b0bad46),
	.w5(32'h3abfe369),
	.w6(32'h3b960251),
	.w7(32'h3acc22a7),
	.w8(32'h3b8127a3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a229744),
	.w1(32'hbb5fd613),
	.w2(32'hbb3a586a),
	.w3(32'hba131581),
	.w4(32'hbb40be68),
	.w5(32'h39ca285f),
	.w6(32'hba88b6da),
	.w7(32'hbb2088be),
	.w8(32'hbb0d0c1f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32015c),
	.w1(32'h3b0133bb),
	.w2(32'hbb535922),
	.w3(32'hbbad9804),
	.w4(32'h3b63e411),
	.w5(32'h3b45360f),
	.w6(32'hbb92d077),
	.w7(32'h3b0e8fb1),
	.w8(32'hba8a4e5e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f6b52),
	.w1(32'h3913b5c0),
	.w2(32'hba3a8c3a),
	.w3(32'hb82a5b5f),
	.w4(32'hb9f16680),
	.w5(32'hb8c0ead5),
	.w6(32'hb7b744e4),
	.w7(32'h3ac4eee9),
	.w8(32'hba74426b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5a712),
	.w1(32'hbae2f1f5),
	.w2(32'hbbc3ee1d),
	.w3(32'h3a8fe0b3),
	.w4(32'h3babd007),
	.w5(32'h3a6f5280),
	.w6(32'h3af6bf36),
	.w7(32'h3b677d9b),
	.w8(32'h39488202),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56cc8d),
	.w1(32'h3a25f56f),
	.w2(32'hbb8c8fa5),
	.w3(32'hbadcda25),
	.w4(32'hba273d59),
	.w5(32'h3a25cb4b),
	.w6(32'hba967300),
	.w7(32'hba543238),
	.w8(32'h3be17cd9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule