module layer_8_featuremap_156(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26687),
	.w1(32'h3b519faf),
	.w2(32'h3b888ac2),
	.w3(32'h3a2fe54d),
	.w4(32'h3c5e4826),
	.w5(32'h3c16ecb1),
	.w6(32'h3bc942cb),
	.w7(32'h3bd59a22),
	.w8(32'hbb8c291c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d7dbc),
	.w1(32'h3b835267),
	.w2(32'hba8b5d72),
	.w3(32'h3a9d0083),
	.w4(32'h3b14281c),
	.w5(32'hbaec1102),
	.w6(32'hbb689b86),
	.w7(32'h3b665ff8),
	.w8(32'h3a55e6ef),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44d97),
	.w1(32'hbbded061),
	.w2(32'hbc91fd68),
	.w3(32'hbac9833c),
	.w4(32'hbc9cbc9b),
	.w5(32'hbca93e53),
	.w6(32'hbbaa5e0d),
	.w7(32'hbca71414),
	.w8(32'hbc7d6d52),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6424b2),
	.w1(32'hbc6d31ec),
	.w2(32'h3c587cb9),
	.w3(32'hbc03821f),
	.w4(32'hbb2fbd58),
	.w5(32'hbbe88c6f),
	.w6(32'hbc225854),
	.w7(32'hbc3fd992),
	.w8(32'h3ca3a14d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb8271),
	.w1(32'h3b9ef378),
	.w2(32'hba813721),
	.w3(32'h3b5eeacc),
	.w4(32'h3ace6745),
	.w5(32'h3bd8c2a0),
	.w6(32'hba99c038),
	.w7(32'h3b91a38a),
	.w8(32'h3a4a0352),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409a06),
	.w1(32'hbbf2f196),
	.w2(32'h3a5b688f),
	.w3(32'hbaf193d3),
	.w4(32'hbbdbb146),
	.w5(32'h3c3eeef3),
	.w6(32'hbc3300f2),
	.w7(32'h3b689b92),
	.w8(32'h3b5abab0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae3e8c),
	.w1(32'hbbf76fe6),
	.w2(32'hbc1e4720),
	.w3(32'hbb18f06f),
	.w4(32'hbbc33a87),
	.w5(32'hbb538b83),
	.w6(32'h3b34f8ea),
	.w7(32'hbc3065ab),
	.w8(32'h3b4c08d7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52e606),
	.w1(32'hbcbb03d3),
	.w2(32'h3aa6b8c0),
	.w3(32'hbb54e747),
	.w4(32'h3bbf4af2),
	.w5(32'hbc03465b),
	.w6(32'h3ad54485),
	.w7(32'hbb0b1a44),
	.w8(32'h3c0022aa),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b979),
	.w1(32'hbb4ca45e),
	.w2(32'h3b00ef41),
	.w3(32'h3b7a6499),
	.w4(32'h3c368a85),
	.w5(32'h3bf4ef79),
	.w6(32'hbc927322),
	.w7(32'h3b87f860),
	.w8(32'h3b21cabc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09f07a),
	.w1(32'h3bc544ea),
	.w2(32'h3bd37542),
	.w3(32'h3bbfc424),
	.w4(32'h3b950957),
	.w5(32'hba802db3),
	.w6(32'h3be8ed0d),
	.w7(32'hbb8dac03),
	.w8(32'h3c813483),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90de73),
	.w1(32'h3994d2dd),
	.w2(32'hba63cd02),
	.w3(32'h3c1afb3e),
	.w4(32'h3c51ecf4),
	.w5(32'hbb8ad2a3),
	.w6(32'h3c07693d),
	.w7(32'h3addca17),
	.w8(32'hbc2fa7da),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9b31e),
	.w1(32'h3bcea6f1),
	.w2(32'h39e79c11),
	.w3(32'h3b1da98a),
	.w4(32'hbb99ad7c),
	.w5(32'hbbe3a3d9),
	.w6(32'h3ac5313d),
	.w7(32'hbc0a159c),
	.w8(32'h3a1dd2d9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbca90),
	.w1(32'hbbca3032),
	.w2(32'h3bc014e7),
	.w3(32'hbc0c1ddc),
	.w4(32'hbae6d289),
	.w5(32'h3abd7604),
	.w6(32'hbca77d5a),
	.w7(32'hbc485b07),
	.w8(32'hbb3ed66f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b992ac9),
	.w1(32'h3aca8c05),
	.w2(32'hbb4a424c),
	.w3(32'h3a51d01d),
	.w4(32'h3a116269),
	.w5(32'hb9991ba3),
	.w6(32'hbac475a6),
	.w7(32'hbadb24c6),
	.w8(32'hbbc80ebc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf5d0f),
	.w1(32'h3c0ddf99),
	.w2(32'hbaaa1b4c),
	.w3(32'hbadeba1b),
	.w4(32'hb91b36e8),
	.w5(32'hbb155ab2),
	.w6(32'hbb8788ed),
	.w7(32'hbaf1431d),
	.w8(32'hbc090d8f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8baa),
	.w1(32'hbb071d87),
	.w2(32'h3d069f0c),
	.w3(32'hbb9e9d64),
	.w4(32'h3bf1badc),
	.w5(32'h3bcf00b4),
	.w6(32'hbbda9230),
	.w7(32'hbb9f0b40),
	.w8(32'h3d24d05c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5ac5f),
	.w1(32'h3c1f3ed0),
	.w2(32'hbb8f39ea),
	.w3(32'hbc0b8c7b),
	.w4(32'h3bbcd2de),
	.w5(32'hbc42e1c5),
	.w6(32'h3ccecbdf),
	.w7(32'h3c4481f0),
	.w8(32'h3c331255),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d9543),
	.w1(32'hbbdccf04),
	.w2(32'h3cbddd88),
	.w3(32'h3b6fb58f),
	.w4(32'h3c6651e5),
	.w5(32'h3c6b0b8c),
	.w6(32'h3c08782c),
	.w7(32'hbb4aca8f),
	.w8(32'h3c67f8eb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d89d),
	.w1(32'hbba84523),
	.w2(32'hbcb252ee),
	.w3(32'h3bb58aca),
	.w4(32'h3bd07f02),
	.w5(32'hbc99793d),
	.w6(32'h3c8d0052),
	.w7(32'hbbeb3a3a),
	.w8(32'hbb41da51),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9be6ac),
	.w1(32'hbc11c240),
	.w2(32'h3b108620),
	.w3(32'h3af96b3e),
	.w4(32'hb9bcb9e2),
	.w5(32'h3c09f3ae),
	.w6(32'h3c9c37ba),
	.w7(32'h3c9f45d2),
	.w8(32'hbcbe6740),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebee74),
	.w1(32'h3cb78b5b),
	.w2(32'h3c6523de),
	.w3(32'hbbe07d7f),
	.w4(32'h3c328ab3),
	.w5(32'h3c3069c3),
	.w6(32'hbc12ae67),
	.w7(32'hbcbaad87),
	.w8(32'hbb9e8706),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b9f90),
	.w1(32'hbb65c361),
	.w2(32'h3ae48a63),
	.w3(32'hbb4a0469),
	.w4(32'hbc8229e6),
	.w5(32'h3b4f962a),
	.w6(32'hbc929776),
	.w7(32'hbc06f0f5),
	.w8(32'hbc331af5),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d818d1a),
	.w1(32'hbc23e1a7),
	.w2(32'h3c28bfef),
	.w3(32'h3ca426ea),
	.w4(32'h3ce7c2e1),
	.w5(32'h3c354afd),
	.w6(32'h3cad751a),
	.w7(32'h3c82f59b),
	.w8(32'h3c9c840a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e90ba),
	.w1(32'h3c17fccb),
	.w2(32'h3bfc0d8f),
	.w3(32'hbaceea72),
	.w4(32'h3b62cae7),
	.w5(32'h3b6524d8),
	.w6(32'h3c61d040),
	.w7(32'h3c448a2c),
	.w8(32'h3ccb28fc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cac61),
	.w1(32'hbbd45015),
	.w2(32'h3b2d1750),
	.w3(32'hbbe6cac7),
	.w4(32'h3b419fb4),
	.w5(32'hbad6ec50),
	.w6(32'h3ae5bdce),
	.w7(32'hbaedfd8b),
	.w8(32'hba95adf3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eed69),
	.w1(32'h3b679974),
	.w2(32'h3ca75519),
	.w3(32'h3b43bf10),
	.w4(32'h3c6effb3),
	.w5(32'h3bd66e8b),
	.w6(32'h3be6117a),
	.w7(32'h3c689184),
	.w8(32'h3c9c167c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3af5b),
	.w1(32'hba9eb7d7),
	.w2(32'h3baba5cf),
	.w3(32'hbc71337d),
	.w4(32'h3b4020b0),
	.w5(32'h3baa552e),
	.w6(32'hbbbf29b2),
	.w7(32'h3c108d5e),
	.w8(32'hbcc5fcde),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26f6e0),
	.w1(32'hbae9b827),
	.w2(32'hbb8e6015),
	.w3(32'h3c62bd33),
	.w4(32'h3cf09c86),
	.w5(32'h3cb29ab4),
	.w6(32'h3cc0e66c),
	.w7(32'h3d113e49),
	.w8(32'h3d0b8b76),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d707c02),
	.w1(32'h3c8fd55a),
	.w2(32'hba0cf5e3),
	.w3(32'hbc6aeeb7),
	.w4(32'hbbeeaeba),
	.w5(32'h3be413ca),
	.w6(32'hbc9fc8c4),
	.w7(32'hbbb69206),
	.w8(32'hbcd0e6c6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6e9f66),
	.w1(32'hbc28a428),
	.w2(32'h3c0900dc),
	.w3(32'h3ba660bd),
	.w4(32'hbade724f),
	.w5(32'hbbe7ee19),
	.w6(32'hbbaf2515),
	.w7(32'hbc691ce3),
	.w8(32'hbb2be496),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a6cd8),
	.w1(32'h3b73efc0),
	.w2(32'hba5c8033),
	.w3(32'hbbf953c4),
	.w4(32'h3a932c42),
	.w5(32'hbae061a8),
	.w6(32'hbbd5753e),
	.w7(32'hbbc00dd4),
	.w8(32'hbbbdf08c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b128d87),
	.w1(32'h3b20d2b0),
	.w2(32'h3d250aef),
	.w3(32'hba8adbae),
	.w4(32'hbbecbd58),
	.w5(32'h3c505e66),
	.w6(32'hbbd608cb),
	.w7(32'hbcb6b26e),
	.w8(32'hbc67ffbe),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4c143e),
	.w1(32'h3c7259b3),
	.w2(32'h3bb7d08a),
	.w3(32'hbbba725d),
	.w4(32'h3c463c1b),
	.w5(32'h3c44fd7e),
	.w6(32'hbc4c85c6),
	.w7(32'h3b282488),
	.w8(32'hbc4919b1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2a496a),
	.w1(32'hbc888dae),
	.w2(32'hbc30c152),
	.w3(32'h3c32bb5b),
	.w4(32'h3c2622dd),
	.w5(32'h3cb536c8),
	.w6(32'h3c80e2a9),
	.w7(32'hbbf99e8a),
	.w8(32'h3c8242c5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd016d61),
	.w1(32'hbc490c16),
	.w2(32'h3a4b88a1),
	.w3(32'h3b84978c),
	.w4(32'hbbe84d3b),
	.w5(32'h3ae22335),
	.w6(32'h3cd31204),
	.w7(32'hbc4f7fd7),
	.w8(32'h3ac64e59),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42a996),
	.w1(32'h3adcb307),
	.w2(32'h3c128b81),
	.w3(32'hbb1293eb),
	.w4(32'hbc99d433),
	.w5(32'hbb5002f2),
	.w6(32'hbb74dc80),
	.w7(32'h38f77315),
	.w8(32'hbc6ac6fd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01ea00),
	.w1(32'h3bd1f39c),
	.w2(32'h3cf67201),
	.w3(32'h3982c473),
	.w4(32'hbc88a621),
	.w5(32'hbc5fa4d5),
	.w6(32'hba0afba6),
	.w7(32'hbca75912),
	.w8(32'hbcd74182),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39f5b1),
	.w1(32'hbc9547ea),
	.w2(32'hbc562a4b),
	.w3(32'hbcadb07d),
	.w4(32'h3c3c66b3),
	.w5(32'h3bfcaa0c),
	.w6(32'hbcad8154),
	.w7(32'h3cc96e43),
	.w8(32'h3ce781c8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b9964),
	.w1(32'h3bf247f4),
	.w2(32'h3cf53de9),
	.w3(32'h3bb77e3b),
	.w4(32'hbc77b48a),
	.w5(32'hbc3c482e),
	.w6(32'h3c5ad471),
	.w7(32'h3ba4a933),
	.w8(32'hbc35ee87),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f2409),
	.w1(32'hbccd2ca8),
	.w2(32'h3bb458d8),
	.w3(32'hbc5e141d),
	.w4(32'hbb28427b),
	.w5(32'h3b06ae12),
	.w6(32'hbc4b313f),
	.w7(32'hbc094265),
	.w8(32'hbbb31929),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88a3ab),
	.w1(32'h3bf87ae9),
	.w2(32'h3c97f6ee),
	.w3(32'h3c4620c1),
	.w4(32'h3a5f486a),
	.w5(32'h3c88f8d7),
	.w6(32'h3bc77bc7),
	.w7(32'hbbefc2af),
	.w8(32'h3d1a0773),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16434),
	.w1(32'h3afb410f),
	.w2(32'h3b54cd7e),
	.w3(32'hbc7faec5),
	.w4(32'h3b8e08ae),
	.w5(32'h3b41bcb2),
	.w6(32'h3beede15),
	.w7(32'hbc02e52c),
	.w8(32'hbc4a4ff7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9c50a),
	.w1(32'h3a0e7e0b),
	.w2(32'hbc84c10e),
	.w3(32'hbbd6e9d1),
	.w4(32'h3c39e23b),
	.w5(32'h3be5f072),
	.w6(32'hbc9efea2),
	.w7(32'hbba95cb0),
	.w8(32'h3cb7fbeb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0013b5),
	.w1(32'hbbaf2177),
	.w2(32'h3c092d05),
	.w3(32'h3c09e979),
	.w4(32'h3bc949a2),
	.w5(32'h3b4868d6),
	.w6(32'h3c983513),
	.w7(32'hbbc860a1),
	.w8(32'h3a86715f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b267),
	.w1(32'h3abc98f2),
	.w2(32'h3b31c592),
	.w3(32'hb93decbd),
	.w4(32'hbc86305a),
	.w5(32'hbc985b97),
	.w6(32'h3b58c663),
	.w7(32'h3cda09fa),
	.w8(32'hbc8c3d25),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08cabe),
	.w1(32'hbbddef1e),
	.w2(32'h3ca30170),
	.w3(32'hbb770cb4),
	.w4(32'hbbcc83de),
	.w5(32'hbbfb87dd),
	.w6(32'hbc80a35c),
	.w7(32'hbb2b57b0),
	.w8(32'h3aea249f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabde1b),
	.w1(32'hbc404d2b),
	.w2(32'hbb5710af),
	.w3(32'hbbda9417),
	.w4(32'hbcb1d015),
	.w5(32'h3b9adc47),
	.w6(32'h3b6eddfc),
	.w7(32'hbc837644),
	.w8(32'hbcf76154),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5e0359),
	.w1(32'h3ca5b326),
	.w2(32'h3cae0ec1),
	.w3(32'hba798058),
	.w4(32'hbb1f7c8b),
	.w5(32'hbc312157),
	.w6(32'h3bb50d9a),
	.w7(32'h3be6c630),
	.w8(32'hbc8ac363),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44d14d),
	.w1(32'hbd0a0c42),
	.w2(32'hbc509203),
	.w3(32'h3b6aaa3a),
	.w4(32'hbbf5b473),
	.w5(32'hbbd5a1c9),
	.w6(32'h3c380e31),
	.w7(32'hbbad07de),
	.w8(32'hbb2ddfba),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccc8d7),
	.w1(32'h3c595eec),
	.w2(32'hbc1ae266),
	.w3(32'h3b4c449e),
	.w4(32'hbd06e7d3),
	.w5(32'hbcc15bbf),
	.w6(32'hbc6e64f7),
	.w7(32'hbb3ee7c2),
	.w8(32'h3c25fb2f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74c782),
	.w1(32'hbca2d5b1),
	.w2(32'hbc664ac8),
	.w3(32'hbd3e0b97),
	.w4(32'h3c62b7db),
	.w5(32'h3bd20c48),
	.w6(32'hbce4717a),
	.w7(32'hbc142f1a),
	.w8(32'h3d61ad6d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd55152b),
	.w1(32'hbc699690),
	.w2(32'hbb8dbd31),
	.w3(32'hbc6d2cb8),
	.w4(32'h3c628030),
	.w5(32'h3b9c4ba6),
	.w6(32'h3d0bf716),
	.w7(32'hbbcd709b),
	.w8(32'hbd342f64),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c42a4),
	.w1(32'hbaa8d2c3),
	.w2(32'hbc87644d),
	.w3(32'h3cea56fb),
	.w4(32'h3c0ca69b),
	.w5(32'h3a6c8326),
	.w6(32'hbc2e2f86),
	.w7(32'h3ba85e45),
	.w8(32'h3c035ba5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb50736),
	.w1(32'h3bac7f57),
	.w2(32'hba91c7c7),
	.w3(32'hbbd3f10f),
	.w4(32'h3b4df54e),
	.w5(32'hbaace8b7),
	.w6(32'hbc23c322),
	.w7(32'hbc0579d4),
	.w8(32'hbbe56189),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d076),
	.w1(32'h3b2db400),
	.w2(32'hba19685c),
	.w3(32'hbb4b1da5),
	.w4(32'hbca1a761),
	.w5(32'hbc5badac),
	.w6(32'hbb66e43a),
	.w7(32'h3cbc8cc6),
	.w8(32'hbc59ceb3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9011d4),
	.w1(32'h3c456695),
	.w2(32'hbc89ab93),
	.w3(32'h3a2b5ca3),
	.w4(32'h3a47e4d9),
	.w5(32'hbc4794ec),
	.w6(32'hbce91813),
	.w7(32'h3b8bbb1b),
	.w8(32'h3c9f0ad5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc639380),
	.w1(32'hbc3953db),
	.w2(32'hbc38e3a7),
	.w3(32'hbc06e6fa),
	.w4(32'hbb765a47),
	.w5(32'hbb9f66e9),
	.w6(32'hbb456baf),
	.w7(32'hbc6b445d),
	.w8(32'hbbe8a449),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139a6b),
	.w1(32'hbb7f2fc3),
	.w2(32'h3b2a1df7),
	.w3(32'h3bdd72b5),
	.w4(32'hbb277e67),
	.w5(32'hbcaf1925),
	.w6(32'h3bc5d2b7),
	.w7(32'h3c1a7cae),
	.w8(32'h3ce55482),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c277),
	.w1(32'hbc270649),
	.w2(32'h3b044f42),
	.w3(32'hbc7f4a4b),
	.w4(32'h3ada5c18),
	.w5(32'hba01479f),
	.w6(32'h3bc596db),
	.w7(32'hbbdc8355),
	.w8(32'hbb17ce38),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab8994),
	.w1(32'h3b755803),
	.w2(32'h3b598281),
	.w3(32'hbac1ef80),
	.w4(32'h3bfe231e),
	.w5(32'hbbeb0762),
	.w6(32'h3ac43112),
	.w7(32'hba85e030),
	.w8(32'h3ccc346c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43f14e),
	.w1(32'h3b53fea8),
	.w2(32'h3b3a9acb),
	.w3(32'hbbf2ad95),
	.w4(32'h3af663ed),
	.w5(32'hbbefda04),
	.w6(32'h3be19b30),
	.w7(32'h3c0b6cae),
	.w8(32'h3cb0286e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad63b3e),
	.w1(32'h3bf2c9b0),
	.w2(32'hbbfce49c),
	.w3(32'hbc97ed78),
	.w4(32'hbb2f718f),
	.w5(32'hbb8c88c0),
	.w6(32'hbc9153d1),
	.w7(32'hbb14f9fc),
	.w8(32'hbba42545),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a61f6),
	.w1(32'hbc14a6cf),
	.w2(32'hbd001d20),
	.w3(32'hbb853cb8),
	.w4(32'h3c18587a),
	.w5(32'h3a3cd81f),
	.w6(32'h3ba48d8c),
	.w7(32'h3d21b822),
	.w8(32'h3c627253),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad45b6),
	.w1(32'h3c163866),
	.w2(32'h3badbf4d),
	.w3(32'h3c63bfd3),
	.w4(32'hbc25afc2),
	.w5(32'hbbd5116c),
	.w6(32'h3a1c7b92),
	.w7(32'hbb99716c),
	.w8(32'hbc366d40),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5bab910),
	.w1(32'h3acec2cf),
	.w2(32'hbc5b1774),
	.w3(32'hbb8b0af2),
	.w4(32'hbc261eb7),
	.w5(32'hbc1fe957),
	.w6(32'hbcdc61fc),
	.w7(32'hbc96940f),
	.w8(32'hba6a3407),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcfea9),
	.w1(32'hbbeb3996),
	.w2(32'hbcdf4046),
	.w3(32'hbc82b4fa),
	.w4(32'h3cb4d484),
	.w5(32'h3c3323e8),
	.w6(32'hbb92a48a),
	.w7(32'h3bdfc1ed),
	.w8(32'h3ccd9e34),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd209d3b),
	.w1(32'hbc0d9f2b),
	.w2(32'hbc8653c3),
	.w3(32'hbbc1709c),
	.w4(32'h3bafa50c),
	.w5(32'hba3e2469),
	.w6(32'h3c9588a3),
	.w7(32'h3ceb076a),
	.w8(32'h3b665bae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce35b37),
	.w1(32'hbc555a5b),
	.w2(32'hbc71d6a5),
	.w3(32'hba108c04),
	.w4(32'h3c4eb174),
	.w5(32'h3c812c05),
	.w6(32'h3c4cccbe),
	.w7(32'hbce7b42e),
	.w8(32'hbc66351f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee97f8),
	.w1(32'h3c18d45e),
	.w2(32'h3b35b80e),
	.w3(32'h3cb00d62),
	.w4(32'hbc8cf7c7),
	.w5(32'hbc3b6362),
	.w6(32'h3b2926e9),
	.w7(32'hbb0aacca),
	.w8(32'hbb4df83a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda7698),
	.w1(32'hbc2ac4f3),
	.w2(32'hbca54f29),
	.w3(32'h3a1ad2e4),
	.w4(32'h3cc4973a),
	.w5(32'h3cb2446e),
	.w6(32'hbbda5d29),
	.w7(32'h3c40b78f),
	.w8(32'h3c48786c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5cc63c),
	.w1(32'hbb8a14be),
	.w2(32'h3bea710e),
	.w3(32'h3c1e2eb1),
	.w4(32'hb80e90c7),
	.w5(32'h3c816355),
	.w6(32'h3ccee6f1),
	.w7(32'hbbcf5e2f),
	.w8(32'h3cc6ed41),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b2f52),
	.w1(32'h3cc6c305),
	.w2(32'hbc00fed1),
	.w3(32'h3cb7fa0c),
	.w4(32'h3b36ae66),
	.w5(32'hb9eb2fa8),
	.w6(32'h3d0da98b),
	.w7(32'h3cb723ac),
	.w8(32'h3ba3e380),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36b409),
	.w1(32'hbc47ca04),
	.w2(32'h3c6f9420),
	.w3(32'hbc782152),
	.w4(32'hbc543c5c),
	.w5(32'h3b190c83),
	.w6(32'hbc594e29),
	.w7(32'hbc377680),
	.w8(32'hbb8b826b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca43ec6),
	.w1(32'h3c7abd42),
	.w2(32'hbd05ac95),
	.w3(32'hbaf622af),
	.w4(32'h3caeeac4),
	.w5(32'h3cd5d244),
	.w6(32'hbc18bd7f),
	.w7(32'hbc71e6c2),
	.w8(32'h3d72716d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd62857b),
	.w1(32'h3cba8a79),
	.w2(32'h3c0f0590),
	.w3(32'h3a262bd3),
	.w4(32'hbc6f1d76),
	.w5(32'hbbd952ab),
	.w6(32'h3d07b2b8),
	.w7(32'hbb442592),
	.w8(32'hbd12381a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4751b2),
	.w1(32'hbc1561eb),
	.w2(32'hbcaa986f),
	.w3(32'h3c26e2cf),
	.w4(32'hba1f4cf5),
	.w5(32'hbc0e2672),
	.w6(32'hbb0c983d),
	.w7(32'h3abbd7f7),
	.w8(32'hbae4b1cb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c9007),
	.w1(32'hbc04d794),
	.w2(32'hbadc9a3a),
	.w3(32'hbbd88c52),
	.w4(32'h39ab7600),
	.w5(32'hba05a75b),
	.w6(32'hbb0ff827),
	.w7(32'h3ae40a53),
	.w8(32'hbb9ca53f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8fd33),
	.w1(32'h3b23d752),
	.w2(32'hbb47672e),
	.w3(32'h3c310b89),
	.w4(32'h3c26cb8a),
	.w5(32'hbb577dab),
	.w6(32'h3c2f5dda),
	.w7(32'h3c5a5aae),
	.w8(32'hbbc44a76),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15addf),
	.w1(32'hbb05ae56),
	.w2(32'h3a9c5128),
	.w3(32'h3a6b0dc0),
	.w4(32'h3ba5898f),
	.w5(32'hbaff421f),
	.w6(32'hbb11bb3c),
	.w7(32'h3b92c313),
	.w8(32'hbba47a34),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db3b5),
	.w1(32'hba14a5e3),
	.w2(32'h3bbe4fed),
	.w3(32'h3af91290),
	.w4(32'h3c0d012a),
	.w5(32'hbb6ce9ee),
	.w6(32'hbb222ab5),
	.w7(32'hbcccf8c1),
	.w8(32'hbad1dc36),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39980bf4),
	.w1(32'hbca8456c),
	.w2(32'hbb4fd058),
	.w3(32'hbc074d0e),
	.w4(32'h3bbace3c),
	.w5(32'h3ba15ec7),
	.w6(32'h3bf69d15),
	.w7(32'hbbbdbd89),
	.w8(32'hbc5d170a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70b644),
	.w1(32'hbadb4259),
	.w2(32'h39745a48),
	.w3(32'h3bfbcaea),
	.w4(32'hbbd93de6),
	.w5(32'hbc40b351),
	.w6(32'h3c47fcf7),
	.w7(32'h3c86ec2a),
	.w8(32'h3d2a14a2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc9c1e4),
	.w1(32'h3cafa897),
	.w2(32'h3b9caca5),
	.w3(32'h3cce543b),
	.w4(32'h3ca4b033),
	.w5(32'h3ac61866),
	.w6(32'h3b9f1b23),
	.w7(32'h3c180d88),
	.w8(32'h3c29e692),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94f9a),
	.w1(32'h3b7cffe4),
	.w2(32'hbc02db19),
	.w3(32'h3c13e1ea),
	.w4(32'hbc1e54c0),
	.w5(32'hbc7353d4),
	.w6(32'h3c503f27),
	.w7(32'h3c952864),
	.w8(32'h3c0ebaa6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91c5d8),
	.w1(32'h3c8635b7),
	.w2(32'h3b19db8e),
	.w3(32'h3ce08996),
	.w4(32'h3d08fd25),
	.w5(32'h3ac9a633),
	.w6(32'h3aa74410),
	.w7(32'h3cdc527b),
	.w8(32'h3cd15802),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dda66),
	.w1(32'hbc16a8f7),
	.w2(32'h3b76ed92),
	.w3(32'h3c07152d),
	.w4(32'h3c2f10f5),
	.w5(32'h3b7bde2c),
	.w6(32'h3cae2888),
	.w7(32'h3c3b7f5d),
	.w8(32'hbc1c02cf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536a09),
	.w1(32'hbb9834f3),
	.w2(32'hbc9baa97),
	.w3(32'hbbb9735a),
	.w4(32'h3c3fb9df),
	.w5(32'h3c6891ff),
	.w6(32'hbacd73bf),
	.w7(32'hbc4edc3c),
	.w8(32'hbbee12c1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c8851),
	.w1(32'hbb9fc95c),
	.w2(32'h3b912609),
	.w3(32'h3ba0e509),
	.w4(32'h3bdd9e97),
	.w5(32'h3b682ffb),
	.w6(32'hbc9cc71c),
	.w7(32'h3bbc238e),
	.w8(32'hbc1642a9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b230e5f),
	.w1(32'hba7b7b87),
	.w2(32'hbab13d8e),
	.w3(32'h3ad20d56),
	.w4(32'h3bc6155c),
	.w5(32'hbb934fa0),
	.w6(32'hbbd49066),
	.w7(32'hbb8991d2),
	.w8(32'h3bcb0ead),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc70a),
	.w1(32'h3c05411e),
	.w2(32'hbc181ede),
	.w3(32'h3baf9d48),
	.w4(32'h3bf41eb7),
	.w5(32'hbbb5288f),
	.w6(32'h39ed8507),
	.w7(32'h3aefd87f),
	.w8(32'h3cb28ded),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c5eb3),
	.w1(32'h3b5253f7),
	.w2(32'hbc82bc9a),
	.w3(32'h3c9d43e9),
	.w4(32'h3b1ed175),
	.w5(32'h3986e10a),
	.w6(32'hbc2994c9),
	.w7(32'h3bab2fb4),
	.w8(32'h3cf7df46),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb657bff),
	.w1(32'h3bdd154c),
	.w2(32'h3cbbdea9),
	.w3(32'hbbef8962),
	.w4(32'hbbd9e703),
	.w5(32'hbc90d0ae),
	.w6(32'hbba64839),
	.w7(32'hbcdff27f),
	.w8(32'h3d2854f8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a000b3f),
	.w1(32'hbcb8605c),
	.w2(32'h3c6e0600),
	.w3(32'h3c6a1a67),
	.w4(32'h3c0b0ee5),
	.w5(32'h3c81a983),
	.w6(32'h3c8952a6),
	.w7(32'h3ca834d7),
	.w8(32'hbba025ff),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2b76c),
	.w1(32'h3c25cd22),
	.w2(32'h3bed039c),
	.w3(32'h3b538371),
	.w4(32'hbb8ef90c),
	.w5(32'h3cc0e6f7),
	.w6(32'h3c8754b4),
	.w7(32'h3a14d366),
	.w8(32'hbd8808eb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ed52a),
	.w1(32'hbcb7e479),
	.w2(32'h3b0048ea),
	.w3(32'hbc9dc107),
	.w4(32'h3b494fd0),
	.w5(32'h38f23a4c),
	.w6(32'h3cdf8206),
	.w7(32'h3bcd6d3f),
	.w8(32'hb9883b50),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e62ac),
	.w1(32'hb95d9777),
	.w2(32'hbb08abbc),
	.w3(32'h3b9831af),
	.w4(32'hbb96ec60),
	.w5(32'hbcb695b8),
	.w6(32'h3ad22817),
	.w7(32'hbc497870),
	.w8(32'hbcb8c979),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e72f),
	.w1(32'hbced8c34),
	.w2(32'hbbc528ce),
	.w3(32'h3ca5e0ad),
	.w4(32'h3c8ad438),
	.w5(32'h3cf5d52d),
	.w6(32'hbae53bd4),
	.w7(32'h3ca70ff8),
	.w8(32'hbcfe6bb0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25fc48),
	.w1(32'h3c8dacf6),
	.w2(32'h3c10bda6),
	.w3(32'hbc057192),
	.w4(32'hbbc336ce),
	.w5(32'hbc0b2f15),
	.w6(32'h3c40e2a0),
	.w7(32'h3c41e48e),
	.w8(32'h3d108214),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce38e53),
	.w1(32'hba4b2daa),
	.w2(32'h3c15a29f),
	.w3(32'h3c460b62),
	.w4(32'h3b8d555b),
	.w5(32'h3a80da97),
	.w6(32'hbc62ce11),
	.w7(32'h3b2da560),
	.w8(32'hbc0ab3c7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95960e),
	.w1(32'h3a25b9ba),
	.w2(32'h3ac0536d),
	.w3(32'h3b097a70),
	.w4(32'h3b629a65),
	.w5(32'h3c13f9a5),
	.w6(32'hbadb3086),
	.w7(32'hbbd5cd8f),
	.w8(32'hbc682126),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6d791),
	.w1(32'h3c005d66),
	.w2(32'h3a854880),
	.w3(32'hbaa4a1c6),
	.w4(32'hbbe857f4),
	.w5(32'hbbf37eeb),
	.w6(32'hbc22f0f7),
	.w7(32'hb9e92869),
	.w8(32'hbb15e92f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80b422),
	.w1(32'h3b2f7f1e),
	.w2(32'hbb95636b),
	.w3(32'hbbfc07b8),
	.w4(32'h3b5703a0),
	.w5(32'h3b5b0635),
	.w6(32'hbae453b6),
	.w7(32'h3b6eaa87),
	.w8(32'hbc3a2df9),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05bed0),
	.w1(32'h3baeaf1c),
	.w2(32'hbbc678ea),
	.w3(32'h3b96e6ae),
	.w4(32'hbb5183bf),
	.w5(32'hbb7c9b52),
	.w6(32'h3c1f39ef),
	.w7(32'h3beddafd),
	.w8(32'hbc131c3d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a69f2),
	.w1(32'hbb30b709),
	.w2(32'hb90b9b59),
	.w3(32'h3c340a43),
	.w4(32'h3c358719),
	.w5(32'h3bcbe78a),
	.w6(32'hbbe8448c),
	.w7(32'h3ba7241a),
	.w8(32'hbb9ae912),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032eb2),
	.w1(32'h3b39c551),
	.w2(32'hba84810e),
	.w3(32'hbb3b90f2),
	.w4(32'hb8f6df67),
	.w5(32'hbc597e12),
	.w6(32'hbb78b089),
	.w7(32'hbbb9a356),
	.w8(32'h3c14e668),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22cd86),
	.w1(32'h3c4d5bbf),
	.w2(32'h3c008f44),
	.w3(32'h3c44a4c5),
	.w4(32'h3cc3c6d2),
	.w5(32'h3bbb0c2a),
	.w6(32'hbb1998fa),
	.w7(32'hbcbd9474),
	.w8(32'h3d7ffa9e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922d65),
	.w1(32'h3b0871b9),
	.w2(32'hbcd99582),
	.w3(32'h3bdeaff7),
	.w4(32'h3c4eaf51),
	.w5(32'h3d05b66c),
	.w6(32'h3c4bea04),
	.w7(32'h3d505aa1),
	.w8(32'hbdbe5663),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7be09b),
	.w1(32'h3bdd9937),
	.w2(32'h3a4bb5f4),
	.w3(32'hbc547bb8),
	.w4(32'h3b15b955),
	.w5(32'h3b0d2796),
	.w6(32'h3c0ad3b2),
	.w7(32'h3b3a470e),
	.w8(32'hbb59311f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e5972),
	.w1(32'hba827937),
	.w2(32'hbab20b55),
	.w3(32'hbba3c9df),
	.w4(32'hbb8b9211),
	.w5(32'h3bafde0a),
	.w6(32'hbb087cef),
	.w7(32'hbb590a3b),
	.w8(32'hbc9fe63b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07ebfe),
	.w1(32'hbbeaa2ab),
	.w2(32'hbc14ee55),
	.w3(32'hbb7ca089),
	.w4(32'h3c0ad481),
	.w5(32'h3cf58576),
	.w6(32'hbc07e1d8),
	.w7(32'h3c3d9907),
	.w8(32'hbd623f2b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc88bdf),
	.w1(32'h3ad50f19),
	.w2(32'h3b271c57),
	.w3(32'hbc02ae4d),
	.w4(32'h3c3b6cf8),
	.w5(32'h3c01f46b),
	.w6(32'h3bf60e96),
	.w7(32'h3c97e424),
	.w8(32'hbc31830f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50453d),
	.w1(32'h3bd6d266),
	.w2(32'h3bb0de14),
	.w3(32'h3c077bd6),
	.w4(32'h3b384171),
	.w5(32'h3cb4e69e),
	.w6(32'hbbc13183),
	.w7(32'h3c0958a0),
	.w8(32'hbc9cc8a3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6eaff),
	.w1(32'h3b0a868a),
	.w2(32'h3b616901),
	.w3(32'hba9b8519),
	.w4(32'hbc6308d4),
	.w5(32'hbc638855),
	.w6(32'h3c7c4884),
	.w7(32'hbcc8406c),
	.w8(32'h3d5811cf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd222d56),
	.w1(32'h3b3e10ae),
	.w2(32'hbc80302e),
	.w3(32'hbc82fd06),
	.w4(32'hbc479196),
	.w5(32'hbc535b30),
	.w6(32'h3b7c3313),
	.w7(32'hbc71b0a9),
	.w8(32'h3c78b8e0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc869dab),
	.w1(32'hbccbc78a),
	.w2(32'h3cc6f8ef),
	.w3(32'hbc0a7b15),
	.w4(32'h3bb3d18c),
	.w5(32'h3b8e4d47),
	.w6(32'hbc311512),
	.w7(32'hbc18c6d7),
	.w8(32'h3b2983f6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8dea6),
	.w1(32'hbb9a1991),
	.w2(32'hbc13c2ac),
	.w3(32'hbbb89b79),
	.w4(32'hbbf024f3),
	.w5(32'hbbdc952f),
	.w6(32'h3ca6d0a4),
	.w7(32'h3c5f3ab2),
	.w8(32'hbb4bc51a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b363),
	.w1(32'hbbd9a78c),
	.w2(32'h3bd29831),
	.w3(32'hbc40015f),
	.w4(32'hbbc36ee3),
	.w5(32'hbcb30b09),
	.w6(32'h3c4ba4be),
	.w7(32'hbb9b2ff1),
	.w8(32'h3c170af5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc60cc6),
	.w1(32'hbb4e9a7e),
	.w2(32'h3aec2bd2),
	.w3(32'h3ba0bf2c),
	.w4(32'h378e54dd),
	.w5(32'h3a1104ef),
	.w6(32'hbb276aba),
	.w7(32'h3a83a71d),
	.w8(32'hbb15c68b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d9abb),
	.w1(32'hbb3350a3),
	.w2(32'hbc6f60c3),
	.w3(32'hb92a34bf),
	.w4(32'hbbc7df90),
	.w5(32'hbb0aab9c),
	.w6(32'hbb0a370f),
	.w7(32'hbb996b04),
	.w8(32'hbcb80b77),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c4b4),
	.w1(32'hbbbf0e0b),
	.w2(32'hbb3d5d1e),
	.w3(32'hbc998575),
	.w4(32'hbb921b88),
	.w5(32'h3a32dd68),
	.w6(32'h3bef5d4d),
	.w7(32'hbc0afa0d),
	.w8(32'hbc12309e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26551f),
	.w1(32'hbc0cea89),
	.w2(32'hbb103f1e),
	.w3(32'h3af292d1),
	.w4(32'h3b6abc9f),
	.w5(32'hbb9ed40f),
	.w6(32'hbbba7c85),
	.w7(32'h3b72cb7c),
	.w8(32'h3c363836),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa10bb),
	.w1(32'hbae68188),
	.w2(32'h3c4ea1c2),
	.w3(32'hba311180),
	.w4(32'hbc054f19),
	.w5(32'hbb61f693),
	.w6(32'h3c3c2238),
	.w7(32'hbbb63d1b),
	.w8(32'hbb729314),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceeb5db),
	.w1(32'hbc425801),
	.w2(32'hbaab8c5b),
	.w3(32'hbc348ed3),
	.w4(32'hbb61ec70),
	.w5(32'hbacb4db3),
	.w6(32'h3c53beea),
	.w7(32'hbb1d3755),
	.w8(32'hbbcac047),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae36572),
	.w1(32'hbb2b0c45),
	.w2(32'hbcd77cf2),
	.w3(32'hba905840),
	.w4(32'hbc3661ad),
	.w5(32'hbc8a5bdc),
	.w6(32'hbb03a8cf),
	.w7(32'h3d006ecc),
	.w8(32'h3d25e815),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6b2e3),
	.w1(32'h3c1e6082),
	.w2(32'hbc2497a2),
	.w3(32'h3c734fb4),
	.w4(32'hbc27ad1c),
	.w5(32'hbc18e3c1),
	.w6(32'hbd8b05af),
	.w7(32'h3a33def1),
	.w8(32'h3cb58a52),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842515),
	.w1(32'h3aa4dfb2),
	.w2(32'h3bff028a),
	.w3(32'h3c3dcc8a),
	.w4(32'h3b74dc6b),
	.w5(32'h3b9e90a1),
	.w6(32'hbcaef445),
	.w7(32'h3bcfd7cb),
	.w8(32'h39921068),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5a6ef),
	.w1(32'h3bab30f9),
	.w2(32'h3bb8fc3b),
	.w3(32'h3b875ebb),
	.w4(32'hbbb58373),
	.w5(32'h3ba589f4),
	.w6(32'h3927332f),
	.w7(32'h3bddf135),
	.w8(32'hbc13847f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeafec),
	.w1(32'hbb2afbca),
	.w2(32'hbaa42ab2),
	.w3(32'hbb46a979),
	.w4(32'hba592ed3),
	.w5(32'hbb7a034e),
	.w6(32'h3c2b506b),
	.w7(32'h3c923ff4),
	.w8(32'hbbe16d38),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule