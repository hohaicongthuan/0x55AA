module layer_10_featuremap_264(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4014f),
	.w1(32'hbc416969),
	.w2(32'hbc2379aa),
	.w3(32'h3c0e9131),
	.w4(32'h3a4f7512),
	.w5(32'h3bac4efc),
	.w6(32'h3baafc19),
	.w7(32'hbb34b0ae),
	.w8(32'h3790e9bf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bae25),
	.w1(32'hbc5985ca),
	.w2(32'hbbd52638),
	.w3(32'h3c8483fe),
	.w4(32'h3b89c1a1),
	.w5(32'hb98170c5),
	.w6(32'hbbec8f68),
	.w7(32'h3c1ecf24),
	.w8(32'hbaaf61ae),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90460e),
	.w1(32'hbb1f0383),
	.w2(32'h3bc5fe8c),
	.w3(32'hbc252a64),
	.w4(32'hbb466e3b),
	.w5(32'hbc0cf0d5),
	.w6(32'hbb424266),
	.w7(32'h3b79a2d3),
	.w8(32'h3c05a599),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0315b5),
	.w1(32'h3bcffbf7),
	.w2(32'h3acbfc3b),
	.w3(32'hbb8a9f2a),
	.w4(32'hbc3ae8e8),
	.w5(32'hbbef8c72),
	.w6(32'h3b6e6c5f),
	.w7(32'hba46702a),
	.w8(32'hbd24d466),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ec8d),
	.w1(32'h3c84304e),
	.w2(32'hbc128c94),
	.w3(32'hb9e6c6b1),
	.w4(32'h3b805897),
	.w5(32'hbbb212db),
	.w6(32'hbd1e0757),
	.w7(32'hbd31c59a),
	.w8(32'hbaf71109),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37c1e6),
	.w1(32'hbc912d09),
	.w2(32'hbc4cc9bf),
	.w3(32'h3beeab57),
	.w4(32'hbb8f85d9),
	.w5(32'h3b56211d),
	.w6(32'hbb4a22c6),
	.w7(32'hbb115ed2),
	.w8(32'hba10f1b1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb697b31),
	.w1(32'hbc4ae516),
	.w2(32'hbbd98432),
	.w3(32'h3beb02af),
	.w4(32'h3b7d6fb3),
	.w5(32'hbc0097cd),
	.w6(32'hbbb54ff7),
	.w7(32'h3b36c0c6),
	.w8(32'hbbba76ac),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7710b1),
	.w1(32'hbc52c371),
	.w2(32'hbc6f2d08),
	.w3(32'h3c427ada),
	.w4(32'h3b63e9b8),
	.w5(32'hbb9da392),
	.w6(32'hbb300a85),
	.w7(32'hba969f6f),
	.w8(32'hbc146108),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fea5d),
	.w1(32'hbcd65a94),
	.w2(32'hbc8a1484),
	.w3(32'h3cdf8a25),
	.w4(32'h3c6cff86),
	.w5(32'hbbf163c9),
	.w6(32'h3c014160),
	.w7(32'h3c0fea4d),
	.w8(32'hb960e8ac),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d7ded),
	.w1(32'hbb56d6bd),
	.w2(32'hba33b61d),
	.w3(32'h3b9b165b),
	.w4(32'hbb5c022f),
	.w5(32'h3c348eed),
	.w6(32'hbc0e3604),
	.w7(32'h3a8ba1bf),
	.w8(32'h3ba9a1cc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189913),
	.w1(32'hbb37a3b4),
	.w2(32'hbaf79f99),
	.w3(32'h3c3b81cf),
	.w4(32'h3ae146eb),
	.w5(32'h3bad4f20),
	.w6(32'hbaf34602),
	.w7(32'hb8681e4b),
	.w8(32'h398e4c24),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60304),
	.w1(32'hbb6bb36e),
	.w2(32'hbb85def3),
	.w3(32'hbb2613e9),
	.w4(32'h3a7888a2),
	.w5(32'h3b22bd4a),
	.w6(32'h3c3d44df),
	.w7(32'h3b820077),
	.w8(32'hbc253399),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc584201),
	.w1(32'hbc2e977b),
	.w2(32'h3b606ed3),
	.w3(32'h3cc6f361),
	.w4(32'h3cb8a710),
	.w5(32'h3c8ae16f),
	.w6(32'hbc258644),
	.w7(32'hbb12dbe3),
	.w8(32'h3acf8f01),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc06d7),
	.w1(32'h3b96812c),
	.w2(32'h3ba47ca1),
	.w3(32'h3c869675),
	.w4(32'h3bd65a06),
	.w5(32'h3b2c1c11),
	.w6(32'h3c321255),
	.w7(32'h3bd6bde6),
	.w8(32'h3bcc9cec),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfad157),
	.w1(32'hbbba95a3),
	.w2(32'h3bb20268),
	.w3(32'h3c242e7a),
	.w4(32'h3bc8a1e6),
	.w5(32'h3c30bd60),
	.w6(32'h3b1cd3ed),
	.w7(32'h39953cc5),
	.w8(32'hbb3f3644),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2184bf),
	.w1(32'hbbbb4592),
	.w2(32'h3a227ec1),
	.w3(32'h3ce21cdd),
	.w4(32'h3c432883),
	.w5(32'h3c9b43df),
	.w6(32'hbbd907e6),
	.w7(32'h3be41f5f),
	.w8(32'hb82e808f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32a680),
	.w1(32'hbce3f973),
	.w2(32'hbc479eb1),
	.w3(32'h3cdd4840),
	.w4(32'h3c5182d4),
	.w5(32'hbbd0b32b),
	.w6(32'hbb85ce2f),
	.w7(32'hbb8e0396),
	.w8(32'h3b467c68),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f633),
	.w1(32'h3bc5554a),
	.w2(32'hbbebc13c),
	.w3(32'hbc691589),
	.w4(32'hbc7ad231),
	.w5(32'hbcd1efd1),
	.w6(32'hbc0d158b),
	.w7(32'hbc46807b),
	.w8(32'hbcc61946),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14dfd6),
	.w1(32'h3ce39197),
	.w2(32'hba76bbeb),
	.w3(32'hbca12d7d),
	.w4(32'hbc7860d9),
	.w5(32'hbbcf0f7a),
	.w6(32'hbc6dfec2),
	.w7(32'hbc43c480),
	.w8(32'hbb811987),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b23dc),
	.w1(32'hb8dd1674),
	.w2(32'hbb886a9f),
	.w3(32'hbc17edbe),
	.w4(32'hbb71565a),
	.w5(32'h3941414c),
	.w6(32'h3c03a0b0),
	.w7(32'hbaaafd2e),
	.w8(32'h3a102576),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b527d),
	.w1(32'hbc06a297),
	.w2(32'hbc71909b),
	.w3(32'h3c7b0ed3),
	.w4(32'h3bad4e9a),
	.w5(32'h3b1bbe7c),
	.w6(32'hba89c053),
	.w7(32'hbb0e6515),
	.w8(32'h3b4eb9cd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bb641),
	.w1(32'h3b959ec6),
	.w2(32'h3b0214d6),
	.w3(32'h3ab0c483),
	.w4(32'hbb68324e),
	.w5(32'hbb139219),
	.w6(32'h3b58cb2f),
	.w7(32'h3b5545c0),
	.w8(32'hba18507f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e6d29),
	.w1(32'hbc7c3fbd),
	.w2(32'hbc9fa767),
	.w3(32'hbc98ba72),
	.w4(32'hbc4aedb0),
	.w5(32'hbc59675f),
	.w6(32'hbca3627e),
	.w7(32'hbba50202),
	.w8(32'hbcb25bb2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35c8c1),
	.w1(32'hbc154ee1),
	.w2(32'h3b896577),
	.w3(32'h3d0bfd7e),
	.w4(32'h3be6e761),
	.w5(32'h3b4fc035),
	.w6(32'hbb75deb3),
	.w7(32'h3c11db44),
	.w8(32'hb9a22eb0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801fd4),
	.w1(32'h3c2260aa),
	.w2(32'h3c404240),
	.w3(32'hbb602d2e),
	.w4(32'h3bc1f498),
	.w5(32'h3c35078a),
	.w6(32'h3c4d77fb),
	.w7(32'hbaa98b9c),
	.w8(32'h3c53e363),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc434),
	.w1(32'hbc2ae507),
	.w2(32'h3b26e876),
	.w3(32'h3c144129),
	.w4(32'hbab4bc24),
	.w5(32'h3b2e3e8f),
	.w6(32'h3ba6de63),
	.w7(32'h3be109ca),
	.w8(32'h3b28a0ed),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13ac9f),
	.w1(32'h3b259e67),
	.w2(32'h3b5b9465),
	.w3(32'h3c16833b),
	.w4(32'h3bb50db1),
	.w5(32'hb9f08f6d),
	.w6(32'h3bf1d197),
	.w7(32'h3b386391),
	.w8(32'hbc11712d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53aa51),
	.w1(32'hbcc9ea0f),
	.w2(32'hbc8f32a7),
	.w3(32'h3c50a502),
	.w4(32'hbb94e9d7),
	.w5(32'h3b8c392f),
	.w6(32'hbb3fe179),
	.w7(32'hbbe81f13),
	.w8(32'h3c097076),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f9cc6),
	.w1(32'h3bbeb00c),
	.w2(32'hbbb1da75),
	.w3(32'hbc21a02d),
	.w4(32'hbb1e5bf5),
	.w5(32'h3bb7ce39),
	.w6(32'h3c5eaa9e),
	.w7(32'hbb83f2dd),
	.w8(32'h3a23ef42),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba62a11),
	.w1(32'hbb039946),
	.w2(32'h3b347bb7),
	.w3(32'h3ca80c7d),
	.w4(32'h3c7ce946),
	.w5(32'h3c823e99),
	.w6(32'hbb30decb),
	.w7(32'h3c23f90f),
	.w8(32'hb97e6111),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69e7f5),
	.w1(32'hba788033),
	.w2(32'hbbb8e382),
	.w3(32'hb820031b),
	.w4(32'h3c1a41b9),
	.w5(32'h3b5d8638),
	.w6(32'hbbb13a68),
	.w7(32'hbbd3a6ac),
	.w8(32'hbc230041),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad77384),
	.w1(32'hbb9da9e2),
	.w2(32'hbbdf2695),
	.w3(32'hbaa6061f),
	.w4(32'hba854a39),
	.w5(32'hb9d7777b),
	.w6(32'h3bb75d29),
	.w7(32'hbcaf3450),
	.w8(32'hbab662b8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926156),
	.w1(32'h3c0f3837),
	.w2(32'h3c325e00),
	.w3(32'hbbfc3260),
	.w4(32'hbbdf7028),
	.w5(32'h3aba189b),
	.w6(32'hbca61bd7),
	.w7(32'hbb655bc1),
	.w8(32'h3b8de8e3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a336),
	.w1(32'h3b924e1c),
	.w2(32'h3bcb97e6),
	.w3(32'hbba2ad64),
	.w4(32'hbc021003),
	.w5(32'hbb991f9b),
	.w6(32'hbad3395c),
	.w7(32'hbb582745),
	.w8(32'h3b43f54c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f8464),
	.w1(32'hbbe22084),
	.w2(32'hbc37e26d),
	.w3(32'hbbe63e69),
	.w4(32'h3b342a09),
	.w5(32'hbb897ab7),
	.w6(32'h3c5da8a7),
	.w7(32'hbb77eed8),
	.w8(32'hbbf8b6da),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2066a2),
	.w1(32'hbbda3a8d),
	.w2(32'hbb6241a2),
	.w3(32'hbb571ac7),
	.w4(32'hbb8c6843),
	.w5(32'h39a79b37),
	.w6(32'hbbd4554e),
	.w7(32'h3a948a80),
	.w8(32'hbbdfce84),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc7e72),
	.w1(32'h3c4aa65d),
	.w2(32'hbbb8c3cc),
	.w3(32'hbcb1ce94),
	.w4(32'h3be2c580),
	.w5(32'hb9c6f218),
	.w6(32'hbc77ad21),
	.w7(32'hbc78b6dd),
	.w8(32'h3bbde04b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f42d2),
	.w1(32'h3c7f8286),
	.w2(32'h3c4fa35a),
	.w3(32'h3a669ee6),
	.w4(32'hbb9d4f7c),
	.w5(32'h3c2dabed),
	.w6(32'h3b89b260),
	.w7(32'h3b63be3c),
	.w8(32'h3c13979f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f71e),
	.w1(32'hbba88ae9),
	.w2(32'hbadbd4a5),
	.w3(32'h3c6514b1),
	.w4(32'h3c04e630),
	.w5(32'hbb5e1e0c),
	.w6(32'h3c56d101),
	.w7(32'hba46d8de),
	.w8(32'h3cac5c09),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce93569),
	.w1(32'h3d821421),
	.w2(32'h3c30b457),
	.w3(32'hbd29954f),
	.w4(32'hbcb15c53),
	.w5(32'h3ad28094),
	.w6(32'hbb59b72c),
	.w7(32'hbc6b9ac1),
	.w8(32'hba833410),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8971a3),
	.w1(32'hbc113e41),
	.w2(32'hbb62b4e1),
	.w3(32'hbb838740),
	.w4(32'hbb666a8a),
	.w5(32'h3a1851ae),
	.w6(32'hbc175b3a),
	.w7(32'hbc1970c7),
	.w8(32'hb9b906b1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf0931),
	.w1(32'hbb85ae7c),
	.w2(32'h3b8b97ae),
	.w3(32'h3c0c7ba3),
	.w4(32'hbb8a284f),
	.w5(32'hbae5753b),
	.w6(32'hbb22a15c),
	.w7(32'h3b886592),
	.w8(32'hba3fe77e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0897d6),
	.w1(32'h3c8c0f47),
	.w2(32'h3acedf4b),
	.w3(32'hbbfd3094),
	.w4(32'hbb20f6b1),
	.w5(32'h3c870379),
	.w6(32'hbc75ec62),
	.w7(32'hbc18cb8f),
	.w8(32'hbac120d3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8248b0),
	.w1(32'hbcc10b01),
	.w2(32'h3bbc19f1),
	.w3(32'h3d0afe58),
	.w4(32'h3ceadc8d),
	.w5(32'hbadfd707),
	.w6(32'hbc2c544f),
	.w7(32'h3c95374a),
	.w8(32'h3c4a36f4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b570f),
	.w1(32'h3d3a9424),
	.w2(32'h3ca5cd3b),
	.w3(32'hbd0cdae2),
	.w4(32'hbcbe3764),
	.w5(32'h3c4a0c5b),
	.w6(32'hbc74b5a8),
	.w7(32'hbc485131),
	.w8(32'h3ba8ad95),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f3dfe),
	.w1(32'h3b8be5b7),
	.w2(32'h3c4d6cc4),
	.w3(32'hbb9c61c3),
	.w4(32'hbb006467),
	.w5(32'h3c689829),
	.w6(32'hbc2ce71e),
	.w7(32'h39acffd9),
	.w8(32'h3c5952b2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc78cf),
	.w1(32'h3cebeba1),
	.w2(32'h3c558882),
	.w3(32'hbcaf71bd),
	.w4(32'hbbabacb2),
	.w5(32'h3c6cd0b0),
	.w6(32'hbae48be7),
	.w7(32'h3ab15c60),
	.w8(32'hbc0d8a30),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1467e),
	.w1(32'hbd101808),
	.w2(32'hbcf1455e),
	.w3(32'h3d1bc931),
	.w4(32'h3c972ec5),
	.w5(32'h3a7f6a47),
	.w6(32'h3b3f591a),
	.w7(32'h3b9e83ff),
	.w8(32'hbbe24d3c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe95ec0),
	.w1(32'hbca07570),
	.w2(32'h3b2df16c),
	.w3(32'h3ce2099a),
	.w4(32'h3c6e4a06),
	.w5(32'h3babe2c6),
	.w6(32'h3c35e690),
	.w7(32'h3c60489a),
	.w8(32'h3ac7053d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137dae),
	.w1(32'h3bc401dc),
	.w2(32'h3b58af3b),
	.w3(32'h3c1b7f8f),
	.w4(32'hbaaeded1),
	.w5(32'h3bb723c4),
	.w6(32'h3b908782),
	.w7(32'hbb63178d),
	.w8(32'h3b0b0dce),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8acd39),
	.w1(32'h3bb52a48),
	.w2(32'hbb016aee),
	.w3(32'h3affb8f0),
	.w4(32'hbb8c7906),
	.w5(32'hbc0f04f4),
	.w6(32'hbb86ce95),
	.w7(32'hbc0d0300),
	.w8(32'hbb989f00),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18a846),
	.w1(32'h3bbeb13e),
	.w2(32'h3c075403),
	.w3(32'hbc353a5e),
	.w4(32'hbb1c4b92),
	.w5(32'h3c04b15c),
	.w6(32'hbc0901f8),
	.w7(32'h3b487c2f),
	.w8(32'hbb367ec3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8891d8),
	.w1(32'h3af36cdd),
	.w2(32'hba8d3b9c),
	.w3(32'hbadf10d2),
	.w4(32'hbbbcf854),
	.w5(32'hbc006ff4),
	.w6(32'h3bf56f0a),
	.w7(32'hba504b8a),
	.w8(32'hbb384e3e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7020d),
	.w1(32'hbc069015),
	.w2(32'hbba19513),
	.w3(32'hbac0e88f),
	.w4(32'h397b6425),
	.w5(32'hbb8c2814),
	.w6(32'hbc541138),
	.w7(32'hbc0c14cd),
	.w8(32'hbb238b06),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1d675),
	.w1(32'h39eba8dc),
	.w2(32'hbbdbdb0d),
	.w3(32'hbc3218af),
	.w4(32'hbb7d7a2e),
	.w5(32'hbc225918),
	.w6(32'h3c0dd822),
	.w7(32'hbb561df3),
	.w8(32'h39f58cbb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43f299),
	.w1(32'h3bd10e68),
	.w2(32'hbad4e1b6),
	.w3(32'hbc16c67f),
	.w4(32'hbc00bb16),
	.w5(32'h3b8c8727),
	.w6(32'h3b41eb5e),
	.w7(32'hbbbd029e),
	.w8(32'h3ab2e765),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3191),
	.w1(32'hbc3b9ed8),
	.w2(32'hbb2e8ee3),
	.w3(32'hbacf8641),
	.w4(32'h3bf2e3cb),
	.w5(32'hbc236aa7),
	.w6(32'hbacc41f9),
	.w7(32'hbb19a45c),
	.w8(32'hba8ad613),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52f34c),
	.w1(32'h3c1e1341),
	.w2(32'h3bf2b3a4),
	.w3(32'h3b944daa),
	.w4(32'h3b183fbe),
	.w5(32'h3b968ef7),
	.w6(32'hbc5c3813),
	.w7(32'hbb355e13),
	.w8(32'h3af9dc69),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6e08d),
	.w1(32'hbb1d1508),
	.w2(32'hba2b2fd5),
	.w3(32'h3c0b220c),
	.w4(32'h3b289844),
	.w5(32'hba44d415),
	.w6(32'h3bac3988),
	.w7(32'h3a313cec),
	.w8(32'h3bc9ba61),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a1117),
	.w1(32'h3d049975),
	.w2(32'h3b98be78),
	.w3(32'hbd0e593c),
	.w4(32'hbc9681f7),
	.w5(32'hb8e981f2),
	.w6(32'h3bd8e3f0),
	.w7(32'hbb673476),
	.w8(32'hba277cc3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7883),
	.w1(32'hbbb2c7e2),
	.w2(32'hbb8c64f2),
	.w3(32'h3b857918),
	.w4(32'h3bc74d9c),
	.w5(32'h3ab8715c),
	.w6(32'hba7ad14d),
	.w7(32'hbbb05aa6),
	.w8(32'hbbe18729),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d87e8),
	.w1(32'hbc207202),
	.w2(32'hbc1ed9ac),
	.w3(32'h3c6f2371),
	.w4(32'hbc511799),
	.w5(32'hbc218194),
	.w6(32'hbc048d09),
	.w7(32'hbbe3c4ef),
	.w8(32'hbca1e229),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5f246),
	.w1(32'h3b914bb7),
	.w2(32'hbb16c398),
	.w3(32'hb9f5d87e),
	.w4(32'h3befb589),
	.w5(32'h3a11562f),
	.w6(32'h3a01dad9),
	.w7(32'hbbf2bf07),
	.w8(32'hbab51cf9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8fca),
	.w1(32'hba2ceb37),
	.w2(32'h3b0524af),
	.w3(32'hbb5d4f67),
	.w4(32'h3bba8927),
	.w5(32'hbb8c4eef),
	.w6(32'hbbeeacfc),
	.w7(32'hbc00e6fb),
	.w8(32'hbb4e110b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2d07b),
	.w1(32'h3b90f6f6),
	.w2(32'hbc33a66d),
	.w3(32'hbb3e0706),
	.w4(32'hbad79d6e),
	.w5(32'hbb42e84c),
	.w6(32'hb9025438),
	.w7(32'hbbcbc38b),
	.w8(32'h3b24f4e7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c8e2),
	.w1(32'h3c57c3b5),
	.w2(32'hba8e37e9),
	.w3(32'hbc42582c),
	.w4(32'hbc0f1283),
	.w5(32'hbc327a25),
	.w6(32'h3c9a7293),
	.w7(32'hb7520dd7),
	.w8(32'hbc81e314),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc60d0b),
	.w1(32'hbcb262eb),
	.w2(32'hbbd935d4),
	.w3(32'h3c9711d4),
	.w4(32'h3c51e448),
	.w5(32'h3abf834a),
	.w6(32'h39a1fbbc),
	.w7(32'h3b766799),
	.w8(32'hbbe8dfba),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbd24c),
	.w1(32'hbd0fd1a4),
	.w2(32'hbbf4de3b),
	.w3(32'h3cf787cc),
	.w4(32'h3cad7e5f),
	.w5(32'h3c2ef616),
	.w6(32'hbb644ea0),
	.w7(32'h3c91afd8),
	.w8(32'h3c62e16f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90dc117),
	.w1(32'hbc2b04f3),
	.w2(32'hbc38bf77),
	.w3(32'h3b27c3b9),
	.w4(32'hbc2865a3),
	.w5(32'hbbbfe215),
	.w6(32'hbc8f8f0b),
	.w7(32'hbbdad0c3),
	.w8(32'hbc107f46),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc667bb1),
	.w1(32'hbad5e63c),
	.w2(32'h3c7e5fe5),
	.w3(32'h3c203792),
	.w4(32'hb9da6580),
	.w5(32'h3c8705ca),
	.w6(32'hbc0ca434),
	.w7(32'h3bc33c1d),
	.w8(32'h3c723fc9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5d288),
	.w1(32'h3c605fb5),
	.w2(32'h3b41107a),
	.w3(32'hbbd76a4f),
	.w4(32'h3b1ec2b7),
	.w5(32'hbae9b70b),
	.w6(32'hbc076e88),
	.w7(32'hbba33d59),
	.w8(32'hbbc0c3d9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe3591),
	.w1(32'hbcad0c09),
	.w2(32'hbb8082e5),
	.w3(32'h3ca67d09),
	.w4(32'h3c351a45),
	.w5(32'h3b001bd6),
	.w6(32'h3b7cead7),
	.w7(32'h3af6203e),
	.w8(32'hbbfc0da2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66e095),
	.w1(32'hbc8f4155),
	.w2(32'hbbd87876),
	.w3(32'h3c2decb2),
	.w4(32'h3b28ada9),
	.w5(32'hbb37ee6d),
	.w6(32'h3b8e3002),
	.w7(32'h3c22c42a),
	.w8(32'h3bfd9077),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb85df9),
	.w1(32'h3c4bb8d0),
	.w2(32'h3b7bdec4),
	.w3(32'hbb922b28),
	.w4(32'h39984ece),
	.w5(32'hbb9dc466),
	.w6(32'hbc03f4e7),
	.w7(32'hbbc6b53a),
	.w8(32'hbc840404),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5aaa23),
	.w1(32'hbc92e5d5),
	.w2(32'hbbda686b),
	.w3(32'h3cb6f052),
	.w4(32'h3b787972),
	.w5(32'hbb1a6c7e),
	.w6(32'hba113969),
	.w7(32'hbaa67b5e),
	.w8(32'hbaaf43d2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9848a45),
	.w1(32'h3aac5e7b),
	.w2(32'hbba7944f),
	.w3(32'hbc486309),
	.w4(32'hb9993168),
	.w5(32'hbc409616),
	.w6(32'hbbda7b20),
	.w7(32'hbc3237e4),
	.w8(32'hbc2089b5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21d5e3),
	.w1(32'hbc137333),
	.w2(32'hbb77e76c),
	.w3(32'hbc74436e),
	.w4(32'hbb173698),
	.w5(32'hbcba00c6),
	.w6(32'hbb148243),
	.w7(32'hbba3f8be),
	.w8(32'hbc7e3d74),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b6de),
	.w1(32'h3d18e997),
	.w2(32'h3c43528d),
	.w3(32'hbc91ac97),
	.w4(32'hbbfe274c),
	.w5(32'h3ade14c1),
	.w6(32'h3b44731e),
	.w7(32'h3b72a8ec),
	.w8(32'h3c9e2c17),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b934b72),
	.w1(32'h3cc3790d),
	.w2(32'h38c32d28),
	.w3(32'hbce8110c),
	.w4(32'hbc5f72b6),
	.w5(32'h3b084d96),
	.w6(32'h3c04ae69),
	.w7(32'h3b81aed6),
	.w8(32'hbc0d8b65),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf391a0),
	.w1(32'hbd2b8860),
	.w2(32'hbc95710f),
	.w3(32'h3d16244f),
	.w4(32'h3c6e57cb),
	.w5(32'h3c499faa),
	.w6(32'h3ba5df0c),
	.w7(32'h3c21fb55),
	.w8(32'h3c5ce249),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96aa2b),
	.w1(32'h3cbac77c),
	.w2(32'h3b26abd3),
	.w3(32'hbc5bee38),
	.w4(32'h3b079f8a),
	.w5(32'h3b439498),
	.w6(32'hbb81606a),
	.w7(32'h3b0a2f19),
	.w8(32'hb8d114dc),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeb823),
	.w1(32'h3c0c900a),
	.w2(32'hbade462a),
	.w3(32'hbb4a4cdb),
	.w4(32'hbad2aafa),
	.w5(32'hbb9deb76),
	.w6(32'hbb418918),
	.w7(32'hbbb570e7),
	.w8(32'hbb2cd49b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a128e06),
	.w1(32'h3b7db04c),
	.w2(32'h3bc37037),
	.w3(32'h3b2ca862),
	.w4(32'hba63c752),
	.w5(32'hbc1b2c3d),
	.w6(32'hb914a0de),
	.w7(32'h3b96f7fb),
	.w8(32'hbc560a8c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6b0d3),
	.w1(32'hbb93f62e),
	.w2(32'hba999a97),
	.w3(32'h3c8f4ace),
	.w4(32'hbb785158),
	.w5(32'hbbbefdb2),
	.w6(32'hbbaa4544),
	.w7(32'h3b02a9c3),
	.w8(32'h3b2fa4a7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f903f),
	.w1(32'hbadbf807),
	.w2(32'hbb6846ad),
	.w3(32'hbc17c431),
	.w4(32'hba838fd7),
	.w5(32'h3b801e22),
	.w6(32'h3b94a43a),
	.w7(32'h3b67adaa),
	.w8(32'hbb957e14),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1019),
	.w1(32'hbb939e6b),
	.w2(32'h3ba966fc),
	.w3(32'hb8a96d30),
	.w4(32'h3b8100eb),
	.w5(32'h3b6d4a4d),
	.w6(32'hbc239b9e),
	.w7(32'hbac0b504),
	.w8(32'h3b904407),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91fb55),
	.w1(32'hb9184d85),
	.w2(32'h3bbed430),
	.w3(32'h3c24b124),
	.w4(32'hbad90621),
	.w5(32'hbb1e4eea),
	.w6(32'hbb32ebdb),
	.w7(32'hbb482e48),
	.w8(32'hbc11ff11),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a3f5),
	.w1(32'hba72587e),
	.w2(32'hbb7be59e),
	.w3(32'hbb6633fa),
	.w4(32'hb91e3ecb),
	.w5(32'h3b192513),
	.w6(32'h3c3e157e),
	.w7(32'hbba18e6a),
	.w8(32'hbb5080a2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2377fb),
	.w1(32'hbc892ff0),
	.w2(32'hbc1a7610),
	.w3(32'h3c86162b),
	.w4(32'h3c413ab2),
	.w5(32'h3bf23108),
	.w6(32'hba83931b),
	.w7(32'h3b09787b),
	.w8(32'hbb679537),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b1d18),
	.w1(32'hbce9df86),
	.w2(32'hbcd05201),
	.w3(32'h3c77661a),
	.w4(32'hbba739c7),
	.w5(32'hbc1aa76f),
	.w6(32'hbc203476),
	.w7(32'hbc1d4a74),
	.w8(32'hbc979d37),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bf376),
	.w1(32'hbcb2ce9b),
	.w2(32'hbb64f562),
	.w3(32'h3c89cddf),
	.w4(32'hbbb3e236),
	.w5(32'hb9709f13),
	.w6(32'hb9e17b1b),
	.w7(32'h3a32230b),
	.w8(32'hbb0080c3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dae0f),
	.w1(32'h3c2a32bb),
	.w2(32'hba5daf8e),
	.w3(32'h3b7a0905),
	.w4(32'h3bce3c2b),
	.w5(32'hbb831784),
	.w6(32'hbbff76a1),
	.w7(32'hbb09ff0b),
	.w8(32'hbbf5d56f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06b1b2),
	.w1(32'h3c079862),
	.w2(32'h3c819102),
	.w3(32'h3b204de2),
	.w4(32'h3c094d9a),
	.w5(32'h3b0ebc89),
	.w6(32'hbba45cff),
	.w7(32'hbbb30658),
	.w8(32'h3b972c5d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc030636),
	.w1(32'hbbcac1d2),
	.w2(32'h3b258e5b),
	.w3(32'hbc1a4411),
	.w4(32'h3932fab7),
	.w5(32'hbbda4c29),
	.w6(32'hbbc5e30b),
	.w7(32'h3b9ca3b8),
	.w8(32'hbc1af737),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38cb97),
	.w1(32'h3bf04805),
	.w2(32'h39fb45a2),
	.w3(32'h3c07f3f6),
	.w4(32'hbb85942c),
	.w5(32'hbbbbce7a),
	.w6(32'hbbc085d8),
	.w7(32'hbba3d28b),
	.w8(32'hbc08801c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee3f7),
	.w1(32'h3c9a0b74),
	.w2(32'h3c80a601),
	.w3(32'hbc83aeb6),
	.w4(32'hbb2caaa2),
	.w5(32'hbaf63452),
	.w6(32'hbc076784),
	.w7(32'hbc20f4e9),
	.w8(32'h3c7a3888),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb22a8),
	.w1(32'h3d6311d1),
	.w2(32'h3c7c1738),
	.w3(32'hbd37fd46),
	.w4(32'hbcb709b3),
	.w5(32'h3af5b429),
	.w6(32'h3c4e16ad),
	.w7(32'hbb33b7d4),
	.w8(32'h3bd8f76f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bfef3),
	.w1(32'h3b18cc6f),
	.w2(32'h3be760fd),
	.w3(32'h3bb3776d),
	.w4(32'hbb123d7a),
	.w5(32'h3b43457c),
	.w6(32'hbc4a5269),
	.w7(32'h39e0ed0f),
	.w8(32'hbb2425a1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb1aba),
	.w1(32'hbbafe6ad),
	.w2(32'hb9c7fb20),
	.w3(32'hbba0de71),
	.w4(32'hbb89277b),
	.w5(32'h3774d257),
	.w6(32'hbbca6a26),
	.w7(32'hbbef12ee),
	.w8(32'hbae2464b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd274ba),
	.w1(32'hbba89844),
	.w2(32'hbc30fbb9),
	.w3(32'hbbaa24d9),
	.w4(32'hbbc31173),
	.w5(32'hbc933944),
	.w6(32'hbbdea286),
	.w7(32'hbbd46f27),
	.w8(32'hbc68936e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd34e50),
	.w1(32'hbc0ded4d),
	.w2(32'hbaafd7b2),
	.w3(32'hbb3b2b4f),
	.w4(32'h3a63fb1b),
	.w5(32'h3c41f3f6),
	.w6(32'h3a539a0d),
	.w7(32'hb9277e90),
	.w8(32'h3bc57342),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab10e3b),
	.w1(32'h3c135202),
	.w2(32'h3c06b538),
	.w3(32'h3b232158),
	.w4(32'h3c4a5f97),
	.w5(32'h3ca15355),
	.w6(32'hbbf3e100),
	.w7(32'h3bacd560),
	.w8(32'h3c617dd3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a36ed),
	.w1(32'hbbbe0544),
	.w2(32'hbbe1050a),
	.w3(32'hbb07f7ba),
	.w4(32'hba30398f),
	.w5(32'hbc04c8f1),
	.w6(32'hbb698c08),
	.w7(32'h3972b83c),
	.w8(32'hbc2b0c4d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349275),
	.w1(32'hb99eda51),
	.w2(32'h3992fcb3),
	.w3(32'hba07b586),
	.w4(32'h3adbb71c),
	.w5(32'h3b538d63),
	.w6(32'hbb01bb1f),
	.w7(32'h3a9297b5),
	.w8(32'h3b52adbb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf09ca3),
	.w1(32'hbc22155e),
	.w2(32'hbca0df84),
	.w3(32'hbc2cd04f),
	.w4(32'hbc2b117a),
	.w5(32'hbca1dd10),
	.w6(32'hbbe3729d),
	.w7(32'hbc0c82fe),
	.w8(32'hbc574fd2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffe3ad),
	.w1(32'hbb0bdc94),
	.w2(32'h3b82fe7c),
	.w3(32'h3a2657a3),
	.w4(32'hbad7bd4c),
	.w5(32'h3bc417e2),
	.w6(32'hba631f01),
	.w7(32'h394c95b3),
	.w8(32'h3c0786d9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404917),
	.w1(32'h39388c5b),
	.w2(32'h3a7e35e3),
	.w3(32'h3ade8406),
	.w4(32'hb9d80040),
	.w5(32'hba640bda),
	.w6(32'h3a847cf0),
	.w7(32'hbafe9719),
	.w8(32'h39c3ae0e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a7fdf),
	.w1(32'h3b4e6b12),
	.w2(32'h3b31d56c),
	.w3(32'h3b181370),
	.w4(32'h3b19d818),
	.w5(32'hbadafc90),
	.w6(32'h3b0cc6ff),
	.w7(32'h3b459fc7),
	.w8(32'hbac8db72),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06d0a8),
	.w1(32'h3ba6c29f),
	.w2(32'h3b807bfb),
	.w3(32'h3b304e62),
	.w4(32'h3c0ff8a6),
	.w5(32'h3be5611a),
	.w6(32'hbb192bf3),
	.w7(32'h3b8f69b4),
	.w8(32'h3b274ee3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8d388),
	.w1(32'h3b7cf7e8),
	.w2(32'h3bdff8b4),
	.w3(32'hb8dfaea4),
	.w4(32'h3bfeffcc),
	.w5(32'h3c0e30bc),
	.w6(32'hbbcca9e2),
	.w7(32'h3bae2efa),
	.w8(32'h3bbdb234),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc35ae),
	.w1(32'hbc0b2424),
	.w2(32'hbbf83234),
	.w3(32'hbbff0121),
	.w4(32'hbb99790a),
	.w5(32'h3b17c26f),
	.w6(32'hbbd4594e),
	.w7(32'hbb8054fb),
	.w8(32'h3ae03e78),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2f834),
	.w1(32'h3a85871c),
	.w2(32'h3b95e0b3),
	.w3(32'h391a6f23),
	.w4(32'h3a4f09f6),
	.w5(32'h3bbcc167),
	.w6(32'hbaf6b874),
	.w7(32'h3b2e8ec6),
	.w8(32'h3bb44389),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40fe1b),
	.w1(32'h3a469eea),
	.w2(32'h3b085f59),
	.w3(32'h3a7fcaa2),
	.w4(32'h3b3ec7aa),
	.w5(32'h3a3c5c54),
	.w6(32'h3a3b6473),
	.w7(32'h3abf793d),
	.w8(32'hb9b23655),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a8e23),
	.w1(32'h3acfb549),
	.w2(32'hba735a0b),
	.w3(32'hba971c7a),
	.w4(32'h3b43f7b8),
	.w5(32'h3b05808d),
	.w6(32'hbab73d85),
	.w7(32'h3a741f1a),
	.w8(32'hbabd244b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b0457),
	.w1(32'h3b55ef13),
	.w2(32'h3bcae3d8),
	.w3(32'h3b02f2d8),
	.w4(32'h3b85d5bf),
	.w5(32'h3c0eb8ef),
	.w6(32'hb84479c6),
	.w7(32'h3ba3306a),
	.w8(32'h3ba1c548),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb512e63d),
	.w1(32'h39f89cfc),
	.w2(32'h3a4af754),
	.w3(32'h3aff3989),
	.w4(32'h39adb30c),
	.w5(32'h3b8df261),
	.w6(32'hba0103e1),
	.w7(32'hb53a21aa),
	.w8(32'h3b8185fe),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba746d0),
	.w1(32'h3b8e8476),
	.w2(32'h3b349bf2),
	.w3(32'h3b2c552f),
	.w4(32'h3ac6691a),
	.w5(32'hbb1ed596),
	.w6(32'h3b582a69),
	.w7(32'h3ae3cdd2),
	.w8(32'hbaf2c354),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52520b),
	.w1(32'hbae822aa),
	.w2(32'hbb03b733),
	.w3(32'hb9009cf2),
	.w4(32'hb9e560ef),
	.w5(32'hbb2d90f0),
	.w6(32'hbb0fa83a),
	.w7(32'hb905309f),
	.w8(32'hbb574780),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb258d21),
	.w1(32'hbb27ade5),
	.w2(32'hbac77a18),
	.w3(32'hbb0618ec),
	.w4(32'hba64c19d),
	.w5(32'hbb840120),
	.w6(32'hbb62721e),
	.w7(32'hbb35f010),
	.w8(32'hbb91187d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63d083),
	.w1(32'h3b1c558c),
	.w2(32'h3b8dab99),
	.w3(32'hbb4a79ca),
	.w4(32'h3b67014c),
	.w5(32'h3ca12622),
	.w6(32'hbbbcf3b6),
	.w7(32'h3a63330b),
	.w8(32'h3c67a117),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ad68),
	.w1(32'h3af4c632),
	.w2(32'h3b3efe41),
	.w3(32'h3b9333de),
	.w4(32'h3b02cdaf),
	.w5(32'h3b03a91a),
	.w6(32'h3b644f9c),
	.w7(32'h3b21249c),
	.w8(32'h3b78edb4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cb610),
	.w1(32'hba7d810f),
	.w2(32'hbbcfd4df),
	.w3(32'hba28216c),
	.w4(32'hbb6bc004),
	.w5(32'h3af795bc),
	.w6(32'h3aefe7ec),
	.w7(32'hbb8f904c),
	.w8(32'h39f1460d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b75ce),
	.w1(32'hbac8066b),
	.w2(32'hba0fe1bf),
	.w3(32'h3be8de50),
	.w4(32'h3c0853f6),
	.w5(32'h3bad32c2),
	.w6(32'hbb382983),
	.w7(32'h3b593de5),
	.w8(32'h3bc772c1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a760c),
	.w1(32'h383f57b7),
	.w2(32'hbb1f092e),
	.w3(32'hbb6c1aaf),
	.w4(32'hbb90108e),
	.w5(32'h3a9a4ca4),
	.w6(32'hbab7b43f),
	.w7(32'hbb716039),
	.w8(32'h3a07a8dd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f268f),
	.w1(32'hbb70b6a7),
	.w2(32'hbb2949af),
	.w3(32'h3b94787a),
	.w4(32'h3b2bec1a),
	.w5(32'h3b50d140),
	.w6(32'h39dfc2a7),
	.w7(32'h3b097eba),
	.w8(32'h3aafc070),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5185f),
	.w1(32'h3b5f11c2),
	.w2(32'h3b0a7c13),
	.w3(32'h3bb640ef),
	.w4(32'h3be9d17d),
	.w5(32'hb92fe3ce),
	.w6(32'h3aa6b07d),
	.w7(32'h3b3d25bf),
	.w8(32'h3aba7895),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4c29),
	.w1(32'h3ae52d8c),
	.w2(32'h3a16ade8),
	.w3(32'h3b29f16d),
	.w4(32'h3ad8d6a3),
	.w5(32'h3b2358f3),
	.w6(32'h3abc76ef),
	.w7(32'h3a92e7d7),
	.w8(32'h3a3f7af4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a623e53),
	.w1(32'h3b76635c),
	.w2(32'h3b5f5ebd),
	.w3(32'h3a70c629),
	.w4(32'h3b3639a1),
	.w5(32'h3b3c3a2f),
	.w6(32'hba56627f),
	.w7(32'h3ac69f29),
	.w8(32'h3a8c1b23),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987c102),
	.w1(32'h3b89e43d),
	.w2(32'h3bccb8f7),
	.w3(32'h3b2a67a7),
	.w4(32'h3bfc7314),
	.w5(32'h3ba64a1e),
	.w6(32'hba0c2916),
	.w7(32'h3bf6fffd),
	.w8(32'h3ae69744),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53d727),
	.w1(32'hbb3f4e90),
	.w2(32'hbb8f820f),
	.w3(32'hbad1367b),
	.w4(32'hbad3a918),
	.w5(32'hba6d91ea),
	.w6(32'hbb410a40),
	.w7(32'hbadf1a95),
	.w8(32'h3a12f3e1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b66375),
	.w1(32'hbaf3d2fc),
	.w2(32'h39ede6dc),
	.w3(32'hbaad1ad4),
	.w4(32'hb9a98366),
	.w5(32'hbaf16762),
	.w6(32'hb908e8c6),
	.w7(32'hbb2040f8),
	.w8(32'hba5664c7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c1b5c),
	.w1(32'hb95b57a7),
	.w2(32'hba23ae0f),
	.w3(32'hba8ba2c0),
	.w4(32'hba9316fc),
	.w5(32'h3b2e0740),
	.w6(32'hbb3e873c),
	.w7(32'hbad180cd),
	.w8(32'h3b8827d2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba66ed0),
	.w1(32'h3c091411),
	.w2(32'h3bfe51b8),
	.w3(32'h3b86811f),
	.w4(32'h3bf28bfe),
	.w5(32'hba8a596d),
	.w6(32'h3b6ffa81),
	.w7(32'h3c13b4c9),
	.w8(32'hbb21c022),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6e5d7),
	.w1(32'h3a3f3da4),
	.w2(32'hba9d2760),
	.w3(32'hbb157e48),
	.w4(32'hba969a9d),
	.w5(32'hbab04ad5),
	.w6(32'hbb351ad1),
	.w7(32'hbb220ca4),
	.w8(32'hbb4b1a06),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905176),
	.w1(32'hbb9974e7),
	.w2(32'hbbfeb342),
	.w3(32'hbb67f34d),
	.w4(32'hbb888515),
	.w5(32'hba9147f4),
	.w6(32'hbc03a33f),
	.w7(32'hbbeac7df),
	.w8(32'hbb903845),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f8a3),
	.w1(32'h3ba1c710),
	.w2(32'h3bdb928a),
	.w3(32'h3b77fcd1),
	.w4(32'h3c066560),
	.w5(32'h3c1a932b),
	.w6(32'h3a13e63d),
	.w7(32'h3bb69f6e),
	.w8(32'h3bd80f28),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a085935),
	.w1(32'h3b248cd4),
	.w2(32'h3b23cfbb),
	.w3(32'hbac712ba),
	.w4(32'h3a797e1e),
	.w5(32'hbb052cf3),
	.w6(32'hba76f2f2),
	.w7(32'h3a199f74),
	.w8(32'hbb9d6e2a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3604a),
	.w1(32'hbbd6892d),
	.w2(32'hbc07bd86),
	.w3(32'hbbb5f754),
	.w4(32'hbba0e252),
	.w5(32'hbbc8b5bb),
	.w6(32'hbc083396),
	.w7(32'hbb9ce6f7),
	.w8(32'hbbafd769),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380941de),
	.w1(32'hb9be7c5d),
	.w2(32'hbb222f75),
	.w3(32'hbaa07897),
	.w4(32'hb886a662),
	.w5(32'hbade0b0a),
	.w6(32'hbb2976d4),
	.w7(32'hba672319),
	.w8(32'hbaea75f7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f7ccc),
	.w1(32'hbb03d011),
	.w2(32'hbb0d6f76),
	.w3(32'hbb5844b0),
	.w4(32'hba3d1ac8),
	.w5(32'h3b12bc83),
	.w6(32'hbb5f8e16),
	.w7(32'hbafb8b01),
	.w8(32'h3a365c0b),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb445922),
	.w1(32'hb992b485),
	.w2(32'h3b4da7e6),
	.w3(32'h3a8a6433),
	.w4(32'h3ba38f18),
	.w5(32'h3ba52b74),
	.w6(32'hbade7e46),
	.w7(32'h3b641537),
	.w8(32'h3b6d7fa7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b2327),
	.w1(32'h3bd48736),
	.w2(32'h3c6ba9d7),
	.w3(32'h3be90848),
	.w4(32'h3c6eb739),
	.w5(32'h3b9dba2b),
	.w6(32'h3ba8f7bf),
	.w7(32'h3c8c4039),
	.w8(32'h3b8a8c17),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaab53),
	.w1(32'hbbfb746f),
	.w2(32'hbc156302),
	.w3(32'hbbfde7d2),
	.w4(32'hbbf90649),
	.w5(32'hbbfe3f68),
	.w6(32'hbc0d3895),
	.w7(32'hbc0c86cf),
	.w8(32'hbc284940),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb653871),
	.w1(32'hbaea7f36),
	.w2(32'h3a21c5f4),
	.w3(32'h3946d222),
	.w4(32'h3b74c22c),
	.w5(32'h3a90d50c),
	.w6(32'hbb479346),
	.w7(32'h3b43addf),
	.w8(32'h3aef6c7c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa7fd),
	.w1(32'hb9a53ed1),
	.w2(32'hb8689c63),
	.w3(32'h3ac3389a),
	.w4(32'h39eb6c35),
	.w5(32'hba9ceb6f),
	.w6(32'h3a92ed31),
	.w7(32'h3ac4892d),
	.w8(32'hb9926017),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa3b81),
	.w1(32'h38ffbb92),
	.w2(32'h3af9553a),
	.w3(32'hbaa9c64c),
	.w4(32'hba08a0f7),
	.w5(32'h3b042e4d),
	.w6(32'h398b9c00),
	.w7(32'hb92b29fc),
	.w8(32'h3b0ce2c4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7154e6),
	.w1(32'hbba19e12),
	.w2(32'hbb463edf),
	.w3(32'hbbb2a982),
	.w4(32'hbb045723),
	.w5(32'h3a55efb0),
	.w6(32'hbc0f5125),
	.w7(32'hbb1bf19d),
	.w8(32'hbb37e0ad),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f507),
	.w1(32'h3c12f8aa),
	.w2(32'h3c64e8bd),
	.w3(32'h3bf17dc5),
	.w4(32'h3c4657e9),
	.w5(32'h3c4fa394),
	.w6(32'h3ae9a550),
	.w7(32'h3bf29512),
	.w8(32'h3c0a1968),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6712d98),
	.w1(32'h39f65e0a),
	.w2(32'h3b587c08),
	.w3(32'h3b047a28),
	.w4(32'h3bd1dea3),
	.w5(32'h3ad065b7),
	.w6(32'hb959a1b8),
	.w7(32'h3bd5bb26),
	.w8(32'h3af2980d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a663f87),
	.w1(32'h3b9972b6),
	.w2(32'h3b897341),
	.w3(32'h3aee1a9a),
	.w4(32'h3b63d7f0),
	.w5(32'h3c1b3d7d),
	.w6(32'hba7e020b),
	.w7(32'h3b1c515d),
	.w8(32'h3b987141),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d1a00),
	.w1(32'h3ba1cabb),
	.w2(32'h3ba12243),
	.w3(32'h3b2a1e77),
	.w4(32'h3bdb9989),
	.w5(32'h3b35115e),
	.w6(32'hba5b71d0),
	.w7(32'h3b4dc087),
	.w8(32'hbb1a4cc4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9689a),
	.w1(32'h39c89c62),
	.w2(32'h3b89265d),
	.w3(32'h3a577966),
	.w4(32'h3bcee75d),
	.w5(32'hbb67c915),
	.w6(32'hbb618932),
	.w7(32'h3bfddb1d),
	.w8(32'hbba56cbb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077692),
	.w1(32'h3b4e82b1),
	.w2(32'h3c004c57),
	.w3(32'hba9ce146),
	.w4(32'h3b32946c),
	.w5(32'h3c0cc62b),
	.w6(32'hbba42a98),
	.w7(32'hba734993),
	.w8(32'h3be3b426),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51d425),
	.w1(32'hb7eefc31),
	.w2(32'hba64b6ba),
	.w3(32'h3877c7fc),
	.w4(32'hbb01377d),
	.w5(32'hbb333bab),
	.w6(32'h3a29a993),
	.w7(32'hbaad3cdb),
	.w8(32'hba4f9ecd),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7b1d),
	.w1(32'h3a9e8e4c),
	.w2(32'hbafb2bc1),
	.w3(32'h3aadc8c7),
	.w4(32'hb98febab),
	.w5(32'h3ade519d),
	.w6(32'h3b019e0d),
	.w7(32'hb967fd38),
	.w8(32'h3b5e92f1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba873d8c),
	.w1(32'h3b6347af),
	.w2(32'h3ba857e5),
	.w3(32'h3a06baa2),
	.w4(32'h3be5ba20),
	.w5(32'h3a8e34b6),
	.w6(32'hba71b3e7),
	.w7(32'h3bdda609),
	.w8(32'hb9b8459d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ba4ee),
	.w1(32'hbbac5f03),
	.w2(32'hbb868e23),
	.w3(32'hbb8d67aa),
	.w4(32'hbb813a66),
	.w5(32'h3b43d445),
	.w6(32'hbb8f5e9f),
	.w7(32'hbbbb53f3),
	.w8(32'h3bd8d648),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d653),
	.w1(32'h3bb40d1c),
	.w2(32'h3b0d323c),
	.w3(32'h3bbfe1ae),
	.w4(32'h3a692c15),
	.w5(32'h3b4b09a8),
	.w6(32'h3bf41862),
	.w7(32'h3a1f9cf8),
	.w8(32'h3b9bbf6e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dbd61),
	.w1(32'h3c0b2e32),
	.w2(32'h3b8582f0),
	.w3(32'h3b277ab9),
	.w4(32'h3b8ddfc7),
	.w5(32'h3b6df005),
	.w6(32'h3bb51bdb),
	.w7(32'h3b9e6ef4),
	.w8(32'h3b2dd75a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933046),
	.w1(32'h3b8bd627),
	.w2(32'h3bc61513),
	.w3(32'h3bce445f),
	.w4(32'h3b89ef98),
	.w5(32'hba9caa38),
	.w6(32'h3c01b95e),
	.w7(32'h3bd2d0f2),
	.w8(32'hbaf649a2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e96ea),
	.w1(32'hbb005607),
	.w2(32'hbb16cf7b),
	.w3(32'hbb8cd438),
	.w4(32'hbb29fd59),
	.w5(32'hbb1df095),
	.w6(32'hbba8ffe2),
	.w7(32'hbb5e9737),
	.w8(32'hbb790c85),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c1342),
	.w1(32'hbb05823b),
	.w2(32'hbaf7fb7e),
	.w3(32'hbb0bbf1a),
	.w4(32'hba69d68e),
	.w5(32'h3afcf817),
	.w6(32'hbb12ebed),
	.w7(32'hba1a3bfd),
	.w8(32'h3a1cd270),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98f41e),
	.w1(32'h3b67cc34),
	.w2(32'h3bc83ab9),
	.w3(32'h3b1185a1),
	.w4(32'h3bb8016c),
	.w5(32'h3b1dc7f5),
	.w6(32'hbb0db519),
	.w7(32'h3b9a0f21),
	.w8(32'h3b06eb7f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5ad31),
	.w1(32'hba0fc1ab),
	.w2(32'hbaa0a767),
	.w3(32'hbb17f456),
	.w4(32'h39b16ddc),
	.w5(32'h396bd18f),
	.w6(32'hbb52178b),
	.w7(32'hb964a796),
	.w8(32'h3a2f39d7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f4afc),
	.w1(32'h3b4b3f64),
	.w2(32'h3a2ee622),
	.w3(32'h3b4b074a),
	.w4(32'h3b84539c),
	.w5(32'h3b4c4cd4),
	.w6(32'h3be840b0),
	.w7(32'h3b8c162c),
	.w8(32'h3ba5978c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b250444),
	.w1(32'h3ab76149),
	.w2(32'hb9dc7c27),
	.w3(32'h3a2d799d),
	.w4(32'hb9a23be1),
	.w5(32'hba2eaec8),
	.w6(32'h3a390658),
	.w7(32'h39e013c4),
	.w8(32'h3aacd4a9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b127a9f),
	.w1(32'h3b950bd1),
	.w2(32'h3b30c467),
	.w3(32'hbb3b33be),
	.w4(32'hbafd2659),
	.w5(32'h39f45b16),
	.w6(32'hb866750a),
	.w7(32'h3a8387aa),
	.w8(32'h3a48d4af),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ccc39),
	.w1(32'hbad8e66d),
	.w2(32'hbb0b436e),
	.w3(32'hb892b567),
	.w4(32'hba0428d9),
	.w5(32'h3a2f6116),
	.w6(32'hbad73a40),
	.w7(32'hbb396b7f),
	.w8(32'hbac33960),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb9fbb),
	.w1(32'hbb884762),
	.w2(32'hbbcd6d6b),
	.w3(32'hbbeff359),
	.w4(32'hba0642ba),
	.w5(32'h3b1a0b4e),
	.w6(32'hbc224e27),
	.w7(32'hbba17ee6),
	.w8(32'hbb7ba4dc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e107e),
	.w1(32'h3a74888c),
	.w2(32'hba0181de),
	.w3(32'h3b3f0949),
	.w4(32'h3a6f14b3),
	.w5(32'h3b67e836),
	.w6(32'h3b939b04),
	.w7(32'h3a898229),
	.w8(32'h3bb6edec),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e8e9),
	.w1(32'h3b97ca22),
	.w2(32'h3bb2278c),
	.w3(32'h3b5a3e0d),
	.w4(32'h3bf8538f),
	.w5(32'h3bf0c185),
	.w6(32'h3a99ec8b),
	.w7(32'h3bf0d1b3),
	.w8(32'h3ba1a933),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf94eec),
	.w1(32'hb9f3fa70),
	.w2(32'hbb0b907f),
	.w3(32'hbaaac394),
	.w4(32'hbb41eae7),
	.w5(32'hbb83a318),
	.w6(32'hbad43043),
	.w7(32'hba9718cd),
	.w8(32'hbb8a21b0),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf0ae3),
	.w1(32'hbb720b55),
	.w2(32'hbb4845aa),
	.w3(32'hbc055ed4),
	.w4(32'hbb2589b2),
	.w5(32'h3b81e70b),
	.w6(32'hbbdc193c),
	.w7(32'hbbb1419e),
	.w8(32'h3b03ad34),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06063a),
	.w1(32'h3b28b905),
	.w2(32'h3b61617f),
	.w3(32'h3a7930b5),
	.w4(32'h3b364067),
	.w5(32'hbb8f8cbb),
	.w6(32'h3a3ee912),
	.w7(32'h3a9a72ef),
	.w8(32'hbbb21383),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7f90e),
	.w1(32'hbaeab5fe),
	.w2(32'hbb9d2d02),
	.w3(32'hbb849623),
	.w4(32'hba458e66),
	.w5(32'h3bf2ddb6),
	.w6(32'hbc0288b8),
	.w7(32'hbb8462fb),
	.w8(32'h3add16b5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e61e),
	.w1(32'h3a76b420),
	.w2(32'hba0b4001),
	.w3(32'h3aa8940c),
	.w4(32'h3a96f44c),
	.w5(32'hbb080968),
	.w6(32'h3a9e612c),
	.w7(32'h3a9b8404),
	.w8(32'hbaedade7),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce0d43),
	.w1(32'hbb84e843),
	.w2(32'hbb116bb0),
	.w3(32'hbb7dec78),
	.w4(32'hba16c2c3),
	.w5(32'h3b83bca4),
	.w6(32'hbba5c686),
	.w7(32'hbaf56aee),
	.w8(32'h3ae36123),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d4560),
	.w1(32'h3b251981),
	.w2(32'hb99002af),
	.w3(32'h3b0b5380),
	.w4(32'hba277db7),
	.w5(32'h3ac558c1),
	.w6(32'h3b6fad59),
	.w7(32'hb9ef542b),
	.w8(32'h38119437),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbf44c),
	.w1(32'h3a4af33b),
	.w2(32'h3b479d06),
	.w3(32'h3ae7ec7b),
	.w4(32'h3b19cf79),
	.w5(32'hb97556f3),
	.w6(32'hb83f5fe8),
	.w7(32'h3b4ce67b),
	.w8(32'h3a5da77f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeec27),
	.w1(32'hba2c5d42),
	.w2(32'hba5cd91c),
	.w3(32'hb8093354),
	.w4(32'h39f7f3ae),
	.w5(32'h396c956b),
	.w6(32'hbb033272),
	.w7(32'h3a406455),
	.w8(32'hb879bcba),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40b217),
	.w1(32'h3b0bc0d9),
	.w2(32'h3b311703),
	.w3(32'hba1d29b4),
	.w4(32'h3a9855ae),
	.w5(32'h3bcb3b0a),
	.w6(32'hbb140f1f),
	.w7(32'h390be728),
	.w8(32'h3b92bab8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15335a),
	.w1(32'h3b02194a),
	.w2(32'h39cd0db6),
	.w3(32'h3af6ba34),
	.w4(32'h3adbdc58),
	.w5(32'hbabf5386),
	.w6(32'h3b8bc535),
	.w7(32'hb9f9fc0f),
	.w8(32'hbaa62940),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa60612),
	.w1(32'hbb08b063),
	.w2(32'hbb35d352),
	.w3(32'hba9e4e2e),
	.w4(32'hbad087be),
	.w5(32'h3b038f64),
	.w6(32'hbb316f1f),
	.w7(32'hbb16072a),
	.w8(32'h3a78857f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea128e),
	.w1(32'h3ab6d5e2),
	.w2(32'h3bbcf118),
	.w3(32'h3b98eb8c),
	.w4(32'h3bc2e49f),
	.w5(32'h3b0f7af0),
	.w6(32'h3ad2fb0d),
	.w7(32'h3bcd7049),
	.w8(32'h3a8440bd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070e2b),
	.w1(32'h383be283),
	.w2(32'h3bc1003a),
	.w3(32'h3b1c3507),
	.w4(32'h3b42b269),
	.w5(32'h3bf2434e),
	.w6(32'h398910d6),
	.w7(32'h3b68c8cf),
	.w8(32'h3bb29737),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3df9de),
	.w1(32'h3b04a494),
	.w2(32'h392b17f4),
	.w3(32'h3b192cd5),
	.w4(32'h3a1715cf),
	.w5(32'h3a67218d),
	.w6(32'h3ad6e670),
	.w7(32'h396e19fe),
	.w8(32'h3b15bd23),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d132f),
	.w1(32'hb90e40f5),
	.w2(32'hbb225dc6),
	.w3(32'h3b338756),
	.w4(32'hba96c3a6),
	.w5(32'hbb29c1a8),
	.w6(32'h3b89726b),
	.w7(32'hbab03fbf),
	.w8(32'hbb62aaf4),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8d377),
	.w1(32'h3b43ee9b),
	.w2(32'h3b7eaeb1),
	.w3(32'h3ac569b7),
	.w4(32'h3c388ca2),
	.w5(32'h3c2a7ac4),
	.w6(32'hbb722a18),
	.w7(32'h3bf35730),
	.w8(32'h3c3eddb9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038c5a),
	.w1(32'h3ba23b45),
	.w2(32'h3b831b5e),
	.w3(32'hbad1fb3d),
	.w4(32'hba79315a),
	.w5(32'h3b289a65),
	.w6(32'h3b416363),
	.w7(32'h3b2b346f),
	.w8(32'h3abe18b7),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0797),
	.w1(32'h39628cb3),
	.w2(32'hb9c442de),
	.w3(32'h3abe8d9c),
	.w4(32'h3a9d7b9a),
	.w5(32'h3b61a5f2),
	.w6(32'h3a33f2bc),
	.w7(32'h3a3245ce),
	.w8(32'h3b805d36),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2e9f),
	.w1(32'h3bcf3bcf),
	.w2(32'h3baf49a8),
	.w3(32'h3b0c126a),
	.w4(32'h3a70fc22),
	.w5(32'h39e35873),
	.w6(32'h3b5f638b),
	.w7(32'h3b50f10b),
	.w8(32'h3a6cd90f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edbf92),
	.w1(32'h3abbc4ed),
	.w2(32'h3b15caa0),
	.w3(32'h3a93bc4e),
	.w4(32'h3b502e30),
	.w5(32'h3ac5e665),
	.w6(32'h3b05e59b),
	.w7(32'h3b7da8d4),
	.w8(32'h3b1a71f9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2946ed),
	.w1(32'h3b182068),
	.w2(32'h3abe0311),
	.w3(32'h3b38159d),
	.w4(32'h3a1f8e9f),
	.w5(32'h39fd10ed),
	.w6(32'h3b464222),
	.w7(32'h3b0c1f9d),
	.w8(32'hb9dbf7d0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d462e9),
	.w1(32'hbaae2469),
	.w2(32'hbb13f5e8),
	.w3(32'hb9c0bf1d),
	.w4(32'hbb1be62e),
	.w5(32'h3afc2abf),
	.w6(32'hbb6d0d0d),
	.w7(32'hbb66cf18),
	.w8(32'h3afd4ff1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb401b),
	.w1(32'hbb43db22),
	.w2(32'hbc005d84),
	.w3(32'hbb04cf3a),
	.w4(32'hbb40d2d6),
	.w5(32'hbbdc4891),
	.w6(32'hbac787bf),
	.w7(32'hbb7ed23a),
	.w8(32'hbbe2f5eb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb600558),
	.w1(32'h3a94e40e),
	.w2(32'h3b5bfc13),
	.w3(32'hbb6fb5a8),
	.w4(32'h3b7d1e14),
	.w5(32'h3c117bcb),
	.w6(32'hbbece9a5),
	.w7(32'hb92d2640),
	.w8(32'h3b90b926),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba968435),
	.w1(32'hb9d42073),
	.w2(32'h3a0ac05f),
	.w3(32'hbaea45e3),
	.w4(32'hba923cc7),
	.w5(32'hba428c55),
	.w6(32'hbae85977),
	.w7(32'hba2b1300),
	.w8(32'hb98b75af),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69fddd),
	.w1(32'h3b4b4921),
	.w2(32'h3b13b7e4),
	.w3(32'h3971f730),
	.w4(32'h3b0478b2),
	.w5(32'h3c04f91c),
	.w6(32'hbb430c4a),
	.w7(32'h3b57c4bd),
	.w8(32'h3bcb8479),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b644b48),
	.w1(32'h3af312cc),
	.w2(32'h3b10b112),
	.w3(32'h3a5ecb5f),
	.w4(32'h3a8cfb80),
	.w5(32'h3a96a391),
	.w6(32'h3a1d025f),
	.w7(32'h3a92e698),
	.w8(32'h3a552d7b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cd14e),
	.w1(32'hba94e55d),
	.w2(32'h3b52d64c),
	.w3(32'hbb48c6a6),
	.w4(32'hb78db2e1),
	.w5(32'hbb77d40a),
	.w6(32'hbb8d2c08),
	.w7(32'h3a2cff3b),
	.w8(32'hbb63d58e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb466e9a),
	.w1(32'hbadff594),
	.w2(32'hba928671),
	.w3(32'hbbd4d44b),
	.w4(32'hbba14c7d),
	.w5(32'hbac364d5),
	.w6(32'hbbd058ca),
	.w7(32'hbb71431e),
	.w8(32'hbad2f9ea),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac15567),
	.w1(32'hb7ae1e2f),
	.w2(32'hbaf89312),
	.w3(32'hba8f0971),
	.w4(32'hba90dbb0),
	.w5(32'h3ab987b3),
	.w6(32'hba37e12c),
	.w7(32'hbb103ff3),
	.w8(32'h3b21f318),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aec2e),
	.w1(32'hbac73a39),
	.w2(32'hbb21375b),
	.w3(32'h3b10d432),
	.w4(32'h39eaef7e),
	.w5(32'h3a8a93ff),
	.w6(32'hbb96c0a4),
	.w7(32'hbb3db55c),
	.w8(32'hbac14b2e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad02623),
	.w1(32'hba27f0e1),
	.w2(32'h3ad262ad),
	.w3(32'h3a80616b),
	.w4(32'h3b170fa2),
	.w5(32'h3933ca18),
	.w6(32'h3a3ed9cd),
	.w7(32'h3a9dc324),
	.w8(32'h3a27ed1e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bffe5),
	.w1(32'h3ba4f4f3),
	.w2(32'h3b9c134d),
	.w3(32'h3b36f8dc),
	.w4(32'h3bcb4103),
	.w5(32'h3b68ac4e),
	.w6(32'h39888da5),
	.w7(32'h3b904d03),
	.w8(32'h39d6f9e5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a7372),
	.w1(32'hba81c98e),
	.w2(32'hb9e58996),
	.w3(32'h39249dc5),
	.w4(32'hba91d50b),
	.w5(32'hbb93b444),
	.w6(32'hb91cba9e),
	.w7(32'hb979d429),
	.w8(32'hbb88fe97),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56d52d),
	.w1(32'hbaf01c3d),
	.w2(32'h3b99da9a),
	.w3(32'hbafd4310),
	.w4(32'h3b8af339),
	.w5(32'h3bdc48cf),
	.w6(32'hbbae830a),
	.w7(32'h3abbbe12),
	.w8(32'h3b6d81ff),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba566f92),
	.w1(32'h3a28c5af),
	.w2(32'h395e44d0),
	.w3(32'h3a1f0aaf),
	.w4(32'h3b578c22),
	.w5(32'h3c3cfc07),
	.w6(32'hbb875acc),
	.w7(32'h3b0d8886),
	.w8(32'h3bf95404),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ec16),
	.w1(32'h3c27088c),
	.w2(32'h3c80daa6),
	.w3(32'h3b7ee5b4),
	.w4(32'h3c367967),
	.w5(32'h3c4e205e),
	.w6(32'hbad2551f),
	.w7(32'h3c133285),
	.w8(32'h3c25fdaf),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d3fb),
	.w1(32'hba0c6a7a),
	.w2(32'hb9a9bf50),
	.w3(32'hbaa0bf6b),
	.w4(32'hb989ca07),
	.w5(32'h3b889b47),
	.w6(32'hbacd8bca),
	.w7(32'h38cf179c),
	.w8(32'h3b53bb1c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5d11),
	.w1(32'h3b0e6f2a),
	.w2(32'hb9a1233c),
	.w3(32'h3b84e879),
	.w4(32'h3b16b994),
	.w5(32'h3b204f61),
	.w6(32'h3afaed44),
	.w7(32'h3946d123),
	.w8(32'hb892dea8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e387ad),
	.w1(32'hba982657),
	.w2(32'h3ac03ddc),
	.w3(32'hbb81d617),
	.w4(32'h3b22f865),
	.w5(32'h3c3d95d8),
	.w6(32'hbc1be879),
	.w7(32'hbb8e9d86),
	.w8(32'h3bc882d4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd65cc0),
	.w1(32'h39dac2ef),
	.w2(32'hbb7b11b2),
	.w3(32'h3ac01afb),
	.w4(32'h3bcecc2b),
	.w5(32'h3b9c5933),
	.w6(32'hbc0176e5),
	.w7(32'hbb30851e),
	.w8(32'hbb5351cd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a28928),
	.w1(32'h3c0d5eea),
	.w2(32'h3c20217c),
	.w3(32'h3b793968),
	.w4(32'h3c01e3b4),
	.w5(32'h3bd80c2b),
	.w6(32'hbaf16513),
	.w7(32'h3bb1928f),
	.w8(32'h3b1c995a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f474ea),
	.w1(32'hbabd01a3),
	.w2(32'hbabc2c61),
	.w3(32'hbaa3d2b5),
	.w4(32'hba41b9f7),
	.w5(32'h3b276065),
	.w6(32'h3a68213f),
	.w7(32'hb98b701e),
	.w8(32'h3b36d60c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddd8a9),
	.w1(32'h3bc6b045),
	.w2(32'h3b6504e1),
	.w3(32'h3b9a31ff),
	.w4(32'h3bb8f81c),
	.w5(32'h39bcd581),
	.w6(32'h3b2026ff),
	.w7(32'h3b405d21),
	.w8(32'h3a357bb2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a9fd9),
	.w1(32'hb9d09dd0),
	.w2(32'hbac45d17),
	.w3(32'hba127a62),
	.w4(32'hba901d11),
	.w5(32'hbb2eb1b6),
	.w6(32'hb9a7188f),
	.w7(32'hb9d0df0f),
	.w8(32'h38975293),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1eed8),
	.w1(32'hbc02858b),
	.w2(32'hbc05957c),
	.w3(32'hbbaa3f1f),
	.w4(32'hbbe86fc8),
	.w5(32'hbb6f7c14),
	.w6(32'hbbb33bb4),
	.w7(32'hbbdee16b),
	.w8(32'hbb4ed66e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc131aae),
	.w1(32'hbc0bdacf),
	.w2(32'hbbe0cb21),
	.w3(32'hba830aa4),
	.w4(32'hbb1743bd),
	.w5(32'hbb484121),
	.w6(32'hbb403fb1),
	.w7(32'hbb5bf159),
	.w8(32'hba09a25e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afacd93),
	.w1(32'hbad492a9),
	.w2(32'hbbafeda8),
	.w3(32'hbacb837e),
	.w4(32'hbb1b98c4),
	.w5(32'h39d570f2),
	.w6(32'h38b1f908),
	.w7(32'hbaaf2db3),
	.w8(32'hbae6554f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c280),
	.w1(32'h3ba34946),
	.w2(32'h3c0ee9bf),
	.w3(32'h3b971048),
	.w4(32'h3adab5af),
	.w5(32'h388a679e),
	.w6(32'h3be3f582),
	.w7(32'h3ba5bb2e),
	.w8(32'hbb2b53d4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54f883),
	.w1(32'hba93d914),
	.w2(32'h3af0e3dd),
	.w3(32'hba89153b),
	.w4(32'h3a9632ba),
	.w5(32'h3ba5b2da),
	.w6(32'hbb927aaa),
	.w7(32'hbad005dc),
	.w8(32'h3b4d6fb3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4d883),
	.w1(32'hba51061c),
	.w2(32'hba1abce6),
	.w3(32'h3a49440b),
	.w4(32'hba9849e4),
	.w5(32'h3aaf7a10),
	.w6(32'hb9e1bf68),
	.w7(32'hba9dae8f),
	.w8(32'h3b0cb7c1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d4f65),
	.w1(32'h3aa5b638),
	.w2(32'h3a894a44),
	.w3(32'h3ab68ab2),
	.w4(32'h3a4ec364),
	.w5(32'hbb8686b0),
	.w6(32'h3a90f577),
	.w7(32'h3ac4403e),
	.w8(32'hbbc1e447),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cee42),
	.w1(32'hbb82a0c0),
	.w2(32'hba98eb9c),
	.w3(32'hbb5ebf5c),
	.w4(32'h39ed866b),
	.w5(32'h3b9fd8d3),
	.w6(32'hbbcad558),
	.w7(32'hbb0869f4),
	.w8(32'h3b6bf36b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babdee3),
	.w1(32'h3c014dde),
	.w2(32'h3be3bbc4),
	.w3(32'h3b9d49e0),
	.w4(32'h3bdedb47),
	.w5(32'hba3a0a29),
	.w6(32'h3bc2d51c),
	.w7(32'h3bec62ff),
	.w8(32'hba966f7e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c6c0e),
	.w1(32'hbaa63b20),
	.w2(32'hb9091da3),
	.w3(32'h38232451),
	.w4(32'h3a18be0b),
	.w5(32'hbb07e08f),
	.w6(32'hba821a1c),
	.w7(32'hb9121764),
	.w8(32'hbae06137),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8866),
	.w1(32'hbab9a00c),
	.w2(32'h391e199a),
	.w3(32'hbb8d8ee1),
	.w4(32'hb936552d),
	.w5(32'h3b01499e),
	.w6(32'hbc021d6f),
	.w7(32'hbb82e7a2),
	.w8(32'h3a41b45f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace4378),
	.w1(32'h3a917069),
	.w2(32'h3b3fd3d2),
	.w3(32'h37bddc28),
	.w4(32'h3b457c88),
	.w5(32'h3b1e7836),
	.w6(32'h397694bc),
	.w7(32'h3b4223c9),
	.w8(32'h3a3a6c01),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b9c5f),
	.w1(32'hba96d7c9),
	.w2(32'hbaaccce8),
	.w3(32'hbb22e2e0),
	.w4(32'hbb01d84c),
	.w5(32'h38edebe4),
	.w6(32'hb9b1af35),
	.w7(32'hbabf0ad1),
	.w8(32'hb983e919),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd06d06),
	.w1(32'hbbdd0332),
	.w2(32'hbbf005ce),
	.w3(32'hba61e7e6),
	.w4(32'hbb3fdef2),
	.w5(32'hbc17fc13),
	.w6(32'hbb8f5fab),
	.w7(32'hbb99ff1f),
	.w8(32'hbc0ccf4f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dbcc7),
	.w1(32'hbb589e53),
	.w2(32'hbb1d76f4),
	.w3(32'hbb8dade8),
	.w4(32'hbadfb87e),
	.w5(32'h391415ac),
	.w6(32'hbb898ce1),
	.w7(32'hbb05f418),
	.w8(32'hbb2866e3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9468094),
	.w1(32'hb9c67461),
	.w2(32'h39fe7444),
	.w3(32'hba60182c),
	.w4(32'hb9b39aea),
	.w5(32'hba1abfc1),
	.w6(32'hba4b5f4d),
	.w7(32'hbb0bbaff),
	.w8(32'hba26f6db),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5164fd),
	.w1(32'hbad643eb),
	.w2(32'hbb32a33d),
	.w3(32'hb9fb7a4f),
	.w4(32'hb8155bd4),
	.w5(32'hba466c3e),
	.w6(32'hbb1280ef),
	.w7(32'h39eea0c4),
	.w8(32'hbaed7f21),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72ce5a),
	.w1(32'hb94c040f),
	.w2(32'h39791f53),
	.w3(32'hba615f1e),
	.w4(32'hbad5ee70),
	.w5(32'hb98cd0c4),
	.w6(32'hba482047),
	.w7(32'hbac667aa),
	.w8(32'hb9da8fe2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3975fd),
	.w1(32'h3a8be440),
	.w2(32'h3a82d192),
	.w3(32'h3900cfab),
	.w4(32'h3a31f40b),
	.w5(32'hbb1048e2),
	.w6(32'hb8f265bc),
	.w7(32'h39f70002),
	.w8(32'hbb194a11),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb026c86),
	.w1(32'hbb1bad15),
	.w2(32'hbb031f87),
	.w3(32'hbb1f4219),
	.w4(32'hbb1ea040),
	.w5(32'hbab823fd),
	.w6(32'hbb671fd4),
	.w7(32'hbb2f8c33),
	.w8(32'hba88f6cc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3819a6e2),
	.w1(32'h3a367a57),
	.w2(32'h39bbd173),
	.w3(32'hba2b5c81),
	.w4(32'hba01f15f),
	.w5(32'h39f99f32),
	.w6(32'hb93b88a5),
	.w7(32'hb83c41d2),
	.w8(32'h39a7e2a0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d3161),
	.w1(32'hb8770bac),
	.w2(32'h3aacaae0),
	.w3(32'hbb1bb294),
	.w4(32'hba4c48ca),
	.w5(32'h39c5dad3),
	.w6(32'hba3fa867),
	.w7(32'hba200d07),
	.w8(32'h3a227af9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad684ba),
	.w1(32'h3ba125f7),
	.w2(32'h3b88f515),
	.w3(32'h3977715a),
	.w4(32'h3bc96163),
	.w5(32'h3c1a7a88),
	.w6(32'hbb3eea97),
	.w7(32'h3b94ad82),
	.w8(32'h3b985ccf),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50405b),
	.w1(32'h39b0fd1a),
	.w2(32'h3b16db61),
	.w3(32'hb9ce3174),
	.w4(32'h3ade72f6),
	.w5(32'h3b971df7),
	.w6(32'hbb2aff37),
	.w7(32'h3aa2ffc3),
	.w8(32'h3a24397e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c7680),
	.w1(32'h3ad73b53),
	.w2(32'h3a704377),
	.w3(32'h3ae73cb7),
	.w4(32'h3b92523d),
	.w5(32'h3b383783),
	.w6(32'hba8b853b),
	.w7(32'h3a990949),
	.w8(32'h3a2c447f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba598838),
	.w1(32'hb9693d80),
	.w2(32'h3aa1d4e7),
	.w3(32'hb8c40f2b),
	.w4(32'h3b01421b),
	.w5(32'hba33ebf2),
	.w6(32'hb9bb0d14),
	.w7(32'h3adc16b7),
	.w8(32'hbaa7ea79),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62f705),
	.w1(32'h3a5365dd),
	.w2(32'h3934f47a),
	.w3(32'hbac36047),
	.w4(32'hba84c9ef),
	.w5(32'h3a4631a6),
	.w6(32'hb9c5b100),
	.w7(32'hb9e3675c),
	.w8(32'h3a166495),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a496c05),
	.w1(32'h3a8c4a84),
	.w2(32'h3ad524cd),
	.w3(32'h3a70c2a7),
	.w4(32'h3a5ac6b2),
	.w5(32'h3a8c0de4),
	.w6(32'h3a588572),
	.w7(32'h3abf6284),
	.w8(32'hba145572),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad94b4f),
	.w1(32'h3b165b3e),
	.w2(32'h3b33cf4f),
	.w3(32'h3a85574b),
	.w4(32'hba2e5606),
	.w5(32'hb9a41a52),
	.w6(32'h39cb4078),
	.w7(32'h3a58d87f),
	.w8(32'hba650c0f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19e3c8),
	.w1(32'hbbe6f3ce),
	.w2(32'hbbb032d1),
	.w3(32'hbbfa9b36),
	.w4(32'hbb74697e),
	.w5(32'hbc0c69e3),
	.w6(32'hbc0f5b1d),
	.w7(32'hbbb89760),
	.w8(32'hbc362dac),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5133d),
	.w1(32'hbbc14682),
	.w2(32'hbb5ee3d5),
	.w3(32'hbbab26c8),
	.w4(32'hbb992a29),
	.w5(32'hba9ccd0a),
	.w6(32'hbbf27025),
	.w7(32'hbb891c91),
	.w8(32'hba390f0e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae41fa5),
	.w1(32'h3a2a11da),
	.w2(32'h3a08763b),
	.w3(32'h3b017cb3),
	.w4(32'h3a20b32f),
	.w5(32'h3a7587d3),
	.w6(32'h3aa7b8c6),
	.w7(32'h3a07ad85),
	.w8(32'h3a6e8273),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acad811),
	.w1(32'h3a123eb6),
	.w2(32'hbaaa10d0),
	.w3(32'h3a9f0943),
	.w4(32'hb882739b),
	.w5(32'h3aa0c2fe),
	.w6(32'h3abf3533),
	.w7(32'h3921674c),
	.w8(32'h3a7c0c86),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99d293),
	.w1(32'hb974489e),
	.w2(32'h392f3d56),
	.w3(32'h3a06fa76),
	.w4(32'h39945d35),
	.w5(32'hba42422c),
	.w6(32'h3a52ed26),
	.w7(32'h39f48a29),
	.w8(32'h391e3a7b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f829d),
	.w1(32'hb9cea902),
	.w2(32'hb9f3ff86),
	.w3(32'hb9317d61),
	.w4(32'h3aa9b511),
	.w5(32'h3af39586),
	.w6(32'hb91bbafe),
	.w7(32'h39c7dfaf),
	.w8(32'h3ab2f830),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8852a5),
	.w1(32'h3a9ebc07),
	.w2(32'h3a80552a),
	.w3(32'h3a1fa6da),
	.w4(32'h3834997e),
	.w5(32'hba01166d),
	.w6(32'h3a2e1899),
	.w7(32'h39781376),
	.w8(32'hba669637),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74f94),
	.w1(32'hbbb0316b),
	.w2(32'hbc08c883),
	.w3(32'hbb2d49f5),
	.w4(32'hbb22f7e6),
	.w5(32'hbbdf694a),
	.w6(32'hbb472dd4),
	.w7(32'hbb4432b6),
	.w8(32'hbbfe870e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9822ea3),
	.w1(32'hb9dbb99f),
	.w2(32'h3874e574),
	.w3(32'hba071cd0),
	.w4(32'h38313c02),
	.w5(32'h390d03a9),
	.w6(32'h393924eb),
	.w7(32'h38affd3d),
	.w8(32'h39390843),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fbef7),
	.w1(32'hbb31de42),
	.w2(32'h3b41a63e),
	.w3(32'hbb4f7f05),
	.w4(32'hbaded66d),
	.w5(32'hb9fb18d6),
	.w6(32'hbb708fe2),
	.w7(32'hbb4dd90e),
	.w8(32'hbac5d743),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule