module layer_8_featuremap_52(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f83eb),
	.w1(32'h39da14fc),
	.w2(32'h3a4e828d),
	.w3(32'h3b04058f),
	.w4(32'hba1369ac),
	.w5(32'hb8bdeefc),
	.w6(32'h3aa9486c),
	.w7(32'hba16ec25),
	.w8(32'hb97c4448),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3f13f),
	.w1(32'h37ac88f4),
	.w2(32'hb9dea4b6),
	.w3(32'hba0e53b3),
	.w4(32'h38c758d0),
	.w5(32'hb972eee7),
	.w6(32'hba800800),
	.w7(32'hb89efbd5),
	.w8(32'h38835609),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb163997),
	.w1(32'hbab9ea07),
	.w2(32'hba7b26ae),
	.w3(32'hbaf28229),
	.w4(32'hba9e3f43),
	.w5(32'hba921b6d),
	.w6(32'hbb0b2fdb),
	.w7(32'hbaaf09b8),
	.w8(32'hba3cc180),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcdcff),
	.w1(32'hba5729bd),
	.w2(32'h3ae48d24),
	.w3(32'h3b31380b),
	.w4(32'hba22aab8),
	.w5(32'h3a87c1f8),
	.w6(32'h3b3e9adf),
	.w7(32'h3b04a50e),
	.w8(32'h3b05be45),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc7beb),
	.w1(32'h393710de),
	.w2(32'h3a0914e8),
	.w3(32'h3a5e57a6),
	.w4(32'h3a0d021c),
	.w5(32'h3a34537a),
	.w6(32'h3a80876a),
	.w7(32'h3a275ef2),
	.w8(32'h3abf3184),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d037),
	.w1(32'hb96111fb),
	.w2(32'h3b2c8b1a),
	.w3(32'h3a06ccb0),
	.w4(32'hb99b2197),
	.w5(32'h3a34ec7b),
	.w6(32'h395cb045),
	.w7(32'h3ac44f27),
	.w8(32'h39a660fd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65705f1),
	.w1(32'h3893265c),
	.w2(32'hb7627026),
	.w3(32'h3904806f),
	.w4(32'h375f20d0),
	.w5(32'hb946f189),
	.w6(32'h376d10a2),
	.w7(32'h392e067a),
	.w8(32'h38a45ef1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3661e),
	.w1(32'hba11d872),
	.w2(32'hbad76556),
	.w3(32'hba44b2c6),
	.w4(32'h3a972154),
	.w5(32'hb910aced),
	.w6(32'hba2b4f2f),
	.w7(32'hba50633b),
	.w8(32'hbaec967e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08ac69),
	.w1(32'hb8b51fc2),
	.w2(32'hba08d90f),
	.w3(32'h3a00a8ea),
	.w4(32'hb8f12de1),
	.w5(32'hb98006ef),
	.w6(32'h3865ea86),
	.w7(32'hb9157e06),
	.w8(32'hba2328c6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403582),
	.w1(32'hba596218),
	.w2(32'hba6d08cc),
	.w3(32'hbb428839),
	.w4(32'hbaadfd17),
	.w5(32'hb9de260e),
	.w6(32'h38e35049),
	.w7(32'hbb2dec74),
	.w8(32'hbb03eebb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8103605),
	.w1(32'hba64d701),
	.w2(32'hb9cde285),
	.w3(32'h3b19aeb7),
	.w4(32'hba7b6e88),
	.w5(32'hbb0efe97),
	.w6(32'h3a08c43c),
	.w7(32'hb792f2cb),
	.w8(32'hba41ae81),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b77a2b),
	.w1(32'h3a9f4922),
	.w2(32'h3a98eca8),
	.w3(32'h3af363f3),
	.w4(32'h3b1c6184),
	.w5(32'h3b0cd716),
	.w6(32'h3a0866d0),
	.w7(32'h38252076),
	.w8(32'h39e196ec),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b6a47),
	.w1(32'h3a337cda),
	.w2(32'h3a3b5244),
	.w3(32'hba57b546),
	.w4(32'h3912e3b8),
	.w5(32'h39f9ca01),
	.w6(32'hba377ba8),
	.w7(32'h37284e14),
	.w8(32'h3abee77c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b7007),
	.w1(32'h3a5680ba),
	.w2(32'h3a6e53da),
	.w3(32'h3a8f3582),
	.w4(32'h3a214156),
	.w5(32'h39d96cfd),
	.w6(32'h3a4c7c68),
	.w7(32'h3a61ebf3),
	.w8(32'h39e56912),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8373f),
	.w1(32'h39c756dc),
	.w2(32'h39c56385),
	.w3(32'h3a03a380),
	.w4(32'h398fa213),
	.w5(32'h38df0274),
	.w6(32'h39b5d9d4),
	.w7(32'h39eaf4c4),
	.w8(32'hb886c8ba),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ffe8e4),
	.w1(32'hb9319261),
	.w2(32'hb7d40347),
	.w3(32'hb60be2c8),
	.w4(32'hb9051372),
	.w5(32'hb6f34f63),
	.w6(32'hb969a332),
	.w7(32'hb99c411d),
	.w8(32'hb92d6625),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bb9f5),
	.w1(32'hbad1bf88),
	.w2(32'hbaa52c3c),
	.w3(32'hba67fb44),
	.w4(32'hb99c7944),
	.w5(32'h38918895),
	.w6(32'hbad084f6),
	.w7(32'hba62d290),
	.w8(32'hb9f68f02),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d368e),
	.w1(32'h3a768aed),
	.w2(32'hb72f8390),
	.w3(32'hba9041aa),
	.w4(32'h393a3ea8),
	.w5(32'h3a05e65c),
	.w6(32'hba499144),
	.w7(32'hba16815a),
	.w8(32'h3a58c8c9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb191120),
	.w1(32'hbb1200f0),
	.w2(32'h39c028f8),
	.w3(32'h3bfdbd60),
	.w4(32'h3a90c523),
	.w5(32'h3aca2031),
	.w6(32'hba3654da),
	.w7(32'hbb14d0e5),
	.w8(32'hba2148f9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71d5b2),
	.w1(32'h3bc00333),
	.w2(32'h3b2c8e25),
	.w3(32'h3b1c5fbf),
	.w4(32'h3ab82602),
	.w5(32'h3ade2594),
	.w6(32'h3b9bdfbc),
	.w7(32'h3b1cf74d),
	.w8(32'h3b0c0c32),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2d76b),
	.w1(32'h39a8b54e),
	.w2(32'hb95f1a82),
	.w3(32'h3a90f6ca),
	.w4(32'hb9a31bef),
	.w5(32'hba63fc0a),
	.w6(32'hbaf0f2db),
	.w7(32'hba025aa8),
	.w8(32'h3a8d3994),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a182d9),
	.w1(32'hba077537),
	.w2(32'hba53601a),
	.w3(32'hbaab9ccf),
	.w4(32'hba861773),
	.w5(32'hba821a53),
	.w6(32'hbb0f064f),
	.w7(32'hbac83b9d),
	.w8(32'hbaa7e17d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9af5b3),
	.w1(32'h3b94be43),
	.w2(32'h3b89e8db),
	.w3(32'h3b8b6fc2),
	.w4(32'h3b47e839),
	.w5(32'h3ab6467d),
	.w6(32'h3abe12a2),
	.w7(32'h3a2d5096),
	.w8(32'h3a12700f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a300d38),
	.w1(32'h39d97e14),
	.w2(32'hb9672f5c),
	.w3(32'hb97b0b15),
	.w4(32'hb9c19c31),
	.w5(32'hba51c696),
	.w6(32'hb9bad171),
	.w7(32'hb9a43dd5),
	.w8(32'hbab32db4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a45e3),
	.w1(32'hba20992a),
	.w2(32'hba6fa956),
	.w3(32'hbab4c831),
	.w4(32'hbaa68cb7),
	.w5(32'hba3454e3),
	.w6(32'hbaa428c6),
	.w7(32'hba888e9d),
	.w8(32'hb8fbb816),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2f5b0),
	.w1(32'h39495b76),
	.w2(32'h3b2204ad),
	.w3(32'h3b497f33),
	.w4(32'h3b38e327),
	.w5(32'h3b712a09),
	.w6(32'h3ab8fd05),
	.w7(32'h3a95d446),
	.w8(32'h3adfb9b7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b69344),
	.w1(32'hba184df6),
	.w2(32'hb934db2d),
	.w3(32'hb911329a),
	.w4(32'hb973fddc),
	.w5(32'h393f92ec),
	.w6(32'hb9ea6c01),
	.w7(32'hb921f0f9),
	.w8(32'hba1bb3b7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4843f1),
	.w1(32'hb94f32b6),
	.w2(32'hbbdd54f0),
	.w3(32'h3c6ff1ff),
	.w4(32'h3c8ae11d),
	.w5(32'hbbaa4058),
	.w6(32'hbc0d0c3c),
	.w7(32'hb951971e),
	.w8(32'h3ad6e5e1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae29ac),
	.w1(32'hba89210f),
	.w2(32'h3a96e3f6),
	.w3(32'h39a1b2a7),
	.w4(32'hb9f46107),
	.w5(32'h3a834ed7),
	.w6(32'h3aaedd83),
	.w7(32'h3990d834),
	.w8(32'h3a35b666),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9195c3b),
	.w1(32'h37c1ca7d),
	.w2(32'hb8cbc979),
	.w3(32'h37ac60a3),
	.w4(32'h38faa26e),
	.w5(32'hb8a86dba),
	.w6(32'hb85c0125),
	.w7(32'h399b5edd),
	.w8(32'hb9fee787),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf093b),
	.w1(32'hba9b63cb),
	.w2(32'hbade6b4f),
	.w3(32'hbab2acd4),
	.w4(32'hbaa24f69),
	.w5(32'hbab0e535),
	.w6(32'hbaa84340),
	.w7(32'hbaa02e3c),
	.w8(32'hba8b8521),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4c04c),
	.w1(32'hba00493a),
	.w2(32'hb8d942dc),
	.w3(32'h3a94a470),
	.w4(32'h39cbcd57),
	.w5(32'h3a2462f0),
	.w6(32'hba5a6cc8),
	.w7(32'h39dd31ec),
	.w8(32'h3ae1ca2a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cffb42),
	.w1(32'hba406518),
	.w2(32'hba348cb8),
	.w3(32'hba273287),
	.w4(32'hba05f90b),
	.w5(32'hb9edb5ea),
	.w6(32'hb7791d76),
	.w7(32'hb9716635),
	.w8(32'hb6c652d0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c12be),
	.w1(32'h390f4cce),
	.w2(32'hb4c3adac),
	.w3(32'hba2a1b7a),
	.w4(32'hba252a6b),
	.w5(32'h3954b9dc),
	.w6(32'hb9c16946),
	.w7(32'hba812bd2),
	.w8(32'h3a713445),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c09c0),
	.w1(32'h3b18739b),
	.w2(32'h3ac296ce),
	.w3(32'h390876a9),
	.w4(32'h3a47ca6c),
	.w5(32'h39d91caa),
	.w6(32'hba1e8995),
	.w7(32'hb7550be3),
	.w8(32'hb95e9c05),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca11ec),
	.w1(32'hba8a9c45),
	.w2(32'hbac2255e),
	.w3(32'h3a0e0fa4),
	.w4(32'h3992384c),
	.w5(32'hb8caaa1b),
	.w6(32'hba655430),
	.w7(32'hbab927fa),
	.w8(32'hbacaf666),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa1040),
	.w1(32'hba38d4bf),
	.w2(32'hb9fddd68),
	.w3(32'hba2c18f5),
	.w4(32'hba01b2f2),
	.w5(32'hb992eced),
	.w6(32'hba68b839),
	.w7(32'hba3620da),
	.w8(32'hb89f9752),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb636a4f3),
	.w1(32'h3998170d),
	.w2(32'h399313a4),
	.w3(32'h3a0de217),
	.w4(32'h3a4389c7),
	.w5(32'h39a84a84),
	.w6(32'h390462e4),
	.w7(32'h3a3ead02),
	.w8(32'h3ac31ad7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57b838),
	.w1(32'h3a431d16),
	.w2(32'h3a31a636),
	.w3(32'h3a66693b),
	.w4(32'h3a08bfb5),
	.w5(32'h39894565),
	.w6(32'h3a01648a),
	.w7(32'h3a50bf17),
	.w8(32'hb9fa3a75),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b6ea95),
	.w1(32'hba02630a),
	.w2(32'hb98ae301),
	.w3(32'hb990dde1),
	.w4(32'hba3b94a8),
	.w5(32'hb9a32e83),
	.w6(32'hba34c94c),
	.w7(32'hb9618271),
	.w8(32'hb88f441c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47fe83),
	.w1(32'h3aef2b50),
	.w2(32'h3bdde382),
	.w3(32'h3b3a0d68),
	.w4(32'h3adff8c1),
	.w5(32'h3b955eb6),
	.w6(32'h3b7dcd5e),
	.w7(32'h3ae83fa9),
	.w8(32'h3bc35d49),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eeea4),
	.w1(32'hbb9ae44d),
	.w2(32'h3978716e),
	.w3(32'hba9a692c),
	.w4(32'h3b33b040),
	.w5(32'hb9db1056),
	.w6(32'h3b12b5fc),
	.w7(32'h3b4cf3fa),
	.w8(32'hbca45c55),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0257),
	.w1(32'h3bfc4e64),
	.w2(32'h3bc915ae),
	.w3(32'h3b00ebda),
	.w4(32'hbcf28148),
	.w5(32'hbcc3dd27),
	.w6(32'hbc5dce53),
	.w7(32'h3c37b57d),
	.w8(32'h3b9c446b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcab5bb),
	.w1(32'hbbb98126),
	.w2(32'hbbc6afb5),
	.w3(32'hba884085),
	.w4(32'h3a3a526b),
	.w5(32'hbb564ba1),
	.w6(32'h3af11aa0),
	.w7(32'h3b3be604),
	.w8(32'h3a87dff8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed8b3f),
	.w1(32'hbb277925),
	.w2(32'h3a3ee1ed),
	.w3(32'hbb7b5921),
	.w4(32'h37862807),
	.w5(32'hbb523069),
	.w6(32'h3b0755d0),
	.w7(32'h3b48cbf3),
	.w8(32'hbb8a8e8c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fcb89),
	.w1(32'h3b7acb66),
	.w2(32'hbbbacae0),
	.w3(32'hbaa270c2),
	.w4(32'hbb723ff4),
	.w5(32'hbb4517f5),
	.w6(32'hbb34aad4),
	.w7(32'hbb605b08),
	.w8(32'hbcc7a26f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d847c),
	.w1(32'h3d28911b),
	.w2(32'h3a92881e),
	.w3(32'h3b95acb6),
	.w4(32'hbc29368e),
	.w5(32'hba95e29f),
	.w6(32'h3cb22007),
	.w7(32'h3b9cdb77),
	.w8(32'hbaf6ee2d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec8af6),
	.w1(32'h3ab84877),
	.w2(32'h3a8fb69e),
	.w3(32'hbc67a0c8),
	.w4(32'hbb0fc8c5),
	.w5(32'hbbf16356),
	.w6(32'hbc1a624f),
	.w7(32'hbbb345dc),
	.w8(32'hbc38fbf4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e01e),
	.w1(32'hbb0b510e),
	.w2(32'h3c49fa07),
	.w3(32'h3c2d2277),
	.w4(32'h3c352d03),
	.w5(32'h3cbf7667),
	.w6(32'hbc5065d1),
	.w7(32'hbb9c1f76),
	.w8(32'h3aae79ee),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf24b4d),
	.w1(32'hbb4a9919),
	.w2(32'h3b0a2a7c),
	.w3(32'hbae907e8),
	.w4(32'h3ad58874),
	.w5(32'h3a1866f6),
	.w6(32'h3be7413d),
	.w7(32'h3b979c2a),
	.w8(32'h3b669247),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd46e3),
	.w1(32'hbab42d95),
	.w2(32'hbaa69abc),
	.w3(32'hbbd3643b),
	.w4(32'hba499c4c),
	.w5(32'hb7c2b6ae),
	.w6(32'hbb5d1f06),
	.w7(32'h3ad63859),
	.w8(32'h3c1e5651),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc259b0e),
	.w1(32'hbbce978c),
	.w2(32'hbb83a365),
	.w3(32'hbaaf1d6e),
	.w4(32'hba6c933b),
	.w5(32'hbb9bd838),
	.w6(32'h3ba9ba97),
	.w7(32'h3b7afbb2),
	.w8(32'h3c62b075),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e25b4),
	.w1(32'h3d1c5ad5),
	.w2(32'h3ad3c576),
	.w3(32'hbc430863),
	.w4(32'h39b6eaa5),
	.w5(32'hbaa79749),
	.w6(32'hbcd26723),
	.w7(32'hbbc4a952),
	.w8(32'hbafc1e39),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85a4fc),
	.w1(32'hbaa7f252),
	.w2(32'h3a8849f7),
	.w3(32'hb922293a),
	.w4(32'h3ad33bf3),
	.w5(32'h3bf9c250),
	.w6(32'hb95ba4af),
	.w7(32'hbb95facf),
	.w8(32'hbcb151b2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c092ccc),
	.w1(32'h3c5ad509),
	.w2(32'hbc6e9241),
	.w3(32'hbad8cb3d),
	.w4(32'hbca4aacf),
	.w5(32'hbc987890),
	.w6(32'h3accc65c),
	.w7(32'hbbc75d92),
	.w8(32'hbbdd68ce),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcdd51),
	.w1(32'hbb335193),
	.w2(32'hbc4d3bb2),
	.w3(32'hbb342a23),
	.w4(32'hbbae1ef2),
	.w5(32'hbb1796ba),
	.w6(32'hbc1cfa90),
	.w7(32'hbcb3849a),
	.w8(32'hbaa557a6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c20c),
	.w1(32'hbc2a98b6),
	.w2(32'hbbe43cd6),
	.w3(32'hbc2fc032),
	.w4(32'h3b923c3a),
	.w5(32'h3a5c239f),
	.w6(32'h3a0d738a),
	.w7(32'hbc182521),
	.w8(32'h3b38efe9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d93b),
	.w1(32'hbb778a72),
	.w2(32'hbb7df53e),
	.w3(32'hbb024368),
	.w4(32'hb9fb178c),
	.w5(32'hbc22d83a),
	.w6(32'hbb8191e9),
	.w7(32'hbb9e3ddd),
	.w8(32'hbb2d05e1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5af9ff),
	.w1(32'hbb518dd9),
	.w2(32'h3ba72282),
	.w3(32'h3c17877c),
	.w4(32'h3bc0f86f),
	.w5(32'h3c3b4bf9),
	.w6(32'hbc11af2f),
	.w7(32'h3a315b99),
	.w8(32'h3b47b784),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8512ca),
	.w1(32'h3bcec4cb),
	.w2(32'hbb409629),
	.w3(32'hbc84771b),
	.w4(32'hbc31bb98),
	.w5(32'hbbf1ade0),
	.w6(32'h3b47d123),
	.w7(32'hbb26262d),
	.w8(32'hbc435929),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b62d4),
	.w1(32'h3d4826ec),
	.w2(32'h3c90d917),
	.w3(32'h3c2be30c),
	.w4(32'h3ce7b4d7),
	.w5(32'hbc092ef8),
	.w6(32'hbd18f0d8),
	.w7(32'h3bb00634),
	.w8(32'hbc4fbc06),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba917a07),
	.w1(32'hbb827a74),
	.w2(32'hbc120779),
	.w3(32'hbc20f396),
	.w4(32'hbbb3c315),
	.w5(32'hbc0e2bb6),
	.w6(32'hbbb487e6),
	.w7(32'hbc5778a2),
	.w8(32'h3b6963e3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a763),
	.w1(32'hbb43a049),
	.w2(32'hba2fb5d1),
	.w3(32'hbafd2383),
	.w4(32'h3b6c3f14),
	.w5(32'h3ad9b254),
	.w6(32'h3bc03cf5),
	.w7(32'h3bbfad50),
	.w8(32'h3bdb8b5d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598624),
	.w1(32'h3c8e041e),
	.w2(32'hbbc9c1a9),
	.w3(32'hbc46dcc4),
	.w4(32'hba6d3d3c),
	.w5(32'hbaa15129),
	.w6(32'h3c6a9b34),
	.w7(32'h3c1636ac),
	.w8(32'h398b3c74),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1389),
	.w1(32'hbb31c21d),
	.w2(32'hbaa39582),
	.w3(32'hbb874e97),
	.w4(32'hba413518),
	.w5(32'hbb1e3a8f),
	.w6(32'h3afebf1a),
	.w7(32'h3ba732ce),
	.w8(32'h3b27536b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79b3b8),
	.w1(32'hbb62a9dc),
	.w2(32'hbb67a475),
	.w3(32'hbaef72dc),
	.w4(32'hba85363b),
	.w5(32'hbb3bb3be),
	.w6(32'hba46d1c3),
	.w7(32'hb910a3b0),
	.w8(32'h3a66d6cf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6612c2),
	.w1(32'hbab7cbbf),
	.w2(32'hbab5c954),
	.w3(32'hbb209f78),
	.w4(32'hbae57469),
	.w5(32'hbb213ae3),
	.w6(32'hb9e41603),
	.w7(32'h3ae8c89a),
	.w8(32'hbb8fe671),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7ffc),
	.w1(32'h3cb6f722),
	.w2(32'h3c9c56c3),
	.w3(32'hbc23cb42),
	.w4(32'hb98482e0),
	.w5(32'hbbd0ff12),
	.w6(32'hbc3ea23f),
	.w7(32'hbbc68c32),
	.w8(32'h3abb7fac),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f27a),
	.w1(32'hbaf00833),
	.w2(32'h3a82a45b),
	.w3(32'hbba3c600),
	.w4(32'hb85e597c),
	.w5(32'hbaa9d32c),
	.w6(32'h3b02b818),
	.w7(32'h3b102817),
	.w8(32'h3c627def),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4466f),
	.w1(32'hba6fcf31),
	.w2(32'hbadeec7e),
	.w3(32'h3c30c9ff),
	.w4(32'hba91a920),
	.w5(32'hbbf69639),
	.w6(32'h3ae928cb),
	.w7(32'h3bba3150),
	.w8(32'h3b824d7e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae3ca),
	.w1(32'hbb844436),
	.w2(32'hba3260e7),
	.w3(32'hbaf3dfd9),
	.w4(32'h3ac01453),
	.w5(32'hbaa698cf),
	.w6(32'h3ba573c8),
	.w7(32'h3bd93941),
	.w8(32'h3abb761f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc63eb),
	.w1(32'hbb1d2f71),
	.w2(32'h3b0c6f02),
	.w3(32'hbb5a77f2),
	.w4(32'h3a1807ff),
	.w5(32'hba26f43b),
	.w6(32'h3b649ca2),
	.w7(32'h3b603427),
	.w8(32'h3bc39ddd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7d86),
	.w1(32'hbb5717ff),
	.w2(32'h39e1301f),
	.w3(32'hbb66ae30),
	.w4(32'h3733c5b9),
	.w5(32'hbb37553a),
	.w6(32'h3bbefbcd),
	.w7(32'h3c025c5b),
	.w8(32'h3cb98ce5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e56a0),
	.w1(32'h3d281755),
	.w2(32'h3c3329a0),
	.w3(32'hba841d72),
	.w4(32'h3b9ab586),
	.w5(32'h3be216d5),
	.w6(32'h3c964149),
	.w7(32'hbca881bf),
	.w8(32'h3b97f086),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8727eb),
	.w1(32'h3b74c779),
	.w2(32'h3b8a8ad8),
	.w3(32'hbb93ca64),
	.w4(32'hbb4bcebf),
	.w5(32'hbbbb8f58),
	.w6(32'h3b775c0b),
	.w7(32'h3b927c44),
	.w8(32'h3b5aded2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba56092),
	.w1(32'hbb754f0e),
	.w2(32'hbb8deb5e),
	.w3(32'hb9c3aa6a),
	.w4(32'h3ac3937c),
	.w5(32'hbae93414),
	.w6(32'h3b5fff02),
	.w7(32'h3b8c5813),
	.w8(32'h3b7d060f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f5f9),
	.w1(32'hbb631a3b),
	.w2(32'hbaeb09d0),
	.w3(32'hbb6ff40f),
	.w4(32'h39c02d02),
	.w5(32'hbb3e65de),
	.w6(32'h3b9ffe59),
	.w7(32'h3b291491),
	.w8(32'h3c76f087),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc99b87),
	.w1(32'hba8bf3c2),
	.w2(32'hbb1678f3),
	.w3(32'h3c309c16),
	.w4(32'h3a546631),
	.w5(32'hbb612d03),
	.w6(32'h3b462da7),
	.w7(32'h3c10220c),
	.w8(32'h3c68de60),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79db09),
	.w1(32'hb94e9e41),
	.w2(32'hbba45832),
	.w3(32'h3b263328),
	.w4(32'h3b3cfa93),
	.w5(32'hbb3b44ac),
	.w6(32'h3c009287),
	.w7(32'h3bbbc4aa),
	.w8(32'h3afa919a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006327),
	.w1(32'h3bac49b6),
	.w2(32'hbaa91661),
	.w3(32'hbb25ea35),
	.w4(32'hbb2b2879),
	.w5(32'h3985ff95),
	.w6(32'h3ac4993e),
	.w7(32'hbaedb66c),
	.w8(32'hba389027),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e54ee),
	.w1(32'h3d71d5df),
	.w2(32'h3ca1761c),
	.w3(32'hbc4e85b5),
	.w4(32'h3cadff37),
	.w5(32'h3bbef675),
	.w6(32'hba998a73),
	.w7(32'h3c09ca1f),
	.w8(32'hbb3c41c0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb893b76),
	.w1(32'hbbb2f2d7),
	.w2(32'hbb146932),
	.w3(32'hbbea7918),
	.w4(32'hbba1bb67),
	.w5(32'hbbfd2300),
	.w6(32'h3b1b80dc),
	.w7(32'hbad56a22),
	.w8(32'hb9d62a8a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99566b),
	.w1(32'h3ba6b2b7),
	.w2(32'hbb77ba40),
	.w3(32'hbb226ff2),
	.w4(32'hbb072e9b),
	.w5(32'hbb87ebcd),
	.w6(32'h3c250a3a),
	.w7(32'hb89509ef),
	.w8(32'h3c8a1fbf),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63dc34),
	.w1(32'h3ca0fae6),
	.w2(32'h3d25dd20),
	.w3(32'hbc5c8869),
	.w4(32'h3cabd228),
	.w5(32'h3ca53e61),
	.w6(32'h3c805256),
	.w7(32'h3c2ebb5d),
	.w8(32'h3b81bf97),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c07a),
	.w1(32'h3afdcde2),
	.w2(32'h3b7a8b1c),
	.w3(32'h3b97a453),
	.w4(32'h3ab87b8f),
	.w5(32'h3b8c2508),
	.w6(32'h3b50ba7a),
	.w7(32'hb95cd956),
	.w8(32'h3b4241d0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe390b7),
	.w1(32'hbb08c0a2),
	.w2(32'h3b8ff8ab),
	.w3(32'hbb657b2b),
	.w4(32'h3a22dc83),
	.w5(32'hbaa050b4),
	.w6(32'h3c1a1766),
	.w7(32'h3bf6e7be),
	.w8(32'hbc7282e6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa1f1d),
	.w1(32'hbac8812f),
	.w2(32'h3c907d66),
	.w3(32'h3c7dd946),
	.w4(32'h3c81a284),
	.w5(32'h3d0414f2),
	.w6(32'hbc7d7f69),
	.w7(32'hbbb09321),
	.w8(32'h3b59f1b8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94409a),
	.w1(32'hbb9088ac),
	.w2(32'hbb39a5a2),
	.w3(32'hbc1e8214),
	.w4(32'hbac00f29),
	.w5(32'hbb95e0b0),
	.w6(32'hbb29bd24),
	.w7(32'h3bd82e10),
	.w8(32'hbb0991b1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5de9b),
	.w1(32'hbaad83d1),
	.w2(32'h3a637a73),
	.w3(32'hbc720ddc),
	.w4(32'hbc3d1212),
	.w5(32'hb9bc4ccb),
	.w6(32'hbb96cf4a),
	.w7(32'h3b97b535),
	.w8(32'hbc6f0759),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafa316),
	.w1(32'hba9ea3b1),
	.w2(32'h3c8850fd),
	.w3(32'h3c7646fc),
	.w4(32'h3c7706be),
	.w5(32'h3cf9f0f3),
	.w6(32'hbc60b0b7),
	.w7(32'hbb9b1ce2),
	.w8(32'hbc49bba6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb276d2),
	.w1(32'h3a36d547),
	.w2(32'h3c80d3d5),
	.w3(32'h3c6181f4),
	.w4(32'h3c614cd6),
	.w5(32'h3cdbd269),
	.w6(32'hbc39093f),
	.w7(32'hbb7ca167),
	.w8(32'hba9d3c07),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5b0f8),
	.w1(32'hbb2cf09a),
	.w2(32'h3aa39403),
	.w3(32'h39f0bfcc),
	.w4(32'hbb185732),
	.w5(32'h3ab56390),
	.w6(32'hba64e98c),
	.w7(32'hb98231f5),
	.w8(32'h3b28fb60),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81e7f5),
	.w1(32'h3c8cd10b),
	.w2(32'h3c712ae2),
	.w3(32'hbb9f7a18),
	.w4(32'hbc9d78fc),
	.w5(32'hbb620296),
	.w6(32'h3bc860a9),
	.w7(32'hbc9080b8),
	.w8(32'h3b04135b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f5382),
	.w1(32'hbb075149),
	.w2(32'hbb553ed1),
	.w3(32'hbab7ee54),
	.w4(32'hba7090a7),
	.w5(32'hbb31f03e),
	.w6(32'h3aa5baf4),
	.w7(32'h3a81e2eb),
	.w8(32'hbb129b71),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e64bc),
	.w1(32'hbcbd919c),
	.w2(32'hbc5b5975),
	.w3(32'h3ac39d1d),
	.w4(32'h3c85ce07),
	.w5(32'hba3f9f0b),
	.w6(32'h3b8bb878),
	.w7(32'hbc143883),
	.w8(32'hbb568dc6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bcb6c),
	.w1(32'hbc970c01),
	.w2(32'hbc177bfc),
	.w3(32'hbab820ae),
	.w4(32'h3a2dea81),
	.w5(32'h3be27d9c),
	.w6(32'h3a9baf47),
	.w7(32'hb92cd265),
	.w8(32'h3c0d1ee1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9766),
	.w1(32'hbc1a0a3f),
	.w2(32'hb8c9cd89),
	.w3(32'h3c9cf720),
	.w4(32'h3c6cc748),
	.w5(32'h3c7c81eb),
	.w6(32'h3c4fce47),
	.w7(32'h3b8f9321),
	.w8(32'h3c2b96a9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc527422),
	.w1(32'hbb6c4c75),
	.w2(32'h3a778501),
	.w3(32'h3c84de53),
	.w4(32'h3bbe39aa),
	.w5(32'h3bde883a),
	.w6(32'h3d1f884b),
	.w7(32'h3c6ea400),
	.w8(32'h3c58c508),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9acb4),
	.w1(32'hba7c2af3),
	.w2(32'hbb350b50),
	.w3(32'h3bc56881),
	.w4(32'hba8122a9),
	.w5(32'hbb59936e),
	.w6(32'h3b0fef76),
	.w7(32'h3bef3c65),
	.w8(32'h3ac82d3e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77840d),
	.w1(32'hbb8d7b82),
	.w2(32'hbb131a27),
	.w3(32'hbbf7b35e),
	.w4(32'h375bfbeb),
	.w5(32'hbb7544f3),
	.w6(32'h3aacc9bc),
	.w7(32'h3b351855),
	.w8(32'hbb4d2874),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fcf35),
	.w1(32'h3c7440fe),
	.w2(32'hbc15526d),
	.w3(32'hbc413b85),
	.w4(32'hbaefbfc3),
	.w5(32'hbc0849d3),
	.w6(32'h3b09994a),
	.w7(32'hbb235f45),
	.w8(32'h3ad49fa7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16c8c),
	.w1(32'hbb427a27),
	.w2(32'hbbb76e13),
	.w3(32'hbb86989d),
	.w4(32'hbb693aae),
	.w5(32'hbba7bb01),
	.w6(32'hb9b4a984),
	.w7(32'h3adb1b37),
	.w8(32'h3cdc2395),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a544a),
	.w1(32'hbb962419),
	.w2(32'hbc12b982),
	.w3(32'h3b79f0f2),
	.w4(32'h3b646c60),
	.w5(32'hbc03c748),
	.w6(32'h3cb32b13),
	.w7(32'h3c481672),
	.w8(32'hbaf798b2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39d56),
	.w1(32'hbb0eadf0),
	.w2(32'h3b36477f),
	.w3(32'hbb19dd18),
	.w4(32'hbb5d72b5),
	.w5(32'hba1e9c15),
	.w6(32'hba74beb6),
	.w7(32'hb9a7125e),
	.w8(32'hbbda34d9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac58d3a),
	.w1(32'hba4b051e),
	.w2(32'h3bc1eac1),
	.w3(32'h3b963395),
	.w4(32'h3ba6e07b),
	.w5(32'h3c3452cf),
	.w6(32'hbbcf26cb),
	.w7(32'hbb30cf84),
	.w8(32'h3b099f0a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34faaa),
	.w1(32'hbb8acabc),
	.w2(32'hbb3aee81),
	.w3(32'hbb6f3c30),
	.w4(32'hbb497394),
	.w5(32'hbc15e55d),
	.w6(32'hb990743c),
	.w7(32'h3b299b4a),
	.w8(32'h3cbda6cb),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c69a5f8),
	.w1(32'hbba532fd),
	.w2(32'h3b7bf3da),
	.w3(32'h3b79804e),
	.w4(32'hbca78022),
	.w5(32'h3c604d96),
	.w6(32'h3c40d970),
	.w7(32'hbc9591a0),
	.w8(32'hba42fc69),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c18a9),
	.w1(32'hba8fb196),
	.w2(32'hba91095c),
	.w3(32'h3b24131a),
	.w4(32'h3c040f42),
	.w5(32'hba3331fe),
	.w6(32'hbc43b657),
	.w7(32'hbacde1ca),
	.w8(32'h3b3af4f8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cafe4),
	.w1(32'h3a6c3f9b),
	.w2(32'h3a8986f1),
	.w3(32'hbc3b9711),
	.w4(32'hbbe9d733),
	.w5(32'hbc24bb39),
	.w6(32'hba6a1de9),
	.w7(32'h3befbc70),
	.w8(32'h3c695b0c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b271b7a),
	.w1(32'h3b0bc68c),
	.w2(32'h3b825c8f),
	.w3(32'hbbe754ef),
	.w4(32'hbca25ee5),
	.w5(32'hbc27ca39),
	.w6(32'h3be0ede3),
	.w7(32'h3c55dbfc),
	.w8(32'h3be25489),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b613b3b),
	.w1(32'hbb975cca),
	.w2(32'hbc1e774c),
	.w3(32'hbc94c64e),
	.w4(32'hbb1a033a),
	.w5(32'hbb84015d),
	.w6(32'hbc404c2b),
	.w7(32'hbcc60b7b),
	.w8(32'hb9ed8282),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33ba70),
	.w1(32'hbb1b33c9),
	.w2(32'h3c1ae03c),
	.w3(32'hbbc172dd),
	.w4(32'hbc342d56),
	.w5(32'h39be2e16),
	.w6(32'hb9ac92ec),
	.w7(32'h3c8ea6d4),
	.w8(32'h3c716314),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc63b3),
	.w1(32'h3a8a8998),
	.w2(32'hba1d545d),
	.w3(32'hbc451547),
	.w4(32'hbc98a9f4),
	.w5(32'hbb8071c5),
	.w6(32'h3d1edd29),
	.w7(32'h3c591d48),
	.w8(32'h3b437b02),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20785f),
	.w1(32'hba8f1e67),
	.w2(32'h38cf3f27),
	.w3(32'hbc537c69),
	.w4(32'hbc30a9d8),
	.w5(32'hbc3a1cf2),
	.w6(32'hba716999),
	.w7(32'h3c0dd152),
	.w8(32'hbacd7962),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd4084),
	.w1(32'h3b0528c1),
	.w2(32'h3b18f08b),
	.w3(32'h3ae676d7),
	.w4(32'h3b8336ee),
	.w5(32'h3aa8c9cf),
	.w6(32'hbbb41300),
	.w7(32'hb904b6b3),
	.w8(32'hbaff1f27),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec42f),
	.w1(32'h3a9a0854),
	.w2(32'h398af199),
	.w3(32'h3b8aadf9),
	.w4(32'h3c299dc7),
	.w5(32'hba54e978),
	.w6(32'hbc76bbca),
	.w7(32'hbb335dde),
	.w8(32'hbccb762f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06c8ef),
	.w1(32'h3c65890e),
	.w2(32'hbaab7181),
	.w3(32'h3c74dcf7),
	.w4(32'hbc225216),
	.w5(32'hbc991cd1),
	.w6(32'h3b889ba4),
	.w7(32'hbbe5a45c),
	.w8(32'h3d068e87),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c9ff),
	.w1(32'h3bda249a),
	.w2(32'h3bb450f3),
	.w3(32'hbcc913d6),
	.w4(32'hbd140df2),
	.w5(32'hbca9fb6a),
	.w6(32'h3d42bbe9),
	.w7(32'h3d02350d),
	.w8(32'h3c30a44c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f078a),
	.w1(32'hbc35c609),
	.w2(32'h3c5b4814),
	.w3(32'hbc57bac0),
	.w4(32'h3b079784),
	.w5(32'h3c94d936),
	.w6(32'hbccf2ef4),
	.w7(32'hbc8e058b),
	.w8(32'h3c035383),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d7d79),
	.w1(32'h3bc80c98),
	.w2(32'h3c9bbf91),
	.w3(32'h3c07f7f6),
	.w4(32'h3cbd674d),
	.w5(32'hbaa369a8),
	.w6(32'h3b8c291e),
	.w7(32'h3c6352e3),
	.w8(32'h3a3a1daa),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953e332),
	.w1(32'hbc058849),
	.w2(32'hbaf10233),
	.w3(32'hbb9af696),
	.w4(32'hbbcb6593),
	.w5(32'h3b89d7ba),
	.w6(32'hbb792131),
	.w7(32'hbb6add39),
	.w8(32'h3bd57354),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1a320),
	.w1(32'hbc89ff72),
	.w2(32'hbbf5186a),
	.w3(32'h3c1e060f),
	.w4(32'hbc85c24c),
	.w5(32'hbb268fe2),
	.w6(32'h3b1f2889),
	.w7(32'h3b881ef9),
	.w8(32'hbc829997),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc138212),
	.w1(32'hb9d3554f),
	.w2(32'hbb96f0d3),
	.w3(32'h3c44160e),
	.w4(32'h3cc826b8),
	.w5(32'h3c503ed9),
	.w6(32'hbc31420d),
	.w7(32'hbc2aeddd),
	.w8(32'h3c783cbd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9671d7),
	.w1(32'h3b86dcdd),
	.w2(32'hbc08d2de),
	.w3(32'hbc0c392d),
	.w4(32'hbcc3b2fe),
	.w5(32'hbbda7171),
	.w6(32'h3cb5cefa),
	.w7(32'h3b1eded6),
	.w8(32'h3b8c5035),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6fe19),
	.w1(32'h3c0dec92),
	.w2(32'hbc4ed97a),
	.w3(32'hbb846d7c),
	.w4(32'hbb12703c),
	.w5(32'h3c8c2671),
	.w6(32'h3c0300b6),
	.w7(32'hbcb8302b),
	.w8(32'h3c41704c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc469889),
	.w1(32'hbc7106b2),
	.w2(32'hbc636881),
	.w3(32'hbc82deb0),
	.w4(32'hbccfd485),
	.w5(32'hbc90dcdf),
	.w6(32'h3b845864),
	.w7(32'h3bae3105),
	.w8(32'h3ae05673),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d516),
	.w1(32'h3b940ca5),
	.w2(32'hb9cb34c4),
	.w3(32'hbbaefe8a),
	.w4(32'hbb2c4b62),
	.w5(32'hbc40004e),
	.w6(32'hba8c3d59),
	.w7(32'h3ab0a127),
	.w8(32'hbc4e94c6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f11d2),
	.w1(32'h3b489e04),
	.w2(32'hbc46aff8),
	.w3(32'hbb065fbb),
	.w4(32'hbbd95fae),
	.w5(32'hbc99101e),
	.w6(32'hbb9cc0d1),
	.w7(32'hbaa23de5),
	.w8(32'hbb0683f9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule