module layer_8_featuremap_97(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb41ae6),
	.w1(32'hbb89b4cd),
	.w2(32'h3a847a58),
	.w3(32'h3c073420),
	.w4(32'hbc01a330),
	.w5(32'hbc22de57),
	.w6(32'hbbfc4694),
	.w7(32'hbcf01107),
	.w8(32'h3c9dbe7a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c516e),
	.w1(32'hbbb4635b),
	.w2(32'hbc482735),
	.w3(32'h3ca072c2),
	.w4(32'h3b7758a8),
	.w5(32'hbc89f757),
	.w6(32'h3cbec591),
	.w7(32'hbc1d65ab),
	.w8(32'hbb63a844),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65ed50),
	.w1(32'hbbe62857),
	.w2(32'h3ba59240),
	.w3(32'hbc00e5bb),
	.w4(32'hbc0a669d),
	.w5(32'h3c2b0f9b),
	.w6(32'h3c90cec6),
	.w7(32'hbc385cec),
	.w8(32'h3bae9689),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc710ccd),
	.w1(32'hb99b3c01),
	.w2(32'hba33631e),
	.w3(32'hb92e1cc5),
	.w4(32'h3c8ae9a2),
	.w5(32'h3b8f3aeb),
	.w6(32'hbaa5b42b),
	.w7(32'h3cddaa20),
	.w8(32'hbc68f1e1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc943dd6),
	.w1(32'h3bad8bc8),
	.w2(32'h3b49ce14),
	.w3(32'h3b70b2ad),
	.w4(32'h3b2c5f47),
	.w5(32'h3ce2eda8),
	.w6(32'hbbcbc501),
	.w7(32'h3d213ce1),
	.w8(32'hbc93ef6e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc8731),
	.w1(32'h3aa5a2a9),
	.w2(32'h3c0570b3),
	.w3(32'h3ca34871),
	.w4(32'hbb90b9db),
	.w5(32'hbb3ab7e8),
	.w6(32'h3b1b97b8),
	.w7(32'h3c4aa259),
	.w8(32'hbbb0da31),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fcee2),
	.w1(32'h3b9c994f),
	.w2(32'hbcd0486a),
	.w3(32'hbc8b4c83),
	.w4(32'hbb24b7d8),
	.w5(32'hbbf5d2ba),
	.w6(32'h3bb841a4),
	.w7(32'h3b661929),
	.w8(32'hbbf07c4a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c0990),
	.w1(32'hbbb9a2d8),
	.w2(32'hbd0c6a9e),
	.w3(32'h3adbb10b),
	.w4(32'hbbe2b23b),
	.w5(32'hbc92c82d),
	.w6(32'h3ca6276a),
	.w7(32'hbbe7393a),
	.w8(32'hbd267c25),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf21ad5),
	.w1(32'h3c389468),
	.w2(32'hbb8cddf2),
	.w3(32'h3b409d61),
	.w4(32'h3b0a4059),
	.w5(32'hba7f27f9),
	.w6(32'h3c8c065b),
	.w7(32'h3b98796c),
	.w8(32'hbbddbb8a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e8168),
	.w1(32'h3bd4b618),
	.w2(32'hbb24c15f),
	.w3(32'h3bef9f6d),
	.w4(32'h3b0354a6),
	.w5(32'h3b2b35e8),
	.w6(32'h3ba2f0f1),
	.w7(32'hbaf3e62e),
	.w8(32'h3b708448),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc509bfd),
	.w1(32'h3bd7b8ca),
	.w2(32'h3b664556),
	.w3(32'h3b69866f),
	.w4(32'h3cf40cff),
	.w5(32'hbb9b15f3),
	.w6(32'h3bacb96d),
	.w7(32'h3b2de94a),
	.w8(32'hbcc8270a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97035),
	.w1(32'h3af18edc),
	.w2(32'h3b60ffec),
	.w3(32'hbbed11aa),
	.w4(32'h3c2f61bd),
	.w5(32'hbb82fca8),
	.w6(32'hbbf1e7f0),
	.w7(32'h3cad63e9),
	.w8(32'hbc96639b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c1dec),
	.w1(32'h3b10ae27),
	.w2(32'hbaa4e0ab),
	.w3(32'h3b817551),
	.w4(32'hb9b1217c),
	.w5(32'hba688570),
	.w6(32'h3c910548),
	.w7(32'h3a837905),
	.w8(32'hb9e42900),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b6de),
	.w1(32'h3a68c1ac),
	.w2(32'h3a9ce31c),
	.w3(32'h3ad742c0),
	.w4(32'h3a8fb477),
	.w5(32'h3a2f058e),
	.w6(32'h3a598dce),
	.w7(32'h3a1813b4),
	.w8(32'h39f5efcd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b14a12),
	.w1(32'hb727360a),
	.w2(32'hb83743f6),
	.w3(32'h392ea63d),
	.w4(32'h38f827b3),
	.w5(32'h3859149e),
	.w6(32'h397e9e3f),
	.w7(32'h396c68e5),
	.w8(32'h3925aa82),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb3f74),
	.w1(32'h3a92fce5),
	.w2(32'h3aa2834d),
	.w3(32'h3ade5cfb),
	.w4(32'h3ae65431),
	.w5(32'h3adffe9b),
	.w6(32'h3aa1c565),
	.w7(32'h3aaf18f4),
	.w8(32'h3ae20d59),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacda878),
	.w1(32'hbac0a75e),
	.w2(32'hba8dc1e8),
	.w3(32'hbab8f535),
	.w4(32'h39154bf9),
	.w5(32'h3ae158a1),
	.w6(32'hb978b266),
	.w7(32'h3b62ccc8),
	.w8(32'h3b80cf50),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d24468),
	.w1(32'hb9448d2b),
	.w2(32'hbb1c322f),
	.w3(32'h3b80eef0),
	.w4(32'h3b6d65d8),
	.w5(32'h3a4b4556),
	.w6(32'h3b94ab5e),
	.w7(32'h3b41ff8e),
	.w8(32'hba1cfc1b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc21c22),
	.w1(32'h3c4927ff),
	.w2(32'hbb8d3e23),
	.w3(32'h3cb7aa86),
	.w4(32'h3d15f0fa),
	.w5(32'h3c4034fc),
	.w6(32'h3a92fd37),
	.w7(32'h3c0d082d),
	.w8(32'hbc3f666a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af5c28),
	.w1(32'h3b9fbf22),
	.w2(32'h3c22a0db),
	.w3(32'h3ac196fc),
	.w4(32'h3c177abe),
	.w5(32'h3c38ba53),
	.w6(32'hbb86426f),
	.w7(32'h3b2d8feb),
	.w8(32'h3bd76bf3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be70286),
	.w1(32'h3be27e3a),
	.w2(32'h3c01b604),
	.w3(32'hbb21e711),
	.w4(32'h3a34a6d7),
	.w5(32'h3bf3eaa0),
	.w6(32'hbc2d33d0),
	.w7(32'hbbf2ca43),
	.w8(32'h3b20dc33),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb644d96),
	.w1(32'hbc267d86),
	.w2(32'hbbc07243),
	.w3(32'hbb4eba7b),
	.w4(32'hbc41ca72),
	.w5(32'hbbe1d5d2),
	.w6(32'hba31f781),
	.w7(32'hbbd55263),
	.w8(32'hbae5d8e0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc853261),
	.w1(32'hbacc1602),
	.w2(32'hbbaffae0),
	.w3(32'hbc17027d),
	.w4(32'h3cab2475),
	.w5(32'h3c26b1bf),
	.w6(32'hbc04ff44),
	.w7(32'h3c32f2d8),
	.w8(32'h3ae267b7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e1ad),
	.w1(32'hb9f7a81c),
	.w2(32'hb9e8bd6b),
	.w3(32'hba261127),
	.w4(32'h3838c080),
	.w5(32'h3a53d9c5),
	.w6(32'hbaf026ab),
	.w7(32'h3a8bd236),
	.w8(32'h3b2d8a0b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd27a),
	.w1(32'h3bb975cf),
	.w2(32'h3c05213a),
	.w3(32'h398ce585),
	.w4(32'h39ad7f0e),
	.w5(32'h3b84dcaf),
	.w6(32'h3aeec569),
	.w7(32'h399c53c7),
	.w8(32'h3bf9b979),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104303),
	.w1(32'hbb85db1a),
	.w2(32'hbb311937),
	.w3(32'hbb494152),
	.w4(32'h3c028f3b),
	.w5(32'h3bf660b9),
	.w6(32'hbc1254d4),
	.w7(32'h3a8019d2),
	.w8(32'h3adc5cfd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24005a),
	.w1(32'hbaf863f2),
	.w2(32'hba8647bb),
	.w3(32'hbb495c1a),
	.w4(32'hba9cbbd8),
	.w5(32'hb9ae9e90),
	.w6(32'hbb38dac7),
	.w7(32'hba843bdf),
	.w8(32'hba064780),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c1f92),
	.w1(32'h3cb4239f),
	.w2(32'h3c96cefc),
	.w3(32'hba9cdecb),
	.w4(32'h3d31fa68),
	.w5(32'h3da4759a),
	.w6(32'hbc6e9127),
	.w7(32'h3cc16b22),
	.w8(32'h3d170768),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46a784),
	.w1(32'h39f8878f),
	.w2(32'h3a2bda8d),
	.w3(32'h3b5364e6),
	.w4(32'h3beefdb4),
	.w5(32'h3bb233f3),
	.w6(32'hb9d1b859),
	.w7(32'h3b1ad777),
	.w8(32'h3a9a8514),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82941c),
	.w1(32'h396069c2),
	.w2(32'h3a558d51),
	.w3(32'h3a80e77d),
	.w4(32'h3a96bde9),
	.w5(32'h3ad1c676),
	.w6(32'h3a989829),
	.w7(32'h3a352c6a),
	.w8(32'h3b0cc742),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81b49f),
	.w1(32'hbb828e66),
	.w2(32'hba520360),
	.w3(32'hbbe186be),
	.w4(32'hbbf5917a),
	.w5(32'hbbb81ea6),
	.w6(32'hbc04b96a),
	.w7(32'hbbf26629),
	.w8(32'hbbba9b8e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9f805),
	.w1(32'hba0b041c),
	.w2(32'h3b195042),
	.w3(32'hbaf2e73e),
	.w4(32'hbad872df),
	.w5(32'h3b33a7df),
	.w6(32'hbb1fe7ee),
	.w7(32'hbab5dd14),
	.w8(32'h3b05cfda),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968b185),
	.w1(32'h3958a209),
	.w2(32'h3847d197),
	.w3(32'h3859fa64),
	.w4(32'h38f3989f),
	.w5(32'h37886498),
	.w6(32'h3842952c),
	.w7(32'h3920de71),
	.w8(32'h38d7cb30),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d9e23),
	.w1(32'h38efe2eb),
	.w2(32'hb83f5ee0),
	.w3(32'h384de4ad),
	.w4(32'h39040643),
	.w5(32'hb857cfce),
	.w6(32'h3819d89c),
	.w7(32'h38a4931a),
	.w8(32'hb89c6620),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6d5e7),
	.w1(32'hba7b738a),
	.w2(32'h3aeb46d9),
	.w3(32'hbb7f4732),
	.w4(32'hbc0b9c4a),
	.w5(32'hbb9c79ea),
	.w6(32'hbb2dcc63),
	.w7(32'hbbc71683),
	.w8(32'hbb13d5a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b9cd0),
	.w1(32'h3bef77c0),
	.w2(32'h3b983326),
	.w3(32'h3bc70a5a),
	.w4(32'h3c424dbe),
	.w5(32'h3c2fd9ea),
	.w6(32'h3b0a7994),
	.w7(32'h3b82bee6),
	.w8(32'h3b887a4c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395313fc),
	.w1(32'hb89a8f77),
	.w2(32'h39354fab),
	.w3(32'h39236f5b),
	.w4(32'h3a37e88e),
	.w5(32'h3abaf166),
	.w6(32'h3a05a0fc),
	.w7(32'h3a5704fc),
	.w8(32'h3a74941d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f38df),
	.w1(32'hbba1ef96),
	.w2(32'hbb5727ad),
	.w3(32'hbb38ae16),
	.w4(32'hbb9fcd9f),
	.w5(32'hbb4cfe53),
	.w6(32'hbb7b56c1),
	.w7(32'hbba8a467),
	.w8(32'hbb820694),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9622ba8),
	.w1(32'h37c9f796),
	.w2(32'hb8d4777d),
	.w3(32'hb94dec08),
	.w4(32'h390859b1),
	.w5(32'h37b0ed9c),
	.w6(32'h37baf7c4),
	.w7(32'h3987695f),
	.w8(32'h39709874),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57cf74),
	.w1(32'hba743896),
	.w2(32'hba3c3fdd),
	.w3(32'hbafa7797),
	.w4(32'hbaa5afd2),
	.w5(32'hbabf4184),
	.w6(32'hbabaf605),
	.w7(32'hb9c050eb),
	.w8(32'hba251246),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13c84e),
	.w1(32'h3c7a2c91),
	.w2(32'h3cc282d2),
	.w3(32'h3cb986b3),
	.w4(32'h3cd195f4),
	.w5(32'h3d001253),
	.w6(32'h3c5eb754),
	.w7(32'h3c430cb0),
	.w8(32'h3cb0a97d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6a37),
	.w1(32'h3afe26f8),
	.w2(32'hbadcfb19),
	.w3(32'h3b5c891f),
	.w4(32'h3b6059c7),
	.w5(32'h39a95d38),
	.w6(32'h3a181b07),
	.w7(32'h3a1f5237),
	.w8(32'hbaa8b108),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9809b81),
	.w1(32'hba124c04),
	.w2(32'h365b5846),
	.w3(32'hb9bef5b9),
	.w4(32'hba180e08),
	.w5(32'h393e5cd0),
	.w6(32'hba610a47),
	.w7(32'hba821bd5),
	.w8(32'hba322f32),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55ed58),
	.w1(32'h3b8f6d33),
	.w2(32'h3b9289fe),
	.w3(32'h3baace24),
	.w4(32'h3c0a1346),
	.w5(32'h3c14a2c0),
	.w6(32'h3b8f280c),
	.w7(32'h3bd2e7a3),
	.w8(32'h3bce125f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02cf0),
	.w1(32'hbb1ecab2),
	.w2(32'hbbb20b7f),
	.w3(32'h3b22f12e),
	.w4(32'h3c22afb1),
	.w5(32'h3af0f8ec),
	.w6(32'hbb3e7c01),
	.w7(32'h3b552fba),
	.w8(32'hbb2f2d78),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f57a),
	.w1(32'h3b7f9b99),
	.w2(32'h36ad71f0),
	.w3(32'h3b1413fb),
	.w4(32'h3b2e371b),
	.w5(32'hba899b43),
	.w6(32'hbacaabf3),
	.w7(32'hbb26c2db),
	.w8(32'hbb7b91a5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65a5008),
	.w1(32'h378268c1),
	.w2(32'hb8234ffe),
	.w3(32'h3803d5ba),
	.w4(32'h3853487a),
	.w5(32'hb7cb3640),
	.w6(32'h386eefc3),
	.w7(32'h38887147),
	.w8(32'hb768d9a9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49fd57),
	.w1(32'h3b7cfb05),
	.w2(32'h3b9ea577),
	.w3(32'h3b32abe5),
	.w4(32'h3c7d66a9),
	.w5(32'h3c464cbb),
	.w6(32'hbab9b2ef),
	.w7(32'h3bde1dfe),
	.w8(32'h3ac23448),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71575),
	.w1(32'h3a33fa8a),
	.w2(32'hb885f5c7),
	.w3(32'h3b41cf1d),
	.w4(32'h3ae075a2),
	.w5(32'h3acb1db6),
	.w6(32'h3b0c8273),
	.w7(32'h3a6f3ea8),
	.w8(32'h3a41cb16),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806629),
	.w1(32'hb957f4c8),
	.w2(32'hbab2531e),
	.w3(32'h3b868f01),
	.w4(32'h3bc32aff),
	.w5(32'h3b6ec4e9),
	.w6(32'hb96f77b5),
	.w7(32'h3b1a2721),
	.w8(32'h3a7bbb2d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53ebd2),
	.w1(32'hbc6ea6a5),
	.w2(32'hbbea2f91),
	.w3(32'hbc3f4b54),
	.w4(32'hbc8a640e),
	.w5(32'hbc28b088),
	.w6(32'hbc61dbde),
	.w7(32'hbca2153a),
	.w8(32'hbc47edb2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2843b4),
	.w1(32'hbb8334f1),
	.w2(32'h3a71d778),
	.w3(32'h3c9233c9),
	.w4(32'h3ce3d101),
	.w5(32'h3c776acc),
	.w6(32'h3c4e02d2),
	.w7(32'h3cd5f0cc),
	.w8(32'h3c1e8917),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb54938),
	.w1(32'hbba8db08),
	.w2(32'hbb2c63c8),
	.w3(32'h3b15a4b4),
	.w4(32'h3c0666b0),
	.w5(32'h3bc8cffe),
	.w6(32'h3b0b35d1),
	.w7(32'h3c092003),
	.w8(32'h3ba184d2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92bd6c),
	.w1(32'h3c3616a4),
	.w2(32'h3c17b363),
	.w3(32'h3b90440e),
	.w4(32'h3c0f31b6),
	.w5(32'h3bb2f3dd),
	.w6(32'h3b23b875),
	.w7(32'h3b33f78f),
	.w8(32'hbadcf6f4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728a6b7),
	.w1(32'h3919666a),
	.w2(32'h36b311dc),
	.w3(32'h38f394c0),
	.w4(32'h39886625),
	.w5(32'h390463d2),
	.w6(32'h38a21009),
	.w7(32'h3954cf75),
	.w8(32'h38b29d94),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7027af),
	.w1(32'h3c1018f6),
	.w2(32'h3bcb9a92),
	.w3(32'hbb8c4c0b),
	.w4(32'h3c2d08d4),
	.w5(32'h3c2e48d1),
	.w6(32'hbb7d7301),
	.w7(32'hbb41b673),
	.w8(32'hbbf96025),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b903897),
	.w1(32'h385da33d),
	.w2(32'hb99ea243),
	.w3(32'hbb38fa3c),
	.w4(32'hbba7bbee),
	.w5(32'hbba29199),
	.w6(32'hbb693ea7),
	.w7(32'hbaf2c53d),
	.w8(32'hba65f586),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982a54a),
	.w1(32'hbbb0d966),
	.w2(32'hbc016594),
	.w3(32'h3c014813),
	.w4(32'h3bfe632c),
	.w5(32'h3a88bd5a),
	.w6(32'h3c223406),
	.w7(32'h3c098ee0),
	.w8(32'h3aeb55c7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefa77),
	.w1(32'hb9c242ce),
	.w2(32'hb901063b),
	.w3(32'hba72c51a),
	.w4(32'h3ba0d118),
	.w5(32'h3b48ddb2),
	.w6(32'h3a4db273),
	.w7(32'h3bb39ac8),
	.w8(32'h3b67740a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fbea6),
	.w1(32'h39a90fec),
	.w2(32'h3b69bd47),
	.w3(32'h3811e9f5),
	.w4(32'h3b3f6e9d),
	.w5(32'h3b9af1d4),
	.w6(32'h3b400109),
	.w7(32'h3b856659),
	.w8(32'h3bb72505),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd0cd),
	.w1(32'h3ace8be6),
	.w2(32'h3af925e8),
	.w3(32'h3aafc62d),
	.w4(32'h3b221bee),
	.w5(32'h3b8df9f4),
	.w6(32'h3b3386ae),
	.w7(32'h3b2aebeb),
	.w8(32'h3b9688eb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de42f),
	.w1(32'hba1e6e5c),
	.w2(32'hb98dea7b),
	.w3(32'hba82de6b),
	.w4(32'hb9d48691),
	.w5(32'hb9becab8),
	.w6(32'hba80f311),
	.w7(32'hb914e1b3),
	.w8(32'hba0f404a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b449b27),
	.w1(32'h3c14bd7d),
	.w2(32'h3c27c408),
	.w3(32'h3c38c91c),
	.w4(32'h3c834a32),
	.w5(32'h3c852f29),
	.w6(32'h3ae5d565),
	.w7(32'h3b9434dc),
	.w8(32'h3bd87489),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7cbaa),
	.w1(32'h3acbb44f),
	.w2(32'h3a901452),
	.w3(32'h3acdfc3a),
	.w4(32'h3b7b80e3),
	.w5(32'h3b0f4d19),
	.w6(32'h3b9c1816),
	.w7(32'h3bfe0d6f),
	.w8(32'h3b627bdd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64818e),
	.w1(32'hbb2199b3),
	.w2(32'hbb0edc8f),
	.w3(32'hbb32b85b),
	.w4(32'hba6021ca),
	.w5(32'hb9af5945),
	.w6(32'hbb185895),
	.w7(32'hba063407),
	.w8(32'hba1c5dd8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a539aff),
	.w1(32'hba2abfb0),
	.w2(32'hbb6aa571),
	.w3(32'h3b29820d),
	.w4(32'h3b513287),
	.w5(32'h3afd33c4),
	.w6(32'h3ab192a1),
	.w7(32'h3aff39cb),
	.w8(32'h3af22d5e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eea57),
	.w1(32'h38664c3a),
	.w2(32'h3af74cca),
	.w3(32'h3b1c3ab5),
	.w4(32'h3ba5e11d),
	.w5(32'h3b64ee51),
	.w6(32'h3bc13c87),
	.w7(32'h3b8395cd),
	.w8(32'h3b94b366),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba072fc6),
	.w1(32'h38b471fe),
	.w2(32'h3b5b213f),
	.w3(32'hbb0c9d73),
	.w4(32'h3b582373),
	.w5(32'h3bef1e52),
	.w6(32'hbba08e86),
	.w7(32'hbb1f283e),
	.w8(32'h3aad2bd8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7a162),
	.w1(32'hba462eb3),
	.w2(32'hba0b074a),
	.w3(32'hbadf0b98),
	.w4(32'h39fac2ee),
	.w5(32'h3a7d7674),
	.w6(32'hba296a5b),
	.w7(32'h3a49a84f),
	.w8(32'h388887a2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a8c24),
	.w1(32'hbb0824f3),
	.w2(32'h3a5c3712),
	.w3(32'hbc07bbfd),
	.w4(32'h3c87640d),
	.w5(32'h3c94a442),
	.w6(32'hbae6ae2f),
	.w7(32'h3c882cbc),
	.w8(32'h3c853cbf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6208),
	.w1(32'hbabcf4e9),
	.w2(32'hba844ebc),
	.w3(32'hbb0d4a2d),
	.w4(32'hbafd211f),
	.w5(32'hbac45404),
	.w6(32'hbb057ac0),
	.w7(32'hbad46e3a),
	.w8(32'hbaa72f9b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b75139),
	.w1(32'h3a961ea2),
	.w2(32'h3a854742),
	.w3(32'h3a014164),
	.w4(32'h3b98c812),
	.w5(32'h3bb64887),
	.w6(32'hb8ee8a64),
	.w7(32'h3b91cee8),
	.w8(32'h3ba195bf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1bbf),
	.w1(32'hbad08fcd),
	.w2(32'hbac70bd6),
	.w3(32'hbaaad72d),
	.w4(32'h3983d306),
	.w5(32'hb894ca05),
	.w6(32'hb98456d2),
	.w7(32'h3953683c),
	.w8(32'hba8ae1d1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897f7e),
	.w1(32'h3b6faca3),
	.w2(32'h3b5ebbc0),
	.w3(32'h3b9095b6),
	.w4(32'h3b7526fb),
	.w5(32'h3c380ff5),
	.w6(32'h3b84a0c5),
	.w7(32'hba395355),
	.w8(32'h3b3d8a05),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f27fb1),
	.w1(32'h386bc9ac),
	.w2(32'h380f2ec7),
	.w3(32'h3712a256),
	.w4(32'h38068a92),
	.w5(32'h376589cf),
	.w6(32'hb7db7a37),
	.w7(32'hb70c99a9),
	.w8(32'h3684657a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a113f),
	.w1(32'hbb4e788c),
	.w2(32'hbb3188c5),
	.w3(32'hbb1d0bcf),
	.w4(32'hba205ea7),
	.w5(32'h39a2326f),
	.w6(32'hbb7bb4da),
	.w7(32'hba831d94),
	.w8(32'h3a875fbe),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927c0f3),
	.w1(32'hb697d492),
	.w2(32'h3a3cf186),
	.w3(32'hb7b8f4b6),
	.w4(32'h3b66796b),
	.w5(32'h3b4c1561),
	.w6(32'hb85acc90),
	.w7(32'h3be7d29f),
	.w8(32'h3b11bcae),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc021152),
	.w1(32'hbb2d9e1e),
	.w2(32'h3c143e65),
	.w3(32'h3c5652a4),
	.w4(32'h3cb71d78),
	.w5(32'h3c272933),
	.w6(32'h3b5117b5),
	.w7(32'h3c0ee561),
	.w8(32'h3abf9cfa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba286ea),
	.w1(32'hbbb6bd92),
	.w2(32'h3ba9b913),
	.w3(32'h3c23742b),
	.w4(32'h3b91ab23),
	.w5(32'h3ba90f73),
	.w6(32'h3aebddb9),
	.w7(32'h3a6b51f0),
	.w8(32'hb9cc33df),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fde8a),
	.w1(32'hbc41368e),
	.w2(32'hbbbee32c),
	.w3(32'h3bb1fe52),
	.w4(32'h3bebaf58),
	.w5(32'hbc7a621d),
	.w6(32'hbbadd610),
	.w7(32'hbbe2197c),
	.w8(32'hbc610e49),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8927f),
	.w1(32'h3bff79d9),
	.w2(32'h3d3fdfc3),
	.w3(32'hbc7225e7),
	.w4(32'hbcc7bb4c),
	.w5(32'hbd22e0c0),
	.w6(32'h3c2849f6),
	.w7(32'hbbf690c1),
	.w8(32'hbc4c6b57),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d43bb3e),
	.w1(32'h3c1d015c),
	.w2(32'h3cae369f),
	.w3(32'hbc83f0e1),
	.w4(32'hbb8567ff),
	.w5(32'h3c88afc6),
	.w6(32'hbbe7d435),
	.w7(32'h3cb9b881),
	.w8(32'h3b8b6bbe),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c453271),
	.w1(32'h3c1d5d30),
	.w2(32'h3ca01e5d),
	.w3(32'hbb4c03db),
	.w4(32'h3c8a4acf),
	.w5(32'h3b986dde),
	.w6(32'hbb7e77c3),
	.w7(32'h3a0420ed),
	.w8(32'h3b821f8f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4becb),
	.w1(32'h3ca36283),
	.w2(32'h3ce94cff),
	.w3(32'h3c977971),
	.w4(32'hbc1150af),
	.w5(32'h3cbccafe),
	.w6(32'h3c9e3995),
	.w7(32'hbc4ea1c7),
	.w8(32'h3d2237ec),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdba71),
	.w1(32'h3baed920),
	.w2(32'hbc8f7917),
	.w3(32'h3c4cef1c),
	.w4(32'h3d197931),
	.w5(32'h3d14fc0d),
	.w6(32'h3ccb4749),
	.w7(32'h3c840287),
	.w8(32'h3c8e6b37),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87602f),
	.w1(32'hbb5952dc),
	.w2(32'hbc19d99e),
	.w3(32'h3cd9a09e),
	.w4(32'hbc1a054e),
	.w5(32'hbc8ad39b),
	.w6(32'h3a2bd4cf),
	.w7(32'h3b625e1d),
	.w8(32'h3c64d334),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15f7d8),
	.w1(32'h3d020e38),
	.w2(32'hbc7dbb39),
	.w3(32'hbbb344f6),
	.w4(32'hbb956ebe),
	.w5(32'hbaa9cab0),
	.w6(32'h3c8f2968),
	.w7(32'hbc62e603),
	.w8(32'h3bd5426a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb618c12),
	.w1(32'hbc7324c0),
	.w2(32'h3b598b15),
	.w3(32'h3bb7dbab),
	.w4(32'hbc14d8d3),
	.w5(32'h3a795432),
	.w6(32'h3c009486),
	.w7(32'hbb0c0923),
	.w8(32'h3ae5e3a4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c788ad6),
	.w1(32'h3c0330df),
	.w2(32'h3b0dcd84),
	.w3(32'hbc27618a),
	.w4(32'hbb378efc),
	.w5(32'hbc275cb2),
	.w6(32'hbc22fa28),
	.w7(32'hbc31d933),
	.w8(32'hbb65b060),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a986d54),
	.w1(32'h3c039b74),
	.w2(32'h3c95426c),
	.w3(32'hbba4fffc),
	.w4(32'hbbb51472),
	.w5(32'hbcc190a7),
	.w6(32'h3c030c1c),
	.w7(32'hbb85ff5c),
	.w8(32'h3c92a004),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d40b87c),
	.w1(32'h3c5e03f2),
	.w2(32'hbca5e465),
	.w3(32'h3b1597e9),
	.w4(32'h3c3e6a11),
	.w5(32'h3c901947),
	.w6(32'h3c8f139b),
	.w7(32'hbc0db386),
	.w8(32'h3c128759),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbad799),
	.w1(32'hbbbcb8a7),
	.w2(32'hbcda983e),
	.w3(32'h3ca130b2),
	.w4(32'hbbbbb3ae),
	.w5(32'h3c7f1c6e),
	.w6(32'hbba7794f),
	.w7(32'hbc64b74f),
	.w8(32'hbbe06afe),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f2462),
	.w1(32'hbab3dfe2),
	.w2(32'h3c368213),
	.w3(32'h3cddd2bc),
	.w4(32'h3a9b3c3e),
	.w5(32'hbc0c1584),
	.w6(32'h3cbf9edf),
	.w7(32'hbc13a8f8),
	.w8(32'hbad52e49),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be16f17),
	.w1(32'h3cb7ab2b),
	.w2(32'hbbd956b5),
	.w3(32'hb9c4dd68),
	.w4(32'h3c225905),
	.w5(32'hbafed28f),
	.w6(32'h3c3cc439),
	.w7(32'hbbd36bfd),
	.w8(32'h3be2c74b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb1f1),
	.w1(32'h3acb3d2f),
	.w2(32'hba5c48b0),
	.w3(32'hbb63d3a1),
	.w4(32'h3bfa2a74),
	.w5(32'h3c0e8d56),
	.w6(32'h3b3a0174),
	.w7(32'hb8ffa5f1),
	.w8(32'h3b49196b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba543c2b),
	.w1(32'hbbbe2a6d),
	.w2(32'hbce1af77),
	.w3(32'h3b5ec25b),
	.w4(32'hbcb4c110),
	.w5(32'hbb185f72),
	.w6(32'hbbbf9209),
	.w7(32'hbc498c5a),
	.w8(32'hbc22c15c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca60c1f),
	.w1(32'h3ccd8ca1),
	.w2(32'h3c731577),
	.w3(32'h3cf9117a),
	.w4(32'h3c7a9bdd),
	.w5(32'h3b8a1aa6),
	.w6(32'h3ca073ad),
	.w7(32'h3c4b1ccd),
	.w8(32'hbb8157e5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4bc71),
	.w1(32'hbabf8af7),
	.w2(32'h3cabe643),
	.w3(32'hbc81d39d),
	.w4(32'h3b90cd95),
	.w5(32'hbc1f4ed7),
	.w6(32'hbcda4aef),
	.w7(32'h3c286e70),
	.w8(32'h3bff1126),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e56f9),
	.w1(32'h3c98bba9),
	.w2(32'h3a694d03),
	.w3(32'hbd07d8f7),
	.w4(32'h3d01e6d2),
	.w5(32'h3cc3d3f6),
	.w6(32'hbbfc40dd),
	.w7(32'h3cb4a696),
	.w8(32'h3c28f3f4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4df5d7),
	.w1(32'hbcd4f254),
	.w2(32'hbc9f3397),
	.w3(32'h3c337f51),
	.w4(32'h3bdf2b8c),
	.w5(32'h3c804599),
	.w6(32'hbbceaac2),
	.w7(32'h3b77a75b),
	.w8(32'hbb114941),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5c1cf),
	.w1(32'hbc8ba152),
	.w2(32'hbd12f2e5),
	.w3(32'h3cbdba81),
	.w4(32'hbbde23b4),
	.w5(32'h3c02fb98),
	.w6(32'hbb8530a2),
	.w7(32'hbcf498b0),
	.w8(32'h3bf73712),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55435d),
	.w1(32'h3c128059),
	.w2(32'h3d06dd6f),
	.w3(32'h3c7ba68f),
	.w4(32'hbc5559d1),
	.w5(32'hbd186540),
	.w6(32'h3cfbb22c),
	.w7(32'h3bc7b6b2),
	.w8(32'hbc6435fb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d038166),
	.w1(32'h3c7419ae),
	.w2(32'hbba0a8b8),
	.w3(32'hbd1da2a5),
	.w4(32'hbbda81f9),
	.w5(32'hbca91456),
	.w6(32'hbc0ce5bd),
	.w7(32'hbc8c4293),
	.w8(32'h3ba8879a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9ae47),
	.w1(32'h3cd71cf2),
	.w2(32'hbc0b93f8),
	.w3(32'hbc1540c2),
	.w4(32'hbbc66cc6),
	.w5(32'h3b17c402),
	.w6(32'h3cdc4b69),
	.w7(32'hb8a3c5bf),
	.w8(32'h3c6aabf7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb327468),
	.w1(32'h3b93d6e0),
	.w2(32'hb92f91a5),
	.w3(32'h3ba7d8cf),
	.w4(32'hbbd5464f),
	.w5(32'hbc560b6e),
	.w6(32'h3c9a4e89),
	.w7(32'hbcc61125),
	.w8(32'hbcc04e0e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f59ff),
	.w1(32'h3c1a9708),
	.w2(32'hbd1af787),
	.w3(32'hbbaf2c2b),
	.w4(32'h3d1390e2),
	.w5(32'h3d7a6ed4),
	.w6(32'h3bfcc830),
	.w7(32'h3c969614),
	.w8(32'h3cd11db7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3945b9),
	.w1(32'hbc9fe4fd),
	.w2(32'h3c99e5b5),
	.w3(32'h3d134ea9),
	.w4(32'h3ba6f61e),
	.w5(32'hbc250b06),
	.w6(32'hba1ce5e0),
	.w7(32'h3bec6dd1),
	.w8(32'hbb916f22),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08a8df),
	.w1(32'h3bd2ac5c),
	.w2(32'h3b1ec306),
	.w3(32'hbb56be14),
	.w4(32'h3ba2ab0d),
	.w5(32'h3b5555f7),
	.w6(32'hbc79759e),
	.w7(32'h3b82f1ca),
	.w8(32'h39b14ff1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc200b16),
	.w1(32'hbc3b5896),
	.w2(32'h3b8c8869),
	.w3(32'hbb357cf5),
	.w4(32'hbc97b913),
	.w5(32'hbcd0d1e0),
	.w6(32'hbbe1898c),
	.w7(32'hbc1abdc7),
	.w8(32'hbb611435),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc33876),
	.w1(32'h3cbe3bdc),
	.w2(32'hbb45ea65),
	.w3(32'h3c41cb12),
	.w4(32'h3c52dc02),
	.w5(32'h3c83f4d8),
	.w6(32'h3bed78a5),
	.w7(32'h3c5627ec),
	.w8(32'h3b77a8d1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc503218),
	.w1(32'hbc27ad5d),
	.w2(32'h3b69dd9c),
	.w3(32'h3bbc660e),
	.w4(32'h3af6e998),
	.w5(32'h3c5554f3),
	.w6(32'h3a19bd49),
	.w7(32'hbd23cb33),
	.w8(32'hbc4dbc5b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25778f),
	.w1(32'h3ca396ac),
	.w2(32'h3c1f97de),
	.w3(32'h3c859ee2),
	.w4(32'hbc813bbb),
	.w5(32'hbcd64080),
	.w6(32'h3cc8eee0),
	.w7(32'h3c47de36),
	.w8(32'h3c2a4e0e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25740b),
	.w1(32'h3cacb65a),
	.w2(32'hbccefb45),
	.w3(32'h39123534),
	.w4(32'hbcc80556),
	.w5(32'hbc6ee2b3),
	.w6(32'h3b97816f),
	.w7(32'hbc22683b),
	.w8(32'hbb4966fb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc956894),
	.w1(32'h3d076b92),
	.w2(32'hbbfe6b21),
	.w3(32'hba414ce9),
	.w4(32'hbd9606b1),
	.w5(32'hbd75e585),
	.w6(32'h3ca18a96),
	.w7(32'hbd516680),
	.w8(32'hbc68f2b4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d165240),
	.w1(32'h3da84dd8),
	.w2(32'h3d0deb82),
	.w3(32'hbca4726e),
	.w4(32'h3ba75df3),
	.w5(32'h3b55bceb),
	.w6(32'h3d26f00f),
	.w7(32'h3cbbf6df),
	.w8(32'h3c4ccc9d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8471a5),
	.w1(32'h3b8c9c2c),
	.w2(32'hbbf35fbe),
	.w3(32'hbd12e47e),
	.w4(32'h3c34e08b),
	.w5(32'h3c38ce88),
	.w6(32'hbccc7644),
	.w7(32'h3a6b28cf),
	.w8(32'hbc6257f0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1b42),
	.w1(32'hbc1599ca),
	.w2(32'h3c9c263a),
	.w3(32'h3c4016d8),
	.w4(32'hbbbd1e9b),
	.w5(32'h3b8bf7ba),
	.w6(32'h3b5d2616),
	.w7(32'h3c597b36),
	.w8(32'hbc6df75d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178dc2),
	.w1(32'h3c4946c8),
	.w2(32'h3aa3e3fb),
	.w3(32'h3b0350d8),
	.w4(32'h3c4265f2),
	.w5(32'h3c282210),
	.w6(32'h3a24787b),
	.w7(32'h3bb19564),
	.w8(32'h3b7322a4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a11b9),
	.w1(32'hbbf307ed),
	.w2(32'h3b9913b7),
	.w3(32'h3bc4b419),
	.w4(32'hbbedc7cf),
	.w5(32'hbb4088e8),
	.w6(32'h3ae41c02),
	.w7(32'hbcd3ab6e),
	.w8(32'hbbd3467c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41d441),
	.w1(32'h3bc5df59),
	.w2(32'h3ba07c17),
	.w3(32'hbc5653dc),
	.w4(32'hbcd9adaf),
	.w5(32'hbcadd661),
	.w6(32'h3c127e41),
	.w7(32'hbc456a32),
	.w8(32'hbbbc5b75),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5a056),
	.w1(32'h3cb9fecf),
	.w2(32'hbbac2e80),
	.w3(32'hbcd62cea),
	.w4(32'hbc60d2ec),
	.w5(32'hbba62e52),
	.w6(32'hb9c8c952),
	.w7(32'hbbc5c0ee),
	.w8(32'hb9f5b41f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb36ab9),
	.w1(32'hbbc6d1cc),
	.w2(32'h3ce2057d),
	.w3(32'h3aea53cf),
	.w4(32'h3be19873),
	.w5(32'hbb9277a2),
	.w6(32'hbb952639),
	.w7(32'hbae9b5c4),
	.w8(32'hbc28a225),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10e77b),
	.w1(32'h3beb211d),
	.w2(32'h3a30dcbc),
	.w3(32'hbd157715),
	.w4(32'h3ba7a306),
	.w5(32'h3b3ec817),
	.w6(32'hbcf6d268),
	.w7(32'h3b6635ca),
	.w8(32'hbaf04d1d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58ccc),
	.w1(32'hbc01ed71),
	.w2(32'hbb801994),
	.w3(32'h398a478d),
	.w4(32'hbc2e44ad),
	.w5(32'hbb675bf8),
	.w6(32'hbb097e60),
	.w7(32'hbb7f52c5),
	.w8(32'h3ca116a0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c519008),
	.w1(32'hbb6eff15),
	.w2(32'h3c02e510),
	.w3(32'h3c611ab8),
	.w4(32'hbc27903e),
	.w5(32'h3b8a98ae),
	.w6(32'h3c1a8a9e),
	.w7(32'hbb8e5059),
	.w8(32'h3bbfb197),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59f63d),
	.w1(32'hbb1fc0c7),
	.w2(32'h3bbaa42f),
	.w3(32'h3bfa5263),
	.w4(32'hbcc54df7),
	.w5(32'hbc83be81),
	.w6(32'hbc012f92),
	.w7(32'hbc8e8d5e),
	.w8(32'hbc486c17),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42b42e),
	.w1(32'h3c3e6c3e),
	.w2(32'h3c4cd46d),
	.w3(32'hbbbed42f),
	.w4(32'hbc56f878),
	.w5(32'hbc857349),
	.w6(32'hbbb69af2),
	.w7(32'hbc482342),
	.w8(32'h3a8107d7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c871eca),
	.w1(32'h3c572ad0),
	.w2(32'h3bcba1d0),
	.w3(32'h3bb2fc99),
	.w4(32'hb889af69),
	.w5(32'h3b751aa2),
	.w6(32'h3c023b7a),
	.w7(32'h388b84ed),
	.w8(32'h3aeb6e06),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule