module layer_10_featuremap_223(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911289),
	.w1(32'hbb85e5e7),
	.w2(32'h3b805f3c),
	.w3(32'hbacc6059),
	.w4(32'hbb2c1688),
	.w5(32'hbabdb804),
	.w6(32'h3c0ca5a7),
	.w7(32'h3c0dddc8),
	.w8(32'hbbf7a65b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d87b),
	.w1(32'hbbfd0da3),
	.w2(32'h3b117fa7),
	.w3(32'h3c61b4eb),
	.w4(32'h3bc5732b),
	.w5(32'hbaa94af3),
	.w6(32'h3c707746),
	.w7(32'hb9c0bf53),
	.w8(32'h3c3a1022),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ffcf3),
	.w1(32'hbbb4a5f0),
	.w2(32'hbd0044ef),
	.w3(32'h3b2b40df),
	.w4(32'hb98449c8),
	.w5(32'h3c9575e3),
	.w6(32'hbb23bc52),
	.w7(32'h3ac23d2f),
	.w8(32'hbc388048),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44dcab),
	.w1(32'hbbcdab9a),
	.w2(32'hbb4853e6),
	.w3(32'hbb7525fa),
	.w4(32'hbbdfd66d),
	.w5(32'h3bef9587),
	.w6(32'h3c24d17b),
	.w7(32'hbc54ad40),
	.w8(32'hbc363182),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ad962),
	.w1(32'h3b0507a8),
	.w2(32'hbbfb4bdc),
	.w3(32'h3b9cf5ea),
	.w4(32'hbbb123c7),
	.w5(32'hb9ee5271),
	.w6(32'hbc9b4219),
	.w7(32'h3b783da9),
	.w8(32'hbaaa3443),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc249c68),
	.w1(32'hbaedd81e),
	.w2(32'hbc1d89c9),
	.w3(32'hbb862aa3),
	.w4(32'h3a83ac00),
	.w5(32'hbcafcee2),
	.w6(32'hbb27a386),
	.w7(32'hbb1277ac),
	.w8(32'hbabab955),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789ec8),
	.w1(32'h3ba9b58f),
	.w2(32'hbc2dc04b),
	.w3(32'hbca1a27c),
	.w4(32'h3b985e79),
	.w5(32'hbacb2573),
	.w6(32'hbbc40663),
	.w7(32'hbca8deec),
	.w8(32'hbb40e100),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f1e89),
	.w1(32'hba2af8bd),
	.w2(32'hb9bde92e),
	.w3(32'hbbf4b959),
	.w4(32'hbb59d27b),
	.w5(32'hbac9b8b7),
	.w6(32'hbbf50876),
	.w7(32'hbc28318c),
	.w8(32'h3b0de6ca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4c09),
	.w1(32'hbc5e4393),
	.w2(32'hbc23a3e3),
	.w3(32'hbabf7e77),
	.w4(32'hbc0d82b3),
	.w5(32'hbb866c5b),
	.w6(32'hbc1178de),
	.w7(32'hbb74ce24),
	.w8(32'h3a810b42),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78cfc1),
	.w1(32'hb9bb0bd7),
	.w2(32'h3d25a732),
	.w3(32'h3be4bc02),
	.w4(32'hbc18d93a),
	.w5(32'hbbe96660),
	.w6(32'hbb53f41c),
	.w7(32'h3a6a176f),
	.w8(32'h3cc9a50c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3cd26),
	.w1(32'h3c8bbc6b),
	.w2(32'h3c5872bc),
	.w3(32'hbc07874a),
	.w4(32'hbbdefeb1),
	.w5(32'h3a6a92ae),
	.w6(32'h3a9b5c23),
	.w7(32'hbc1159c5),
	.w8(32'h3b5eeb47),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39969f8c),
	.w1(32'hbb8f4ba9),
	.w2(32'hbb904f7f),
	.w3(32'hbb53cf4e),
	.w4(32'hbb42f862),
	.w5(32'hb88b7f0c),
	.w6(32'hbbe72095),
	.w7(32'hb7dcba49),
	.w8(32'hbc2419d1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a7ec8),
	.w1(32'hbbe62bc0),
	.w2(32'hbaa6600b),
	.w3(32'hbb1a2149),
	.w4(32'hbc0ff384),
	.w5(32'h3cef47f6),
	.w6(32'hbb5f45ef),
	.w7(32'hbcacf6f8),
	.w8(32'hbb01c65d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e602),
	.w1(32'h3a89851b),
	.w2(32'hbd238f0b),
	.w3(32'hbbf3a6e2),
	.w4(32'h3b07c1c9),
	.w5(32'h3a2b9dd3),
	.w6(32'h3c4178db),
	.w7(32'h3ac201d2),
	.w8(32'hbb81c214),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914340),
	.w1(32'h3be297c5),
	.w2(32'hbbaedb9c),
	.w3(32'hbc02c0e5),
	.w4(32'h3bbfb8e9),
	.w5(32'h3c4712ba),
	.w6(32'h3c63dd2e),
	.w7(32'h3b14b922),
	.w8(32'hba990303),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878bd1),
	.w1(32'hbbe8afac),
	.w2(32'h3bd81df4),
	.w3(32'hba152f00),
	.w4(32'h3b89ee1e),
	.w5(32'hbb710933),
	.w6(32'hbab2a11d),
	.w7(32'hbaf88d5c),
	.w8(32'h3b2b0d49),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2caa),
	.w1(32'hba9881b6),
	.w2(32'h3b1b48cc),
	.w3(32'h3a6f802c),
	.w4(32'h38e365d0),
	.w5(32'hbc3ab925),
	.w6(32'h3a96e719),
	.w7(32'h3bc4a66b),
	.w8(32'hbbd06c5d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34f128),
	.w1(32'hbb89ea18),
	.w2(32'hbc4e69d6),
	.w3(32'h3bc7ab32),
	.w4(32'hbb1457ea),
	.w5(32'hb996bb24),
	.w6(32'h3bdca75f),
	.w7(32'h3b1e4be5),
	.w8(32'hbbedb2d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab7a58),
	.w1(32'hbb3b3099),
	.w2(32'hbb9a525d),
	.w3(32'h3c61bf4b),
	.w4(32'hbb1d9222),
	.w5(32'hbbe75be6),
	.w6(32'hbb87af0a),
	.w7(32'hbb028990),
	.w8(32'hbbcc1167),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0f58),
	.w1(32'hbc1b7b4f),
	.w2(32'hbb756918),
	.w3(32'h3b48bd49),
	.w4(32'hbbf3ab8c),
	.w5(32'h3be6f76e),
	.w6(32'hbc15c328),
	.w7(32'hbb57134b),
	.w8(32'hbb3a03d2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ceeaf4),
	.w1(32'hbbbb3252),
	.w2(32'hbb52eb33),
	.w3(32'hbb7adbdb),
	.w4(32'hbc2e2004),
	.w5(32'h3b471d9c),
	.w6(32'h3ac44392),
	.w7(32'hbc3677ca),
	.w8(32'h3a2e669a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97404b),
	.w1(32'hbbfc5247),
	.w2(32'hbbde59c9),
	.w3(32'h3abbc8bd),
	.w4(32'hbb35edf3),
	.w5(32'hbba792aa),
	.w6(32'h3b8207c3),
	.w7(32'h37c51df1),
	.w8(32'h3c6e0e73),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a8636),
	.w1(32'hba2cfb47),
	.w2(32'hbc388b86),
	.w3(32'hbc087cbc),
	.w4(32'h3c06ba14),
	.w5(32'hbb712400),
	.w6(32'h3abbea7e),
	.w7(32'hbbb4f8bd),
	.w8(32'h393e0b7a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fd8a4),
	.w1(32'hba47950b),
	.w2(32'hbb080475),
	.w3(32'hba4d451e),
	.w4(32'h3ac01ade),
	.w5(32'hbc8bf4ef),
	.w6(32'hbb0ea3dc),
	.w7(32'hbc51d6b5),
	.w8(32'h3c6e5fb7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7e91),
	.w1(32'hbb236966),
	.w2(32'h39d9bd57),
	.w3(32'h3b9d5c25),
	.w4(32'h3b44399d),
	.w5(32'h3cc7ab03),
	.w6(32'hbae52aa0),
	.w7(32'hbb962ab0),
	.w8(32'hbab35b03),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc344231),
	.w1(32'h3b66dac9),
	.w2(32'h3968bfd1),
	.w3(32'h3c714816),
	.w4(32'hbc8ac7f9),
	.w5(32'hbb8df9a5),
	.w6(32'hbb91cb05),
	.w7(32'h39ed21cf),
	.w8(32'h3bee3251),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20c2a6),
	.w1(32'hbba000c3),
	.w2(32'hb9330186),
	.w3(32'h3c779205),
	.w4(32'h3aa74123),
	.w5(32'hbb768565),
	.w6(32'h3ca7dfdf),
	.w7(32'hbbbbe3ae),
	.w8(32'h3ac10a71),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe579c0),
	.w1(32'hbc1e7ddb),
	.w2(32'h3a89eeab),
	.w3(32'hbba6cce8),
	.w4(32'hbc7ffe4e),
	.w5(32'hbb4ef538),
	.w6(32'hb9895e71),
	.w7(32'h3c71c1ec),
	.w8(32'hba970673),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa6e53),
	.w1(32'h3a0c52c2),
	.w2(32'hbc9168e5),
	.w3(32'hbb0e3317),
	.w4(32'h3a024b99),
	.w5(32'h3a76c901),
	.w6(32'h3b9d14a8),
	.w7(32'h3aba92e5),
	.w8(32'h3bb13756),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb2225),
	.w1(32'hbb9e6bf2),
	.w2(32'h3baef686),
	.w3(32'hba038db6),
	.w4(32'h3cbff0d5),
	.w5(32'hbc30533f),
	.w6(32'h3bf2894c),
	.w7(32'h3b6c3f76),
	.w8(32'hbb39832a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5845e),
	.w1(32'hbb16b25b),
	.w2(32'hbb2eb9d1),
	.w3(32'hbc73712e),
	.w4(32'h3b819d7c),
	.w5(32'h3b9af7cb),
	.w6(32'h3b0beb61),
	.w7(32'hba3004e6),
	.w8(32'hbc3eb31d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc92cb3),
	.w1(32'hbbb49d06),
	.w2(32'hbb47f043),
	.w3(32'h3b566789),
	.w4(32'hbbabf3da),
	.w5(32'hba638ebc),
	.w6(32'hbbc67e01),
	.w7(32'h3a70fce7),
	.w8(32'hbcad66d1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d53c2a),
	.w1(32'hbb95b217),
	.w2(32'hbb087ac9),
	.w3(32'hbb431d09),
	.w4(32'h3be8effc),
	.w5(32'hba1e4cb4),
	.w6(32'hbba1cb8f),
	.w7(32'hbc25068e),
	.w8(32'hbb2127c1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3e88),
	.w1(32'hbd08e17d),
	.w2(32'h3c3b7fef),
	.w3(32'hbb899001),
	.w4(32'h3b3f9a1d),
	.w5(32'hbb24ddfa),
	.w6(32'hba4e6391),
	.w7(32'hbb128d49),
	.w8(32'hb9dbf967),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae15964),
	.w1(32'hbb9d0eb1),
	.w2(32'hbb9f3034),
	.w3(32'h3b0886a0),
	.w4(32'hbb9c90e9),
	.w5(32'hba8803c6),
	.w6(32'hbbe9bcc1),
	.w7(32'h3aaa344d),
	.w8(32'h3cdb0c2a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea04a8),
	.w1(32'hbac2da51),
	.w2(32'hbbe9f47f),
	.w3(32'hbba0ead0),
	.w4(32'hbb5fee3b),
	.w5(32'hbb59717f),
	.w6(32'hbb81861a),
	.w7(32'hbb023494),
	.w8(32'h39eeed72),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1426),
	.w1(32'hbc3a9305),
	.w2(32'h3c13d7ed),
	.w3(32'h3ac95bcd),
	.w4(32'hbc582293),
	.w5(32'hba93cb98),
	.w6(32'h3a63fb12),
	.w7(32'h3a2b65c4),
	.w8(32'hba4cacb6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985286c),
	.w1(32'h3a899cc6),
	.w2(32'h3b0e0000),
	.w3(32'hbbea08e5),
	.w4(32'hbd138e4e),
	.w5(32'h39a6ebf8),
	.w6(32'hbbfd0a02),
	.w7(32'h3be6d044),
	.w8(32'h3b1a3b99),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda55f5),
	.w1(32'h3b0045f3),
	.w2(32'h3c250f22),
	.w3(32'h3c4a002f),
	.w4(32'hbbef8d9b),
	.w5(32'hbbabceab),
	.w6(32'hbb1aff59),
	.w7(32'hbb1c5dd0),
	.w8(32'hbc109554),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd35db8),
	.w1(32'hbbbde528),
	.w2(32'h3ab61576),
	.w3(32'h3c120370),
	.w4(32'h3b9dbe1f),
	.w5(32'hbb1511c9),
	.w6(32'hbcf90a74),
	.w7(32'h3b90a257),
	.w8(32'hbc70498a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ec99d6),
	.w1(32'hbafb0b5a),
	.w2(32'h3ba92159),
	.w3(32'hbcae8638),
	.w4(32'hbbd3edc1),
	.w5(32'hbb610b8e),
	.w6(32'hba348fe0),
	.w7(32'h3a49089a),
	.w8(32'hba85556a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf803f),
	.w1(32'hbadab842),
	.w2(32'h3c236a89),
	.w3(32'hbbc23e67),
	.w4(32'hbca2aa15),
	.w5(32'hbb32c4d3),
	.w6(32'h3afc1d0b),
	.w7(32'h3c00b57e),
	.w8(32'h3d3575cc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9047a9),
	.w1(32'h3b839ae9),
	.w2(32'hbb58fd33),
	.w3(32'hbc11086f),
	.w4(32'h3bb0035f),
	.w5(32'hb8d82500),
	.w6(32'h3b8a31ca),
	.w7(32'h3a32e6e7),
	.w8(32'h3bff7172),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bed84),
	.w1(32'h39d9ba53),
	.w2(32'hbb778de7),
	.w3(32'hbb02a711),
	.w4(32'hbaab6692),
	.w5(32'h3af3f778),
	.w6(32'hbbdfc93a),
	.w7(32'h3b13af94),
	.w8(32'hbb29e071),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0323f),
	.w1(32'hbce05769),
	.w2(32'hbb515277),
	.w3(32'h3a35adfe),
	.w4(32'hbbbe1ee5),
	.w5(32'hb92e46bf),
	.w6(32'h3bbaf1f2),
	.w7(32'h3b55ef09),
	.w8(32'h374db38c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba851409),
	.w1(32'hbba60cf4),
	.w2(32'hbb575f88),
	.w3(32'h3a0aca20),
	.w4(32'hba541193),
	.w5(32'h3c004928),
	.w6(32'hbbaff63f),
	.w7(32'hbbe6ce5c),
	.w8(32'hb8c806e6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18a4f9),
	.w1(32'hbb4b1015),
	.w2(32'h3bf50d13),
	.w3(32'hbc296d31),
	.w4(32'hbb9bfe46),
	.w5(32'hbc60c6ca),
	.w6(32'h39b2fb65),
	.w7(32'h3b941cb1),
	.w8(32'h3a89988a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe101e8),
	.w1(32'h3b351cd2),
	.w2(32'hbb7c66a3),
	.w3(32'hbbbf4937),
	.w4(32'hbbe0c6d8),
	.w5(32'hbbdb683f),
	.w6(32'hbc12c9c5),
	.w7(32'hbaca85d4),
	.w8(32'h3c0368d7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a062b98),
	.w1(32'h3bf8e432),
	.w2(32'h3b910083),
	.w3(32'hbbc1576a),
	.w4(32'h393de937),
	.w5(32'hbb709f4c),
	.w6(32'h3aac4afb),
	.w7(32'hb892eca6),
	.w8(32'h3a51914c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08250),
	.w1(32'h3c56987a),
	.w2(32'hbaea6868),
	.w3(32'h3c30c2a8),
	.w4(32'h3c90eddb),
	.w5(32'hbc0b89a8),
	.w6(32'h3b7cba8e),
	.w7(32'h398593b1),
	.w8(32'hbb919ea7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b2129),
	.w1(32'h3a47f8d0),
	.w2(32'h39c1bb16),
	.w3(32'h3b583682),
	.w4(32'hba903351),
	.w5(32'hb8c14691),
	.w6(32'hbaba283c),
	.w7(32'hbbb8f84a),
	.w8(32'h3a813803),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8234369),
	.w1(32'h3cab0d02),
	.w2(32'h3b7db5a6),
	.w3(32'hbcde7d44),
	.w4(32'hbcbd4abe),
	.w5(32'hbb0521b5),
	.w6(32'hbac370bd),
	.w7(32'h3a47eca6),
	.w8(32'hbb87498d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb42f09),
	.w1(32'hbbfd18b2),
	.w2(32'hbb43a494),
	.w3(32'hb86311c8),
	.w4(32'hbb731b34),
	.w5(32'hbb33401c),
	.w6(32'h3b5afa8f),
	.w7(32'h3a84154f),
	.w8(32'h3d29e896),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf9811),
	.w1(32'h3afad807),
	.w2(32'h3af69da8),
	.w3(32'h3a42b08e),
	.w4(32'hbb84bb27),
	.w5(32'hbc5d567a),
	.w6(32'h3aefcfcf),
	.w7(32'hbc0e806e),
	.w8(32'hbc739747),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977242),
	.w1(32'hba9785b0),
	.w2(32'hbb3148a6),
	.w3(32'h3bcc7e64),
	.w4(32'hbaed1e69),
	.w5(32'h3b51cce2),
	.w6(32'hbaee0c05),
	.w7(32'h38730649),
	.w8(32'hbb57afac),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65479c),
	.w1(32'hbc8da6b1),
	.w2(32'hbc919793),
	.w3(32'hbc9226f3),
	.w4(32'hbc2159f7),
	.w5(32'hbbe3e9d4),
	.w6(32'hbacc0a1f),
	.w7(32'h3a7bac14),
	.w8(32'h3b2ef641),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73dfa1),
	.w1(32'h3a83c083),
	.w2(32'hbc363edd),
	.w3(32'hbb02bde8),
	.w4(32'hbc6aeac9),
	.w5(32'h3b2bb920),
	.w6(32'hbc1e2e07),
	.w7(32'h3bbeb76e),
	.w8(32'hbb63c391),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a1e20),
	.w1(32'hbbeab892),
	.w2(32'h3d0bd647),
	.w3(32'h3a353cb3),
	.w4(32'hbb9eb79a),
	.w5(32'hbc4989c1),
	.w6(32'h3a80c972),
	.w7(32'hbc3f0ab9),
	.w8(32'hbabe83f2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c31ee),
	.w1(32'h3b997dec),
	.w2(32'hbc0b32fb),
	.w3(32'hbbfdac9a),
	.w4(32'hbc73f2a3),
	.w5(32'hbc092961),
	.w6(32'hbb8137bf),
	.w7(32'h3b607e6b),
	.w8(32'hbc2a13b1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba20c4),
	.w1(32'h3c99bdf0),
	.w2(32'hbba4958f),
	.w3(32'h3b709aec),
	.w4(32'hbc2e1dd3),
	.w5(32'hbc7bdbcf),
	.w6(32'hbc31e36b),
	.w7(32'hbc941127),
	.w8(32'hbc1256aa),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c4fa6),
	.w1(32'hbc09c620),
	.w2(32'hbc33baab),
	.w3(32'hbc269833),
	.w4(32'hbc3f4c4f),
	.w5(32'hbb9a4458),
	.w6(32'hbb0b0488),
	.w7(32'hbc01c4b8),
	.w8(32'hbb63c18f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4df31d),
	.w1(32'hba8563a8),
	.w2(32'h3bc297f7),
	.w3(32'hbb946cb6),
	.w4(32'hbb94705e),
	.w5(32'h3b5b22d1),
	.w6(32'hbc59d7f8),
	.w7(32'hbbc91e9f),
	.w8(32'hbc721e80),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc946f6b),
	.w1(32'hbb4c43ca),
	.w2(32'h3c0b64e4),
	.w3(32'hba6ab634),
	.w4(32'hbb704149),
	.w5(32'hbba0fcd0),
	.w6(32'h3bb258e3),
	.w7(32'hbc40b4a1),
	.w8(32'hbab6c401),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a8b7e),
	.w1(32'h3c1a8da6),
	.w2(32'h3bd81e5b),
	.w3(32'h3b255bb7),
	.w4(32'hba2cc79c),
	.w5(32'h3c339cb8),
	.w6(32'hbcd29460),
	.w7(32'hbc9b0143),
	.w8(32'hbba24347),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a7f9a),
	.w1(32'h3b433bcd),
	.w2(32'h3aa00175),
	.w3(32'hbb99905f),
	.w4(32'hbc0be863),
	.w5(32'hbc17ec7b),
	.w6(32'hbba2e912),
	.w7(32'hbb63e351),
	.w8(32'hba81af5c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9362f4),
	.w1(32'hbc8e864f),
	.w2(32'hbb3196b0),
	.w3(32'hbc006a30),
	.w4(32'hbc3873cc),
	.w5(32'hbb65dea9),
	.w6(32'h3c9376c3),
	.w7(32'h3b293abc),
	.w8(32'h3a04e8b0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e48d3),
	.w1(32'hbb2b3e91),
	.w2(32'hbcb270a2),
	.w3(32'hbb598e15),
	.w4(32'hbb0eed07),
	.w5(32'hbc147c40),
	.w6(32'hb94320f3),
	.w7(32'hbc2e2baf),
	.w8(32'h3c018f45),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98384e4),
	.w1(32'hbb5354fb),
	.w2(32'h3b98a645),
	.w3(32'h3b811867),
	.w4(32'hbbd84e1a),
	.w5(32'hbbd482b5),
	.w6(32'hba430953),
	.w7(32'hbc0a563e),
	.w8(32'hbb0442b9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57be57),
	.w1(32'h3c66763c),
	.w2(32'h393311f9),
	.w3(32'hbb60c163),
	.w4(32'hb92522b3),
	.w5(32'h3b95b61b),
	.w6(32'hbb9fcf50),
	.w7(32'h3abe7d45),
	.w8(32'hbcc2c911),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83b265),
	.w1(32'hbbf5f00e),
	.w2(32'h3a87be8c),
	.w3(32'h3b8a32ff),
	.w4(32'hbc747a74),
	.w5(32'h3b944ee7),
	.w6(32'hbc83a2a6),
	.w7(32'hbc2fd5f7),
	.w8(32'hba60f93d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6756a),
	.w1(32'h3b8e3f8f),
	.w2(32'h3aafde13),
	.w3(32'h3989b5fb),
	.w4(32'hbc0bc826),
	.w5(32'hbc43d78e),
	.w6(32'h3bb6cd62),
	.w7(32'hbc6fca37),
	.w8(32'h39abcd7c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c0028),
	.w1(32'hbbe4b7e1),
	.w2(32'h3be41a64),
	.w3(32'h3bc161c4),
	.w4(32'hbbca8be3),
	.w5(32'hbad7480e),
	.w6(32'hbc9812c1),
	.w7(32'hbc158530),
	.w8(32'hbc7d6bbf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e85c2),
	.w1(32'hbbc7d8ab),
	.w2(32'hbc2376bd),
	.w3(32'hbad5f484),
	.w4(32'hbb9b36d7),
	.w5(32'hbb86b0b2),
	.w6(32'hbc366381),
	.w7(32'h3a64f16b),
	.w8(32'hbbc91512),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b626992),
	.w1(32'h377af9a4),
	.w2(32'hbc427780),
	.w3(32'hbc667b8e),
	.w4(32'hbc0aa22c),
	.w5(32'hbbb8250f),
	.w6(32'h3906c592),
	.w7(32'hbc1aebef),
	.w8(32'hbc75d788),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26e045),
	.w1(32'hbb560b50),
	.w2(32'hb8bb442b),
	.w3(32'h3bdef13e),
	.w4(32'h3c1a20e3),
	.w5(32'hbb8a76d7),
	.w6(32'hbb201f87),
	.w7(32'hbbfdd0a4),
	.w8(32'h3bb1f972),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb610d4a),
	.w1(32'hbc1322d1),
	.w2(32'hbb5b3c5b),
	.w3(32'hbac84543),
	.w4(32'hbbbd1551),
	.w5(32'hbc54274e),
	.w6(32'hbb816074),
	.w7(32'hbbad0bde),
	.w8(32'hbb4103b0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc370224),
	.w1(32'hbb8f0a0c),
	.w2(32'hbb28678d),
	.w3(32'hbbcdc847),
	.w4(32'h3bd2db75),
	.w5(32'hbc6259f8),
	.w6(32'hbc50cc71),
	.w7(32'h3bc9ccc6),
	.w8(32'hbab3e583),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c3a0),
	.w1(32'hbba2eca1),
	.w2(32'hbc6f29f5),
	.w3(32'hbbbb5e5c),
	.w4(32'hbbc94ccd),
	.w5(32'hbc508f45),
	.w6(32'hbc2fb0c6),
	.w7(32'h3c0d0914),
	.w8(32'h3c7fcc50),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034285),
	.w1(32'hba8b32d9),
	.w2(32'hbab79ab6),
	.w3(32'hbabf58d4),
	.w4(32'hb91b735b),
	.w5(32'hbbcf35cf),
	.w6(32'hbc516b0d),
	.w7(32'hbb2c46f0),
	.w8(32'hbbfdc9c7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb7a9),
	.w1(32'hbbffacc1),
	.w2(32'hbc94d58e),
	.w3(32'h3af6a0c5),
	.w4(32'hbc42e9cb),
	.w5(32'hbb72fc81),
	.w6(32'h3945d119),
	.w7(32'hbbcf0c7d),
	.w8(32'h3ab9743a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb062da),
	.w1(32'hbb20201d),
	.w2(32'h388c30d1),
	.w3(32'hbb9780a9),
	.w4(32'h3bea2e9e),
	.w5(32'hbc3acfb0),
	.w6(32'hbba7fbe8),
	.w7(32'hbb1f970c),
	.w8(32'h399593ab),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d2af6),
	.w1(32'hbbc27721),
	.w2(32'hbc3a0f58),
	.w3(32'hbc38aedc),
	.w4(32'hbc59f3d7),
	.w5(32'h3b2afb93),
	.w6(32'hbb88afa5),
	.w7(32'hbb4a2cc7),
	.w8(32'hbb806a5e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31f0f2),
	.w1(32'hbad0414d),
	.w2(32'hbc143977),
	.w3(32'h3b59ce83),
	.w4(32'hbb302d7f),
	.w5(32'hbc749349),
	.w6(32'hbbcdab78),
	.w7(32'hbac106a8),
	.w8(32'hbbe3d173),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d0900),
	.w1(32'hbc119e24),
	.w2(32'hbae5e793),
	.w3(32'h3b0d0436),
	.w4(32'hbb6e912a),
	.w5(32'hbb05a654),
	.w6(32'hba307889),
	.w7(32'hbb46796f),
	.w8(32'h3ac066e1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55aa20),
	.w1(32'h3c381d84),
	.w2(32'hbb9efa81),
	.w3(32'h3ca377c0),
	.w4(32'hbb97d6bb),
	.w5(32'hbb5b4e8c),
	.w6(32'hbb02c464),
	.w7(32'hbbcd2919),
	.w8(32'h3c2412fd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b690260),
	.w1(32'hbb41fd2d),
	.w2(32'hbc92096f),
	.w3(32'hbb97f627),
	.w4(32'hba1763b4),
	.w5(32'hbbfe2089),
	.w6(32'hbc346307),
	.w7(32'hbbb6724c),
	.w8(32'h3b2cf37d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b7523),
	.w1(32'hbbdd6a9f),
	.w2(32'hbc6d429e),
	.w3(32'h3baf2e2f),
	.w4(32'hba61155e),
	.w5(32'hbbb69d97),
	.w6(32'hbafd6a75),
	.w7(32'hbad1325b),
	.w8(32'hbc781959),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe9c75),
	.w1(32'h3c89b972),
	.w2(32'h3bd88d63),
	.w3(32'h3b884c97),
	.w4(32'h3a6770b6),
	.w5(32'h3b282f90),
	.w6(32'hba2ebc03),
	.w7(32'hbba643b7),
	.w8(32'hbbcfcdcb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1a9a6),
	.w1(32'h3a043637),
	.w2(32'hbb0b7eb8),
	.w3(32'h3b1b39f4),
	.w4(32'hbaede3d0),
	.w5(32'hbb8caf2f),
	.w6(32'hbba8bd3d),
	.w7(32'hbc1cfe46),
	.w8(32'hbc547001),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb501798),
	.w1(32'h3c1fdc70),
	.w2(32'h3b718cad),
	.w3(32'hbc667a30),
	.w4(32'hbc55c991),
	.w5(32'h3cbd5f03),
	.w6(32'hbc48b70a),
	.w7(32'h3c6655d6),
	.w8(32'hbbc988cd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c044f06),
	.w1(32'h3badb43d),
	.w2(32'hbbca89cb),
	.w3(32'h391c3b4b),
	.w4(32'h3c919989),
	.w5(32'hba6f4384),
	.w6(32'hbc09092f),
	.w7(32'h3a9a9321),
	.w8(32'hbb030b9a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9582d4),
	.w1(32'hb9603cfc),
	.w2(32'h3bc48533),
	.w3(32'hbb09badd),
	.w4(32'h3c2dc3ec),
	.w5(32'hbbc9dfa5),
	.w6(32'hbbad2f7d),
	.w7(32'hb986f38d),
	.w8(32'hbc08273f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98db650),
	.w1(32'hbae8e90d),
	.w2(32'h3bf7b46a),
	.w3(32'hb9ac8953),
	.w4(32'hbb21bfab),
	.w5(32'hbbba923e),
	.w6(32'hbc4d700f),
	.w7(32'hbcad3d3e),
	.w8(32'hbc3e7c30),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3597a1),
	.w1(32'hbb823b0b),
	.w2(32'h39445801),
	.w3(32'h3b956fd8),
	.w4(32'h3c26c80e),
	.w5(32'hbc723194),
	.w6(32'hbcb82e01),
	.w7(32'hbb869bf6),
	.w8(32'h3bc628ce),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d84d8),
	.w1(32'h3aa51c06),
	.w2(32'hb9b20edd),
	.w3(32'hbb4869da),
	.w4(32'h3a941757),
	.w5(32'hbc0e16de),
	.w6(32'h385120a3),
	.w7(32'h3b834506),
	.w8(32'hbbb267b0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06cdcb),
	.w1(32'hbc689fc8),
	.w2(32'hbbac779a),
	.w3(32'h3b678c01),
	.w4(32'h3cc1be9c),
	.w5(32'h3a402504),
	.w6(32'h3caf1297),
	.w7(32'h3b3c0dec),
	.w8(32'hbb7d3040),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2464bf),
	.w1(32'hbb81961c),
	.w2(32'h3b20048c),
	.w3(32'hbb9f04de),
	.w4(32'hbb3cf39c),
	.w5(32'hbc24f09e),
	.w6(32'h3a9df49c),
	.w7(32'hbab5d317),
	.w8(32'hba41d608),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8946ec),
	.w1(32'hbc6123ae),
	.w2(32'h3c026f56),
	.w3(32'h3b672046),
	.w4(32'h3baa8fa5),
	.w5(32'h3c3fdd53),
	.w6(32'hbcfdff47),
	.w7(32'hbc5622f0),
	.w8(32'hbad8a6ec),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d474f),
	.w1(32'hbb28f6ab),
	.w2(32'h3bf82ac4),
	.w3(32'hbc3ac100),
	.w4(32'hbb0c91b4),
	.w5(32'h3c1631c4),
	.w6(32'h3b36c621),
	.w7(32'h3a684abd),
	.w8(32'h3ad9d186),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9854),
	.w1(32'hbbe32f23),
	.w2(32'hbc20758b),
	.w3(32'hbba203b5),
	.w4(32'hbc5f955c),
	.w5(32'h3add8b38),
	.w6(32'h3b09e6f6),
	.w7(32'h3b5145cd),
	.w8(32'h3be7a0ac),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cef82ed),
	.w1(32'hbc424290),
	.w2(32'h3c2c5c7c),
	.w3(32'hba441761),
	.w4(32'hbb51f8c5),
	.w5(32'h395a4975),
	.w6(32'h3b67f72d),
	.w7(32'hbb77fd4b),
	.w8(32'h3c35ea32),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1317e6),
	.w1(32'hbb63de59),
	.w2(32'hba741950),
	.w3(32'h3b08932e),
	.w4(32'hbb1b916c),
	.w5(32'hba92b650),
	.w6(32'hbbfadabf),
	.w7(32'h3c5936cb),
	.w8(32'hbae57026),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db006),
	.w1(32'h3bcb7c85),
	.w2(32'h3c41e4d9),
	.w3(32'h3b0fbc6d),
	.w4(32'hb99cc465),
	.w5(32'hbc017f06),
	.w6(32'hbaf9f4d2),
	.w7(32'hbbd08712),
	.w8(32'hbbd03371),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eed9d),
	.w1(32'h3bbe9ccb),
	.w2(32'hbc195b8b),
	.w3(32'h3ae8fce1),
	.w4(32'hbc6a39c1),
	.w5(32'h3b2de1f6),
	.w6(32'hbb856a09),
	.w7(32'hbbf67467),
	.w8(32'h3a5f0165),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d4400),
	.w1(32'h3ba11714),
	.w2(32'hbb56f8a4),
	.w3(32'h3c5cf58c),
	.w4(32'hba56e4c8),
	.w5(32'h3bd5c0ab),
	.w6(32'h3b40356a),
	.w7(32'h3c120353),
	.w8(32'h38ab8a1c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb2d88),
	.w1(32'hbc2dd2a3),
	.w2(32'h38ee6f16),
	.w3(32'h3a3bf7df),
	.w4(32'h3c1402ed),
	.w5(32'h3b48be5d),
	.w6(32'hbb8e61b8),
	.w7(32'hba0db90c),
	.w8(32'hbb06bab2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a231cff),
	.w1(32'hbbf4b158),
	.w2(32'h3bd3b954),
	.w3(32'hbc0a406f),
	.w4(32'h3a9d77d9),
	.w5(32'h3c2d526b),
	.w6(32'h3bfd622c),
	.w7(32'hbbddea6b),
	.w8(32'h387fee20),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b975406),
	.w1(32'h3c5cd855),
	.w2(32'h389cad64),
	.w3(32'hba264a75),
	.w4(32'hb92abbe4),
	.w5(32'h3b3e9054),
	.w6(32'hbc1ef5c3),
	.w7(32'h3a23448b),
	.w8(32'h3c4dfb3c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd66e8),
	.w1(32'h3bb51e3c),
	.w2(32'h3b9c7c13),
	.w3(32'hbc87e7b1),
	.w4(32'hbc8021c3),
	.w5(32'h3c63f881),
	.w6(32'hba3a9948),
	.w7(32'hba21b93b),
	.w8(32'h3c84fc35),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf16aed),
	.w1(32'h3c4df349),
	.w2(32'hbb2de923),
	.w3(32'hbc1ec16b),
	.w4(32'hbc181eec),
	.w5(32'hbb6aa836),
	.w6(32'h3bd93f52),
	.w7(32'hbc3ffde9),
	.w8(32'hbb368f6b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52eec7),
	.w1(32'h3be31240),
	.w2(32'hbbda554b),
	.w3(32'h3a94ad64),
	.w4(32'hbc5ef033),
	.w5(32'hbc54f77d),
	.w6(32'hbc14fc95),
	.w7(32'h3a4a8fe8),
	.w8(32'h3bcbb324),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99dab0),
	.w1(32'hbd03c59c),
	.w2(32'hbc2dddcf),
	.w3(32'hbbe7d1fb),
	.w4(32'hbc7bf426),
	.w5(32'h3b9ac9e1),
	.w6(32'h3c6a3a08),
	.w7(32'h3c08154b),
	.w8(32'hbb8159fc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5196),
	.w1(32'hba71b2de),
	.w2(32'h3bdbf555),
	.w3(32'h3afa43c0),
	.w4(32'hbb43cdb1),
	.w5(32'hbb56174f),
	.w6(32'h3ba36e61),
	.w7(32'hbbc6392d),
	.w8(32'h3b7220a2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d3592),
	.w1(32'hbc6825db),
	.w2(32'h3c6ea46f),
	.w3(32'h3c3916d5),
	.w4(32'h3bbc0af2),
	.w5(32'h3b5d001a),
	.w6(32'hbb7ed306),
	.w7(32'h3c2d8ec1),
	.w8(32'hbb380810),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c421930),
	.w1(32'h3b3b28ec),
	.w2(32'hbc11693c),
	.w3(32'hbba29ba1),
	.w4(32'hbc00f110),
	.w5(32'h3c24e50f),
	.w6(32'h3b051a0b),
	.w7(32'hbb962512),
	.w8(32'h3c7eded4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3030ca),
	.w1(32'h3c90e5ef),
	.w2(32'hbc01f5a8),
	.w3(32'hba99345e),
	.w4(32'h3bd0b544),
	.w5(32'hbc684a93),
	.w6(32'h3c432075),
	.w7(32'hbafeab14),
	.w8(32'h3c8db1a2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851d35),
	.w1(32'hbb5c3206),
	.w2(32'h3b76c916),
	.w3(32'hbc756e92),
	.w4(32'hbc90df4e),
	.w5(32'h3d20976a),
	.w6(32'h3c119227),
	.w7(32'hbbe168ff),
	.w8(32'h3bc64073),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6306),
	.w1(32'h3c1ad282),
	.w2(32'hbbf5d6d9),
	.w3(32'hb98c14b0),
	.w4(32'hbc69e850),
	.w5(32'hbbec6a02),
	.w6(32'hbc558d59),
	.w7(32'h381531b8),
	.w8(32'hbb58ef3d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a43ae),
	.w1(32'hba15e6cd),
	.w2(32'h3c0faeff),
	.w3(32'hbc7eb446),
	.w4(32'hbb870eec),
	.w5(32'hbbd55e18),
	.w6(32'h3c74dba0),
	.w7(32'h3aa4c3e1),
	.w8(32'hbc60c7b6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fdc45),
	.w1(32'hbb2c9431),
	.w2(32'h3cccb391),
	.w3(32'hbbd0403a),
	.w4(32'hbb244097),
	.w5(32'h3b1e5e82),
	.w6(32'h3a4b0870),
	.w7(32'h3c365456),
	.w8(32'hbc0d9627),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a5020),
	.w1(32'h3c0997a6),
	.w2(32'hb9fd9dd0),
	.w3(32'h3d39ada2),
	.w4(32'h3c985318),
	.w5(32'hbb891a39),
	.w6(32'hbc4cc52b),
	.w7(32'h3b504524),
	.w8(32'h3c3374b8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7186e9),
	.w1(32'hbbabe0ce),
	.w2(32'hbca57447),
	.w3(32'h3c5c91b1),
	.w4(32'hbb50c24e),
	.w5(32'h3bd1df1f),
	.w6(32'hbbb0c5e1),
	.w7(32'h3aabe68a),
	.w8(32'hb8aa6df3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376d10),
	.w1(32'h3ad3bfc1),
	.w2(32'h3ab26a80),
	.w3(32'h3b9e8c04),
	.w4(32'hbb1247c3),
	.w5(32'h3c8620c7),
	.w6(32'h3c8454c3),
	.w7(32'hbabfcf37),
	.w8(32'h3c0ffded),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839b32),
	.w1(32'h3c1a7f7c),
	.w2(32'h3cb6e3da),
	.w3(32'hb9a5c2aa),
	.w4(32'h3cb7c40a),
	.w5(32'hbb47cf11),
	.w6(32'hbb8a0665),
	.w7(32'h3c6cbd4c),
	.w8(32'h3cb64d59),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cfd4b),
	.w1(32'hbb47c827),
	.w2(32'h3c818c62),
	.w3(32'h3c1cd60c),
	.w4(32'hbbf24c72),
	.w5(32'hbc3bed7e),
	.w6(32'h3be34ee2),
	.w7(32'h3b7a1b09),
	.w8(32'hbbbd3435),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be08665),
	.w1(32'hb73c95cd),
	.w2(32'h3b8b85be),
	.w3(32'h3ae9556a),
	.w4(32'h3c07f202),
	.w5(32'hbc998a3a),
	.w6(32'hbb8c024c),
	.w7(32'hba0af4c9),
	.w8(32'h3bb27f54),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bd9bc),
	.w1(32'hbc640f79),
	.w2(32'h3c56ada0),
	.w3(32'hbc4ef8ca),
	.w4(32'hbc5489a8),
	.w5(32'h3bda0055),
	.w6(32'hbbae48d0),
	.w7(32'hbcac09f7),
	.w8(32'hbc168b8d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e7a25),
	.w1(32'h3c16416c),
	.w2(32'h3b11e247),
	.w3(32'hbbb8b37c),
	.w4(32'h3b6a4ed9),
	.w5(32'h3bc66b95),
	.w6(32'hbc17d7a8),
	.w7(32'h3c3bc803),
	.w8(32'hbc2e1383),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c492634),
	.w1(32'hbbeda7bf),
	.w2(32'hbbb43d9f),
	.w3(32'h3bfc8f35),
	.w4(32'h3baf785a),
	.w5(32'hb9b7fc7e),
	.w6(32'h3b035f2a),
	.w7(32'h3bfda6a0),
	.w8(32'hbaf523bb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49e892),
	.w1(32'hbaef1f30),
	.w2(32'h3ca340a4),
	.w3(32'hbacbd289),
	.w4(32'h3bba704e),
	.w5(32'h3bc97145),
	.w6(32'h3b2860fa),
	.w7(32'hbb955e2d),
	.w8(32'h3c9e867d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1b81b),
	.w1(32'hbb8aadb3),
	.w2(32'hbb51b7d7),
	.w3(32'h3bfaa12f),
	.w4(32'hbb233cc0),
	.w5(32'hbc164192),
	.w6(32'h383cab54),
	.w7(32'hba92b652),
	.w8(32'h3bff4ef5),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e9ae5),
	.w1(32'h3c171957),
	.w2(32'hbb7bd9f7),
	.w3(32'h3cadb481),
	.w4(32'h3b633a86),
	.w5(32'h3cb78da3),
	.w6(32'h3aba351f),
	.w7(32'hba58d99d),
	.w8(32'h3c5c2054),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a0bb2),
	.w1(32'h3a71eadf),
	.w2(32'hbc4929fe),
	.w3(32'h3c5264df),
	.w4(32'h396f3e24),
	.w5(32'h3c5f329c),
	.w6(32'h3be03bcd),
	.w7(32'h3b6f81f2),
	.w8(32'h3c00f24e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27764c),
	.w1(32'h3b1c5916),
	.w2(32'h3b3d5d34),
	.w3(32'h3bb6d0d0),
	.w4(32'h3a903ff3),
	.w5(32'h3c8e4de4),
	.w6(32'h3a1fd746),
	.w7(32'h3bf088d0),
	.w8(32'hbc0daccc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26dfb),
	.w1(32'hba6dc186),
	.w2(32'hbbcbeaba),
	.w3(32'h3a94b02f),
	.w4(32'h3c92b42a),
	.w5(32'h3ca0c3c2),
	.w6(32'h3aaa2a35),
	.w7(32'hbc7f6190),
	.w8(32'hbb39120a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9aed9),
	.w1(32'hb980b4e8),
	.w2(32'h3c28f985),
	.w3(32'h3c1232d0),
	.w4(32'hbba7f46c),
	.w5(32'h3c17773b),
	.w6(32'h3c2afa42),
	.w7(32'hbb4e2455),
	.w8(32'hbc43272a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445a2e),
	.w1(32'hba2a2bce),
	.w2(32'hbbe553ba),
	.w3(32'hb90a486c),
	.w4(32'h3ba79420),
	.w5(32'h3be61ab1),
	.w6(32'hbbd72006),
	.w7(32'hbbea1f3c),
	.w8(32'hbc1c4a3d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e648),
	.w1(32'h3bf78ed0),
	.w2(32'hbc13b79e),
	.w3(32'hbc0f8a4f),
	.w4(32'hbb1b717d),
	.w5(32'hbba245a3),
	.w6(32'hbc7c18db),
	.w7(32'hbc363e77),
	.w8(32'h3bff82ba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f3576),
	.w1(32'h3b1ec1e9),
	.w2(32'hbbafe860),
	.w3(32'hbc36f675),
	.w4(32'h3d31b612),
	.w5(32'hbbd2fbff),
	.w6(32'h3b7d8881),
	.w7(32'hbba14452),
	.w8(32'hbc037271),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a2cef),
	.w1(32'h3c02840b),
	.w2(32'hbc8f86ad),
	.w3(32'hbcbdb654),
	.w4(32'h3b6bb845),
	.w5(32'hbcbb336a),
	.w6(32'h3d53fb9b),
	.w7(32'h39741c74),
	.w8(32'hbb2d0af2),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39b384),
	.w1(32'h3c2b982d),
	.w2(32'h3c30bf94),
	.w3(32'h3b857421),
	.w4(32'h3bd9c248),
	.w5(32'hbbe064b2),
	.w6(32'hbc11a802),
	.w7(32'h3c451c19),
	.w8(32'hba1cc7d6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c845fc6),
	.w1(32'h3c9d6c56),
	.w2(32'hbc232575),
	.w3(32'hba88f3a3),
	.w4(32'h3c6158e0),
	.w5(32'hbbab1ace),
	.w6(32'hbc1752dd),
	.w7(32'hbc0da970),
	.w8(32'h3c4481bc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd41577),
	.w1(32'hbb90b22e),
	.w2(32'h3ca2a410),
	.w3(32'h3c9e8850),
	.w4(32'hbbf2c014),
	.w5(32'h3b7ecdf1),
	.w6(32'hbc34a5d8),
	.w7(32'hbc3129b6),
	.w8(32'hbc93d733),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20c4bc),
	.w1(32'h3d21c8db),
	.w2(32'hbcd55cba),
	.w3(32'h3aebed16),
	.w4(32'hbc971e70),
	.w5(32'h3ad688ed),
	.w6(32'hbba3eb71),
	.w7(32'hbc14b62f),
	.w8(32'hbbbbcbf1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd623b6),
	.w1(32'h3c51e479),
	.w2(32'h3c5801ef),
	.w3(32'h3d175803),
	.w4(32'hbc908ae0),
	.w5(32'h3c1d6a37),
	.w6(32'hbc0b1cc7),
	.w7(32'h3b387691),
	.w8(32'h3c3633ce),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fa840),
	.w1(32'h3c9957ff),
	.w2(32'h3c9e7d23),
	.w3(32'h3c444128),
	.w4(32'h3ca61ed4),
	.w5(32'h3ce71138),
	.w6(32'h3d0bff3e),
	.w7(32'h3cadfecc),
	.w8(32'h3a2706b0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc82ca1),
	.w1(32'hbccece81),
	.w2(32'h3cb75e14),
	.w3(32'hbc5e8816),
	.w4(32'h3c449d3a),
	.w5(32'hbc3a84ce),
	.w6(32'hbcb62c5e),
	.w7(32'h3c8ce158),
	.w8(32'h3bd714b4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d10d9),
	.w1(32'h3b128bc3),
	.w2(32'hbb439504),
	.w3(32'hbc768249),
	.w4(32'h3c8684c1),
	.w5(32'hbc3d5ecf),
	.w6(32'h3bba9996),
	.w7(32'hbbc4b9fc),
	.w8(32'hbb412c10),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd514be),
	.w1(32'hbc86acd0),
	.w2(32'hbcd99e5c),
	.w3(32'hbc5368e6),
	.w4(32'hbb3cd6b3),
	.w5(32'hbb1e630e),
	.w6(32'hbc18f128),
	.w7(32'h3d7833eb),
	.w8(32'hbadb14ab),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a521),
	.w1(32'h3cc44dce),
	.w2(32'hbc11068a),
	.w3(32'h3b9320b4),
	.w4(32'hbcfdfae2),
	.w5(32'hbc3cd678),
	.w6(32'hbd505d0a),
	.w7(32'h3d10b56f),
	.w8(32'h3cc4f62d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb630e),
	.w1(32'h3cda6764),
	.w2(32'h3cbc323e),
	.w3(32'h3ca8384c),
	.w4(32'hbc29bce7),
	.w5(32'h3ca43c97),
	.w6(32'hba6d4735),
	.w7(32'hbc96bbb9),
	.w8(32'h3c72b288),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6a3fd),
	.w1(32'h3cf154fb),
	.w2(32'hbb320431),
	.w3(32'h3bdf612d),
	.w4(32'h3c02060b),
	.w5(32'h3b81a4b1),
	.w6(32'hbc352e09),
	.w7(32'hb94caf64),
	.w8(32'h3c7846fa),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc275630),
	.w1(32'h3d423521),
	.w2(32'hbcbeef3b),
	.w3(32'h3d72ddad),
	.w4(32'h3c9255e8),
	.w5(32'h3a04008b),
	.w6(32'h3ca888a8),
	.w7(32'h3c0d8432),
	.w8(32'hbb2305dc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7913),
	.w1(32'h3c300aed),
	.w2(32'hbb29f8ac),
	.w3(32'h3c7b755a),
	.w4(32'h3be6bf43),
	.w5(32'h39325ac4),
	.w6(32'hbb9263ad),
	.w7(32'hbbc337d6),
	.w8(32'hbc5803ea),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fc5ce),
	.w1(32'h3cad21f3),
	.w2(32'hbb7bb250),
	.w3(32'h3c134406),
	.w4(32'hbc80edcb),
	.w5(32'h3bc1a384),
	.w6(32'h3ce3e771),
	.w7(32'h3c6c6967),
	.w8(32'h3c59e888),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f3714),
	.w1(32'h3ba32bdc),
	.w2(32'hbc1553ec),
	.w3(32'hbb7fb981),
	.w4(32'h3b2ebaab),
	.w5(32'hbc72799c),
	.w6(32'h3bcfd0e0),
	.w7(32'hbc50b197),
	.w8(32'hbc19c482),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a846ca1),
	.w1(32'hbc30c7c5),
	.w2(32'h3c5c9cba),
	.w3(32'h3b2437c6),
	.w4(32'hbc5fe116),
	.w5(32'h3d0003f7),
	.w6(32'hbba8b1f3),
	.w7(32'h3c2947d9),
	.w8(32'h3c8cef2c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c529c66),
	.w1(32'hbca3e192),
	.w2(32'hbb1961d7),
	.w3(32'hbc488881),
	.w4(32'h3c696b56),
	.w5(32'hbce8c9c0),
	.w6(32'h3cd26ae9),
	.w7(32'h3bd72f19),
	.w8(32'h3ab80994),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4537),
	.w1(32'h3c871937),
	.w2(32'h3678f630),
	.w3(32'h3a53a57f),
	.w4(32'h3c05917f),
	.w5(32'h3c50bff2),
	.w6(32'h3ccfe5c9),
	.w7(32'hbb4acc0b),
	.w8(32'hbbc94e1c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d24f9),
	.w1(32'h3ca594e6),
	.w2(32'hbc302b8e),
	.w3(32'hb9adcf19),
	.w4(32'h3c96d119),
	.w5(32'h3c7a9ede),
	.w6(32'hbbfaa9cb),
	.w7(32'hbc4f4bc0),
	.w8(32'h3bac943a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51de8d),
	.w1(32'h3baa18ed),
	.w2(32'h3c14211c),
	.w3(32'hbab7c862),
	.w4(32'hbc8697da),
	.w5(32'h3b8297c0),
	.w6(32'h3caf668c),
	.w7(32'hbc5df98c),
	.w8(32'h3c30f853),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9640ef),
	.w1(32'h3c822335),
	.w2(32'h3b9685b3),
	.w3(32'hbb8835ae),
	.w4(32'h3c53a86b),
	.w5(32'hbb9c5e4c),
	.w6(32'h3b369b8a),
	.w7(32'h3c7ea432),
	.w8(32'h3c9766df),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d59fa),
	.w1(32'hbd06e05d),
	.w2(32'h39950dfa),
	.w3(32'hb950eb44),
	.w4(32'hbcb28aee),
	.w5(32'hbb1a6030),
	.w6(32'h3cf5c110),
	.w7(32'h3c4690f5),
	.w8(32'hbcc4e739),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5350),
	.w1(32'h3bf53cf2),
	.w2(32'h3bb04505),
	.w3(32'hbb98166f),
	.w4(32'h3c043829),
	.w5(32'hb6e90896),
	.w6(32'hbbbd8acb),
	.w7(32'h3bb016be),
	.w8(32'hbaefd1d6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb68adb),
	.w1(32'h3c36c359),
	.w2(32'h3c2965f5),
	.w3(32'h3c1a5c8b),
	.w4(32'h3c009e93),
	.w5(32'h3b8d1caf),
	.w6(32'h3d172e34),
	.w7(32'h3a435da5),
	.w8(32'hbbc55b1a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14d46e),
	.w1(32'hbc5dbb08),
	.w2(32'hbc93579d),
	.w3(32'h3bb5105d),
	.w4(32'h3bda67a8),
	.w5(32'hbc617854),
	.w6(32'h3afa4f7f),
	.w7(32'hbcd0fc82),
	.w8(32'hbcccda49),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c677e),
	.w1(32'h3a53240d),
	.w2(32'h3ccf6d38),
	.w3(32'h3c92bb48),
	.w4(32'hbcbe7b05),
	.w5(32'h3c08b465),
	.w6(32'h3c35f3f9),
	.w7(32'hbaa2824a),
	.w8(32'h3d090f6e),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2879e7),
	.w1(32'hbc1cd8cd),
	.w2(32'hbdcb4e2f),
	.w3(32'h3ab52ac1),
	.w4(32'hbca6bdec),
	.w5(32'h3adfa1e8),
	.w6(32'h3d01f96d),
	.w7(32'hbd6888be),
	.w8(32'h3d5702c1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b4a75),
	.w1(32'h3bdb6851),
	.w2(32'hbc1093f7),
	.w3(32'hbbdfc666),
	.w4(32'h3ca7c89a),
	.w5(32'h3b63e36a),
	.w6(32'hbd6e2a2e),
	.w7(32'hbadf1213),
	.w8(32'h3b5dbf8a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef580e),
	.w1(32'hbbd8a7bf),
	.w2(32'h3aef6770),
	.w3(32'h399dacb3),
	.w4(32'h3b6a2c67),
	.w5(32'h3a904384),
	.w6(32'hbc293fbe),
	.w7(32'hbc300e17),
	.w8(32'hbb7c1131),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5925e1),
	.w1(32'hbb96a4b0),
	.w2(32'hbb14455c),
	.w3(32'hbb1f2632),
	.w4(32'h3abbf71d),
	.w5(32'h3b438530),
	.w6(32'h3a1798bb),
	.w7(32'hbbe1d568),
	.w8(32'h3bb4e5cf),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123d3e),
	.w1(32'hbb1a4e2c),
	.w2(32'h3d5d5bf1),
	.w3(32'h3a191359),
	.w4(32'h3ae20797),
	.w5(32'hbacf48a3),
	.w6(32'h3b466a61),
	.w7(32'hbc12b2da),
	.w8(32'hbb9e8e62),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925251),
	.w1(32'h3bc7f5e8),
	.w2(32'h3c0185e1),
	.w3(32'hbba2b262),
	.w4(32'h3b30a2dc),
	.w5(32'h3aed5e46),
	.w6(32'h3c1aa76d),
	.w7(32'hbba77932),
	.w8(32'h3bd95baa),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec9241),
	.w1(32'hbc01f744),
	.w2(32'h3b69304d),
	.w3(32'hbc3b00d6),
	.w4(32'hbbc5450a),
	.w5(32'h3a95fedb),
	.w6(32'h3c115c9c),
	.w7(32'hbc254f6b),
	.w8(32'h3c116c2a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b62be),
	.w1(32'h3bc94bea),
	.w2(32'h3ba3361b),
	.w3(32'hbbdcd93d),
	.w4(32'h3b566493),
	.w5(32'hbc869a94),
	.w6(32'h3bb5afc3),
	.w7(32'hbb8289b3),
	.w8(32'hbb972763),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c134474),
	.w1(32'hb97b6dd6),
	.w2(32'hbaadf184),
	.w3(32'hbc3cc29c),
	.w4(32'hbb200e8c),
	.w5(32'h3b8fe7d5),
	.w6(32'hbb570512),
	.w7(32'h3beb1ac5),
	.w8(32'hbc84cf48),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc875c44),
	.w1(32'hbbcae8a7),
	.w2(32'hbbd886d3),
	.w3(32'hbba3cc2d),
	.w4(32'hbc4e5586),
	.w5(32'h3b75cc93),
	.w6(32'hbb6ebe11),
	.w7(32'h3b2a94ac),
	.w8(32'hbb22885d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5233bd),
	.w1(32'h3bad0041),
	.w2(32'hbc03f950),
	.w3(32'hbbee22c2),
	.w4(32'h3b82de37),
	.w5(32'h3b333b5c),
	.w6(32'hbbf8c9d9),
	.w7(32'h3c3a3970),
	.w8(32'hbb8e425d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31e85a),
	.w1(32'hbbcf07f7),
	.w2(32'hbb1cca1c),
	.w3(32'hb9ced020),
	.w4(32'hbbc687e3),
	.w5(32'h3bdd9a47),
	.w6(32'hbb5d9a0d),
	.w7(32'h3c1a66e5),
	.w8(32'hba0731cf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf8caa),
	.w1(32'h3c1704b4),
	.w2(32'hbc9f7d4d),
	.w3(32'hb9f498a2),
	.w4(32'h3aa45b16),
	.w5(32'hbba9b298),
	.w6(32'h3b2f5ca3),
	.w7(32'hbbc4e822),
	.w8(32'hbb441d8f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39571a21),
	.w1(32'hbc8dae72),
	.w2(32'hbb9a3592),
	.w3(32'hbb7555e0),
	.w4(32'hbb9b9395),
	.w5(32'hb9bede71),
	.w6(32'h3c2fc9aa),
	.w7(32'hbc50822c),
	.w8(32'hbb94b59d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc8b60),
	.w1(32'h3bf1f3a0),
	.w2(32'h3b2a976b),
	.w3(32'h3bc29125),
	.w4(32'h3b537304),
	.w5(32'hbb1d0a13),
	.w6(32'hbaaa26aa),
	.w7(32'h3bd39b92),
	.w8(32'hba734e3d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1832b),
	.w1(32'h3b2ffef3),
	.w2(32'h3c4fb23f),
	.w3(32'h3b9b2f53),
	.w4(32'hba784c0b),
	.w5(32'h3acef97d),
	.w6(32'hb7cb625f),
	.w7(32'hbbc1d332),
	.w8(32'h3b63d29f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56458c),
	.w1(32'h39defa4a),
	.w2(32'hbd8d3f58),
	.w3(32'h3bb0d6df),
	.w4(32'hbbfc7619),
	.w5(32'h3a2b08a1),
	.w6(32'hbafcaa9f),
	.w7(32'hbb23a628),
	.w8(32'h3a6111ef),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd539e1),
	.w1(32'hba37dcfa),
	.w2(32'hbc505b35),
	.w3(32'h39cfb911),
	.w4(32'hbb3b016f),
	.w5(32'h393aea0e),
	.w6(32'hbbd085e2),
	.w7(32'hb966ad82),
	.w8(32'hbc03a934),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22d206),
	.w1(32'hbb098031),
	.w2(32'hbb7eb0b5),
	.w3(32'hbc60debc),
	.w4(32'hbb6030b5),
	.w5(32'h3c3a2fba),
	.w6(32'h39732977),
	.w7(32'hb9ae0cb3),
	.w8(32'hba1d575a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd638),
	.w1(32'hbb33486d),
	.w2(32'hbb75b0f5),
	.w3(32'hbb681d4c),
	.w4(32'hbbfd93c3),
	.w5(32'hb95b02ee),
	.w6(32'hbb370a43),
	.w7(32'hbd8a3ba9),
	.w8(32'hbb473e4c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85aa13),
	.w1(32'hbb1f049a),
	.w2(32'hbb8b6496),
	.w3(32'h37cbe4be),
	.w4(32'h3b05d4ac),
	.w5(32'h3a27ebeb),
	.w6(32'hbb93971b),
	.w7(32'hbb1c28b4),
	.w8(32'hbaebc64c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d63b188),
	.w1(32'hbb4c47d1),
	.w2(32'hba3270ab),
	.w3(32'hbbda90ea),
	.w4(32'hba7359cd),
	.w5(32'hbc217be7),
	.w6(32'hbbf266d0),
	.w7(32'hbb4586eb),
	.w8(32'hbb186049),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc58dcf),
	.w1(32'h3b81b347),
	.w2(32'h3bf6fbd2),
	.w3(32'hba809329),
	.w4(32'hbc4cc7dd),
	.w5(32'hbb82ba7a),
	.w6(32'hbc4db38d),
	.w7(32'hbbba38ff),
	.w8(32'hba8c9952),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20dd3b),
	.w1(32'h3a677748),
	.w2(32'hbb16545d),
	.w3(32'h3ab0f643),
	.w4(32'hbbacfe7e),
	.w5(32'h3b034b39),
	.w6(32'hba127b2d),
	.w7(32'h3a7bba7f),
	.w8(32'hbc2d215b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebf1ac),
	.w1(32'hbc9c0b79),
	.w2(32'hbb42774c),
	.w3(32'h3be5c003),
	.w4(32'hbb123a7e),
	.w5(32'hbaa9469d),
	.w6(32'hbacf793e),
	.w7(32'h3c0b0275),
	.w8(32'hbcb93db9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc733f49),
	.w1(32'hbb220df4),
	.w2(32'h3b948373),
	.w3(32'hbab8c682),
	.w4(32'hbbc471ab),
	.w5(32'hbbf1a65f),
	.w6(32'hb8b6c83c),
	.w7(32'h3a8d6433),
	.w8(32'hba95116e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68629c),
	.w1(32'hbc676929),
	.w2(32'hbc87ac92),
	.w3(32'h3a8754f7),
	.w4(32'h3cb537db),
	.w5(32'h3b8989c2),
	.w6(32'hbb0b515e),
	.w7(32'h3b40fb02),
	.w8(32'h3a37f480),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34a1a3),
	.w1(32'h3bb8857a),
	.w2(32'hbb63312e),
	.w3(32'hba26cbaf),
	.w4(32'h3b700dd2),
	.w5(32'hbb037cce),
	.w6(32'hbd1eca70),
	.w7(32'h3b02436c),
	.w8(32'h3bb71f90),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17cd28),
	.w1(32'h3a2b85e1),
	.w2(32'hbc4a0d8c),
	.w3(32'h3c27ddb5),
	.w4(32'h3a909ba6),
	.w5(32'hbba891b4),
	.w6(32'hbb533556),
	.w7(32'hbcb3c444),
	.w8(32'h3bb1993e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb760e1b),
	.w1(32'h3c12b0b7),
	.w2(32'hbb074b1c),
	.w3(32'hbc760e3d),
	.w4(32'hbb58669e),
	.w5(32'hba90e42d),
	.w6(32'hba99a654),
	.w7(32'h3b5fec34),
	.w8(32'hbb284103),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c5f0d),
	.w1(32'h3b3004e3),
	.w2(32'hbb686ed4),
	.w3(32'hbb1106fb),
	.w4(32'hbad3ba08),
	.w5(32'hbbd7be82),
	.w6(32'hbb7ff01d),
	.w7(32'hbbe8eedb),
	.w8(32'hbb3fcfaf),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cbcb1),
	.w1(32'h3c90aebb),
	.w2(32'h3bbea881),
	.w3(32'h3b285b01),
	.w4(32'hbbc4b09f),
	.w5(32'hbb8112b2),
	.w6(32'hbc1733c8),
	.w7(32'hbb60ee06),
	.w8(32'hba7476a9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e0606),
	.w1(32'hbb8cdacb),
	.w2(32'hbbc465d1),
	.w3(32'h3a48bfe1),
	.w4(32'h3bfe5b85),
	.w5(32'hbace5a8e),
	.w6(32'hbbc543f1),
	.w7(32'h3825644a),
	.w8(32'h3bb0ba3c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79a437),
	.w1(32'hbba6f024),
	.w2(32'hbb313f9c),
	.w3(32'hbbf274d4),
	.w4(32'h3b2036c7),
	.w5(32'hbaad5e37),
	.w6(32'h3b354fad),
	.w7(32'h3be3e428),
	.w8(32'hb9a3c168),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc132927),
	.w1(32'hbbb469e4),
	.w2(32'h3bdc26cc),
	.w3(32'hbb9e4614),
	.w4(32'hbbc38b4d),
	.w5(32'h3beca377),
	.w6(32'hbbbb0f92),
	.w7(32'h38ca91a8),
	.w8(32'h3ae36dab),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe54b42),
	.w1(32'hbbd9277b),
	.w2(32'hbaa6b95e),
	.w3(32'hba48c183),
	.w4(32'hbc09f33a),
	.w5(32'hbc17d22c),
	.w6(32'hbb366705),
	.w7(32'h3ccc9ff6),
	.w8(32'hbc21822d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001f14),
	.w1(32'hbc53385e),
	.w2(32'hbc5f4277),
	.w3(32'h3b3230f0),
	.w4(32'hbbd4d608),
	.w5(32'h3b6a2c7c),
	.w6(32'hbc04d402),
	.w7(32'h3b25f354),
	.w8(32'hb9e73b5a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046e45),
	.w1(32'hbb0ef8d5),
	.w2(32'hbb38220f),
	.w3(32'h3bc5fe9a),
	.w4(32'hbb511ccf),
	.w5(32'h3aa832df),
	.w6(32'hbb14c396),
	.w7(32'hb9989dc7),
	.w8(32'h3b7ed26a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82e69),
	.w1(32'hb92910a2),
	.w2(32'h39d5b012),
	.w3(32'h39fa89a9),
	.w4(32'hbc7d4025),
	.w5(32'hbb820818),
	.w6(32'h3ba9c248),
	.w7(32'hbbed0e48),
	.w8(32'hbab54b6f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dc505),
	.w1(32'hbc42ef34),
	.w2(32'hba9b673d),
	.w3(32'hbc2bef3f),
	.w4(32'hbb3527e5),
	.w5(32'h3c03bca2),
	.w6(32'h3b18d6f3),
	.w7(32'h3ce3a231),
	.w8(32'h3b212426),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826b07),
	.w1(32'h3b230cd3),
	.w2(32'hbac7b0ee),
	.w3(32'h3a2cf2b1),
	.w4(32'h3b2d9b18),
	.w5(32'h3d1507c4),
	.w6(32'hba6b05fc),
	.w7(32'hbc62807b),
	.w8(32'hbb8ac36c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba808a98),
	.w1(32'h3bfed9ad),
	.w2(32'hbac17e83),
	.w3(32'h3b4d6460),
	.w4(32'h39a82938),
	.w5(32'h3b546f8f),
	.w6(32'hbb25813b),
	.w7(32'h3ce400d2),
	.w8(32'h3c3711d2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f578),
	.w1(32'h3ba77082),
	.w2(32'hbbb998b1),
	.w3(32'hbb773b74),
	.w4(32'h38c114e4),
	.w5(32'hbb142b17),
	.w6(32'hbb9b87cb),
	.w7(32'hbaeae66e),
	.w8(32'h3b20b387),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc4011),
	.w1(32'h3b5d1bbc),
	.w2(32'h35ad916d),
	.w3(32'hbb55128a),
	.w4(32'hbbe0922e),
	.w5(32'hbb80c7a5),
	.w6(32'h3c034e63),
	.w7(32'hbb6dd3c1),
	.w8(32'hb7850d45),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0188a2),
	.w1(32'hb88bcaf3),
	.w2(32'hbb8b59d3),
	.w3(32'hbc5ffd4f),
	.w4(32'hbad0ed5d),
	.w5(32'h3bd8cb27),
	.w6(32'hba31d2b1),
	.w7(32'hbbd0f76c),
	.w8(32'hbc049a10),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46c533),
	.w1(32'hbc3c5e71),
	.w2(32'h3a8a561d),
	.w3(32'hbb0db223),
	.w4(32'h3b97a662),
	.w5(32'h3b81669d),
	.w6(32'hbab1e26f),
	.w7(32'h3ad9c442),
	.w8(32'h3bd9bcf5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9652df),
	.w1(32'h3abb0dda),
	.w2(32'hbb547484),
	.w3(32'h39ad6358),
	.w4(32'h38b5d0d6),
	.w5(32'h3aa2ffe0),
	.w6(32'hbc597cdb),
	.w7(32'hbc372a82),
	.w8(32'hbb7e816d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72cbb4),
	.w1(32'hbac0f434),
	.w2(32'h3bf111a6),
	.w3(32'hbab206d1),
	.w4(32'h3a1b8106),
	.w5(32'hbbade826),
	.w6(32'h3ad0d609),
	.w7(32'hbb8fc07d),
	.w8(32'hbc051f1f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ed1b7),
	.w1(32'hbb5ce4ca),
	.w2(32'hbc45f6b3),
	.w3(32'hbc5b5ed8),
	.w4(32'hbba3e467),
	.w5(32'hbc15e319),
	.w6(32'hbb780a42),
	.w7(32'hb7e1ec20),
	.w8(32'hbbc61845),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75e26),
	.w1(32'h3cc63e13),
	.w2(32'h3bd67e70),
	.w3(32'h3a25625a),
	.w4(32'h3c385e43),
	.w5(32'hbc400417),
	.w6(32'hbaab8086),
	.w7(32'h3a0beb42),
	.w8(32'hb95130bd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd5345),
	.w1(32'h3c041088),
	.w2(32'hbc03e4e8),
	.w3(32'hbb11bd02),
	.w4(32'hbb6dd752),
	.w5(32'hbab317d4),
	.w6(32'h3c4948b1),
	.w7(32'hbcad91fb),
	.w8(32'hbb4112ab),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b164c20),
	.w1(32'hbb39796f),
	.w2(32'hbbe0915a),
	.w3(32'h3b57cc83),
	.w4(32'hbb4278fe),
	.w5(32'h3ba95760),
	.w6(32'h3c8b028c),
	.w7(32'h3c7d7b3e),
	.w8(32'hba00d5d6),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bf3dd),
	.w1(32'h3bf10e99),
	.w2(32'h3b8508ef),
	.w3(32'h3b97907a),
	.w4(32'hbb0e41e8),
	.w5(32'hbc828289),
	.w6(32'hbc0cea55),
	.w7(32'h3ae75da3),
	.w8(32'hbac63a49),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43265),
	.w1(32'hbabdd2b8),
	.w2(32'h37f64916),
	.w3(32'hbbd8c22c),
	.w4(32'hbb6f7544),
	.w5(32'hbaa061a4),
	.w6(32'hba1ea8b7),
	.w7(32'hbb17931e),
	.w8(32'h3b12067a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf30c5f),
	.w1(32'hba0e293a),
	.w2(32'h3b150e14),
	.w3(32'hbac0d1fa),
	.w4(32'hb9e21d56),
	.w5(32'h3b380c44),
	.w6(32'hb990d973),
	.w7(32'hbab0ed1e),
	.w8(32'h3b6a35d1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2fd36),
	.w1(32'hbb1fe19e),
	.w2(32'h3bbbfe90),
	.w3(32'hba371705),
	.w4(32'h398a922d),
	.w5(32'h3c6e8ec3),
	.w6(32'hbbf1a23e),
	.w7(32'hba7dfbe6),
	.w8(32'h3b883ae9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac823b0),
	.w1(32'hbc32626f),
	.w2(32'h3a3da653),
	.w3(32'hbbf6b366),
	.w4(32'hbc4bd302),
	.w5(32'hbbab5a8f),
	.w6(32'hba87b5aa),
	.w7(32'h3cb157fc),
	.w8(32'hbc42bac1),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9d3ca),
	.w1(32'hbb77fa5b),
	.w2(32'hbb8382b4),
	.w3(32'h3c268e69),
	.w4(32'h3bb11c53),
	.w5(32'hbb9a9a08),
	.w6(32'h3c0da0e3),
	.w7(32'hbc84a6e2),
	.w8(32'hbb929e52),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeb6ad),
	.w1(32'hbb96777d),
	.w2(32'h3b568af0),
	.w3(32'h3bc1fda2),
	.w4(32'hbbb2d917),
	.w5(32'h3cf1a9c8),
	.w6(32'hbbaf0e5d),
	.w7(32'hbbd9df60),
	.w8(32'h3ae42f66),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18053a),
	.w1(32'h3baf257b),
	.w2(32'hbc364ae0),
	.w3(32'hbc333863),
	.w4(32'h3b6b2a37),
	.w5(32'hbc7aa936),
	.w6(32'h3a466f60),
	.w7(32'h3b9f4a21),
	.w8(32'hba1f378f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbabf0e),
	.w1(32'h3b3f660b),
	.w2(32'h3b098217),
	.w3(32'hbab6da30),
	.w4(32'h3c005e56),
	.w5(32'hbb866f6a),
	.w6(32'h3a2cba28),
	.w7(32'h3bfbeb2f),
	.w8(32'hbc453895),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf34b7f),
	.w1(32'hbc2d9deb),
	.w2(32'hbc732a76),
	.w3(32'hbc594cc2),
	.w4(32'hbb2d5064),
	.w5(32'h3b86777a),
	.w6(32'h3b6482c1),
	.w7(32'h3c479c19),
	.w8(32'h3b7ad4c8),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ecf1f),
	.w1(32'hba00acb1),
	.w2(32'hba9b33ba),
	.w3(32'hbbb2df9a),
	.w4(32'hb8b6f896),
	.w5(32'hbb8cf702),
	.w6(32'hbb427c74),
	.w7(32'hbab53bd4),
	.w8(32'h3b361d8b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a7dc2),
	.w1(32'hbb207f3d),
	.w2(32'hbc9aedb3),
	.w3(32'hbb77e3a4),
	.w4(32'h3b34a864),
	.w5(32'h3bdac97e),
	.w6(32'hbc749c93),
	.w7(32'hbb1f4659),
	.w8(32'hbbe48bf7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ae21e),
	.w1(32'hba8521dc),
	.w2(32'h3b51615a),
	.w3(32'hbbbaf998),
	.w4(32'h3abd28bc),
	.w5(32'hbc45a9f5),
	.w6(32'hb90775dd),
	.w7(32'h3c276019),
	.w8(32'h3b0e8d48),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a4aa8),
	.w1(32'hbaea9b71),
	.w2(32'hb946c9cc),
	.w3(32'hbbee74d2),
	.w4(32'h3a821032),
	.w5(32'h3b3c6978),
	.w6(32'hbb9bf980),
	.w7(32'h3b230860),
	.w8(32'h3ba5a98f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae77d0e),
	.w1(32'h3c6b075f),
	.w2(32'h3be7d419),
	.w3(32'h3b836c91),
	.w4(32'hbbf353fc),
	.w5(32'hba2990c4),
	.w6(32'h3b5e06c2),
	.w7(32'h3b6a98e9),
	.w8(32'hbcbedd0c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50b935),
	.w1(32'hbbb79fc8),
	.w2(32'h3c0c1a18),
	.w3(32'hbbad6ea7),
	.w4(32'hbc7387ae),
	.w5(32'h3c8acb19),
	.w6(32'h3b0a4eb3),
	.w7(32'hbbf76cf2),
	.w8(32'hbba18eea),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a6b6),
	.w1(32'h3a98832c),
	.w2(32'hbc297ee3),
	.w3(32'hbc3eb1c5),
	.w4(32'hbbaa3887),
	.w5(32'hbb636069),
	.w6(32'hbb08ae38),
	.w7(32'hbb0ea196),
	.w8(32'h3b51fda2),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e02e9),
	.w1(32'h3b87a80d),
	.w2(32'h3c43ec16),
	.w3(32'hba95a49e),
	.w4(32'hbaf5d18f),
	.w5(32'hbc061c3c),
	.w6(32'hbba66c58),
	.w7(32'h3aec1783),
	.w8(32'h39391ec9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6ff5f),
	.w1(32'h3c7c69a7),
	.w2(32'hbc2af4e8),
	.w3(32'h3b385315),
	.w4(32'h3bed2962),
	.w5(32'hbad04745),
	.w6(32'hbc071cc3),
	.w7(32'h3bc11b92),
	.w8(32'hbc10f75c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8aa2d),
	.w1(32'hbb9d676b),
	.w2(32'hbc1fc28c),
	.w3(32'h3afb5b6e),
	.w4(32'h39d34cf2),
	.w5(32'hbc258ed4),
	.w6(32'h3b908ebc),
	.w7(32'hbabde544),
	.w8(32'h3c2313a6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d9c4),
	.w1(32'h3a12c593),
	.w2(32'hbbfffb15),
	.w3(32'hb90f6ff1),
	.w4(32'h3c1c0f9b),
	.w5(32'h3bce0cb6),
	.w6(32'hbc347dfa),
	.w7(32'h3b7dd80f),
	.w8(32'h3c43e4b4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f997c),
	.w1(32'h3cbaf1b2),
	.w2(32'h3d179b54),
	.w3(32'h3b48e6e3),
	.w4(32'hbc1d2d15),
	.w5(32'hbcd3b759),
	.w6(32'h3c66fa8e),
	.w7(32'h3c944ca0),
	.w8(32'hbc3bed54),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64efd),
	.w1(32'hbbcd858b),
	.w2(32'hbbd07ddb),
	.w3(32'h3aa9f46b),
	.w4(32'h3bbd7f2e),
	.w5(32'hbbcc0f6a),
	.w6(32'hbbdcfca0),
	.w7(32'hbbde90a1),
	.w8(32'h3ab80bda),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d045b),
	.w1(32'hbc3adaba),
	.w2(32'hbb81bb38),
	.w3(32'hbb648751),
	.w4(32'h3b877447),
	.w5(32'h3afc1b61),
	.w6(32'h3a84eff5),
	.w7(32'hbb168b90),
	.w8(32'hba9586da),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00c84),
	.w1(32'hbb89170e),
	.w2(32'hba88ce5a),
	.w3(32'hba67c275),
	.w4(32'hbc3f1d7c),
	.w5(32'h3b957ff2),
	.w6(32'h3c02f838),
	.w7(32'hbb66afeb),
	.w8(32'h3b8f792b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3650114c),
	.w1(32'h3c03201a),
	.w2(32'hbc6d8030),
	.w3(32'hbabc944e),
	.w4(32'hbb4917d7),
	.w5(32'hbb9a92ba),
	.w6(32'h3c64a927),
	.w7(32'h3c6c091a),
	.w8(32'hbb103f69),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeedb02),
	.w1(32'h36aa49fa),
	.w2(32'hbba49a46),
	.w3(32'h3c0ab971),
	.w4(32'hbbc3c03e),
	.w5(32'h3b2db87e),
	.w6(32'hbc19c55d),
	.w7(32'h3a8c3d5f),
	.w8(32'h3b162706),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c75af),
	.w1(32'h3cecef19),
	.w2(32'hbb359632),
	.w3(32'h3bdb1a04),
	.w4(32'hbac27e25),
	.w5(32'h3c2b52f5),
	.w6(32'h3b287ee5),
	.w7(32'hbc3da742),
	.w8(32'hbc890696),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d530a),
	.w1(32'hbbf7764e),
	.w2(32'h3b75ec29),
	.w3(32'h3b0c3d12),
	.w4(32'h3bb8457a),
	.w5(32'h3b47be4a),
	.w6(32'hbac32cbf),
	.w7(32'hbb4c534b),
	.w8(32'h3b04b645),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ab2b6),
	.w1(32'hbb234690),
	.w2(32'hb9d3b409),
	.w3(32'h3c402c27),
	.w4(32'h3c1874e4),
	.w5(32'h3c4c1215),
	.w6(32'hbb9609c0),
	.w7(32'hb9686540),
	.w8(32'hbc965204),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a8b5),
	.w1(32'h391b3fdb),
	.w2(32'hba294c86),
	.w3(32'hb94513bc),
	.w4(32'h3a708993),
	.w5(32'hbb4108ea),
	.w6(32'hbba83982),
	.w7(32'hbc167832),
	.w8(32'h398e95eb),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a129174),
	.w1(32'h3b85d5d1),
	.w2(32'h3a90074e),
	.w3(32'h3b5c47a5),
	.w4(32'h3b339bc5),
	.w5(32'hbc0711ed),
	.w6(32'hbb756be1),
	.w7(32'hbae00b95),
	.w8(32'hbaf04737),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6265f),
	.w1(32'h38d5b154),
	.w2(32'hbc01cab9),
	.w3(32'h3c118a50),
	.w4(32'h3bc7829e),
	.w5(32'h3be52234),
	.w6(32'hbc0f8d52),
	.w7(32'hba313223),
	.w8(32'h3a458875),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8c83b),
	.w1(32'h3a82a2e6),
	.w2(32'h3af500fc),
	.w3(32'hbba6f900),
	.w4(32'h3bcffa03),
	.w5(32'hba955d59),
	.w6(32'hbb642fcd),
	.w7(32'h3b9054f6),
	.w8(32'h3c573a68),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3499ca),
	.w1(32'h3bcd4f3e),
	.w2(32'h3c3b19f9),
	.w3(32'h3b2bbfb7),
	.w4(32'h3b8412e5),
	.w5(32'h3a960e78),
	.w6(32'hbc4e43c5),
	.w7(32'h3b83f932),
	.w8(32'hbca9e67f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192390),
	.w1(32'hba832be9),
	.w2(32'h3b18adc5),
	.w3(32'hbc2a114a),
	.w4(32'hba1009d4),
	.w5(32'hbb9ba648),
	.w6(32'hbc4bd598),
	.w7(32'hbac86954),
	.w8(32'hbb68272f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8e0d3),
	.w1(32'h3bd91284),
	.w2(32'hbab3f618),
	.w3(32'hb998a43b),
	.w4(32'h3c015ced),
	.w5(32'h3c25a67e),
	.w6(32'h3c26dbd0),
	.w7(32'h3bbdaf5b),
	.w8(32'hba8d5331),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule