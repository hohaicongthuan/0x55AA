module layer_8_featuremap_170(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061305),
	.w1(32'hbcc2be75),
	.w2(32'h3bce7dac),
	.w3(32'hbc050170),
	.w4(32'hbc554c26),
	.w5(32'hbc47195a),
	.w6(32'hbc93bc0d),
	.w7(32'h3d065995),
	.w8(32'h3bc4af8f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdf70d),
	.w1(32'h3afe2812),
	.w2(32'h395ffc8e),
	.w3(32'h3cccbdba),
	.w4(32'h3a468df5),
	.w5(32'hba066e3c),
	.w6(32'h3bdd9827),
	.w7(32'h38cdc2de),
	.w8(32'hbb6b7097),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d95a0),
	.w1(32'hbb6b0ee7),
	.w2(32'h3c1f3890),
	.w3(32'hba6a7af6),
	.w4(32'h39d92886),
	.w5(32'hbc1580a5),
	.w6(32'h3b8c9aa4),
	.w7(32'h3c80215e),
	.w8(32'hbc132a02),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4ad37),
	.w1(32'hbc884b62),
	.w2(32'h3c8140f0),
	.w3(32'h3bbbdd6c),
	.w4(32'hbbc7795d),
	.w5(32'hbb878735),
	.w6(32'hbb5d5550),
	.w7(32'h3c1dd455),
	.w8(32'hba07e1c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1058c),
	.w1(32'h3c159499),
	.w2(32'h3b7cf4e0),
	.w3(32'h3caa6340),
	.w4(32'h3bf3da2f),
	.w5(32'h3b9261c6),
	.w6(32'h3c2a710a),
	.w7(32'h3bc241ab),
	.w8(32'h3be2a7cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219b2c),
	.w1(32'hbc4c248b),
	.w2(32'hbbcd9641),
	.w3(32'hbae6da93),
	.w4(32'hbba83653),
	.w5(32'h3c00c087),
	.w6(32'hbc87df73),
	.w7(32'hbc363885),
	.w8(32'hbc3bee5f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd2bd0),
	.w1(32'h3aa168de),
	.w2(32'hbb62a9bc),
	.w3(32'hbb4bb0e1),
	.w4(32'hb990bd1e),
	.w5(32'hbb214330),
	.w6(32'h3a815891),
	.w7(32'hb9f00822),
	.w8(32'h3b1a21a8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3654c4),
	.w1(32'hbbcd87d0),
	.w2(32'h3c0cf439),
	.w3(32'h38323868),
	.w4(32'hbb86f65c),
	.w5(32'h3c65129d),
	.w6(32'h3bf45ecb),
	.w7(32'h3c28fa8a),
	.w8(32'hbca381bd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf4443),
	.w1(32'h3c49459d),
	.w2(32'hbb2f9fcb),
	.w3(32'h3bf76383),
	.w4(32'h3c9f172c),
	.w5(32'hbbd5730a),
	.w6(32'h3c85f5e8),
	.w7(32'h3b6d10a4),
	.w8(32'h3a3fe1c1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba221b),
	.w1(32'h3c2ed450),
	.w2(32'hbc3a1673),
	.w3(32'hbb31d363),
	.w4(32'hb752ca48),
	.w5(32'hbb9a4d3d),
	.w6(32'hbbabc14b),
	.w7(32'h3afe962b),
	.w8(32'h3ca0757c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63d777),
	.w1(32'hbbefef6b),
	.w2(32'h3d09dd07),
	.w3(32'hbc57fdb1),
	.w4(32'hbc6638da),
	.w5(32'h3bcf3da8),
	.w6(32'h3c19003c),
	.w7(32'h3bf369f8),
	.w8(32'hbc648208),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc15d91),
	.w1(32'hbb8e9e0f),
	.w2(32'hbc78fe64),
	.w3(32'h3cba6bd1),
	.w4(32'hbba29ec2),
	.w5(32'hbbe0d966),
	.w6(32'h3b1d209b),
	.w7(32'hbb15dba3),
	.w8(32'hba90f89b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf993d),
	.w1(32'h3bcc5940),
	.w2(32'hbb5ed540),
	.w3(32'hbb708a0b),
	.w4(32'h3c0aaf84),
	.w5(32'hbb3dc561),
	.w6(32'h3bad36eb),
	.w7(32'hbc1c3e34),
	.w8(32'h3b8d786c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52c561),
	.w1(32'hbce2170e),
	.w2(32'hbca50cd7),
	.w3(32'hba8bcf70),
	.w4(32'hbbcf5fb3),
	.w5(32'hbce1fba7),
	.w6(32'hbcf9267b),
	.w7(32'h3b5f0c9d),
	.w8(32'h3ca1f392),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25ddb2),
	.w1(32'h3c06dcc0),
	.w2(32'hb9c3866d),
	.w3(32'h3c2d36ad),
	.w4(32'h3bef9273),
	.w5(32'h3a904b20),
	.w6(32'h3b5945a3),
	.w7(32'hbaad8c24),
	.w8(32'h3a9de428),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b18ee8),
	.w1(32'hbad37b29),
	.w2(32'hbcba751f),
	.w3(32'h3a491ab0),
	.w4(32'h39ad6692),
	.w5(32'hbc993da2),
	.w6(32'hbc46aff5),
	.w7(32'hbb5c7a77),
	.w8(32'hbb48d044),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1dc1),
	.w1(32'h3cf64219),
	.w2(32'h3d870bf9),
	.w3(32'hba81664c),
	.w4(32'hbc04a833),
	.w5(32'h3d678aa6),
	.w6(32'h3cfbf45b),
	.w7(32'hbccea862),
	.w8(32'h3d08411a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c238078),
	.w1(32'hbb777895),
	.w2(32'hbbe52106),
	.w3(32'h3c9fc689),
	.w4(32'h3c118c23),
	.w5(32'hbc916a35),
	.w6(32'h3bf14f07),
	.w7(32'h3c6860cc),
	.w8(32'h3c2b8865),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2f37a5),
	.w1(32'h3c751297),
	.w2(32'h3981a8e1),
	.w3(32'h3c6a3d17),
	.w4(32'h3c17e628),
	.w5(32'h3c34d7fd),
	.w6(32'h3c461954),
	.w7(32'hbb5a8be8),
	.w8(32'h3adb4903),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99fe39),
	.w1(32'h3c962461),
	.w2(32'h3c420ea8),
	.w3(32'h3c142209),
	.w4(32'h3c0b31c4),
	.w5(32'h3bc5a7fa),
	.w6(32'h3c855bf1),
	.w7(32'h3c14961d),
	.w8(32'h3b7b2b81),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17bdb3),
	.w1(32'hbb60b51d),
	.w2(32'hbca8ca23),
	.w3(32'hbc381af6),
	.w4(32'hbb9f9faa),
	.w5(32'hbc975626),
	.w6(32'hba29d0dc),
	.w7(32'hbc3170ca),
	.w8(32'hbbccd122),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbce9a2),
	.w1(32'h3b966080),
	.w2(32'h3c1ba867),
	.w3(32'hbc463acc),
	.w4(32'hbbb7cca9),
	.w5(32'h3c31a125),
	.w6(32'h3aa27304),
	.w7(32'hbc4bbebd),
	.w8(32'hbc706b2a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1bbb5a),
	.w1(32'h3cc4cac4),
	.w2(32'h3b032190),
	.w3(32'hbb4a913d),
	.w4(32'h3c8fb76a),
	.w5(32'h3c2b4fa1),
	.w6(32'h3c9d401c),
	.w7(32'hbbe57a8c),
	.w8(32'h3b3069a2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb289a4a),
	.w1(32'h3c37f0f2),
	.w2(32'h3bebf8ba),
	.w3(32'hbbd018d0),
	.w4(32'hb9c725fa),
	.w5(32'h3c9ba744),
	.w6(32'h3b8e8403),
	.w7(32'hba079339),
	.w8(32'hbc0e2cb5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01d1fd),
	.w1(32'h3c864b9c),
	.w2(32'h3b68d4d4),
	.w3(32'hbc21641a),
	.w4(32'h3c1ae843),
	.w5(32'h3b3ccafd),
	.w6(32'h3c7dc5ce),
	.w7(32'hbabf5731),
	.w8(32'hbbc6ab61),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3609),
	.w1(32'hbb839475),
	.w2(32'h3bfdbd12),
	.w3(32'h3b09b930),
	.w4(32'h3b9c799b),
	.w5(32'hbbf018e6),
	.w6(32'hbc076d78),
	.w7(32'h3ca6a92a),
	.w8(32'h3bca7e73),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81488e),
	.w1(32'h3c47a52a),
	.w2(32'h3c2d61bd),
	.w3(32'hbbea62b1),
	.w4(32'h3bf51ec4),
	.w5(32'h3c00cbb7),
	.w6(32'hbb216da1),
	.w7(32'h3be7fdde),
	.w8(32'hbb8ff9da),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caea90f),
	.w1(32'h3b5398e2),
	.w2(32'h3d3382c1),
	.w3(32'h3cde14b2),
	.w4(32'hbb894d91),
	.w5(32'hbc4b2a0f),
	.w6(32'h3cb2f4ef),
	.w7(32'h3d005736),
	.w8(32'h3c138295),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4c4de),
	.w1(32'h3c15733f),
	.w2(32'hbb8a18d5),
	.w3(32'h3c822fb3),
	.w4(32'h3bd70060),
	.w5(32'hbb294757),
	.w6(32'h3bb520e8),
	.w7(32'hbb2068f8),
	.w8(32'hbbac3f0c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecd849),
	.w1(32'h3ab66fc0),
	.w2(32'hbba5bdd5),
	.w3(32'hbc2d8356),
	.w4(32'hbc0f4b48),
	.w5(32'hbc82d017),
	.w6(32'h3aec8cbc),
	.w7(32'hbafc4548),
	.w8(32'h3c88bac5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb34799),
	.w1(32'h3a74aaae),
	.w2(32'hbb0c2acd),
	.w3(32'hba8b08a0),
	.w4(32'h3a551603),
	.w5(32'hbbbe718c),
	.w6(32'hbb01f16c),
	.w7(32'h399161d4),
	.w8(32'h3a122c24),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad324a),
	.w1(32'h3c8b91ed),
	.w2(32'h3b4ae2ee),
	.w3(32'h3a9fd22e),
	.w4(32'h3b18cfcb),
	.w5(32'h3c087742),
	.w6(32'h3c3f5184),
	.w7(32'h3bae49ab),
	.w8(32'h3b9a7b9a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ebd6a),
	.w1(32'hbc2f910a),
	.w2(32'h3c0f8c6b),
	.w3(32'hbc066adb),
	.w4(32'hb984ad19),
	.w5(32'hbc67ac0b),
	.w6(32'hbc28ac1d),
	.w7(32'h3b66fec9),
	.w8(32'h398224b6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2acb6),
	.w1(32'hbc1184c1),
	.w2(32'hbbafe0a2),
	.w3(32'h3ca23867),
	.w4(32'hbb8722cb),
	.w5(32'hbc8c6d57),
	.w6(32'hbc00c3f0),
	.w7(32'hbb64705b),
	.w8(32'h3b3849d7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee988f),
	.w1(32'h3c041d9f),
	.w2(32'h3c258156),
	.w3(32'h3b9c44cf),
	.w4(32'h3bf4101b),
	.w5(32'h3c22e8f1),
	.w6(32'h3c373727),
	.w7(32'h3bc00363),
	.w8(32'h3bd93baf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb959ef),
	.w1(32'h3ca6c686),
	.w2(32'h3c58d0d7),
	.w3(32'hba661e7f),
	.w4(32'h3b1eb7a9),
	.w5(32'h3c0cf672),
	.w6(32'h3c2c53e2),
	.w7(32'h3c54ab86),
	.w8(32'hbbf4a6a6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ff6dd),
	.w1(32'h3bec0831),
	.w2(32'h3b86fbdc),
	.w3(32'hbc1758cc),
	.w4(32'h3b564174),
	.w5(32'h3c04f86f),
	.w6(32'h3b56321b),
	.w7(32'hb99cff4b),
	.w8(32'hbaf0214c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2aa48),
	.w1(32'h3c518f26),
	.w2(32'h3babb194),
	.w3(32'h3a46c759),
	.w4(32'h3c5e07f6),
	.w5(32'h3b1b8d16),
	.w6(32'h3bb68efb),
	.w7(32'h391a584b),
	.w8(32'h3b104d37),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b055fc8),
	.w1(32'h3c24aa99),
	.w2(32'h3b02416a),
	.w3(32'h3b7dcb94),
	.w4(32'h3b3bfad1),
	.w5(32'h3baaa915),
	.w6(32'h3c04d064),
	.w7(32'hbba465fa),
	.w8(32'hbc266dd8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf93830),
	.w1(32'hba65e8f7),
	.w2(32'h3c0b521a),
	.w3(32'h3b52c19f),
	.w4(32'hbbfbb561),
	.w5(32'h3bd2ab3d),
	.w6(32'h3b76d1d7),
	.w7(32'hbbd18b71),
	.w8(32'hbbe8b74e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48e1d),
	.w1(32'h3abc3cbf),
	.w2(32'h3a35b172),
	.w3(32'h3bec31fd),
	.w4(32'h3b855413),
	.w5(32'h3b034d6c),
	.w6(32'h3c6e8dea),
	.w7(32'h3b1d78cf),
	.w8(32'h3b2b1f35),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8dc4b),
	.w1(32'h3a64df91),
	.w2(32'hbba65154),
	.w3(32'h3b0faf80),
	.w4(32'h3be0da8a),
	.w5(32'hbbc5fd4c),
	.w6(32'h3bc4b9da),
	.w7(32'h3b5acb8a),
	.w8(32'hbc62a0ab),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba6c70),
	.w1(32'hbb8658af),
	.w2(32'h3bfdd5a0),
	.w3(32'hba9a2d72),
	.w4(32'hbae78060),
	.w5(32'h3addc897),
	.w6(32'hbb36ab3c),
	.w7(32'hbaccd0ea),
	.w8(32'hbbb3ce9a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91a84c),
	.w1(32'h3b8c4481),
	.w2(32'hbc9277e4),
	.w3(32'h3c1ce8da),
	.w4(32'h3c32d75c),
	.w5(32'hbc2a3c89),
	.w6(32'h3bd6303e),
	.w7(32'hbb4e9702),
	.w8(32'h3c029fd6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b420e),
	.w1(32'hbb92ec71),
	.w2(32'h3c6a2027),
	.w3(32'h3afe7881),
	.w4(32'hbc2e749d),
	.w5(32'h3b36c437),
	.w6(32'hbc62a76c),
	.w7(32'hbc64fca2),
	.w8(32'hbcc6414b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5762ea),
	.w1(32'h3adb6d1f),
	.w2(32'hbb8a24d8),
	.w3(32'hb6ad0114),
	.w4(32'hba87f71f),
	.w5(32'hbb672eb0),
	.w6(32'h3b228f94),
	.w7(32'hbb1790fb),
	.w8(32'h390a4cec),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7fc2d),
	.w1(32'hbb1da598),
	.w2(32'hbc4b3029),
	.w3(32'hbbc350c5),
	.w4(32'h3b2fc4d9),
	.w5(32'hbc02a791),
	.w6(32'h3ba043af),
	.w7(32'hbc17c832),
	.w8(32'hbb8887cc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52c714),
	.w1(32'h3c98db93),
	.w2(32'h3c4f9b75),
	.w3(32'h3b0877ae),
	.w4(32'h3afa7d8d),
	.w5(32'h3c86d59f),
	.w6(32'h3cb2bdcf),
	.w7(32'hba210036),
	.w8(32'hbcf7957b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0acff3),
	.w1(32'h3c2d5767),
	.w2(32'h3c32c2af),
	.w3(32'hbb2e9978),
	.w4(32'hbbd9bc8e),
	.w5(32'hbc13fce5),
	.w6(32'h3c6249c6),
	.w7(32'hbb9fa7d6),
	.w8(32'hbd0c2426),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2d0671),
	.w1(32'hb9fa46bc),
	.w2(32'hbc9e698d),
	.w3(32'hbc854f68),
	.w4(32'hbb1419e2),
	.w5(32'hbc57a981),
	.w6(32'h3a299a2c),
	.w7(32'hbbd3d07c),
	.w8(32'h3aec417b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc9e56c),
	.w1(32'hbbe93182),
	.w2(32'hbbae43b0),
	.w3(32'hbbafcf5d),
	.w4(32'hbba4e1a5),
	.w5(32'hbb6af07c),
	.w6(32'hb99ada88),
	.w7(32'hbc17d49e),
	.w8(32'hbb6f3040),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806710),
	.w1(32'h3c82f88c),
	.w2(32'h3c8ae3b9),
	.w3(32'h3c99d865),
	.w4(32'h3be1f0a2),
	.w5(32'h3c63a3f3),
	.w6(32'h3ca4e411),
	.w7(32'h3bbb1867),
	.w8(32'hbb5035f4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31522e),
	.w1(32'h3bcdc841),
	.w2(32'hbb9989b9),
	.w3(32'h3c7d321e),
	.w4(32'h3b72d700),
	.w5(32'hbbb9a56d),
	.w6(32'h3c5d3e21),
	.w7(32'hbb38d7f6),
	.w8(32'hbb185df3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfb59a),
	.w1(32'hbb85638b),
	.w2(32'hbc644ecc),
	.w3(32'h3b795d2c),
	.w4(32'h3b7684fd),
	.w5(32'hbc09ffd7),
	.w6(32'hbad084b3),
	.w7(32'hbc17f9b1),
	.w8(32'h3b081dd7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895daa),
	.w1(32'h3c29640d),
	.w2(32'hbc7c0ee0),
	.w3(32'h3a8ff734),
	.w4(32'h3bb3b5e0),
	.w5(32'hbbc9dcc2),
	.w6(32'h3bc86424),
	.w7(32'hbb956906),
	.w8(32'h3c12374d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79acfc),
	.w1(32'hbc562953),
	.w2(32'hbc8c3fc1),
	.w3(32'h3a0cbc1d),
	.w4(32'h3b5450a7),
	.w5(32'hbd083127),
	.w6(32'hbb6bb6e4),
	.w7(32'h3c3b0a9f),
	.w8(32'h3a2ba0ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfddc7e),
	.w1(32'hbaa52c3e),
	.w2(32'hbcb4d09d),
	.w3(32'h3a1dd6c9),
	.w4(32'hbb26a960),
	.w5(32'hbc4dc645),
	.w6(32'h3b944255),
	.w7(32'hbc596b34),
	.w8(32'hb917b2ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0499aa),
	.w1(32'h3b05fdae),
	.w2(32'hbba048e1),
	.w3(32'hbba199ac),
	.w4(32'hbb605e2a),
	.w5(32'hbb8395a1),
	.w6(32'h3b895341),
	.w7(32'hbbe9e068),
	.w8(32'hbb00263a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9537054),
	.w1(32'hbb2a3d79),
	.w2(32'hbb8fb9a2),
	.w3(32'h392c3078),
	.w4(32'hbb5e193f),
	.w5(32'hbb951519),
	.w6(32'h3af11204),
	.w7(32'hbb3b4e4f),
	.w8(32'hbbd145cc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7cd23),
	.w1(32'h3c5d1164),
	.w2(32'h3c66f955),
	.w3(32'hbb52a50c),
	.w4(32'h3b880aaa),
	.w5(32'h3c7b392a),
	.w6(32'h3c0937af),
	.w7(32'hbb21c39a),
	.w8(32'hbc9042cf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfeb1e6),
	.w1(32'h3b785ffe),
	.w2(32'h3b58103e),
	.w3(32'h3b17e2b3),
	.w4(32'hba079e8f),
	.w5(32'h3bce86f0),
	.w6(32'hbb0bab13),
	.w7(32'hbb988a94),
	.w8(32'h3ba2b3ea),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7423af),
	.w1(32'h3ba2cb36),
	.w2(32'hbba847a3),
	.w3(32'h3b56e40b),
	.w4(32'h3b8e5832),
	.w5(32'hb9f1a977),
	.w6(32'h3b1fb28f),
	.w7(32'hbc1842fd),
	.w8(32'h3bf76817),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45917d),
	.w1(32'h3c51be13),
	.w2(32'hbb7131cf),
	.w3(32'hba86e531),
	.w4(32'h3b0194d7),
	.w5(32'hbc164130),
	.w6(32'h3c2e8f97),
	.w7(32'h3be7880e),
	.w8(32'h3c3180dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c150831),
	.w1(32'hbbef7bcf),
	.w2(32'hbbc3726c),
	.w3(32'hbbab2571),
	.w4(32'hbb59e042),
	.w5(32'hbb7cca41),
	.w6(32'hbb84b8c3),
	.w7(32'h39f499a4),
	.w8(32'hbbd6a2d6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc369d97),
	.w1(32'hbb01e84a),
	.w2(32'hbb9aadba),
	.w3(32'hbc0cb10a),
	.w4(32'h390ff1e4),
	.w5(32'hbb7b6203),
	.w6(32'hbb8a4cd5),
	.w7(32'hbbe46889),
	.w8(32'hbc057e09),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff0f0b),
	.w1(32'hb997ad02),
	.w2(32'hba6d612e),
	.w3(32'hbbae4c10),
	.w4(32'hbb191476),
	.w5(32'h3c14cb47),
	.w6(32'hbb74ed05),
	.w7(32'hbc114ecb),
	.w8(32'hbc05793c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9033fd),
	.w1(32'hbc614170),
	.w2(32'hbd342d83),
	.w3(32'hbc46cb72),
	.w4(32'hbb8f4355),
	.w5(32'hbcf31f67),
	.w6(32'h3b3a7f68),
	.w7(32'hbc4c486d),
	.w8(32'hbc1c5939),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc969118),
	.w1(32'hbc7f8389),
	.w2(32'hbcc4605b),
	.w3(32'hbccfb9f1),
	.w4(32'hbc149caa),
	.w5(32'hbc8514f1),
	.w6(32'hbc2655ff),
	.w7(32'hbca7c8f3),
	.w8(32'hbc7fe134),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2b06),
	.w1(32'hbc208aad),
	.w2(32'hbaf60665),
	.w3(32'hbc0646ef),
	.w4(32'h3b142c21),
	.w5(32'hbcc7e3a5),
	.w6(32'hbc557af3),
	.w7(32'h3b8e0548),
	.w8(32'h3a949a4b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2b3b10),
	.w1(32'h3cb2b24e),
	.w2(32'h3c297cf4),
	.w3(32'h3cd09c96),
	.w4(32'h3c1120a5),
	.w5(32'h3c6bc603),
	.w6(32'h3ca486fc),
	.w7(32'h3bf77389),
	.w8(32'hbbf17238),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf86d09),
	.w1(32'h3b782ee0),
	.w2(32'hbaa4a89f),
	.w3(32'hbc67ccb8),
	.w4(32'h3ab2716c),
	.w5(32'h37cfb36a),
	.w6(32'hbb174f20),
	.w7(32'hbbbb8f05),
	.w8(32'hbb5328d6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf66e81),
	.w1(32'hba2087d8),
	.w2(32'h3c013d54),
	.w3(32'h3c1648ec),
	.w4(32'h3c11edb1),
	.w5(32'hbbe456d8),
	.w6(32'h3b3f04e2),
	.w7(32'h3c8e473d),
	.w8(32'h3c0941e5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e0063),
	.w1(32'h3c5c52e2),
	.w2(32'h3c6c0f59),
	.w3(32'h3bb23d8c),
	.w4(32'h3b8d976e),
	.w5(32'h3a59ee2a),
	.w6(32'h3c94c390),
	.w7(32'h3bfd620b),
	.w8(32'hbb0dcec3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1b45),
	.w1(32'h3c6032ae),
	.w2(32'h3c0b90e1),
	.w3(32'h3b89b9b4),
	.w4(32'h3c7144f9),
	.w5(32'h3c87a5ff),
	.w6(32'h3c03a9af),
	.w7(32'h3bbd0e6a),
	.w8(32'h3bbe3de0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc013f64),
	.w1(32'h3b831ada),
	.w2(32'hbaacfbc0),
	.w3(32'hba5bf541),
	.w4(32'h3ba3a96c),
	.w5(32'h3c0495c5),
	.w6(32'h3bd5a312),
	.w7(32'hb9940f9d),
	.w8(32'hbb426e50),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf25d63),
	.w1(32'h3c2b4997),
	.w2(32'h3c240334),
	.w3(32'hba18c182),
	.w4(32'h3be1204c),
	.w5(32'h3bd595dd),
	.w6(32'hba232507),
	.w7(32'h3bfab8b5),
	.w8(32'h3b249ac7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1a4a),
	.w1(32'h3b76acfd),
	.w2(32'h3c38fefd),
	.w3(32'hbb51989a),
	.w4(32'h39b82df8),
	.w5(32'h3c18391d),
	.w6(32'hbaef0af6),
	.w7(32'h3a2d384c),
	.w8(32'hbbe16f2e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc02f0f),
	.w1(32'h3b88ef67),
	.w2(32'h3b1c18ca),
	.w3(32'h3b152503),
	.w4(32'hba0fc368),
	.w5(32'hbb3cf498),
	.w6(32'hbab6f7c7),
	.w7(32'hbaa36703),
	.w8(32'hbb29a4fa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b7e97),
	.w1(32'hbbf2c971),
	.w2(32'hba95c482),
	.w3(32'hbbe9269b),
	.w4(32'hbab297b6),
	.w5(32'hbc5ad75b),
	.w6(32'hbbee0f7f),
	.w7(32'h3ba50e64),
	.w8(32'hbb5d249c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91986c),
	.w1(32'hbc784df4),
	.w2(32'h3c4a6033),
	.w3(32'h3c04582d),
	.w4(32'hbbfe8756),
	.w5(32'hbca75bc5),
	.w6(32'hbb7452d2),
	.w7(32'h3cada721),
	.w8(32'hbbd94aa9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90bbb5),
	.w1(32'hbc44b804),
	.w2(32'hbbc373c4),
	.w3(32'h3c75f5b6),
	.w4(32'hbb1edc9f),
	.w5(32'hbc8b55df),
	.w6(32'hbbef32de),
	.w7(32'h3ab97723),
	.w8(32'h3bae3b28),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c3c74),
	.w1(32'hbc6a556d),
	.w2(32'h3a9a118f),
	.w3(32'h3c17a784),
	.w4(32'h3c70ee4e),
	.w5(32'hbc9f972e),
	.w6(32'hbc60827d),
	.w7(32'h3c201bbd),
	.w8(32'h3c0661c3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b52c3),
	.w1(32'h3b2bd41f),
	.w2(32'h3bde97ec),
	.w3(32'h3c9398d4),
	.w4(32'h3b898433),
	.w5(32'h3b2dd2c8),
	.w6(32'h3c1736b7),
	.w7(32'hbb14f1ce),
	.w8(32'hbc0835b0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a559),
	.w1(32'hbbb3ace8),
	.w2(32'h3c1f8496),
	.w3(32'h3c4734e8),
	.w4(32'h3bdbbb09),
	.w5(32'h3ca60c7c),
	.w6(32'hbae66088),
	.w7(32'hbbb6bb4b),
	.w8(32'hbb96e73d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7762e8),
	.w1(32'hbc880f3d),
	.w2(32'hbb8c91a3),
	.w3(32'h3cf55b36),
	.w4(32'h3b80b977),
	.w5(32'hbca1697f),
	.w6(32'h3b150d1e),
	.w7(32'h3cc1f46c),
	.w8(32'h3c39477b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00a118),
	.w1(32'h3b9f2a7d),
	.w2(32'h3cb46dbd),
	.w3(32'h3c7d931b),
	.w4(32'h3c7ba511),
	.w5(32'h3beec5a8),
	.w6(32'h3ac658e8),
	.w7(32'h3c95e027),
	.w8(32'h3c827c32),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9246),
	.w1(32'h3b83ee2f),
	.w2(32'h3b3a9d22),
	.w3(32'hbb72ded1),
	.w4(32'h3a086b08),
	.w5(32'h3b144534),
	.w6(32'hb7f7c389),
	.w7(32'h3afc8b3b),
	.w8(32'hbb6afd20),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a98e5),
	.w1(32'h3b7b1d5f),
	.w2(32'hbb44ec56),
	.w3(32'h3b091c27),
	.w4(32'hbaa65ddd),
	.w5(32'hbbbf9436),
	.w6(32'h3c187ea3),
	.w7(32'hbaa9ce1f),
	.w8(32'hbb94919f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4869ca),
	.w1(32'hbaabd571),
	.w2(32'hbb56ba3a),
	.w3(32'hbbe00863),
	.w4(32'h3b5ccacf),
	.w5(32'h3ad0e199),
	.w6(32'h3a9be53d),
	.w7(32'h3b5efc08),
	.w8(32'h3b14909d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf00485),
	.w1(32'h3c6346aa),
	.w2(32'h3c30e0c9),
	.w3(32'h3aa70a38),
	.w4(32'hb9f7a368),
	.w5(32'h38d084c9),
	.w6(32'h3c20b71b),
	.w7(32'h3ba28ca0),
	.w8(32'hbcb9e4b5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ac4a6),
	.w1(32'h3c21e46e),
	.w2(32'h37c11ac7),
	.w3(32'hbab5a5f1),
	.w4(32'h3c01c04c),
	.w5(32'hba5afc11),
	.w6(32'h3ca095b1),
	.w7(32'h3c3f8fff),
	.w8(32'h3bf6e833),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c2b06),
	.w1(32'hbc590175),
	.w2(32'hbc8e16d9),
	.w3(32'h39be839a),
	.w4(32'hbc0de86a),
	.w5(32'hbc7e3707),
	.w6(32'hbc74ee0e),
	.w7(32'hbbd0a099),
	.w8(32'h3c135ee7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbac354),
	.w1(32'hbaa85adc),
	.w2(32'hbad00706),
	.w3(32'h3b6d5c4a),
	.w4(32'hba81f4a6),
	.w5(32'h398044ed),
	.w6(32'h3bc1baef),
	.w7(32'h3991a3ff),
	.w8(32'hbb177e36),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2d3a7),
	.w1(32'hb9b26aa1),
	.w2(32'hbbda5fca),
	.w3(32'hbb12eaf5),
	.w4(32'hbb06ffc7),
	.w5(32'hbb4957f8),
	.w6(32'h3acdcd32),
	.w7(32'hbbc10e45),
	.w8(32'hbc251ceb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb50ee),
	.w1(32'h3bb71f8e),
	.w2(32'hbc88510d),
	.w3(32'hbbb4bd26),
	.w4(32'hbbf1ed74),
	.w5(32'hbb727b2f),
	.w6(32'hbb4b68a4),
	.w7(32'hbc7e8f91),
	.w8(32'hbbf43600),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc135a30),
	.w1(32'hbb6511d6),
	.w2(32'hbb237566),
	.w3(32'hbc6e5532),
	.w4(32'hb955a701),
	.w5(32'hb9e0b4e2),
	.w6(32'h3aad1e24),
	.w7(32'h3b3b5b04),
	.w8(32'h3b83a348),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5008d0),
	.w1(32'h3c86cce0),
	.w2(32'h3c2abd10),
	.w3(32'h3c44042b),
	.w4(32'h3c2ba4b5),
	.w5(32'h3c47d1c6),
	.w6(32'h3c97879c),
	.w7(32'h3b57133f),
	.w8(32'hbc13e517),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185215),
	.w1(32'h3bf66b0f),
	.w2(32'h3c010dba),
	.w3(32'hbb21d1ac),
	.w4(32'h3b89b7fd),
	.w5(32'h3be3fec9),
	.w6(32'h3bd5306d),
	.w7(32'h3ba8840b),
	.w8(32'hbba16653),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf291bc),
	.w1(32'h3b58658b),
	.w2(32'hbc57a5f0),
	.w3(32'h3bd3511b),
	.w4(32'hbad75807),
	.w5(32'hbbf0fa8e),
	.w6(32'h3c25cd6e),
	.w7(32'hbb3f5f0a),
	.w8(32'hbb17f143),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59238a),
	.w1(32'hbc09d06c),
	.w2(32'h3cdb5981),
	.w3(32'hbbfd2000),
	.w4(32'hbc7d3cd1),
	.w5(32'h3c0e4854),
	.w6(32'hba9c0c37),
	.w7(32'hba8e6cf0),
	.w8(32'hbca60023),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba960f18),
	.w1(32'h3bfc1adc),
	.w2(32'hbd294203),
	.w3(32'h3cd5c730),
	.w4(32'h3cc711e5),
	.w5(32'hbc3409ab),
	.w6(32'hba10d111),
	.w7(32'hbb8d059a),
	.w8(32'h3c7a59fc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0254ae),
	.w1(32'h3b0e7f84),
	.w2(32'h3c1f64f3),
	.w3(32'hbbd0702b),
	.w4(32'h3a5292c1),
	.w5(32'h3bc6a995),
	.w6(32'hbb08c2e8),
	.w7(32'hbc0be27f),
	.w8(32'h3c13ccdc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903b7dd),
	.w1(32'hbcaaf052),
	.w2(32'hbc9dd9f5),
	.w3(32'hbb4b075e),
	.w4(32'h3b33a65a),
	.w5(32'hbcc98564),
	.w6(32'hbc8305b8),
	.w7(32'h3b4a32af),
	.w8(32'h3c9b2fcb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bf5a8),
	.w1(32'h3ca41a50),
	.w2(32'h3c8adc75),
	.w3(32'h3c5b38d7),
	.w4(32'h3b31e9c3),
	.w5(32'h3b89daec),
	.w6(32'h3cec0a26),
	.w7(32'h3c23def9),
	.w8(32'hbc8e4860),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa43af),
	.w1(32'hbc3a3127),
	.w2(32'hbc8d0145),
	.w3(32'hbc1872d5),
	.w4(32'h3be6ba05),
	.w5(32'hbc023148),
	.w6(32'hbb9417a3),
	.w7(32'h3bddd2a3),
	.w8(32'h3a166399),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066160),
	.w1(32'h3be9bff2),
	.w2(32'hbb80059e),
	.w3(32'h3c9b0478),
	.w4(32'h3c2afcc8),
	.w5(32'hbad97d77),
	.w6(32'h3c5455aa),
	.w7(32'h3a7c564c),
	.w8(32'h3b6a544b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf1be),
	.w1(32'h3c650f78),
	.w2(32'h3a0f47d3),
	.w3(32'h3aaeb1bf),
	.w4(32'h3c401277),
	.w5(32'h3c0a58d9),
	.w6(32'h3bc731e9),
	.w7(32'h3be942c0),
	.w8(32'hbb236d2b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bae79),
	.w1(32'h39909ba3),
	.w2(32'hbbe54e18),
	.w3(32'h3b15c8c8),
	.w4(32'h3c2467e4),
	.w5(32'hbb694d13),
	.w6(32'hbb13f3bd),
	.w7(32'h3b209c0b),
	.w8(32'h3c7158d3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd62acd),
	.w1(32'h3aff2058),
	.w2(32'hbc26fac9),
	.w3(32'h3bac57ec),
	.w4(32'hb9a65c55),
	.w5(32'hbb40e638),
	.w6(32'h3bb6e8fb),
	.w7(32'h3bcbca09),
	.w8(32'h3c924a04),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb193ad),
	.w1(32'h3aaef648),
	.w2(32'h39c523eb),
	.w3(32'hb9fa0609),
	.w4(32'h3b630304),
	.w5(32'hba964126),
	.w6(32'h3b41bd50),
	.w7(32'h3bae3c60),
	.w8(32'h3a0ab553),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ebc0),
	.w1(32'hbce4e925),
	.w2(32'hbbc01275),
	.w3(32'h3c0d06c0),
	.w4(32'hba52e483),
	.w5(32'hbcb06bb8),
	.w6(32'hbb7309e1),
	.w7(32'h3b466610),
	.w8(32'h3c1ffe81),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceacb8d),
	.w1(32'h3ba030c2),
	.w2(32'h3a2d5dce),
	.w3(32'h3cd53a49),
	.w4(32'h3b845bc1),
	.w5(32'h3b6dc490),
	.w6(32'h3b6a6d1a),
	.w7(32'hb97a33eb),
	.w8(32'h3ad89ab5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95334f),
	.w1(32'hbaf523f4),
	.w2(32'hbb2b9b23),
	.w3(32'hbbfe72cb),
	.w4(32'hbbc381bd),
	.w5(32'hbbb538ec),
	.w6(32'hbbcad2ce),
	.w7(32'hbbe4912d),
	.w8(32'hbb4a52f5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa59428),
	.w1(32'hbb074ce8),
	.w2(32'h3bb7e5fa),
	.w3(32'hb9832c7c),
	.w4(32'h3c1d478e),
	.w5(32'hbaf81d61),
	.w6(32'h3beaadc2),
	.w7(32'h3c74bf5f),
	.w8(32'hbbc26bf0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31c7ae),
	.w1(32'h39da969b),
	.w2(32'hbb86d05c),
	.w3(32'hbc2f0fa8),
	.w4(32'h3ada77f8),
	.w5(32'hbc02cfce),
	.w6(32'h3a90ba23),
	.w7(32'hb9dba71b),
	.w8(32'hba506a92),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa215cb),
	.w1(32'hbbb0091f),
	.w2(32'hbba1326e),
	.w3(32'h3b38c0ae),
	.w4(32'hbbc2cee8),
	.w5(32'hbbe11e8b),
	.w6(32'hbba18d03),
	.w7(32'hbbfb1f42),
	.w8(32'hbbcef2c0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b16ce),
	.w1(32'h3a4c6207),
	.w2(32'h3b68b4a3),
	.w3(32'hb9eab333),
	.w4(32'h3a9f423a),
	.w5(32'h3bd68850),
	.w6(32'h3baea10e),
	.w7(32'h39dcaad9),
	.w8(32'h3bc8e385),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd827d7),
	.w1(32'hbc2cc3be),
	.w2(32'hbbe646b5),
	.w3(32'h3bba645b),
	.w4(32'hbc13deb8),
	.w5(32'hbc348ef2),
	.w6(32'hbb5729a9),
	.w7(32'hbbe77ee0),
	.w8(32'h38c1c216),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79ae7c),
	.w1(32'hbc225fdc),
	.w2(32'hbc82e107),
	.w3(32'h3a115f64),
	.w4(32'h3b0b7c10),
	.w5(32'hbca43a5d),
	.w6(32'hbca88472),
	.w7(32'h3b1374d8),
	.w8(32'h3b829c4a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f4e8e),
	.w1(32'h3a6b79b2),
	.w2(32'h3a9166d5),
	.w3(32'hba461aa2),
	.w4(32'hbbb0a515),
	.w5(32'h3b10c1e0),
	.w6(32'h3bd78695),
	.w7(32'hba137503),
	.w8(32'hbbedb865),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2bea),
	.w1(32'hbc707157),
	.w2(32'hba9ff052),
	.w3(32'hbb980274),
	.w4(32'hbaa9ddc9),
	.w5(32'hbcd043d8),
	.w6(32'hbc7a17cd),
	.w7(32'h3a405d51),
	.w8(32'h3b87c61a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d237258),
	.w1(32'hbbf1e148),
	.w2(32'h39c4c4fd),
	.w3(32'h3babb156),
	.w4(32'hbb53d449),
	.w5(32'hbbee1fd6),
	.w6(32'hbb812c29),
	.w7(32'hba446761),
	.w8(32'hbc292944),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab14b24),
	.w1(32'h3b257990),
	.w2(32'h394892a7),
	.w3(32'h3b82542b),
	.w4(32'h3b05bb71),
	.w5(32'h3b377479),
	.w6(32'h3bb5104d),
	.w7(32'h3b1adfe9),
	.w8(32'hb98b8df7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf0dc),
	.w1(32'hba1ff016),
	.w2(32'h39c83885),
	.w3(32'hbbb5d398),
	.w4(32'hbba3918c),
	.w5(32'h3bb5f1be),
	.w6(32'hbb4b3cb6),
	.w7(32'hbc45e516),
	.w8(32'hbb904e18),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2ca73),
	.w1(32'h3c5449b7),
	.w2(32'hbcf1bf53),
	.w3(32'h3a96d75b),
	.w4(32'h3c2d478c),
	.w5(32'h3c97a98d),
	.w6(32'hbbef817a),
	.w7(32'hbc2f40bf),
	.w8(32'h3d340e77),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb58fb3),
	.w1(32'h3c2ded12),
	.w2(32'h3c8dee00),
	.w3(32'hbc14bd62),
	.w4(32'h3b944e99),
	.w5(32'h3c6c1204),
	.w6(32'h3cbbecff),
	.w7(32'hbbeb9da3),
	.w8(32'hbd0a741d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd178c8f),
	.w1(32'h3adb8795),
	.w2(32'h3a55e2a0),
	.w3(32'hbc62f6ac),
	.w4(32'h3b0ef97d),
	.w5(32'h3a4aca0c),
	.w6(32'h3a02afc7),
	.w7(32'h3aa37aeb),
	.w8(32'h3a93b140),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e34bbc),
	.w1(32'hbabe7bb7),
	.w2(32'h3bbc30b1),
	.w3(32'h391bfed8),
	.w4(32'hbbc208ce),
	.w5(32'h3b5164f5),
	.w6(32'hbb513d31),
	.w7(32'h3b7f516e),
	.w8(32'hbb3817bc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule