module layer_10_featuremap_218(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17d1ff),
	.w1(32'h3b7eb672),
	.w2(32'h3a75f436),
	.w3(32'h3a1dcd6d),
	.w4(32'h3b3d24dd),
	.w5(32'h3b539a9f),
	.w6(32'h3b10b880),
	.w7(32'h3b7f1a9f),
	.w8(32'h3b743f72),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba570b9),
	.w1(32'hb9fe8f13),
	.w2(32'h39c87940),
	.w3(32'h3b62467b),
	.w4(32'hba8dc715),
	.w5(32'hba1a0794),
	.w6(32'h3a19741d),
	.w7(32'hbaaed933),
	.w8(32'h3a86889e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38880130),
	.w1(32'hb972c12f),
	.w2(32'h3927f413),
	.w3(32'hb7b7fca4),
	.w4(32'hb9af76ac),
	.w5(32'hba48f52d),
	.w6(32'hb9d27c02),
	.w7(32'hba68c125),
	.w8(32'hb8730b83),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c8833),
	.w1(32'h3a94c187),
	.w2(32'h3a90f463),
	.w3(32'h3910d1e6),
	.w4(32'h3adaf705),
	.w5(32'h3aa69278),
	.w6(32'h39c0250e),
	.w7(32'hb9422554),
	.w8(32'hba13bbd3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0e64e),
	.w1(32'h3b19be8d),
	.w2(32'h3ab5c07e),
	.w3(32'h397cafee),
	.w4(32'h3b343227),
	.w5(32'h3adaebb2),
	.w6(32'h3b1dbdfc),
	.w7(32'h3a6477dc),
	.w8(32'h39b1c032),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae29d75),
	.w1(32'h39a466df),
	.w2(32'h3a4e18e9),
	.w3(32'h3a98c155),
	.w4(32'h3a67010f),
	.w5(32'h3a49f158),
	.w6(32'h3a744a2a),
	.w7(32'h3a8bbae6),
	.w8(32'h3aa13470),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a861eb9),
	.w1(32'h3b03fce1),
	.w2(32'h3b31fcbd),
	.w3(32'h3ab89733),
	.w4(32'h3b692f7f),
	.w5(32'h3b73d3d7),
	.w6(32'h3ae25eff),
	.w7(32'h3b1020eb),
	.w8(32'h3b868d1e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8029),
	.w1(32'h3b0df8c4),
	.w2(32'h3ae89f55),
	.w3(32'h3bb3137b),
	.w4(32'h3b64143d),
	.w5(32'h3abe1fbc),
	.w6(32'h3b1cdbb6),
	.w7(32'h39ea37d5),
	.w8(32'h3b15614b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9b1d),
	.w1(32'hba06f509),
	.w2(32'h39ccf8bb),
	.w3(32'hba1fc23e),
	.w4(32'hb986730a),
	.w5(32'h395d9630),
	.w6(32'hb9cfcf6d),
	.w7(32'h39eb2ee8),
	.w8(32'h388a8f95),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24829),
	.w1(32'h3b6e8924),
	.w2(32'h3b9f5cc1),
	.w3(32'h3b912c39),
	.w4(32'h3ab6104c),
	.w5(32'h3b37e8a8),
	.w6(32'h3b66730b),
	.w7(32'h3a6530d7),
	.w8(32'h3b9dbb91),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2696d),
	.w1(32'h3a0f8234),
	.w2(32'h39eb77ed),
	.w3(32'h3ab5a0b4),
	.w4(32'hb8903f61),
	.w5(32'hb9af69af),
	.w6(32'h3a8769fb),
	.w7(32'hb98e34d5),
	.w8(32'h3901f5e3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4c78a),
	.w1(32'hbb193018),
	.w2(32'hb97d7bae),
	.w3(32'h3a8e2082),
	.w4(32'hba7473ae),
	.w5(32'h3adc85ef),
	.w6(32'h3a6e41e8),
	.w7(32'hba4ec105),
	.w8(32'h3b45da2e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82be5c),
	.w1(32'h3ae461e3),
	.w2(32'h3b94d733),
	.w3(32'h3b028455),
	.w4(32'h3ab57c62),
	.w5(32'h3b2f95e1),
	.w6(32'h373a327e),
	.w7(32'hb99a6b65),
	.w8(32'h3b284f16),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9585de4),
	.w1(32'hbad4e914),
	.w2(32'hbae415b1),
	.w3(32'hb9e67a43),
	.w4(32'hbaf82582),
	.w5(32'hbb30c249),
	.w6(32'hbb161419),
	.w7(32'hbb3d1a13),
	.w8(32'hbadf3e89),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d18be),
	.w1(32'h3b857bab),
	.w2(32'h3b6c7996),
	.w3(32'hba718211),
	.w4(32'h3b3144b5),
	.w5(32'h3b0c14d4),
	.w6(32'h3b126630),
	.w7(32'h3a68fc8b),
	.w8(32'h3a48bf8f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4a1a0),
	.w1(32'h3b7a5a80),
	.w2(32'h3b93bd75),
	.w3(32'h3b30a468),
	.w4(32'h3a738442),
	.w5(32'h3a6cf86b),
	.w6(32'h3b8d1e3b),
	.w7(32'h3ae98eca),
	.w8(32'h3add7da4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ed914),
	.w1(32'h3a839e5d),
	.w2(32'h3aeaaf55),
	.w3(32'h3ad557f3),
	.w4(32'h3b0b8f94),
	.w5(32'h3a7bd139),
	.w6(32'h3944d789),
	.w7(32'h3a7a2baf),
	.w8(32'h3a230969),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75a4b1),
	.w1(32'h3b16e700),
	.w2(32'h3bab0dd1),
	.w3(32'h3b7fb6e2),
	.w4(32'h3b23a095),
	.w5(32'h3b96e8b4),
	.w6(32'h3b484486),
	.w7(32'h3b1dfb73),
	.w8(32'h3bac5b0c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b127591),
	.w1(32'h3a559a56),
	.w2(32'h3b46f515),
	.w3(32'h3b0fa737),
	.w4(32'h3a87c2f5),
	.w5(32'h3b16cc58),
	.w6(32'h3955049d),
	.w7(32'h3a2c8aa5),
	.w8(32'h3b289e53),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03bcc4),
	.w1(32'hba297a7c),
	.w2(32'hb88a33a2),
	.w3(32'hba013dce),
	.w4(32'hba519b60),
	.w5(32'hba3bcedf),
	.w6(32'hba4f55d4),
	.w7(32'hba479d8a),
	.w8(32'hba7615b1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59cb1b),
	.w1(32'hb9ccb632),
	.w2(32'hb8747e92),
	.w3(32'hb9e24add),
	.w4(32'hba0dabcd),
	.w5(32'hb91a81cc),
	.w6(32'hb9e2f53a),
	.w7(32'hb885b694),
	.w8(32'hb9684a3a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721e139),
	.w1(32'h395983a0),
	.w2(32'h3a76a683),
	.w3(32'hb91353a3),
	.w4(32'h3aa729ae),
	.w5(32'h3b0d18cd),
	.w6(32'hba4b52fa),
	.w7(32'hba94ba7f),
	.w8(32'h3b120c38),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c481a),
	.w1(32'h3b0c288c),
	.w2(32'h3b7a9264),
	.w3(32'h3be28e74),
	.w4(32'h3a4781eb),
	.w5(32'h3b478cf8),
	.w6(32'h3b64adac),
	.w7(32'h3aa9131a),
	.w8(32'h3b96d207),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e6711),
	.w1(32'h3ae9852f),
	.w2(32'h3ba68545),
	.w3(32'h3ab1d52b),
	.w4(32'hba0bf812),
	.w5(32'h3b28d47a),
	.w6(32'h3b32fc33),
	.w7(32'hb81e4784),
	.w8(32'h3b2f1974),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb66714),
	.w1(32'hb96bce41),
	.w2(32'h3b7fb67f),
	.w3(32'h3b6db393),
	.w4(32'hbb12d145),
	.w5(32'h3abc1d29),
	.w6(32'h3b682f01),
	.w7(32'hbad75186),
	.w8(32'h3954c491),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923c397),
	.w1(32'h3a8e7cd5),
	.w2(32'h3970df6c),
	.w3(32'h3994a315),
	.w4(32'h3a9c15d0),
	.w5(32'hb878c3c6),
	.w6(32'h3a24e648),
	.w7(32'h3ade4319),
	.w8(32'h3a92f5dc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e1dbe),
	.w1(32'hba909259),
	.w2(32'hba2e51e6),
	.w3(32'hb97138da),
	.w4(32'hba979766),
	.w5(32'hbaad15d3),
	.w6(32'hba877084),
	.w7(32'hba8ca2d8),
	.w8(32'hba8b8fe0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa31d29),
	.w1(32'hbb58cc79),
	.w2(32'hb9573814),
	.w3(32'hb92555f5),
	.w4(32'hbb8b65c0),
	.w5(32'hbb08e632),
	.w6(32'hbad859da),
	.w7(32'hbb3cf6e9),
	.w8(32'hbb1f85bf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb19fa),
	.w1(32'hbb7c89b5),
	.w2(32'hbb7320ca),
	.w3(32'h3926c7f7),
	.w4(32'hbb331275),
	.w5(32'hbb3e1f44),
	.w6(32'h3993d2ca),
	.w7(32'hbae5318a),
	.w8(32'hba87875b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397d09),
	.w1(32'h39c9c8e4),
	.w2(32'h3b815e00),
	.w3(32'h3b39d7d2),
	.w4(32'h3a2712c0),
	.w5(32'h3b28971f),
	.w6(32'h3b4d694d),
	.w7(32'h36d559b2),
	.w8(32'h3aac9647),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6d51),
	.w1(32'hba235abf),
	.w2(32'hba2511fc),
	.w3(32'h3a9351e3),
	.w4(32'hba09f1a7),
	.w5(32'hba2f6a45),
	.w6(32'hb9ac0ffc),
	.w7(32'hba1c445f),
	.w8(32'hb99b9004),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff8d61),
	.w1(32'hba140eac),
	.w2(32'hba1902ba),
	.w3(32'hb9cf4a24),
	.w4(32'hba11d053),
	.w5(32'hba53285d),
	.w6(32'hba290710),
	.w7(32'hba2a3f38),
	.w8(32'hb9e6ddb0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9152080),
	.w1(32'h39ccfaa0),
	.w2(32'h3b39a893),
	.w3(32'hba4d3eeb),
	.w4(32'hb8aa9093),
	.w5(32'h3ac46c3d),
	.w6(32'hba3b3486),
	.w7(32'hb9c6bca1),
	.w8(32'h39761303),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71b1bc),
	.w1(32'h38948996),
	.w2(32'h3afc5e53),
	.w3(32'hba3e3967),
	.w4(32'hba3da63e),
	.w5(32'h39c37225),
	.w6(32'h3a969644),
	.w7(32'hb9d8af67),
	.w8(32'hb99f1757),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3abb0c),
	.w1(32'hba657bc5),
	.w2(32'hbab86bb0),
	.w3(32'hb838395a),
	.w4(32'hb931a192),
	.w5(32'hba12d67e),
	.w6(32'h385351bb),
	.w7(32'hb9c553c7),
	.w8(32'h3a10ffda),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdb2d6),
	.w1(32'hb98be322),
	.w2(32'h3a10f1e9),
	.w3(32'h396fed95),
	.w4(32'hb9a499f8),
	.w5(32'h38e3a930),
	.w6(32'hba590d50),
	.w7(32'hba116549),
	.w8(32'hb80b305d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30f36a),
	.w1(32'hbaf1cf8c),
	.w2(32'h3b373eb2),
	.w3(32'h3a88c76f),
	.w4(32'hbb2d0c5a),
	.w5(32'h3ac56c56),
	.w6(32'hbaea7483),
	.w7(32'hbba46151),
	.w8(32'h3b430a3e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2686),
	.w1(32'hbb259f4d),
	.w2(32'hb9003d59),
	.w3(32'h3bd02154),
	.w4(32'hbb895a28),
	.w5(32'hba31913b),
	.w6(32'h3bff1b57),
	.w7(32'hbb296b0c),
	.w8(32'h3af0e70c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd021fe),
	.w1(32'hbb8a35d3),
	.w2(32'hbb0466e1),
	.w3(32'h3bd62359),
	.w4(32'hbb95f8d9),
	.w5(32'hbaa1bf97),
	.w6(32'h3be625df),
	.w7(32'hbb0ead82),
	.w8(32'h3ad2585c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef19c8),
	.w1(32'hba53a3a6),
	.w2(32'h3a4b29c0),
	.w3(32'h3a4f8533),
	.w4(32'hbab0908c),
	.w5(32'hba2fb799),
	.w6(32'h3a602d9e),
	.w7(32'hba2a4ef7),
	.w8(32'hb72d55d1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb968bf29),
	.w1(32'h39a66070),
	.w2(32'h3a118aab),
	.w3(32'hb99b187d),
	.w4(32'h3a187158),
	.w5(32'h3a85be80),
	.w6(32'h3973fa41),
	.w7(32'h3a0c8fd8),
	.w8(32'h38235af9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bf99c),
	.w1(32'hb98bb447),
	.w2(32'hb99d4d74),
	.w3(32'h3a8bf4e4),
	.w4(32'hba5eec65),
	.w5(32'hba98956f),
	.w6(32'hb9f171af),
	.w7(32'hba609ab2),
	.w8(32'hba36bdbf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1918bf),
	.w1(32'hb98e25ed),
	.w2(32'hb9794764),
	.w3(32'h3b0913e4),
	.w4(32'h39f55161),
	.w5(32'h3986e896),
	.w6(32'h3a734487),
	.w7(32'h3983dee0),
	.w8(32'h39cd7b29),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7b35d),
	.w1(32'h3bb4c01f),
	.w2(32'h3bcfe1f5),
	.w3(32'h3bedfbc5),
	.w4(32'h3bd9222c),
	.w5(32'h3bae2f50),
	.w6(32'h3c09fd9f),
	.w7(32'h3bbf7dea),
	.w8(32'h3bd2abea),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00ee95),
	.w1(32'h3b4b1260),
	.w2(32'h3ba5b7d7),
	.w3(32'h3bce83f8),
	.w4(32'h3a91d20c),
	.w5(32'h3b36d460),
	.w6(32'h3b733d1b),
	.w7(32'h39357b53),
	.w8(32'h3b13a67c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be78793),
	.w1(32'h3b58a9ce),
	.w2(32'h3bd3c307),
	.w3(32'h3b8ab728),
	.w4(32'h3a21a9e7),
	.w5(32'h3b4d9543),
	.w6(32'h3b9d4a24),
	.w7(32'hba1530cb),
	.w8(32'h3b04eb8f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62fa6f),
	.w1(32'h3b38ed33),
	.w2(32'h3b82afce),
	.w3(32'h3b00823c),
	.w4(32'h3b13c075),
	.w5(32'h3b814409),
	.w6(32'h3bb56f7e),
	.w7(32'h3ada7beb),
	.w8(32'h3b31a66a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40f283),
	.w1(32'h3a660e69),
	.w2(32'h3b833818),
	.w3(32'h3b5d2d83),
	.w4(32'h3b04d20c),
	.w5(32'h3b0bb6be),
	.w6(32'hba92deca),
	.w7(32'h3902cfd9),
	.w8(32'h3b4d9a87),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbd72d),
	.w1(32'hba09e6b9),
	.w2(32'h39881079),
	.w3(32'hb9fd8c40),
	.w4(32'hb979d023),
	.w5(32'hb94706a2),
	.w6(32'hba2a5ed1),
	.w7(32'hb8cf9da5),
	.w8(32'h371e5c6e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a61b3b),
	.w1(32'h3810f80b),
	.w2(32'hb9ee3cb7),
	.w3(32'h39beb6a6),
	.w4(32'hb91eea07),
	.w5(32'hba4661a7),
	.w6(32'hb9aaaa18),
	.w7(32'hba370f05),
	.w8(32'hba2e42be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95559a6),
	.w1(32'h3a6de584),
	.w2(32'hb93ae6d2),
	.w3(32'h39997254),
	.w4(32'h3a85918b),
	.w5(32'h3a206166),
	.w6(32'h3ab7c7ed),
	.w7(32'h39bd2f05),
	.w8(32'hb8b861eb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4aac25),
	.w1(32'h3b3150e6),
	.w2(32'h3b886b07),
	.w3(32'h3b0d47fa),
	.w4(32'hba1326d1),
	.w5(32'h3b16e951),
	.w6(32'h3adc63f9),
	.w7(32'h3aa51091),
	.w8(32'h3a5122ce),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b016940),
	.w1(32'h3a3d0542),
	.w2(32'h3a940da4),
	.w3(32'h3ade4611),
	.w4(32'h3a26abc8),
	.w5(32'h3a189f0a),
	.w6(32'h3a7047cf),
	.w7(32'hb993d79c),
	.w8(32'h3a13d7c4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1c90),
	.w1(32'h3b2bfb29),
	.w2(32'h3bbcbc97),
	.w3(32'h3bad69a1),
	.w4(32'h3b2f4405),
	.w5(32'h3b63018a),
	.w6(32'h3b434c11),
	.w7(32'h3ab99ff5),
	.w8(32'h3b69faf0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918949d),
	.w1(32'hba9450ba),
	.w2(32'h390ceb78),
	.w3(32'h39c704ae),
	.w4(32'hba0472a3),
	.w5(32'hb91ab6f6),
	.w6(32'h39989bd4),
	.w7(32'h39ebaa9e),
	.w8(32'h39d66902),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b851a6),
	.w1(32'hba8c0b3d),
	.w2(32'h3a5b9ec8),
	.w3(32'h3895ecf6),
	.w4(32'hb9335cb4),
	.w5(32'h39b1fb4a),
	.w6(32'hba560f3b),
	.w7(32'hb8c551e4),
	.w8(32'hb987bbbd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b55cb4),
	.w1(32'hbad8dabd),
	.w2(32'hbad9594f),
	.w3(32'h398226c7),
	.w4(32'hba1784cf),
	.w5(32'hbaa775c1),
	.w6(32'hba9f2e64),
	.w7(32'hbae787d2),
	.w8(32'hbaadfdbd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6d885),
	.w1(32'h3a07d32c),
	.w2(32'hbb07eb20),
	.w3(32'hba913b79),
	.w4(32'h3a7ebdd1),
	.w5(32'hbac617e7),
	.w6(32'h3a05f7ba),
	.w7(32'hbb03c04e),
	.w8(32'hba587bb5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b0873),
	.w1(32'hba4c7ecd),
	.w2(32'hb9a7855c),
	.w3(32'hbabd9399),
	.w4(32'hba6642de),
	.w5(32'hb9824a37),
	.w6(32'h398741e9),
	.w7(32'hb7d9108b),
	.w8(32'h3a167c2b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39516eca),
	.w1(32'h3a2bf4b7),
	.w2(32'h3a415e68),
	.w3(32'hb8560bb4),
	.w4(32'h39e592d2),
	.w5(32'h3a0e4ba4),
	.w6(32'hb8219eee),
	.w7(32'h3a5aeaf7),
	.w8(32'h3a065d8e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4827b8),
	.w1(32'h389ff75a),
	.w2(32'h3ae710cf),
	.w3(32'h3b37db0d),
	.w4(32'h39f2e9ec),
	.w5(32'h39a3d3cd),
	.w6(32'h3ab93cb3),
	.w7(32'hb936f696),
	.w8(32'h3a64b1ad),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c1e2),
	.w1(32'hb8f4858c),
	.w2(32'hb9c494de),
	.w3(32'h3a9dd6d7),
	.w4(32'h3a794f25),
	.w5(32'hb8a692cd),
	.w6(32'h3a3545bb),
	.w7(32'h3a28be42),
	.w8(32'h3991b346),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41405a),
	.w1(32'h3adcf948),
	.w2(32'h3a90231b),
	.w3(32'hba15accc),
	.w4(32'h3ac8eb48),
	.w5(32'h3ad94367),
	.w6(32'hb791dfa0),
	.w7(32'h390571fe),
	.w8(32'hba7fb972),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd2dff),
	.w1(32'h3a22ac44),
	.w2(32'h392599b8),
	.w3(32'hba8b073c),
	.w4(32'h3a8be18b),
	.w5(32'h3a82fda8),
	.w6(32'h3a6cd6ac),
	.w7(32'h3a1101f8),
	.w8(32'h3abb4a33),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb7abb),
	.w1(32'hbac2e3fc),
	.w2(32'hb91a004c),
	.w3(32'h3afcc60d),
	.w4(32'hba869766),
	.w5(32'hba36238d),
	.w6(32'hba83a251),
	.w7(32'hba342936),
	.w8(32'hb8f601e7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fbc7f),
	.w1(32'hbab790fe),
	.w2(32'hba722c1a),
	.w3(32'hba94fadd),
	.w4(32'hbad4066a),
	.w5(32'hba8961b4),
	.w6(32'hbae6b9d9),
	.w7(32'hbaf978be),
	.w8(32'hbb187045),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e18b50),
	.w1(32'h3b1fccf6),
	.w2(32'h3ba51c41),
	.w3(32'h3a5ac70c),
	.w4(32'h3b537e77),
	.w5(32'h3b37b002),
	.w6(32'h3b2ae73d),
	.w7(32'h3b59c53d),
	.w8(32'h3b8aecc6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d772),
	.w1(32'h3accc073),
	.w2(32'h3b78a63c),
	.w3(32'h3b9103e3),
	.w4(32'h3aa326eb),
	.w5(32'h3b613399),
	.w6(32'h3b2343d8),
	.w7(32'hb9f9ccd5),
	.w8(32'h3afe3f60),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eb63a),
	.w1(32'hba1a83ea),
	.w2(32'h3ad1e99e),
	.w3(32'h3aa9e56c),
	.w4(32'hbacdb699),
	.w5(32'h3a982a2a),
	.w6(32'h3b686502),
	.w7(32'hb977e058),
	.w8(32'h3aa0ebdd),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb92913),
	.w1(32'hbb58d538),
	.w2(32'h3b982d84),
	.w3(32'h3b40e649),
	.w4(32'hbbd74b1c),
	.w5(32'hb9efe9e0),
	.w6(32'h3b72c8c2),
	.w7(32'hbbd3edf7),
	.w8(32'h3a3c0cf9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba137389),
	.w1(32'hb9a2eed1),
	.w2(32'hb8881de5),
	.w3(32'hba17de40),
	.w4(32'hb9baf5b4),
	.w5(32'hba102caa),
	.w6(32'hb917e3a9),
	.w7(32'hb982a02a),
	.w8(32'hb98f59bc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a70bd0),
	.w1(32'hb9f07f45),
	.w2(32'hb99d09c0),
	.w3(32'hb99046c5),
	.w4(32'hb9859934),
	.w5(32'hba038a30),
	.w6(32'hb9c73d96),
	.w7(32'hba102eea),
	.w8(32'hb9d0c537),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e42e8),
	.w1(32'h39c0ad91),
	.w2(32'h39eefe4f),
	.w3(32'hb93c7eee),
	.w4(32'h398d094a),
	.w5(32'h39915477),
	.w6(32'h383455d8),
	.w7(32'h394d0188),
	.w8(32'h36d9c05e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28c4a3),
	.w1(32'hba4c3f70),
	.w2(32'hb999489a),
	.w3(32'h3a87de86),
	.w4(32'hba4ca7cf),
	.w5(32'hb9fb8a5e),
	.w6(32'hb9e1832c),
	.w7(32'hba4ee7ab),
	.w8(32'hb9520284),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f86bc),
	.w1(32'hbaae8d4b),
	.w2(32'hba2821d6),
	.w3(32'hba08b884),
	.w4(32'hbab34ef1),
	.w5(32'hba8df1d3),
	.w6(32'hba52c016),
	.w7(32'hb9f45274),
	.w8(32'hba03f835),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c36e1),
	.w1(32'h3a8acc4c),
	.w2(32'h3b22fba0),
	.w3(32'h3a7b2e17),
	.w4(32'hb9d23a70),
	.w5(32'h3a9800d3),
	.w6(32'hba2f4a4a),
	.w7(32'h3a4e8762),
	.w8(32'hba0a02c8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae7b1c),
	.w1(32'h3a62ce75),
	.w2(32'h3ad976b3),
	.w3(32'h3b35f4e6),
	.w4(32'h3a4d184e),
	.w5(32'h3a88765e),
	.w6(32'h3b65cc9b),
	.w7(32'h399a80b4),
	.w8(32'h3b1d4917),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74514e),
	.w1(32'h3af5e2de),
	.w2(32'h3b8649b1),
	.w3(32'h3b1ffb34),
	.w4(32'hb8ddbf08),
	.w5(32'h3a9e8e33),
	.w6(32'h3aa0ea11),
	.w7(32'hb6e66b90),
	.w8(32'h3a709b8d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d912f),
	.w1(32'hba86ed85),
	.w2(32'h3a96f72c),
	.w3(32'h3a0564bc),
	.w4(32'hba24fa0c),
	.w5(32'h39eaa147),
	.w6(32'h3a530f5e),
	.w7(32'h39b5fe85),
	.w8(32'h3ac174a1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d265e8),
	.w1(32'hb9a5574e),
	.w2(32'h3a2b5248),
	.w3(32'h3a172149),
	.w4(32'h38e30e22),
	.w5(32'h39f571ad),
	.w6(32'hb9ed7c25),
	.w7(32'hb9288baf),
	.w8(32'h3a60e15f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae02679),
	.w1(32'h3a59e520),
	.w2(32'h39c01c2f),
	.w3(32'h3a76ac82),
	.w4(32'hb9211e23),
	.w5(32'hba6db16a),
	.w6(32'h3a4730a6),
	.w7(32'hba488de9),
	.w8(32'hba676f63),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8ec9b),
	.w1(32'hb9b7c379),
	.w2(32'h3a6e356f),
	.w3(32'h381dac69),
	.w4(32'h39ef5eaa),
	.w5(32'h3aba5874),
	.w6(32'hb7d300ee),
	.w7(32'hb9d9eaf1),
	.w8(32'h3aaf03a6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9497fc1),
	.w1(32'hba850a91),
	.w2(32'hb9079da0),
	.w3(32'h379f6c44),
	.w4(32'hba6da89a),
	.w5(32'hba22315d),
	.w6(32'hba524703),
	.w7(32'hba5e24fc),
	.w8(32'hba69dff8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f4cdf),
	.w1(32'hb89def5b),
	.w2(32'h399738b5),
	.w3(32'hb98538f5),
	.w4(32'hba128250),
	.w5(32'hb9d1f243),
	.w6(32'h394e51aa),
	.w7(32'h39b22b98),
	.w8(32'h3a13bd74),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924fe77),
	.w1(32'h3a1c05b4),
	.w2(32'hb9782347),
	.w3(32'hb990147b),
	.w4(32'h38ec8fb5),
	.w5(32'hb8c7bc3f),
	.w6(32'h39a5c9a9),
	.w7(32'hba074ffb),
	.w8(32'hb998160d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da5a6a),
	.w1(32'hb9357761),
	.w2(32'h39d43f52),
	.w3(32'hba34ec37),
	.w4(32'h37baf588),
	.w5(32'hb8c0323d),
	.w6(32'h38831a78),
	.w7(32'hb9d2ee7f),
	.w8(32'hb8934fce),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad7b3),
	.w1(32'hbae22924),
	.w2(32'h3ae7c78f),
	.w3(32'h3ae107b6),
	.w4(32'hbb54b9cb),
	.w5(32'hb9cd94c2),
	.w6(32'hb9a6569e),
	.w7(32'hbb0008ce),
	.w8(32'hba6c2ab2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf364cb),
	.w1(32'hba88ebb6),
	.w2(32'hba1bb148),
	.w3(32'hbab4e12c),
	.w4(32'hba5c97d6),
	.w5(32'hba4510c4),
	.w6(32'hb95961dc),
	.w7(32'hba1b0875),
	.w8(32'hba11e0c3),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12b107),
	.w1(32'h3a8ac95f),
	.w2(32'h3b27ba68),
	.w3(32'h3a7aff58),
	.w4(32'hb9f4598b),
	.w5(32'h3aa77204),
	.w6(32'h3ac4c0f2),
	.w7(32'h39359b40),
	.w8(32'h3a888f6f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9410f1),
	.w1(32'h3abffeb6),
	.w2(32'h3a24fe2b),
	.w3(32'h3bbb2237),
	.w4(32'h3ac354ef),
	.w5(32'h3a12050c),
	.w6(32'h3ba8575c),
	.w7(32'h3b09de10),
	.w8(32'h3ab8a7bc),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad61b7c),
	.w1(32'hbad7df23),
	.w2(32'hb9356904),
	.w3(32'h3b18adc0),
	.w4(32'hbb03aaec),
	.w5(32'hb9c78b7e),
	.w6(32'h3abe4611),
	.w7(32'hbafc083e),
	.w8(32'h37f014a2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a729c02),
	.w1(32'h3a99dcc3),
	.w2(32'h3b14cc05),
	.w3(32'h3b0d3d18),
	.w4(32'h38a49ee9),
	.w5(32'h3abc58e2),
	.w6(32'h3a7e1499),
	.w7(32'h3a90727f),
	.w8(32'h3b8c1aa6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a883e57),
	.w1(32'hbb10242c),
	.w2(32'hb59b5245),
	.w3(32'h3b1979c3),
	.w4(32'hbb0caa8e),
	.w5(32'hb9a57627),
	.w6(32'hba279cbc),
	.w7(32'hbb167fd7),
	.w8(32'hb9d267fc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ec206),
	.w1(32'h3841e3ff),
	.w2(32'h3ab8f7ef),
	.w3(32'h39c24167),
	.w4(32'hbb062362),
	.w5(32'hba9ac412),
	.w6(32'h3af4883e),
	.w7(32'hbaa3473a),
	.w8(32'h3a4260ba),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392684b0),
	.w1(32'hba0f7ecd),
	.w2(32'h3b04839a),
	.w3(32'hb9a3e4db),
	.w4(32'hbaff54f7),
	.w5(32'hbade363e),
	.w6(32'hb9d68b63),
	.w7(32'hbaee5249),
	.w8(32'hba2490c7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45eff8),
	.w1(32'hb8e28b83),
	.w2(32'h3b70dcf1),
	.w3(32'h3ad3c9c4),
	.w4(32'hbabe9d00),
	.w5(32'h3b30a07a),
	.w6(32'h3b1a39de),
	.w7(32'hba634968),
	.w8(32'h3b10364b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef060f),
	.w1(32'h3a720e16),
	.w2(32'h3b1abe28),
	.w3(32'h3a83e2d3),
	.w4(32'h3a263bcd),
	.w5(32'h3ac13a1f),
	.w6(32'hba254fe5),
	.w7(32'h3af39f7a),
	.w8(32'h39ae28b8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba0e4),
	.w1(32'h3ad78847),
	.w2(32'h3bacbd5b),
	.w3(32'h3b8c1138),
	.w4(32'h3a975468),
	.w5(32'h3b9b44de),
	.w6(32'h3b0dab95),
	.w7(32'h3afa64ab),
	.w8(32'h3b8ed7f7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984ceda),
	.w1(32'hbb0f982b),
	.w2(32'h3aa35d37),
	.w3(32'h3aacd9fc),
	.w4(32'hbb12fe3c),
	.w5(32'hb9213413),
	.w6(32'hbb0cfecf),
	.w7(32'hbaed8550),
	.w8(32'h3aacfc63),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eb6cb),
	.w1(32'hbaa25315),
	.w2(32'h3b7fc730),
	.w3(32'h3a77d0f6),
	.w4(32'hbaf75407),
	.w5(32'h3b574b3c),
	.w6(32'hbaa6af7d),
	.w7(32'hbb499267),
	.w8(32'h3b2e7889),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b753876),
	.w1(32'hbb353958),
	.w2(32'hba2d004c),
	.w3(32'h3abf5651),
	.w4(32'hbba0d8de),
	.w5(32'hbb2be6b2),
	.w6(32'h3b336a49),
	.w7(32'hbbbe9af5),
	.w8(32'h3a15f72c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce0bc3),
	.w1(32'h3bc6bd48),
	.w2(32'h3c0d75a4),
	.w3(32'h3b8f4127),
	.w4(32'h3b3d9601),
	.w5(32'h3b9a0ab5),
	.w6(32'h3bac719a),
	.w7(32'h3a2dc719),
	.w8(32'h3a8326b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118e70),
	.w1(32'h39d0b868),
	.w2(32'h3b1fd6d0),
	.w3(32'h3aee466f),
	.w4(32'hb8ba4dde),
	.w5(32'h3b193859),
	.w6(32'hbb09ecd3),
	.w7(32'hbaa60ba7),
	.w8(32'h3b6dd7b4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0168be),
	.w1(32'h3a35fa35),
	.w2(32'h3a185f9d),
	.w3(32'h3ab6275f),
	.w4(32'h3a9c8b6c),
	.w5(32'h39837d1b),
	.w6(32'h3a5d1d4d),
	.w7(32'h3a051426),
	.w8(32'h382a2c56),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd767a6),
	.w1(32'h3ac7c87d),
	.w2(32'h3bb21341),
	.w3(32'h3b342804),
	.w4(32'h395418ce),
	.w5(32'h3b9b3330),
	.w6(32'hbaac241c),
	.w7(32'hbaa67758),
	.w8(32'h3b08b9c6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7ba03),
	.w1(32'hba73c2ec),
	.w2(32'h3b2e2487),
	.w3(32'h3a4bc886),
	.w4(32'h39018c72),
	.w5(32'h3b0a2537),
	.w6(32'hbae63814),
	.w7(32'hba8a22e5),
	.w8(32'h3a111abd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba945063),
	.w1(32'hba00d411),
	.w2(32'hb993c5ae),
	.w3(32'hba7d1762),
	.w4(32'hba967e86),
	.w5(32'hba4a72fd),
	.w6(32'hb889da4b),
	.w7(32'hba2f7aec),
	.w8(32'hb8b1cf60),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae7b15),
	.w1(32'hb9d3ce82),
	.w2(32'h393c5359),
	.w3(32'hb9a6a3ba),
	.w4(32'hb99d2b89),
	.w5(32'hb87ee232),
	.w6(32'h3899cc65),
	.w7(32'hb9bfd064),
	.w8(32'hb8c46297),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80df47),
	.w1(32'h3b66a1bf),
	.w2(32'h3b7868a0),
	.w3(32'h3b748762),
	.w4(32'h3b2bf067),
	.w5(32'h3b3d2ddc),
	.w6(32'h3b5c1ef4),
	.w7(32'h3b325bff),
	.w8(32'h3b60f923),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb31e2e),
	.w1(32'h3b9f7317),
	.w2(32'h3bd2ce16),
	.w3(32'h3b900818),
	.w4(32'h3b2f0c2b),
	.w5(32'h3b6e2205),
	.w6(32'h3b624973),
	.w7(32'h3aa0e17f),
	.w8(32'h3b0478d4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ed31),
	.w1(32'h3b0435bb),
	.w2(32'h3b641f84),
	.w3(32'h3b5b40d1),
	.w4(32'h3a53efb4),
	.w5(32'h3b0bc089),
	.w6(32'h3aedb744),
	.w7(32'h3ad1fcf3),
	.w8(32'h3b31c94b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe789f),
	.w1(32'h3ab157f1),
	.w2(32'h3a0f4f5a),
	.w3(32'h3afcf7e7),
	.w4(32'h3a9b7fb1),
	.w5(32'h3afd9fd8),
	.w6(32'h38ec816c),
	.w7(32'h396b0667),
	.w8(32'h3aa81800),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1be07b),
	.w1(32'h39c23434),
	.w2(32'h3a7386ed),
	.w3(32'h3aaecfca),
	.w4(32'h38972dac),
	.w5(32'h3ac34900),
	.w6(32'h3b4bf20a),
	.w7(32'h39e940c3),
	.w8(32'h3ae8ebb4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34e58b),
	.w1(32'h3ab6a506),
	.w2(32'h3b196cb9),
	.w3(32'h3b23c943),
	.w4(32'h3a1aaf6a),
	.w5(32'h3a6fd149),
	.w6(32'h3a082063),
	.w7(32'h3a051198),
	.w8(32'h3971d5ce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21dda5),
	.w1(32'hb9d2a141),
	.w2(32'h3a075e46),
	.w3(32'h3b05f859),
	.w4(32'hba4c5b18),
	.w5(32'hba3f8388),
	.w6(32'h39b5dced),
	.w7(32'hba389f18),
	.w8(32'hba145b35),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd14d),
	.w1(32'hb972f281),
	.w2(32'hb9934d1b),
	.w3(32'hbac06107),
	.w4(32'hb8aab4a0),
	.w5(32'hb928ab79),
	.w6(32'hba1e9283),
	.w7(32'hba121592),
	.w8(32'hb9dd7183),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e6385c),
	.w1(32'hb84d5b9f),
	.w2(32'hb7655924),
	.w3(32'h39aedfe4),
	.w4(32'hb86346a4),
	.w5(32'hb9a3a25a),
	.w6(32'h38760094),
	.w7(32'hb7fb7e8f),
	.w8(32'h3887b28a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccd5ff),
	.w1(32'hb9adfade),
	.w2(32'hb99fb90d),
	.w3(32'h3984ea05),
	.w4(32'hb97978d5),
	.w5(32'hb98864a2),
	.w6(32'hb91690f7),
	.w7(32'hb9195ffa),
	.w8(32'h38ee39bf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0d879),
	.w1(32'hba522c79),
	.w2(32'hbaa7e607),
	.w3(32'h39c8f8f8),
	.w4(32'h3979278a),
	.w5(32'h391fb23e),
	.w6(32'hbad75936),
	.w7(32'hbb17a135),
	.w8(32'hba5954a9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fbd09),
	.w1(32'h3ac38784),
	.w2(32'h3b2666f2),
	.w3(32'h3b108635),
	.w4(32'h39dde59d),
	.w5(32'h3968b98e),
	.w6(32'h3b2a29f9),
	.w7(32'hb917cc06),
	.w8(32'hb7ba549f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9484ea),
	.w1(32'hb94a6c2b),
	.w2(32'hb98628e7),
	.w3(32'hba9ec45f),
	.w4(32'hb9f65033),
	.w5(32'hbaa4deaf),
	.w6(32'hb9f277ae),
	.w7(32'hbaddf6d7),
	.w8(32'hbaa2c34a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4d4cc),
	.w1(32'h39c162a5),
	.w2(32'h3a6c7ce6),
	.w3(32'hb98fcec0),
	.w4(32'h39ac047d),
	.w5(32'h3a419258),
	.w6(32'hba6765fb),
	.w7(32'hb904dbfa),
	.w8(32'h3aaf214f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56856c),
	.w1(32'h3a847e07),
	.w2(32'h3adb5c82),
	.w3(32'h3b3953c0),
	.w4(32'hba40e50b),
	.w5(32'h3a3cf3e5),
	.w6(32'h3b428c51),
	.w7(32'hb899af92),
	.w8(32'h3acacb54),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ae5c6),
	.w1(32'h3b075d25),
	.w2(32'h3a8c6edb),
	.w3(32'h3931e1f2),
	.w4(32'h3aca14cb),
	.w5(32'h3a7624bb),
	.w6(32'h3ab848c3),
	.w7(32'h3a277e99),
	.w8(32'h3a43bd4d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9014c6),
	.w1(32'h3995dcab),
	.w2(32'h3a217866),
	.w3(32'h3aba91dd),
	.w4(32'h39e3dd30),
	.w5(32'h39951ac6),
	.w6(32'h3aa07eea),
	.w7(32'h3a730247),
	.w8(32'h39e2845a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39204c30),
	.w1(32'hbaaf73f9),
	.w2(32'hba82f2c9),
	.w3(32'h3a1eca4a),
	.w4(32'hba8c8e43),
	.w5(32'hba8de4db),
	.w6(32'hba7fb9b3),
	.w7(32'hba9a37e2),
	.w8(32'hba74d7a8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba022b03),
	.w1(32'hb9aaab8d),
	.w2(32'hba8abfe8),
	.w3(32'hb97cf40b),
	.w4(32'h39d0a12d),
	.w5(32'hb7906465),
	.w6(32'h3a4e7215),
	.w7(32'h39dc4c5f),
	.w8(32'h3810e6d6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fa8e7),
	.w1(32'h3a96b981),
	.w2(32'h3a882d46),
	.w3(32'hb9ccb1bc),
	.w4(32'h3a42e001),
	.w5(32'h3ad2ff2d),
	.w6(32'h3a8bf3e0),
	.w7(32'h3a1b1f62),
	.w8(32'h3a0e3f35),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efc52),
	.w1(32'h3a80cfeb),
	.w2(32'h3b99e6ac),
	.w3(32'h3ad3d3ed),
	.w4(32'hb90cefcf),
	.w5(32'h39db4adf),
	.w6(32'h3adb4d1f),
	.w7(32'h39921ffb),
	.w8(32'h3b35953e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a02dec),
	.w1(32'h3a25580f),
	.w2(32'h3ad5c9e2),
	.w3(32'hba7df734),
	.w4(32'hb94deaac),
	.w5(32'h3a3d4c49),
	.w6(32'hb82b4abd),
	.w7(32'h3a1c325d),
	.w8(32'h39703b22),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accc8ec),
	.w1(32'hb8a70c87),
	.w2(32'h3a75ab22),
	.w3(32'h3b11ec52),
	.w4(32'h3910a1d5),
	.w5(32'h3a9d9055),
	.w6(32'h39ca6b63),
	.w7(32'hb9a493cc),
	.w8(32'h398cadbe),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55c8ce),
	.w1(32'h3a7e4254),
	.w2(32'h3b0b9733),
	.w3(32'h3a8c054e),
	.w4(32'hba3beb6f),
	.w5(32'h3a1476a3),
	.w6(32'h3a17ad87),
	.w7(32'h39ccdc53),
	.w8(32'hba0b3f96),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b2caa),
	.w1(32'h3a45b2c6),
	.w2(32'h3a21a525),
	.w3(32'hba3ed671),
	.w4(32'h39501282),
	.w5(32'hb9a9d154),
	.w6(32'h3a896dbe),
	.w7(32'h39e617e4),
	.w8(32'hb92cef02),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5a04),
	.w1(32'h3abc1548),
	.w2(32'h3b379979),
	.w3(32'h3958c2f9),
	.w4(32'hb9bfbe12),
	.w5(32'hb91c0039),
	.w6(32'h3ac17b33),
	.w7(32'h3a991fcc),
	.w8(32'h38b9c3a0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5dd0),
	.w1(32'h3b13bb14),
	.w2(32'h3ba6b177),
	.w3(32'h3a464a19),
	.w4(32'h3aed2bbe),
	.w5(32'h3b8afaef),
	.w6(32'h3af0a590),
	.w7(32'h3b06b2b9),
	.w8(32'h3b70a732),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bb085),
	.w1(32'h39a08722),
	.w2(32'h371f35b7),
	.w3(32'h3afc71b9),
	.w4(32'hba3e5ef0),
	.w5(32'hb972cfbf),
	.w6(32'h3b2f4ea6),
	.w7(32'hb8968a24),
	.w8(32'h3a0cf14e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f8ef),
	.w1(32'h3adbbe17),
	.w2(32'h3b14dd27),
	.w3(32'hb85e373f),
	.w4(32'hba432d6e),
	.w5(32'h3a7d5f3b),
	.w6(32'hb6d88122),
	.w7(32'hb7e601d3),
	.w8(32'h3a9f05a9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af550d5),
	.w1(32'h3a97a01b),
	.w2(32'h3b449522),
	.w3(32'h3a7dfd73),
	.w4(32'hb8e602dc),
	.w5(32'h3adf800d),
	.w6(32'h3ad6d050),
	.w7(32'h3aac9e1d),
	.w8(32'h3a0148fd),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2deeb),
	.w1(32'hbafd00fe),
	.w2(32'hb9e4499a),
	.w3(32'hba4d3a8f),
	.w4(32'hbb0ed138),
	.w5(32'hba04601b),
	.w6(32'hb81b52b0),
	.w7(32'hba61ecad),
	.w8(32'h3ab14488),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a8d4),
	.w1(32'h3a408fcd),
	.w2(32'h3a6c9996),
	.w3(32'h3b1a763e),
	.w4(32'h39fe963d),
	.w5(32'h3a24db3a),
	.w6(32'h3ad9162f),
	.w7(32'h3a855e4d),
	.w8(32'h3ad5b928),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a22cc8),
	.w1(32'hb9d07539),
	.w2(32'hb9bb92b5),
	.w3(32'hba07d846),
	.w4(32'hb9c83c91),
	.w5(32'hb9c060c9),
	.w6(32'h39da4496),
	.w7(32'hba56a59b),
	.w8(32'hb8511946),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86748e),
	.w1(32'hba807980),
	.w2(32'h3abd4061),
	.w3(32'h3b67ca15),
	.w4(32'hbaca600d),
	.w5(32'h3ac6c736),
	.w6(32'h3b9c1d95),
	.w7(32'hb9cd648a),
	.w8(32'h3b088a10),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e663e0),
	.w1(32'hbb1bd084),
	.w2(32'hbad0f2d8),
	.w3(32'h399b7855),
	.w4(32'hbaf25344),
	.w5(32'hbac95ebc),
	.w6(32'hb98b628f),
	.w7(32'hbaad3879),
	.w8(32'h3a500ef7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4776a2),
	.w1(32'h38139067),
	.w2(32'h38a7c76c),
	.w3(32'hbb0fdd84),
	.w4(32'h38de7e7a),
	.w5(32'h39fd1c8f),
	.w6(32'h39c35dd1),
	.w7(32'h3a19eee3),
	.w8(32'hb9046d33),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1aec29),
	.w1(32'h3b7f9cd5),
	.w2(32'h3c07445b),
	.w3(32'hb9f6caf2),
	.w4(32'h3b4cec6e),
	.w5(32'h3beaa1d1),
	.w6(32'h3b2938c4),
	.w7(32'h3ba9725c),
	.w8(32'h3714a947),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa46ee),
	.w1(32'h38b2743c),
	.w2(32'h3aa0b78a),
	.w3(32'h3b7abb65),
	.w4(32'hbabd379b),
	.w5(32'hba89000d),
	.w6(32'h3a3d5d08),
	.w7(32'h39a7010b),
	.w8(32'hb9be10ce),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f762e),
	.w1(32'h39a597c0),
	.w2(32'h3b5d138c),
	.w3(32'hb9c99974),
	.w4(32'hbb11a91c),
	.w5(32'h3ad5cc0f),
	.w6(32'hb93e573e),
	.w7(32'hbac86bb0),
	.w8(32'h3a7b61a5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58a692),
	.w1(32'h39f8d9c1),
	.w2(32'h3b3c0416),
	.w3(32'h3b504ffd),
	.w4(32'hb9cf5fb5),
	.w5(32'h3abcd957),
	.w6(32'h3b29cff2),
	.w7(32'hb8d58748),
	.w8(32'h3b226fb0),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bb6d0),
	.w1(32'hb946b12a),
	.w2(32'hbad59150),
	.w3(32'hba59c6a9),
	.w4(32'h3a48784a),
	.w5(32'h39be8375),
	.w6(32'h3af60849),
	.w7(32'h3a48fac5),
	.w8(32'hb911a75c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b048a24),
	.w1(32'h3ae17e5a),
	.w2(32'h3bd35b38),
	.w3(32'h3ab74ff5),
	.w4(32'h3a74989b),
	.w5(32'h3b61f688),
	.w6(32'h3b0ad37f),
	.w7(32'h3873c50b),
	.w8(32'h3abaee2c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b743c12),
	.w1(32'h3bbae5b7),
	.w2(32'h3be064bd),
	.w3(32'h3ba39600),
	.w4(32'h3a97556c),
	.w5(32'h3b3a75e4),
	.w6(32'h3baaff05),
	.w7(32'h3bc3c313),
	.w8(32'h3adc2da9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae75b8),
	.w1(32'h3aaccb06),
	.w2(32'h3b15d294),
	.w3(32'hbb414ae5),
	.w4(32'h3a503a06),
	.w5(32'h3aff5a17),
	.w6(32'hba1de4f6),
	.w7(32'h39e1236f),
	.w8(32'h3af831a7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95705f3),
	.w1(32'hba86f1df),
	.w2(32'h3b96c9cd),
	.w3(32'hba376ea7),
	.w4(32'hbaeb743d),
	.w5(32'h3b75f1c9),
	.w6(32'h39b1e7d1),
	.w7(32'hbac9730a),
	.w8(32'h39ee45cd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87623f),
	.w1(32'h3aea3755),
	.w2(32'h3b9a784b),
	.w3(32'h3acce0cf),
	.w4(32'h39cf4ac5),
	.w5(32'h3b50f87f),
	.w6(32'h3a8337ed),
	.w7(32'h3aac8591),
	.w8(32'h3a8b1ecd),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7649a9),
	.w1(32'h389af543),
	.w2(32'hb83d5499),
	.w3(32'h3b2a45ae),
	.w4(32'h3a8a10ea),
	.w5(32'h3a956938),
	.w6(32'h3acbb29a),
	.w7(32'h3ade8441),
	.w8(32'h3a9bdb65),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b30a2),
	.w1(32'hbb28d205),
	.w2(32'hbab95d12),
	.w3(32'hb9732853),
	.w4(32'hbb826aa4),
	.w5(32'hbb28f997),
	.w6(32'h38b359cd),
	.w7(32'hbb5ca7eb),
	.w8(32'hbb2df73a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03acf4),
	.w1(32'hb9656adf),
	.w2(32'h3a8fd9b1),
	.w3(32'h39f49c3f),
	.w4(32'hb9d4c467),
	.w5(32'h3b65da3b),
	.w6(32'h3b879d58),
	.w7(32'h3aeb6106),
	.w8(32'h3b52c22a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c007e),
	.w1(32'h3b6fe404),
	.w2(32'h3bce2fb9),
	.w3(32'h3ae2bcde),
	.w4(32'h3b221b58),
	.w5(32'h3bc93c0d),
	.w6(32'h3b22c612),
	.w7(32'h3a4d2937),
	.w8(32'hba965185),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e3867),
	.w1(32'hb79c5138),
	.w2(32'hb9ee44f3),
	.w3(32'h3ba456e0),
	.w4(32'h3a61eb97),
	.w5(32'h3a3d0778),
	.w6(32'h3a657a57),
	.w7(32'h3a00200a),
	.w8(32'h39e4a1c8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e2dd3),
	.w1(32'hba8d44eb),
	.w2(32'hbaaddd4a),
	.w3(32'hb9eb7fd8),
	.w4(32'hba1d656b),
	.w5(32'hba4d121a),
	.w6(32'h392a1013),
	.w7(32'hb96e1800),
	.w8(32'hb97d5404),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a853daf),
	.w1(32'h3aaed84f),
	.w2(32'h3b5dfe8b),
	.w3(32'hb8f35d08),
	.w4(32'h3a5c1c91),
	.w5(32'h3b0020cd),
	.w6(32'h3af76d88),
	.w7(32'h3abb6247),
	.w8(32'h3aa4c4c7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9b39),
	.w1(32'hba8112e5),
	.w2(32'hbb199fe3),
	.w3(32'h39816995),
	.w4(32'hba7c3ede),
	.w5(32'hbad5d768),
	.w6(32'hba8c5913),
	.w7(32'hbb173abc),
	.w8(32'hbab98fdf),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab0e5e),
	.w1(32'hb99134a4),
	.w2(32'h3a96a818),
	.w3(32'hbaf7d10c),
	.w4(32'hbad65bce),
	.w5(32'hba7850b2),
	.w6(32'h3a2e3ddd),
	.w7(32'hb9feed63),
	.w8(32'hbab4a95b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bd8b8),
	.w1(32'hba0402a1),
	.w2(32'hba480c7f),
	.w3(32'hbb0de51a),
	.w4(32'hb9f40792),
	.w5(32'hb9219997),
	.w6(32'h3a108d05),
	.w7(32'h3a27eb6e),
	.w8(32'h3a0c0629),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024cb9),
	.w1(32'hbb09cc2b),
	.w2(32'h39875cb3),
	.w3(32'h3a1e8289),
	.w4(32'hbad430d0),
	.w5(32'hb9e006de),
	.w6(32'hb94c942b),
	.w7(32'hb9e9cc9e),
	.w8(32'h39c9184e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf6926),
	.w1(32'h3aa28ab3),
	.w2(32'h3b1c17bd),
	.w3(32'hba013f5e),
	.w4(32'h3a3e9895),
	.w5(32'h3aedc6c5),
	.w6(32'h3a01b0dd),
	.w7(32'h3aa31750),
	.w8(32'h39006281),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91889a),
	.w1(32'hb7e4d06a),
	.w2(32'hba05231a),
	.w3(32'h3a8c8166),
	.w4(32'h38e53cff),
	.w5(32'hb755b2d6),
	.w6(32'h3a45c4e9),
	.w7(32'h3a0d94a9),
	.w8(32'h39a5e00a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68441a),
	.w1(32'h3915d2ab),
	.w2(32'h3adf4abf),
	.w3(32'hb7bffa6b),
	.w4(32'hba1e525a),
	.w5(32'h3a5e9e5c),
	.w6(32'h3a823ad5),
	.w7(32'h3a22fd64),
	.w8(32'h3accf183),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be66e8b),
	.w1(32'h3b891b1c),
	.w2(32'h3c13738a),
	.w3(32'h3bb34170),
	.w4(32'h3b94b069),
	.w5(32'h3c48c51d),
	.w6(32'h3b7b0332),
	.w7(32'h3b82709a),
	.w8(32'h3aad51f6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2efe1e),
	.w1(32'hbafbbe34),
	.w2(32'hbaf4de77),
	.w3(32'h3ba7c754),
	.w4(32'hbaab65ac),
	.w5(32'hba9de36c),
	.w6(32'h3abbe49c),
	.w7(32'hba0a2e72),
	.w8(32'hba65ee15),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676819),
	.w1(32'h3a8ee27e),
	.w2(32'h3b382146),
	.w3(32'h3b170b15),
	.w4(32'h3954a5e4),
	.w5(32'h3ae34a92),
	.w6(32'h3ac4c773),
	.w7(32'h3986545a),
	.w8(32'h3a31e8a6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9c781),
	.w1(32'h3a827b7c),
	.w2(32'h3b257d72),
	.w3(32'hba693cfb),
	.w4(32'hba7e242e),
	.w5(32'h3a2e57dc),
	.w6(32'h3b4ea231),
	.w7(32'h3b5bb143),
	.w8(32'hba568900),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7137b0),
	.w1(32'h3aa262ce),
	.w2(32'h3bd99964),
	.w3(32'h3aa5168c),
	.w4(32'h3a587ec1),
	.w5(32'h3b7d86aa),
	.w6(32'h3b98a1b6),
	.w7(32'hb98bb812),
	.w8(32'h3b15709a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3f5a6),
	.w1(32'hbac11cdf),
	.w2(32'h3a4c8db7),
	.w3(32'h3a10b6f2),
	.w4(32'hbb084817),
	.w5(32'hba00f98d),
	.w6(32'h3953e953),
	.w7(32'hbb35234d),
	.w8(32'hbaa22ff4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b035faf),
	.w1(32'h3ad2eb33),
	.w2(32'h3b02f4dc),
	.w3(32'h3aecd22f),
	.w4(32'h3b3d4a80),
	.w5(32'h3b79d4ac),
	.w6(32'h3aef89b8),
	.w7(32'h3a9b0f03),
	.w8(32'h3b0b70cc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba624e91),
	.w1(32'h3b0f7529),
	.w2(32'h3b546bec),
	.w3(32'hba01d2b9),
	.w4(32'h3b4b18d5),
	.w5(32'h3b93f4d1),
	.w6(32'h3b15c8c2),
	.w7(32'h3b9376e4),
	.w8(32'h39206153),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02ce96),
	.w1(32'hba2688c3),
	.w2(32'h3ad4de76),
	.w3(32'hb8ee5e47),
	.w4(32'hbabe513e),
	.w5(32'h39699183),
	.w6(32'hba3ccfce),
	.w7(32'hba838c4b),
	.w8(32'hba8c7558),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf2469),
	.w1(32'h398c804a),
	.w2(32'hba000e9a),
	.w3(32'hbab2ef6e),
	.w4(32'h3a04717c),
	.w5(32'h38eeb48e),
	.w6(32'h3a9300ff),
	.w7(32'h3a074709),
	.w8(32'h3a1cb65b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5214e),
	.w1(32'hba19e053),
	.w2(32'h38d530f2),
	.w3(32'h3a0a35ed),
	.w4(32'hba5ed3f8),
	.w5(32'hb7e8955d),
	.w6(32'h399b894e),
	.w7(32'h399d9c39),
	.w8(32'h39e25d39),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83d052),
	.w1(32'hba0511c6),
	.w2(32'hbb714bfc),
	.w3(32'hba96cc04),
	.w4(32'hba490942),
	.w5(32'hba944ebd),
	.w6(32'h39bb883a),
	.w7(32'hbaadbb94),
	.w8(32'hba17ea6e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d3ab9),
	.w1(32'h3b16f096),
	.w2(32'h3bd16039),
	.w3(32'h39dac801),
	.w4(32'h3a610d8d),
	.w5(32'h3b85dc52),
	.w6(32'h3b70aaf9),
	.w7(32'h3b88a792),
	.w8(32'h3b3c9046),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b944),
	.w1(32'hb986bf28),
	.w2(32'h39204afa),
	.w3(32'h3a4c0c50),
	.w4(32'hb9fa8b72),
	.w5(32'hb9c530f3),
	.w6(32'h395e0098),
	.w7(32'h3a5088bc),
	.w8(32'h38cba61c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966eea7),
	.w1(32'h39d0ee6b),
	.w2(32'h3b6d5d05),
	.w3(32'hb9f287a0),
	.w4(32'hb7e22312),
	.w5(32'h3b32c273),
	.w6(32'hb9f59aaa),
	.w7(32'h3b0dab78),
	.w8(32'hba2d5049),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b427c),
	.w1(32'h3b0a47fa),
	.w2(32'h3b04fc49),
	.w3(32'h3ac59229),
	.w4(32'h3b6e98e7),
	.w5(32'h3ba370cb),
	.w6(32'h3b973ea7),
	.w7(32'h3b4942b5),
	.w8(32'h3b31d39c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8130fc),
	.w1(32'hba4fe85e),
	.w2(32'h3afddcf4),
	.w3(32'h3bc5f1ff),
	.w4(32'hba932c75),
	.w5(32'h3acfdb2f),
	.w6(32'h3a18dc18),
	.w7(32'h3adf1f44),
	.w8(32'h3a491c2e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd563a),
	.w1(32'hb804d6ae),
	.w2(32'h3a127ff1),
	.w3(32'h3b40f4ca),
	.w4(32'h39cbf811),
	.w5(32'h3a5f2289),
	.w6(32'hb8829c3b),
	.w7(32'hba059b0b),
	.w8(32'h3a72ed46),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39c62b),
	.w1(32'h39f72bd0),
	.w2(32'h3a2d0ddb),
	.w3(32'hba07a68b),
	.w4(32'h3885aac1),
	.w5(32'h394e175c),
	.w6(32'h3a1ae5ac),
	.w7(32'hba0ea7cb),
	.w8(32'hba9a10a3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff7590),
	.w1(32'h3bb3538a),
	.w2(32'h3c36eda6),
	.w3(32'h3bf52146),
	.w4(32'h3b9fde3a),
	.w5(32'h3bdc2b92),
	.w6(32'h3b9fdb19),
	.w7(32'h3aa5993a),
	.w8(32'h3b18d91f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848dec),
	.w1(32'hb9a3605d),
	.w2(32'h3b523e51),
	.w3(32'h3acab209),
	.w4(32'hbb39360c),
	.w5(32'hba6aeb0a),
	.w6(32'h3a2748ac),
	.w7(32'hbb93e030),
	.w8(32'hbb055a79),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb4564),
	.w1(32'hb98b785c),
	.w2(32'hb9bee913),
	.w3(32'h39ea3e50),
	.w4(32'h3ab09e31),
	.w5(32'h3aa128ca),
	.w6(32'h3a44eb1f),
	.w7(32'h3a7fb008),
	.w8(32'h3ad03764),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6daea),
	.w1(32'h3a5d2c51),
	.w2(32'h391e9ee0),
	.w3(32'h3a1f86b4),
	.w4(32'hba185556),
	.w5(32'hbaf0dc0f),
	.w6(32'h3a882123),
	.w7(32'hbadc7bfd),
	.w8(32'hbaaa12c4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f6ee2),
	.w1(32'h3a48aea2),
	.w2(32'h3aa311d5),
	.w3(32'h3a2dd244),
	.w4(32'hba0fe2a9),
	.w5(32'h38907b95),
	.w6(32'h3ad6425a),
	.w7(32'h3af62a14),
	.w8(32'hba721e6b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba874c98),
	.w1(32'hba1b0bd3),
	.w2(32'hba398ff8),
	.w3(32'hbaed062a),
	.w4(32'hba53e98f),
	.w5(32'hbaa19a2b),
	.w6(32'hba6daa8e),
	.w7(32'hba69b97b),
	.w8(32'hba8fdfd1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abbce),
	.w1(32'hb95f42aa),
	.w2(32'h3a2cbe94),
	.w3(32'hba6e535f),
	.w4(32'h39dcb6d8),
	.w5(32'h3b0177d6),
	.w6(32'hb9ad2ead),
	.w7(32'h3a80a41d),
	.w8(32'h3a22615f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1060b),
	.w1(32'h3b7d23d3),
	.w2(32'h3be64f1d),
	.w3(32'h3ac1e9e6),
	.w4(32'h3b210920),
	.w5(32'h3bc29860),
	.w6(32'h39de2277),
	.w7(32'h3a6ccaf2),
	.w8(32'h3a9ee334),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f88ac),
	.w1(32'h3ba5980d),
	.w2(32'h3c39e422),
	.w3(32'h3c037f85),
	.w4(32'h3b24ecb4),
	.w5(32'h3c3159d6),
	.w6(32'h3bf00d20),
	.w7(32'h3c238bff),
	.w8(32'h3afef745),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ade679),
	.w1(32'hb9be67ed),
	.w2(32'hb7e42a40),
	.w3(32'hb9a77a66),
	.w4(32'hb9a70f14),
	.w5(32'h394614d1),
	.w6(32'h3a8b8db5),
	.w7(32'h3a343b2b),
	.w8(32'h39ba17b2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801342),
	.w1(32'h3b210eb8),
	.w2(32'h3b2a98d7),
	.w3(32'h3b28f10c),
	.w4(32'h3af2ca3b),
	.w5(32'h3af1e0ba),
	.w6(32'h3b2c9b2d),
	.w7(32'h3aa573f8),
	.w8(32'h3b3bacc7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f8e13),
	.w1(32'hb9d0f69c),
	.w2(32'h3a9a622c),
	.w3(32'hb92b49fb),
	.w4(32'hba8834fd),
	.w5(32'h39c1c593),
	.w6(32'h38e3f7a4),
	.w7(32'h39ab2a24),
	.w8(32'hb9021c0e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d937dc),
	.w1(32'h3814d467),
	.w2(32'hb9afb882),
	.w3(32'hba4226f0),
	.w4(32'hb96cc385),
	.w5(32'hb9bc427a),
	.w6(32'h3a0365c5),
	.w7(32'h3995873f),
	.w8(32'hb91000b8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0edbf7),
	.w1(32'h39e92779),
	.w2(32'hb9850add),
	.w3(32'hb78fc9da),
	.w4(32'h397ef2e4),
	.w5(32'hb9ed588c),
	.w6(32'h3a70e5ed),
	.w7(32'h39870fce),
	.w8(32'hb961254e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d6843),
	.w1(32'hbab533dd),
	.w2(32'hbad873ec),
	.w3(32'hb9fdd4b0),
	.w4(32'hba490eb3),
	.w5(32'hba2c6bac),
	.w6(32'h392fab08),
	.w7(32'h3893070f),
	.w8(32'hb996e154),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e354),
	.w1(32'hba2085eb),
	.w2(32'h3a6aefc2),
	.w3(32'h393a7df4),
	.w4(32'hbabe2d68),
	.w5(32'h38bce2da),
	.w6(32'h3aa0eecf),
	.w7(32'hb9e75fb4),
	.w8(32'h395f122e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd914d),
	.w1(32'hbbadaf86),
	.w2(32'hbb64b3f1),
	.w3(32'h38b0e8cc),
	.w4(32'hbbb497a7),
	.w5(32'hbaf3381b),
	.w6(32'h39a47c4b),
	.w7(32'hbb4953fa),
	.w8(32'hba0a3ca2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af58b33),
	.w1(32'h3a0ba52e),
	.w2(32'h3abd28f1),
	.w3(32'h3a893396),
	.w4(32'hb9b50ba7),
	.w5(32'h3a79ea37),
	.w6(32'h3b8acfd1),
	.w7(32'h3b0521c2),
	.w8(32'h3aea819f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d6e1),
	.w1(32'hb9fff6bd),
	.w2(32'hba1d9e16),
	.w3(32'hba8d9e53),
	.w4(32'hba0020cd),
	.w5(32'hba0904d3),
	.w6(32'h39b9b351),
	.w7(32'hbababa1d),
	.w8(32'hbac95a4c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7795f1),
	.w1(32'h3a9753b6),
	.w2(32'h3c23115e),
	.w3(32'h3ae0a37f),
	.w4(32'hbaa79d99),
	.w5(32'h3bc2c5b8),
	.w6(32'h3af02cd5),
	.w7(32'h3bbc7368),
	.w8(32'h3ad0406d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fc4a2),
	.w1(32'h3ad12d6b),
	.w2(32'h3aa1f0e6),
	.w3(32'h3b27920c),
	.w4(32'h3ac673b5),
	.w5(32'h3a98d429),
	.w6(32'h3b5994a2),
	.w7(32'h3a953dee),
	.w8(32'h3a112b0b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b700a3c),
	.w1(32'h3b318d88),
	.w2(32'h3bf90709),
	.w3(32'h3b4ac402),
	.w4(32'h3b618a6d),
	.w5(32'h3c17c43f),
	.w6(32'h3bbd7747),
	.w7(32'h3bc2d727),
	.w8(32'h3b5e65fb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecd7ae),
	.w1(32'h389633bb),
	.w2(32'h39ec6e87),
	.w3(32'h39d1d7d1),
	.w4(32'hb937c239),
	.w5(32'h38eac67d),
	.w6(32'hba402d16),
	.w7(32'hba6290ff),
	.w8(32'hba777a51),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92192be),
	.w1(32'h3a8c3992),
	.w2(32'h3b18d6f5),
	.w3(32'hb8dac8e6),
	.w4(32'h3acf1f2c),
	.w5(32'h3b5c8007),
	.w6(32'h3ab09ff7),
	.w7(32'h3b29c54c),
	.w8(32'h3a925510),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a1cc),
	.w1(32'h3a8b645f),
	.w2(32'h3b482815),
	.w3(32'h3b5ea118),
	.w4(32'hb882a8ea),
	.w5(32'h3b14ceb7),
	.w6(32'h3af09684),
	.w7(32'hba77636e),
	.w8(32'h3a47f57a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93420a),
	.w1(32'h3abfb5e9),
	.w2(32'h3b99cb54),
	.w3(32'h3b36d615),
	.w4(32'hb9ae7446),
	.w5(32'h3b8797bc),
	.w6(32'h3a0f9362),
	.w7(32'h3a6ed619),
	.w8(32'h39f5bb29),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e4e4f),
	.w1(32'h3b81ce92),
	.w2(32'h3bdff8b4),
	.w3(32'h3a3a04ed),
	.w4(32'h3b01edef),
	.w5(32'h3b8f73dd),
	.w6(32'h3b86b998),
	.w7(32'h3a9c09da),
	.w8(32'h3ae33863),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b88bc),
	.w1(32'hba3fdf8f),
	.w2(32'hbaffbf09),
	.w3(32'h3b992857),
	.w4(32'h3a95a692),
	.w5(32'hba923bfc),
	.w6(32'hb9c342d3),
	.w7(32'h3a449f04),
	.w8(32'h39deb151),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa82d8b),
	.w1(32'hb9aec983),
	.w2(32'hba6e522f),
	.w3(32'hba596dcb),
	.w4(32'h39e0c20d),
	.w5(32'h394a5c6f),
	.w6(32'h3a57e97d),
	.w7(32'h39e9e41b),
	.w8(32'h39023ba7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ea135),
	.w1(32'h3a4a01b7),
	.w2(32'h3b36dee5),
	.w3(32'hb891a9c9),
	.w4(32'h39fae042),
	.w5(32'h3b0d9f48),
	.w6(32'hb9456052),
	.w7(32'h3a9a1589),
	.w8(32'hba7c1c42),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96b253),
	.w1(32'hb9f9c3bf),
	.w2(32'h3ab93791),
	.w3(32'h3af0cc58),
	.w4(32'h3b24f78e),
	.w5(32'h3ba24619),
	.w6(32'h3a3c2950),
	.w7(32'h3a8d7f1e),
	.w8(32'h3b6e1411),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83f57b),
	.w1(32'h3b1b21d9),
	.w2(32'h3b88bb56),
	.w3(32'h3b871235),
	.w4(32'h3b3fa002),
	.w5(32'h3b97e115),
	.w6(32'h3b95d1a8),
	.w7(32'h3b03a94e),
	.w8(32'h3b965eb0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39005aa8),
	.w1(32'h3a864e41),
	.w2(32'h3b856c03),
	.w3(32'h397966fd),
	.w4(32'h3a233eb5),
	.w5(32'h3b5b0aa2),
	.w6(32'h38a5986f),
	.w7(32'h3adb8145),
	.w8(32'h3b2c6506),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4d1d7),
	.w1(32'hbaa37922),
	.w2(32'h3b2ccca0),
	.w3(32'h3ac0b20f),
	.w4(32'hbaf02834),
	.w5(32'h3aac256f),
	.w6(32'h3b3043b1),
	.w7(32'h3a738a8e),
	.w8(32'h3a556ddc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb23795),
	.w1(32'h3af5e655),
	.w2(32'h3b33c243),
	.w3(32'h3b647000),
	.w4(32'h3ae41afd),
	.w5(32'h3b977ab5),
	.w6(32'h3bdc1e1d),
	.w7(32'h3b6bf90e),
	.w8(32'h3a380dcd),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023af2),
	.w1(32'h39bd51d3),
	.w2(32'h3a44563a),
	.w3(32'h3988f86b),
	.w4(32'hba084a80),
	.w5(32'hb922c54b),
	.w6(32'hba9382ce),
	.w7(32'hba99c8b5),
	.w8(32'hba739a79),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eac448),
	.w1(32'hba0773fd),
	.w2(32'h375c17b8),
	.w3(32'h390b0d7e),
	.w4(32'hb847558f),
	.w5(32'hb9d82f75),
	.w6(32'h3aac138b),
	.w7(32'h3a320ee8),
	.w8(32'h388c78af),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ee305),
	.w1(32'h3a564b2c),
	.w2(32'h3b6f34f2),
	.w3(32'hb9e9572d),
	.w4(32'hbb179626),
	.w5(32'h3ac8760c),
	.w6(32'h3a9aff8b),
	.w7(32'h3b8ef0a8),
	.w8(32'h3907fa78),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c34282),
	.w1(32'hba1949f9),
	.w2(32'hbaa6d1d9),
	.w3(32'hbb6104dd),
	.w4(32'hbaa6c837),
	.w5(32'hbada48d9),
	.w6(32'hb9d5b05c),
	.w7(32'hba014ecb),
	.w8(32'hba937ed8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75cb1),
	.w1(32'hb9a02eb8),
	.w2(32'h3a33f9e4),
	.w3(32'hbb001fdc),
	.w4(32'hb954c2ca),
	.w5(32'h3a3c1585),
	.w6(32'hbae86c3c),
	.w7(32'hba2b0999),
	.w8(32'hba2b3022),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b693492),
	.w1(32'h3afb248f),
	.w2(32'h3b830c0b),
	.w3(32'h3af01c4d),
	.w4(32'h3a1de649),
	.w5(32'h3b7c034c),
	.w6(32'h3b0954d7),
	.w7(32'h3b0ddb4f),
	.w8(32'h3a776148),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fd5ce),
	.w1(32'hb9d68d02),
	.w2(32'h3a8f8df4),
	.w3(32'h3b1d92e9),
	.w4(32'hbb0f94de),
	.w5(32'hb85c8ecd),
	.w6(32'hba0f1cb6),
	.w7(32'h3aca316c),
	.w8(32'h3adb3ba6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391910d2),
	.w1(32'hbb03f116),
	.w2(32'hbb13c2ae),
	.w3(32'hbacb7813),
	.w4(32'hba82a66d),
	.w5(32'hba484f25),
	.w6(32'hba8d990b),
	.w7(32'hba48bb79),
	.w8(32'hbb31f732),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383420aa),
	.w1(32'h399902f9),
	.w2(32'h3af77b6b),
	.w3(32'h3aa3019c),
	.w4(32'h3aad84f1),
	.w5(32'h3b630f05),
	.w6(32'h3b237144),
	.w7(32'h3b04def0),
	.w8(32'h3b92173f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad1e1),
	.w1(32'h3a241910),
	.w2(32'h3a936529),
	.w3(32'hbac8923c),
	.w4(32'h39727fc7),
	.w5(32'h3a12ea3b),
	.w6(32'h3a57931d),
	.w7(32'h3a261463),
	.w8(32'h3a2cdc98),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e59a7b),
	.w1(32'h36cbc2ce),
	.w2(32'hba25aa49),
	.w3(32'hba141cd2),
	.w4(32'h390b350a),
	.w5(32'hb90ca2e3),
	.w6(32'h3abe158b),
	.w7(32'h3aa2c8ed),
	.w8(32'h39706c9f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba217cfc),
	.w1(32'hb8e7879c),
	.w2(32'h3a5c2ee9),
	.w3(32'hb9891d68),
	.w4(32'h3a2a2462),
	.w5(32'h3a943787),
	.w6(32'h3a4a5f00),
	.w7(32'h3ac6300e),
	.w8(32'h3a5f05bc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba772dd9),
	.w1(32'h3a031578),
	.w2(32'h39e0437a),
	.w3(32'hba6f98e1),
	.w4(32'hb9da5bcc),
	.w5(32'h388c6d4b),
	.w6(32'hbac7a44f),
	.w7(32'hbafe1b6c),
	.w8(32'hbaf1e6f9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed573e),
	.w1(32'hba62ce41),
	.w2(32'hbaeb30df),
	.w3(32'h396c8fe1),
	.w4(32'h38a847ce),
	.w5(32'hb8feecca),
	.w6(32'h3aa18339),
	.w7(32'h3a353cb9),
	.w8(32'h3966dac6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad54ef4),
	.w1(32'hb8e400aa),
	.w2(32'hba169846),
	.w3(32'hbaa5ef82),
	.w4(32'h3906755d),
	.w5(32'hb798d6a9),
	.w6(32'h3ac0dd7f),
	.w7(32'h3a96f1f3),
	.w8(32'h38553920),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9f0bb),
	.w1(32'hba57c7d8),
	.w2(32'hbabbf8f9),
	.w3(32'hba98507d),
	.w4(32'hba93ef47),
	.w5(32'hbabdbd55),
	.w6(32'hba5f338d),
	.w7(32'hbb38440a),
	.w8(32'hbb4a66cd),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0acff0),
	.w1(32'hbaae8061),
	.w2(32'hba83d895),
	.w3(32'hba9588fe),
	.w4(32'hba84b3a8),
	.w5(32'hb8abe48b),
	.w6(32'h3aa404ac),
	.w7(32'h38307626),
	.w8(32'h3a022308),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da0a3),
	.w1(32'h3b449613),
	.w2(32'h3b892277),
	.w3(32'h3ade31ae),
	.w4(32'h3a8e3bf9),
	.w5(32'h3aac516b),
	.w6(32'h3b6e09c4),
	.w7(32'h3a1d7f36),
	.w8(32'h3acf1094),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ce18),
	.w1(32'h3a90f8bc),
	.w2(32'h3b0233ad),
	.w3(32'h3b0a584e),
	.w4(32'h386e4991),
	.w5(32'h3a1d7dd7),
	.w6(32'h3ae74ad1),
	.w7(32'h3a6c9000),
	.w8(32'h3a9685c7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb0627),
	.w1(32'hb9325bfe),
	.w2(32'h3ac0b4db),
	.w3(32'h3ab30764),
	.w4(32'h39385f4f),
	.w5(32'h3a8e2946),
	.w6(32'hba65b7e0),
	.w7(32'hba0fb5b8),
	.w8(32'h3a41b410),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e045),
	.w1(32'hbae207b6),
	.w2(32'hba0e0ec1),
	.w3(32'hbb0a18c1),
	.w4(32'hba879cc1),
	.w5(32'hb985c904),
	.w6(32'hba0d18f7),
	.w7(32'h3a0152a4),
	.w8(32'h3a800cfe),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f76f3),
	.w1(32'h38aadcfa),
	.w2(32'hba4db386),
	.w3(32'h39d73a05),
	.w4(32'h3953d33d),
	.w5(32'hb9100c98),
	.w6(32'h3b14f010),
	.w7(32'h3af3140f),
	.w8(32'h39177a0a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb049556),
	.w1(32'hb9be9f49),
	.w2(32'hba42af8f),
	.w3(32'hbae0728c),
	.w4(32'hb92afbaa),
	.w5(32'hb9d4c8a9),
	.w6(32'h39e63c57),
	.w7(32'h39a2ac42),
	.w8(32'hb90b2cc5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94cd5f),
	.w1(32'hb9b2dbb9),
	.w2(32'hba2917cc),
	.w3(32'hba64f7f4),
	.w4(32'hb95a2b54),
	.w5(32'hb9fffa35),
	.w6(32'h3a651d8c),
	.w7(32'h3a547da8),
	.w8(32'h38d55039),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284ca3),
	.w1(32'h395aee69),
	.w2(32'h3b3c5dd3),
	.w3(32'h390bdc39),
	.w4(32'hba185335),
	.w5(32'h3a15b682),
	.w6(32'h3a363ba3),
	.w7(32'hbae0f262),
	.w8(32'hb9df774b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9f4a),
	.w1(32'hbac5568b),
	.w2(32'hb9809028),
	.w3(32'hba22ae74),
	.w4(32'hbab3ddb5),
	.w5(32'hb5ea6401),
	.w6(32'hbae1116f),
	.w7(32'hb998b2c7),
	.w8(32'hba9cb06b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abb6f),
	.w1(32'hba3816d9),
	.w2(32'h3a8d816d),
	.w3(32'hba8cdbbc),
	.w4(32'hba89bb84),
	.w5(32'h393d20ac),
	.w6(32'h3ab53784),
	.w7(32'h3aae6e3f),
	.w8(32'h3aa991a2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71341),
	.w1(32'h3954ec32),
	.w2(32'h3a27a400),
	.w3(32'h3936cbd4),
	.w4(32'hb9f61f06),
	.w5(32'hb80b7ae4),
	.w6(32'h3a83c8e5),
	.w7(32'h399dfbc1),
	.w8(32'hba0c8031),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfac79),
	.w1(32'hb8fd746a),
	.w2(32'hba35bdbc),
	.w3(32'hba37f360),
	.w4(32'h3969ddf4),
	.w5(32'h37098c73),
	.w6(32'h3a26dc0c),
	.w7(32'h39430405),
	.w8(32'h39063cec),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bda3f3),
	.w1(32'hba2a41b3),
	.w2(32'h3af34edd),
	.w3(32'h3859ccb9),
	.w4(32'hb9d9bcf9),
	.w5(32'hba7a4ffd),
	.w6(32'h3a15be7d),
	.w7(32'hba776f8d),
	.w8(32'hba7fcb7a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39657b29),
	.w1(32'h3a468adb),
	.w2(32'h3b136dab),
	.w3(32'hba24d9b2),
	.w4(32'hb980c341),
	.w5(32'h3a9c13bb),
	.w6(32'h3ac6ef93),
	.w7(32'h3b223648),
	.w8(32'h375f7c87),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec894b),
	.w1(32'h3a55c1d3),
	.w2(32'h3b12ea6b),
	.w3(32'h39e18a59),
	.w4(32'h39f8152c),
	.w5(32'h3ad3794d),
	.w6(32'h3b3a159e),
	.w7(32'h3b0efa54),
	.w8(32'h3a635a37),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac31db0),
	.w1(32'h37a2d453),
	.w2(32'h342b4ad0),
	.w3(32'hba9463b2),
	.w4(32'h37d27255),
	.w5(32'hb5f7cf07),
	.w6(32'hb6b816e0),
	.w7(32'h37f06cc7),
	.w8(32'hb7a53c81),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2f8ef),
	.w1(32'hbb2d6e5c),
	.w2(32'hbb192680),
	.w3(32'hba0b9d6c),
	.w4(32'hbb5781c5),
	.w5(32'hbb32018c),
	.w6(32'h3b5d99d0),
	.w7(32'hbb00c494),
	.w8(32'hb9a9e582),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule