module layer_8_featuremap_128(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc29cb3),
	.w1(32'h3c05c037),
	.w2(32'h3c17c5da),
	.w3(32'hb9eecffe),
	.w4(32'h3bef2bcd),
	.w5(32'h3b9f957c),
	.w6(32'hbc4ca6f6),
	.w7(32'hbba606de),
	.w8(32'hbb9f563b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74591),
	.w1(32'hbc3edcca),
	.w2(32'h3b1ac208),
	.w3(32'hb905519b),
	.w4(32'hbb207ede),
	.w5(32'hbb6b31cc),
	.w6(32'hba7a996f),
	.w7(32'h3a690772),
	.w8(32'h3a429f5e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c602c),
	.w1(32'hbc851f59),
	.w2(32'hbbf0317e),
	.w3(32'hbb68574e),
	.w4(32'h3bd7571e),
	.w5(32'h3bf69a41),
	.w6(32'hbac1bc3a),
	.w7(32'h3bf25a81),
	.w8(32'hb9a41c6d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dde38),
	.w1(32'h3c51a9ff),
	.w2(32'h3beaa457),
	.w3(32'h3b1007b0),
	.w4(32'h3c63288d),
	.w5(32'h3bc4615f),
	.w6(32'h3c1b3142),
	.w7(32'h3c0c1749),
	.w8(32'hbba680fe),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ee108),
	.w1(32'hbb4bcb26),
	.w2(32'hbb6c295d),
	.w3(32'h3a28a844),
	.w4(32'hbb5b5382),
	.w5(32'h3b44fb5d),
	.w6(32'hbc649ae6),
	.w7(32'h3aa74eb1),
	.w8(32'hbba16f21),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c656d),
	.w1(32'hbc01655e),
	.w2(32'hbab0bdca),
	.w3(32'hb97f18f6),
	.w4(32'hbc617d91),
	.w5(32'hbc88eafd),
	.w6(32'hbbe38239),
	.w7(32'h3b9230d1),
	.w8(32'h3c1cd82e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f71c5),
	.w1(32'h3be9313e),
	.w2(32'hbbcc357e),
	.w3(32'h3b136589),
	.w4(32'hbbd57dc8),
	.w5(32'hbb811375),
	.w6(32'hbb85f845),
	.w7(32'hbb0ef937),
	.w8(32'hbc05c2f4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891daa),
	.w1(32'hbbe84677),
	.w2(32'hbba78e35),
	.w3(32'h3b9716f6),
	.w4(32'h3c1d1690),
	.w5(32'hbb9858d3),
	.w6(32'hbb21ee8a),
	.w7(32'h3c1b8931),
	.w8(32'hbbca43c6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d29eb2a),
	.w1(32'h3c9e829f),
	.w2(32'h3b559f61),
	.w3(32'hba9c5415),
	.w4(32'h3c12de8f),
	.w5(32'h3bce4a53),
	.w6(32'h3c1c4314),
	.w7(32'h3c5d1d95),
	.w8(32'h3c33ce31),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35edca),
	.w1(32'h3b912d0e),
	.w2(32'h3c470695),
	.w3(32'hbb86e37d),
	.w4(32'h3c4ec76a),
	.w5(32'h39d8e6c2),
	.w6(32'h3b4a3217),
	.w7(32'h3be580b3),
	.w8(32'hbc4b9b62),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9829b),
	.w1(32'hbb5dca55),
	.w2(32'hbbeb91bd),
	.w3(32'h3c580895),
	.w4(32'h3b396a66),
	.w5(32'hbb143995),
	.w6(32'hbb897693),
	.w7(32'hbc0d18d2),
	.w8(32'hbcb140e5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadafe4),
	.w1(32'h3d2e9561),
	.w2(32'h3c989ef2),
	.w3(32'hbbecb144),
	.w4(32'h3c826c3a),
	.w5(32'h3b99454d),
	.w6(32'h3b8614d8),
	.w7(32'h3c7164ac),
	.w8(32'hbb459d5d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68fc22),
	.w1(32'h3ad667b8),
	.w2(32'h3b8f35dd),
	.w3(32'h3ab74c1b),
	.w4(32'hbaa4a702),
	.w5(32'h3ba09e08),
	.w6(32'h3b950d2e),
	.w7(32'h3c6a0a7c),
	.w8(32'h3ad8f934),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bcc7d),
	.w1(32'hba52669e),
	.w2(32'h3bb1c1f9),
	.w3(32'h3afe201d),
	.w4(32'h3b85845c),
	.w5(32'h3b5c1d3b),
	.w6(32'hbb84f88d),
	.w7(32'hbb221363),
	.w8(32'hbc093359),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36054),
	.w1(32'hbaa3d817),
	.w2(32'h3bed8958),
	.w3(32'h3b9e4d0a),
	.w4(32'h3b989b15),
	.w5(32'h3ba817e8),
	.w6(32'hbb62c7f8),
	.w7(32'h3affce69),
	.w8(32'hbb1a32fe),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c027041),
	.w1(32'h3b3441b8),
	.w2(32'h3b713068),
	.w3(32'h3ba6773f),
	.w4(32'h3c05333a),
	.w5(32'h3c51cd14),
	.w6(32'hb92d08fa),
	.w7(32'h3c27e02f),
	.w8(32'hbc90640c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5c40),
	.w1(32'h3bb04387),
	.w2(32'hbb5dfbc7),
	.w3(32'hbba6d665),
	.w4(32'hbb519918),
	.w5(32'hbbab31f1),
	.w6(32'hba0f56f3),
	.w7(32'h3c06aedc),
	.w8(32'hbc43857b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba36ea),
	.w1(32'hbade45ec),
	.w2(32'hbae3a11a),
	.w3(32'h3aeb153e),
	.w4(32'h3c0fe8e9),
	.w5(32'h3c097c45),
	.w6(32'h3941d9c6),
	.w7(32'h3a960959),
	.w8(32'hbcb46782),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ed721),
	.w1(32'h3c05b055),
	.w2(32'h3a86b3ad),
	.w3(32'h3c9590b6),
	.w4(32'h3d40f79f),
	.w5(32'h3c1d1f80),
	.w6(32'hbbcd56a1),
	.w7(32'hbba74af6),
	.w8(32'h3a0f1b4e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca86bfc),
	.w1(32'h3cafc9c8),
	.w2(32'h3c6eec11),
	.w3(32'h3c2fa646),
	.w4(32'h3c568dd1),
	.w5(32'h3cbe2097),
	.w6(32'hbd0f2464),
	.w7(32'hbc208adc),
	.w8(32'hbb5e1e77),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad98c7),
	.w1(32'h3ab9a498),
	.w2(32'hbcad55ed),
	.w3(32'hbb3b3fb2),
	.w4(32'hbc40b8bf),
	.w5(32'hbbf44263),
	.w6(32'hbbe01519),
	.w7(32'h3c4def43),
	.w8(32'hbb648b66),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d9132),
	.w1(32'h394fc8ce),
	.w2(32'hbce87e99),
	.w3(32'h3bf36db7),
	.w4(32'h3ac69929),
	.w5(32'hbc556023),
	.w6(32'hbc81a567),
	.w7(32'hbcee3824),
	.w8(32'h3d430e36),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ad730),
	.w1(32'h3cb06548),
	.w2(32'h3cc1d712),
	.w3(32'hbcd9e450),
	.w4(32'h3ca81a2f),
	.w5(32'h3d259e2b),
	.w6(32'hbd09fdd8),
	.w7(32'h3caba235),
	.w8(32'hbcf7c3ff),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4eadd),
	.w1(32'hba3cb630),
	.w2(32'h3b1bbb1a),
	.w3(32'h3c110788),
	.w4(32'hb9bdac99),
	.w5(32'h3cb78d6c),
	.w6(32'h3c0ff6c1),
	.w7(32'hbb478a13),
	.w8(32'h3c5edf2e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11089c),
	.w1(32'hbc206e80),
	.w2(32'hbbaa4a43),
	.w3(32'hbb0b5a84),
	.w4(32'hbbd38722),
	.w5(32'hbc01abce),
	.w6(32'hbbb23350),
	.w7(32'hbb026b81),
	.w8(32'hbb04e37e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acace),
	.w1(32'h3a15f94e),
	.w2(32'h3b2c5573),
	.w3(32'hbbcc1300),
	.w4(32'h3bdf1645),
	.w5(32'h3c922c64),
	.w6(32'hbc495a9e),
	.w7(32'hbc451b59),
	.w8(32'h3d4bfd2b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f33f7),
	.w1(32'h3a7978e7),
	.w2(32'h3b6b8b0d),
	.w3(32'hbbfe2682),
	.w4(32'h3b8e71e7),
	.w5(32'hbbd95b5b),
	.w6(32'h3c16fd1c),
	.w7(32'h3c2f05d9),
	.w8(32'hbc3a9a39),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2ab30f),
	.w1(32'h3d1da221),
	.w2(32'h3d22bf56),
	.w3(32'h3ca81465),
	.w4(32'h3cea7011),
	.w5(32'h3dba3128),
	.w6(32'hbd383ca3),
	.w7(32'hbd07743f),
	.w8(32'hbab75605),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65e537),
	.w1(32'h3c56828e),
	.w2(32'h3c89a56f),
	.w3(32'h3af062a4),
	.w4(32'hbc04c214),
	.w5(32'hbbc803bc),
	.w6(32'h3aba40bf),
	.w7(32'hbba4aa74),
	.w8(32'h3d3efb87),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9c051),
	.w1(32'h3c75f4bb),
	.w2(32'h3bd46733),
	.w3(32'hbb059d33),
	.w4(32'hbbd60b2f),
	.w5(32'hbba0070e),
	.w6(32'hba0345fb),
	.w7(32'hbbe7b702),
	.w8(32'h3cb66566),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41efeb),
	.w1(32'h3c529579),
	.w2(32'h3bb81c93),
	.w3(32'hbb9bb76c),
	.w4(32'h3a8a1dda),
	.w5(32'h3b7db73a),
	.w6(32'hbaba454e),
	.w7(32'h3a8a0f28),
	.w8(32'hb7150dd7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b030be5),
	.w1(32'hb89cb5aa),
	.w2(32'h3ada6338),
	.w3(32'h3bade28e),
	.w4(32'hbc2d9654),
	.w5(32'h3c90555b),
	.w6(32'hb9b694f3),
	.w7(32'h3a674778),
	.w8(32'hbc9a8961),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc100db),
	.w1(32'hbac69d94),
	.w2(32'h3c159c48),
	.w3(32'hbb25df0e),
	.w4(32'h3b085d12),
	.w5(32'hbc93fa07),
	.w6(32'hbb40b739),
	.w7(32'h3c845111),
	.w8(32'hbc0d2b2a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf58510),
	.w1(32'hbc9f6292),
	.w2(32'hbbb15551),
	.w3(32'hbbf186f0),
	.w4(32'hbaa4ab9a),
	.w5(32'hbc4dd533),
	.w6(32'hbc8fd1d8),
	.w7(32'hbbf0d0ae),
	.w8(32'hb956f8f1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fcc94),
	.w1(32'hbca1c291),
	.w2(32'hbc398d39),
	.w3(32'h3c64a0ce),
	.w4(32'hbbbbf329),
	.w5(32'hbbe4ec81),
	.w6(32'hbc349a6c),
	.w7(32'hba16e8f1),
	.w8(32'hbbf29c22),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7c9ed),
	.w1(32'h3c5e445d),
	.w2(32'hba418480),
	.w3(32'h3bc714d5),
	.w4(32'h3ccc79ec),
	.w5(32'h3c8c4329),
	.w6(32'h3a398b48),
	.w7(32'hbc36d17f),
	.w8(32'h3c7ffa37),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc466d63),
	.w1(32'h3bb24388),
	.w2(32'hbc78a8e5),
	.w3(32'hbc5c1de0),
	.w4(32'h3c1c9341),
	.w5(32'h3ad992a1),
	.w6(32'h3ce9555f),
	.w7(32'h3c6b0a27),
	.w8(32'hbc1b5265),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17c700),
	.w1(32'hbc32ce10),
	.w2(32'h3c14c0fc),
	.w3(32'h3c236a04),
	.w4(32'hbbbf86c8),
	.w5(32'h3c1cb61e),
	.w6(32'hba3d550b),
	.w7(32'h3b583ac0),
	.w8(32'h3b07018c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba38fd8),
	.w1(32'hba5a4354),
	.w2(32'hbc178dea),
	.w3(32'h3c74f7bc),
	.w4(32'h3b7ae818),
	.w5(32'hbc7ffaaf),
	.w6(32'hbbb41300),
	.w7(32'hbc745241),
	.w8(32'h3d17098f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8343fd),
	.w1(32'h39f33d10),
	.w2(32'hba0ae336),
	.w3(32'hbceb633c),
	.w4(32'hbb68f8a1),
	.w5(32'hbb13c23f),
	.w6(32'h3b10c3f3),
	.w7(32'h3c0686e3),
	.w8(32'h3c01fd3b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ba08),
	.w1(32'h3b15f31e),
	.w2(32'h3c58763a),
	.w3(32'h3beb5134),
	.w4(32'h3c9deb6e),
	.w5(32'h3d0cdab0),
	.w6(32'hbbaf498a),
	.w7(32'h3c1e467b),
	.w8(32'h3ac896f1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e8ea),
	.w1(32'h3cac82cc),
	.w2(32'h3d09f3ba),
	.w3(32'h3aeaf6ca),
	.w4(32'h3c6c6b07),
	.w5(32'h3b562028),
	.w6(32'h3b85e878),
	.w7(32'hbc503ad9),
	.w8(32'hbb2346bc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bec5e),
	.w1(32'h3bda184b),
	.w2(32'hbb45f5e3),
	.w3(32'hbc1d48ae),
	.w4(32'h3bcf166e),
	.w5(32'hbc9b6382),
	.w6(32'h3babb664),
	.w7(32'h3ce23ee8),
	.w8(32'hbb46a603),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccb2bd),
	.w1(32'hbce3a026),
	.w2(32'h3b858256),
	.w3(32'h3c379582),
	.w4(32'h3bda9f25),
	.w5(32'h3c8e8ee8),
	.w6(32'h3b90f263),
	.w7(32'h3bc57d46),
	.w8(32'h3b0af893),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7289c5),
	.w1(32'h3c44c7f5),
	.w2(32'h3c9b55e3),
	.w3(32'h3b7b7b94),
	.w4(32'h3c58d0cc),
	.w5(32'hbb5cd8c1),
	.w6(32'hbc2469b3),
	.w7(32'hbbef1c08),
	.w8(32'h3d259d0d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e53b9),
	.w1(32'h3c8dd268),
	.w2(32'h3c691876),
	.w3(32'hbcbbba80),
	.w4(32'h3ab223df),
	.w5(32'h3ca716c4),
	.w6(32'hbc22b03e),
	.w7(32'hbc9334cf),
	.w8(32'h3c611688),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc2224),
	.w1(32'h3b939278),
	.w2(32'hbc40025e),
	.w3(32'hbaf72f37),
	.w4(32'hbc0f8b79),
	.w5(32'hbc82835e),
	.w6(32'h3c7c0a97),
	.w7(32'hbceba546),
	.w8(32'h3d83710c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75880f),
	.w1(32'h3ca88ac7),
	.w2(32'hbcc9e9d6),
	.w3(32'h3b693b11),
	.w4(32'h3c019823),
	.w5(32'h3c484cf3),
	.w6(32'hbd0ce079),
	.w7(32'hbbe5130b),
	.w8(32'h3d3d42fe),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6aa1f0),
	.w1(32'h3a1fe99e),
	.w2(32'h3acc9298),
	.w3(32'h3bbc159a),
	.w4(32'hbb6e28ad),
	.w5(32'h3b910744),
	.w6(32'hbbb22ced),
	.w7(32'h3c1f7a3e),
	.w8(32'hbd033b0b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd57ff1),
	.w1(32'hbbbce234),
	.w2(32'hbc2a988b),
	.w3(32'hbb908faa),
	.w4(32'hbbd698d1),
	.w5(32'hbc3467e9),
	.w6(32'h3bf9efa4),
	.w7(32'hbc0f1dd4),
	.w8(32'hbba57901),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b1387),
	.w1(32'hbcddebf4),
	.w2(32'h3cceae6c),
	.w3(32'hbcb2cde9),
	.w4(32'hbd03a5c9),
	.w5(32'h3d21d9ce),
	.w6(32'hbc3e7014),
	.w7(32'hbc3788eb),
	.w8(32'hbd5e7458),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36decf),
	.w1(32'h3bdca85a),
	.w2(32'h3c2cfc12),
	.w3(32'h3bcc481d),
	.w4(32'h3c658cb3),
	.w5(32'h3cc004d0),
	.w6(32'hbbab9496),
	.w7(32'h3ca6de16),
	.w8(32'h3c8226d1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a104f),
	.w1(32'h3be76755),
	.w2(32'h3b7c35e5),
	.w3(32'h3b9aac81),
	.w4(32'h3b6f9602),
	.w5(32'h3c6b1414),
	.w6(32'hbc619f49),
	.w7(32'h3c8e8b6b),
	.w8(32'hbc9104de),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca742c5),
	.w1(32'h3c156f1a),
	.w2(32'h3c4f139e),
	.w3(32'h3c0c7f4f),
	.w4(32'h3baf8de2),
	.w5(32'h3c519e8f),
	.w6(32'h3be73f6c),
	.w7(32'h3b709ef2),
	.w8(32'hb96d94a7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab44262),
	.w1(32'hb98b1bb4),
	.w2(32'hbcb95443),
	.w3(32'hb9d0b21b),
	.w4(32'h3c0326d5),
	.w5(32'hbcad1e60),
	.w6(32'hbba75945),
	.w7(32'h3c0a2c46),
	.w8(32'hbcaaaabe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830f0a),
	.w1(32'h3c683249),
	.w2(32'h3c462d4f),
	.w3(32'hbaddf624),
	.w4(32'h3c96ab83),
	.w5(32'h3ce7ee8e),
	.w6(32'hbc219d4a),
	.w7(32'h3c094012),
	.w8(32'h3bd9e69f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ed909),
	.w1(32'h3c352209),
	.w2(32'h3bdae0ca),
	.w3(32'hbc6dd2c0),
	.w4(32'hbc0efc2a),
	.w5(32'hbbe9d0cb),
	.w6(32'hbc27dbd4),
	.w7(32'h3b9f825b),
	.w8(32'hbc4554f5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585587),
	.w1(32'hbc327317),
	.w2(32'hbc3698ad),
	.w3(32'h3c1b64b2),
	.w4(32'h3b8d457b),
	.w5(32'h3cf4843a),
	.w6(32'hbb62fe1f),
	.w7(32'hbc8ccdb0),
	.w8(32'h3cee0be7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b63e),
	.w1(32'h3bd27c25),
	.w2(32'h3b5101dd),
	.w3(32'hbc78b9cd),
	.w4(32'h3bebe351),
	.w5(32'h3c4f71e2),
	.w6(32'h3bfb46d2),
	.w7(32'h3bb1eb8c),
	.w8(32'h39442432),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4155fa),
	.w1(32'h3a3c3648),
	.w2(32'h3b9394ee),
	.w3(32'h3b1433a9),
	.w4(32'hbccef3f2),
	.w5(32'h3cc55063),
	.w6(32'hba676eb3),
	.w7(32'h3cc1cfab),
	.w8(32'hbd292ef8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc930e9),
	.w1(32'hbcdc9120),
	.w2(32'h3ae54178),
	.w3(32'hbc274a36),
	.w4(32'h3c4fb725),
	.w5(32'hbc666e61),
	.w6(32'h3cc1226f),
	.w7(32'hbc58582e),
	.w8(32'h3c506fae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc945567),
	.w1(32'h3c804c3b),
	.w2(32'h3bc34b57),
	.w3(32'hbca98e1c),
	.w4(32'hbc21c508),
	.w5(32'hbc101fce),
	.w6(32'hbc890a2e),
	.w7(32'h3aaf7a15),
	.w8(32'h3bf1c8b3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac14c67),
	.w1(32'h3a7a512e),
	.w2(32'h3cc3bdc3),
	.w3(32'h3c00405f),
	.w4(32'h3c686dd9),
	.w5(32'h3b49ac8e),
	.w6(32'hbb98cbb7),
	.w7(32'h3b34f122),
	.w8(32'h3d2359ef),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82797f),
	.w1(32'hbc3c2a30),
	.w2(32'hbba47cbf),
	.w3(32'h3c2fe373),
	.w4(32'h3bdc1b2c),
	.w5(32'h3bd13dc7),
	.w6(32'hbc1d6ca1),
	.w7(32'hbb5f4888),
	.w8(32'h3c6d0723),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e7326),
	.w1(32'hbb8ee6db),
	.w2(32'h3bdeff16),
	.w3(32'hbbac5112),
	.w4(32'hb969ac13),
	.w5(32'h3c0d9013),
	.w6(32'hbc2a9671),
	.w7(32'hbb19cdfd),
	.w8(32'hbbd2a9a6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a28f5),
	.w1(32'h3a83039c),
	.w2(32'h3c28d7b3),
	.w3(32'h3c0c33fa),
	.w4(32'h3c78160d),
	.w5(32'h3c1bca41),
	.w6(32'h39655ec7),
	.w7(32'h3bcb923a),
	.w8(32'h3b309ae2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247a80),
	.w1(32'hbb2648ad),
	.w2(32'h3c0df049),
	.w3(32'h3c4d99a3),
	.w4(32'hbb93add4),
	.w5(32'hbc9d2c5a),
	.w6(32'h3bdec55d),
	.w7(32'h3c03203e),
	.w8(32'h3d7002b2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9fb33),
	.w1(32'h3c0d56d7),
	.w2(32'hbbf98cd4),
	.w3(32'hbba13f4f),
	.w4(32'h3bfca5f9),
	.w5(32'h3be89428),
	.w6(32'hbd046623),
	.w7(32'hbc50375f),
	.w8(32'h3a94624b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc576456),
	.w1(32'h3baf5f2d),
	.w2(32'hbb938221),
	.w3(32'h3c3e3454),
	.w4(32'h3b3d750f),
	.w5(32'hbc7ef33b),
	.w6(32'h3ba924e7),
	.w7(32'hbc05a99c),
	.w8(32'hbc704fc5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6a005),
	.w1(32'h394b1eb6),
	.w2(32'h3c3c208f),
	.w3(32'hbc1d7db3),
	.w4(32'h3cb75081),
	.w5(32'h3cd6d108),
	.w6(32'hbc00ae97),
	.w7(32'h39ed6361),
	.w8(32'hbbfc2520),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b7541),
	.w1(32'h3adddcba),
	.w2(32'h3c5701b3),
	.w3(32'h3c9f7f3d),
	.w4(32'hbbe31145),
	.w5(32'h3b99d656),
	.w6(32'hbac11827),
	.w7(32'h3d044a06),
	.w8(32'hbcedc720),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9114ef),
	.w1(32'hbb5dd330),
	.w2(32'h3cd6b6ca),
	.w3(32'h3bf5fc7f),
	.w4(32'h3c55d425),
	.w5(32'h3d01e550),
	.w6(32'h3c58913b),
	.w7(32'hbbfc5254),
	.w8(32'h3bd3b24d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118b40),
	.w1(32'hbc235182),
	.w2(32'h3b7457e6),
	.w3(32'hbc186fc3),
	.w4(32'hbc12a9e0),
	.w5(32'h3c080374),
	.w6(32'h3c5637f9),
	.w7(32'h3a0e2a76),
	.w8(32'hbc817661),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc333),
	.w1(32'h3c95591e),
	.w2(32'h3c4afccf),
	.w3(32'h3be2bbfd),
	.w4(32'hbd05ff66),
	.w5(32'h3d32b5e9),
	.w6(32'h3cb2001c),
	.w7(32'h3d625362),
	.w8(32'hbe23fe66),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6a3906),
	.w1(32'hbd337eb4),
	.w2(32'hbc86232c),
	.w3(32'h3c18e8a8),
	.w4(32'hbad104fe),
	.w5(32'hbc8fe191),
	.w6(32'h3d85ff64),
	.w7(32'hbcb0fb55),
	.w8(32'h3d731e7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0cecc),
	.w1(32'hbc59f0dc),
	.w2(32'hba72a978),
	.w3(32'h3a51cc0e),
	.w4(32'h3b4ea6d0),
	.w5(32'h3bc837a5),
	.w6(32'hbd3229af),
	.w7(32'hbc1f10a4),
	.w8(32'hbc82eb97),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cc12),
	.w1(32'h3b8b5d72),
	.w2(32'hbad08c4e),
	.w3(32'hbbbb2221),
	.w4(32'hbb956270),
	.w5(32'h3bb9ae9a),
	.w6(32'h3bd71cb8),
	.w7(32'h3b856ef1),
	.w8(32'hbbea2cb7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4f24),
	.w1(32'h3c2e7018),
	.w2(32'h3c5216f5),
	.w3(32'h3b866021),
	.w4(32'h3c613ebb),
	.w5(32'h3c954f26),
	.w6(32'hbc17e1ba),
	.w7(32'h3b852942),
	.w8(32'h3b329997),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c142bff),
	.w1(32'h3c8be7e3),
	.w2(32'h3ba86094),
	.w3(32'h3b02287b),
	.w4(32'h3b92fac3),
	.w5(32'h3bcd079c),
	.w6(32'h3c1e1dc9),
	.w7(32'hb90b2b17),
	.w8(32'h3b2de41d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd045e9),
	.w1(32'h3bb53348),
	.w2(32'hbb76cdc9),
	.w3(32'h3c195e52),
	.w4(32'h38c08338),
	.w5(32'h3c3cb9e9),
	.w6(32'h3c382836),
	.w7(32'h3c38281e),
	.w8(32'h3b9c7843),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ecdc4),
	.w1(32'h3b6d55ba),
	.w2(32'h3b51c77a),
	.w3(32'hbb34bd9d),
	.w4(32'h3ab8247f),
	.w5(32'hbc627df3),
	.w6(32'hbb4c4052),
	.w7(32'hbc207e18),
	.w8(32'h3b15cb54),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c1c77),
	.w1(32'h3bc16f81),
	.w2(32'hbaa816ed),
	.w3(32'hbadec34e),
	.w4(32'h3ced490f),
	.w5(32'h3c93a7ee),
	.w6(32'h3c9bfc1a),
	.w7(32'h3c89ff13),
	.w8(32'h3c7f3fe9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79da60),
	.w1(32'hbbba4773),
	.w2(32'h3c51c371),
	.w3(32'hbb953855),
	.w4(32'h39e6d0ee),
	.w5(32'h3c88dc54),
	.w6(32'hbbcc5baf),
	.w7(32'hbba35384),
	.w8(32'h3c2d23a4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb0aa5),
	.w1(32'h3c396656),
	.w2(32'h3ce14167),
	.w3(32'h3c107861),
	.w4(32'hbbf9c295),
	.w5(32'hbc32ed7d),
	.w6(32'hbbe0127d),
	.w7(32'hbc50964f),
	.w8(32'hbba89ded),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb94e5),
	.w1(32'h3c0d6053),
	.w2(32'h3ce764ba),
	.w3(32'hbbf8b4dc),
	.w4(32'h3c69af93),
	.w5(32'h3ccaf245),
	.w6(32'hbc246297),
	.w7(32'h3ba347bc),
	.w8(32'h3d818506),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a35e),
	.w1(32'h3b8bcdb6),
	.w2(32'h3aad5a10),
	.w3(32'hbc4cf5be),
	.w4(32'h3be80ddc),
	.w5(32'h3c32d485),
	.w6(32'h3bbe060c),
	.w7(32'h3c812c6d),
	.w8(32'h3b84a488),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce11c5c),
	.w1(32'hbc6f1b06),
	.w2(32'hbc8b3662),
	.w3(32'hbba0d537),
	.w4(32'h3b3e1c40),
	.w5(32'hbb1161f6),
	.w6(32'hbbcfb407),
	.w7(32'hbccd4747),
	.w8(32'hbc088b4a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dcb53),
	.w1(32'hbc2eafb6),
	.w2(32'hbab59bb7),
	.w3(32'hbba865b3),
	.w4(32'h3b946a60),
	.w5(32'h3bc9b962),
	.w6(32'hbb5c176b),
	.w7(32'h3b2b21fe),
	.w8(32'hbbcfe909),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82077e),
	.w1(32'hbab02d77),
	.w2(32'hbb277411),
	.w3(32'h3b30649c),
	.w4(32'h3b3ce0f8),
	.w5(32'hbb762998),
	.w6(32'h3b56bea6),
	.w7(32'hbb9ce8d7),
	.w8(32'hbc10bf97),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49512b),
	.w1(32'hbb9a5f55),
	.w2(32'h3c542708),
	.w3(32'hbc1677bd),
	.w4(32'hbcde5866),
	.w5(32'hbc3bf220),
	.w6(32'hbc58568a),
	.w7(32'h39089787),
	.w8(32'h3d5cc8ac),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3de5d4),
	.w1(32'h3b83efd0),
	.w2(32'h3c164536),
	.w3(32'h3c6c8883),
	.w4(32'h3ad375e8),
	.w5(32'hba6da33a),
	.w6(32'h3d3e881a),
	.w7(32'hb80ad5d0),
	.w8(32'h3cea0496),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4031e),
	.w1(32'hb9f54adf),
	.w2(32'hbc2ebae3),
	.w3(32'hbc4171e8),
	.w4(32'hbd3120ae),
	.w5(32'hbc80c7e2),
	.w6(32'h3c34728b),
	.w7(32'hbd07f406),
	.w8(32'h3d4c0303),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebcbb4),
	.w1(32'hbb17a8c8),
	.w2(32'hbc2bf3a9),
	.w3(32'h3c9b06c0),
	.w4(32'h3c1968c5),
	.w5(32'hbb2525ca),
	.w6(32'h3d01514c),
	.w7(32'hbbe66251),
	.w8(32'hbc4037da),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32d825),
	.w1(32'h3c6589d5),
	.w2(32'hbc44605b),
	.w3(32'h3c315ba4),
	.w4(32'h3c86e476),
	.w5(32'hb9e62ae5),
	.w6(32'h3b1c0ec2),
	.w7(32'hbc94faaa),
	.w8(32'hbd81ae15),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d288d),
	.w1(32'h3c927ce2),
	.w2(32'h3c2e497f),
	.w3(32'hbc615a00),
	.w4(32'h3ba63ac6),
	.w5(32'h3c5b75c7),
	.w6(32'hbc364a22),
	.w7(32'h3be9535f),
	.w8(32'h3c63fb1b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0da82e),
	.w1(32'h3b3b3409),
	.w2(32'hbb457dd4),
	.w3(32'hbafeded7),
	.w4(32'hbb002337),
	.w5(32'h3d1807d0),
	.w6(32'h3b0ef560),
	.w7(32'h3c81956b),
	.w8(32'hbcc08079),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65526e),
	.w1(32'h3d1dc92d),
	.w2(32'hbb9d09c1),
	.w3(32'h3c94ac09),
	.w4(32'h3d2bea6c),
	.w5(32'h3d1e8875),
	.w6(32'hbd06171a),
	.w7(32'h3d009dfd),
	.w8(32'hbcd71f8d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd39c963),
	.w1(32'h3ba00fec),
	.w2(32'h3bb08dd4),
	.w3(32'hbb6dbba7),
	.w4(32'hbace4bb3),
	.w5(32'h3a86c2f7),
	.w6(32'hbd189cec),
	.w7(32'h3c3911bb),
	.w8(32'h3cb817e5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b848ae5),
	.w1(32'hbc89542a),
	.w2(32'h3c0b070e),
	.w3(32'hbc7e5a5c),
	.w4(32'h3b0ae881),
	.w5(32'h3b0994e6),
	.w6(32'h3c383a0c),
	.w7(32'h3bb58cca),
	.w8(32'h3bd97315),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c2279),
	.w1(32'h3bbaf88a),
	.w2(32'hbbf2e1a3),
	.w3(32'h3c6d3cd2),
	.w4(32'h3ccf1e90),
	.w5(32'h3cd7f3d6),
	.w6(32'h3c09c9b6),
	.w7(32'h3b1df826),
	.w8(32'hbc14e257),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73fc44),
	.w1(32'hbbd4da1a),
	.w2(32'hbc293bb3),
	.w3(32'h3ccafd0f),
	.w4(32'hbc258046),
	.w5(32'h3bae5fb6),
	.w6(32'hbcc0b85f),
	.w7(32'h3c21347a),
	.w8(32'h3baedac8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81766d),
	.w1(32'h3bfce953),
	.w2(32'hba4efb49),
	.w3(32'hbc3331b8),
	.w4(32'h3a707ae6),
	.w5(32'h3c881a91),
	.w6(32'hbbb26e84),
	.w7(32'h3c9ff1e4),
	.w8(32'h3c73ab0e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc069c42),
	.w1(32'h3c01786e),
	.w2(32'hbb922f0d),
	.w3(32'hbc3bf400),
	.w4(32'h3c01f5f3),
	.w5(32'hb9c9d24e),
	.w6(32'h3c2a6de7),
	.w7(32'h3b17f712),
	.w8(32'hbbb253dd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73007c),
	.w1(32'h3b936337),
	.w2(32'h3b62112b),
	.w3(32'h3c2f3f2b),
	.w4(32'h3c013f99),
	.w5(32'hbb217a7a),
	.w6(32'h3c0a22dc),
	.w7(32'h3ac7b4d2),
	.w8(32'hbbdbdac1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ea88),
	.w1(32'h3bc040f5),
	.w2(32'h3ad0b5c0),
	.w3(32'hbc1e0a8e),
	.w4(32'hbb8fc643),
	.w5(32'h3b48b3b6),
	.w6(32'hbbd9f7c1),
	.w7(32'h3ac44b28),
	.w8(32'hbc64bd5c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60722c),
	.w1(32'h3c0c508c),
	.w2(32'hbbb9df53),
	.w3(32'hbc011f1e),
	.w4(32'h3c1ec6ab),
	.w5(32'h3c8386fa),
	.w6(32'h3c9748a1),
	.w7(32'hbcffb2b3),
	.w8(32'h3d522b15),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0be994),
	.w1(32'h39d2fd97),
	.w2(32'hb9322c72),
	.w3(32'hbb40c0e6),
	.w4(32'h3cc30bde),
	.w5(32'h3d02f4f0),
	.w6(32'h3bb49d23),
	.w7(32'h3c9a9b89),
	.w8(32'hbce36d5b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1bfbe4),
	.w1(32'h3baf0abc),
	.w2(32'hba7fcce7),
	.w3(32'h3b0df5be),
	.w4(32'hbb2200f7),
	.w5(32'h3c1f0430),
	.w6(32'hbcd9188b),
	.w7(32'h3bb44619),
	.w8(32'hbb7f7bbd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3b7a2),
	.w1(32'h3ae8a7c6),
	.w2(32'hbc8b4843),
	.w3(32'h3b839572),
	.w4(32'hbb9e838e),
	.w5(32'hbc8912e8),
	.w6(32'hb9900945),
	.w7(32'hbd0c4a47),
	.w8(32'hbcc827db),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c023fcc),
	.w1(32'h3c771b74),
	.w2(32'h3bdd3330),
	.w3(32'h3c0e9423),
	.w4(32'h3c831ced),
	.w5(32'h3cddf8b4),
	.w6(32'h3c58492e),
	.w7(32'h3b309842),
	.w8(32'hbb524a46),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a264956),
	.w1(32'hbc0453d9),
	.w2(32'h3b65e2a1),
	.w3(32'h3c7e129e),
	.w4(32'h3c0957f1),
	.w5(32'h3b414d62),
	.w6(32'hbcd4a532),
	.w7(32'hbbbf2b4d),
	.w8(32'hbc48734e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9c7f6),
	.w1(32'h3c9efecd),
	.w2(32'hbba91679),
	.w3(32'h3c89556e),
	.w4(32'h3cb81f23),
	.w5(32'hbc6ade14),
	.w6(32'hbc2fd00f),
	.w7(32'h3c169155),
	.w8(32'hbcb64f8f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48de75),
	.w1(32'h3cb33e8f),
	.w2(32'hbba47720),
	.w3(32'hbcac7d10),
	.w4(32'h3c655443),
	.w5(32'hbc3614b9),
	.w6(32'h3b88f978),
	.w7(32'hbca1d74f),
	.w8(32'h3d1cc9d5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed1036),
	.w1(32'hbcc7be3e),
	.w2(32'hbcf545e5),
	.w3(32'h3b84f9c2),
	.w4(32'h3a93c665),
	.w5(32'h3c2867af),
	.w6(32'h3b9e7b2f),
	.w7(32'hbc89b7dc),
	.w8(32'hbc1b191e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f73df),
	.w1(32'hbbf237fa),
	.w2(32'h3af72952),
	.w3(32'hbca16a71),
	.w4(32'hbb81d44d),
	.w5(32'h3b78d102),
	.w6(32'hbc93b808),
	.w7(32'hbc43a8ce),
	.w8(32'h3cac9b68),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12d779),
	.w1(32'h3c1bff96),
	.w2(32'h3caa0764),
	.w3(32'h3b0c33da),
	.w4(32'hbd0e67c9),
	.w5(32'hbcf483c4),
	.w6(32'h3ba5dbd9),
	.w7(32'h3c273351),
	.w8(32'h3c90ee74),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb33f59),
	.w1(32'h3c92a6d8),
	.w2(32'hbc05becd),
	.w3(32'hbcae79ef),
	.w4(32'hbce2a849),
	.w5(32'h3c5dc1a9),
	.w6(32'h3ce282ba),
	.w7(32'h3c8db085),
	.w8(32'hbac2a7a9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6301),
	.w1(32'h3c5b3c7c),
	.w2(32'h3b1583ba),
	.w3(32'h3b4f96a2),
	.w4(32'hb58b25b6),
	.w5(32'h3c3904a2),
	.w6(32'hbb502fec),
	.w7(32'hb98511eb),
	.w8(32'hba05cf02),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2395db),
	.w1(32'h3ba3dd8a),
	.w2(32'hbae9a62d),
	.w3(32'h3b42e314),
	.w4(32'hbaf8d2d7),
	.w5(32'hbc8d175c),
	.w6(32'h3a9e7d16),
	.w7(32'hbc94809f),
	.w8(32'hbc185375),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b0a28),
	.w1(32'hba643b87),
	.w2(32'hbc154cc4),
	.w3(32'hbc1d7b19),
	.w4(32'hb9fa49d3),
	.w5(32'h3c2bf000),
	.w6(32'hbb049583),
	.w7(32'h3a99e199),
	.w8(32'hbc4ab85d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73162e),
	.w1(32'h3a220b26),
	.w2(32'h3c227cf4),
	.w3(32'hbc0ea2ba),
	.w4(32'hbc0a338f),
	.w5(32'h3bd65e92),
	.w6(32'hbb81772b),
	.w7(32'h3be7f7fb),
	.w8(32'h3ce398af),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8abb00),
	.w1(32'h3c2cb4c6),
	.w2(32'hbb43f105),
	.w3(32'h3c8498d5),
	.w4(32'hbd01b22e),
	.w5(32'hbcf36108),
	.w6(32'h3c3e59fb),
	.w7(32'hbcaa0d7a),
	.w8(32'h3cdd7b5d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00f6bf),
	.w1(32'h3c0eba52),
	.w2(32'h3acb826d),
	.w3(32'h3b3b3ac0),
	.w4(32'hbb2b503f),
	.w5(32'h3c01b9ce),
	.w6(32'h3cd445c8),
	.w7(32'h3a6158e0),
	.w8(32'hbb8fd8b8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8d67),
	.w1(32'hb93a09b5),
	.w2(32'h3c18d889),
	.w3(32'h3b1bb8c0),
	.w4(32'hbc8726e7),
	.w5(32'h3c8364cb),
	.w6(32'h39c16151),
	.w7(32'h3cbea853),
	.w8(32'h3d4eaa69),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aaccd),
	.w1(32'hbca12096),
	.w2(32'hbcd15ec5),
	.w3(32'h3c7f4367),
	.w4(32'hbbc5a900),
	.w5(32'h3ccb050b),
	.w6(32'h3b36c072),
	.w7(32'hbc83650f),
	.w8(32'h3c54c5d9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d540c),
	.w1(32'hbbb70e85),
	.w2(32'h3b3db31c),
	.w3(32'h3ca93d44),
	.w4(32'h3c42c691),
	.w5(32'h3c1ea9c7),
	.w6(32'h3cabf1ac),
	.w7(32'h3a3e40ed),
	.w8(32'hbab8e5b5),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041f72),
	.w1(32'h3bd18faa),
	.w2(32'hbac15684),
	.w3(32'h3bf7f598),
	.w4(32'hbc0f5c54),
	.w5(32'hbb3403e4),
	.w6(32'h3a923f40),
	.w7(32'h3c0e4b9a),
	.w8(32'hbcb8bf5f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0073c),
	.w1(32'h3c86326d),
	.w2(32'hbae059f1),
	.w3(32'hbbba2ae8),
	.w4(32'h3b3409d1),
	.w5(32'h3c1871a7),
	.w6(32'h3c1ea11e),
	.w7(32'h3c197238),
	.w8(32'hbc76efdb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule