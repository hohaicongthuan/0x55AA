module layer_10_featuremap_54(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeee6ef),
	.w1(32'hba9b5858),
	.w2(32'hbbe55d9e),
	.w3(32'hbae80fdf),
	.w4(32'hbb669f57),
	.w5(32'hbbbe2fc3),
	.w6(32'hba8ebf6b),
	.w7(32'hbaf775fc),
	.w8(32'hbb89b86a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d33b5),
	.w1(32'hba7e7810),
	.w2(32'h3ba83ee2),
	.w3(32'hbb2b41e1),
	.w4(32'hbb5b8b71),
	.w5(32'h3a1d4b34),
	.w6(32'hbb38b185),
	.w7(32'hbb4cbb45),
	.w8(32'h3a8c5b65),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c0099),
	.w1(32'hbbde45e4),
	.w2(32'h3a9aafb0),
	.w3(32'h3aab62a0),
	.w4(32'hbbd5b87e),
	.w5(32'h3b15c376),
	.w6(32'hb92e521f),
	.w7(32'hbb9e8bfe),
	.w8(32'h3984c8ee),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2751e9),
	.w1(32'h3b182745),
	.w2(32'h3a04c934),
	.w3(32'hbadda9fd),
	.w4(32'hb7e589a3),
	.w5(32'hbaf2b656),
	.w6(32'hba4b5d75),
	.w7(32'h38edfcd4),
	.w8(32'hba8fe53f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad37a38),
	.w1(32'hbb34d505),
	.w2(32'hbb8a2084),
	.w3(32'hbabbfb26),
	.w4(32'hbb67c8dd),
	.w5(32'hbbc5cd47),
	.w6(32'hba66a8f3),
	.w7(32'hbae05e0a),
	.w8(32'hbbcb5f20),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c094),
	.w1(32'h3b4229a9),
	.w2(32'h3bc62526),
	.w3(32'hbb8adb91),
	.w4(32'h3b8e22a9),
	.w5(32'h3b9ca239),
	.w6(32'hbb8f2183),
	.w7(32'h3c0593ab),
	.w8(32'h3b8aa6a5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c655680),
	.w1(32'h3c0e349a),
	.w2(32'hb95f35ed),
	.w3(32'h3c53c65f),
	.w4(32'h3c26890b),
	.w5(32'hbb8426e0),
	.w6(32'h3c1301bc),
	.w7(32'h3c199388),
	.w8(32'hbbc04cff),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc344),
	.w1(32'hbc552aeb),
	.w2(32'hbbf8766e),
	.w3(32'h3b889d49),
	.w4(32'hbad9cec3),
	.w5(32'hbb8df211),
	.w6(32'hbaf140b4),
	.w7(32'hbbae3955),
	.w8(32'h3a80155d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d14b5),
	.w1(32'hb9a5c377),
	.w2(32'hba932f8e),
	.w3(32'hbb9bce25),
	.w4(32'hbb1edeaf),
	.w5(32'hbaf16338),
	.w6(32'hbb18177c),
	.w7(32'hba32458b),
	.w8(32'hbb45b60f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c718),
	.w1(32'hbb99a3bf),
	.w2(32'hbb827c81),
	.w3(32'h395e4420),
	.w4(32'hbb359af2),
	.w5(32'hbb9c3a64),
	.w6(32'hbaf7e861),
	.w7(32'hbb704091),
	.w8(32'hbb73c0c2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba014e1),
	.w1(32'hbb623e6a),
	.w2(32'hbb214779),
	.w3(32'hbbd2c614),
	.w4(32'hbb90a5ba),
	.w5(32'hbb5f9854),
	.w6(32'hbbc7c0ba),
	.w7(32'hbb81f208),
	.w8(32'hb8a924b4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c19a4),
	.w1(32'h39833835),
	.w2(32'h3c2bf118),
	.w3(32'h3bc2a5ce),
	.w4(32'h3b0d27b4),
	.w5(32'h3c013b57),
	.w6(32'h399c7920),
	.w7(32'h3b861210),
	.w8(32'h3bf64cfb),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb193a),
	.w1(32'h3b72fc34),
	.w2(32'h3b7c1549),
	.w3(32'h3c2737d6),
	.w4(32'h3bada54d),
	.w5(32'hbae95690),
	.w6(32'h3c2e04b8),
	.w7(32'h3bf8ad01),
	.w8(32'h3ad7107e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6278b),
	.w1(32'hb9d87562),
	.w2(32'hbb599e78),
	.w3(32'h3a50075e),
	.w4(32'hba25572f),
	.w5(32'hbbd17f97),
	.w6(32'hbb37dab5),
	.w7(32'hbb22d448),
	.w8(32'hbbb7b6d0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39044b6f),
	.w1(32'hbb0bca39),
	.w2(32'h3b9062ee),
	.w3(32'hbb12eca2),
	.w4(32'hbb3f6966),
	.w5(32'h3ba4dc6e),
	.w6(32'hbb0bf4da),
	.w7(32'hbae3cf5b),
	.w8(32'h3b6c862b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ecb7f),
	.w1(32'h3ba95630),
	.w2(32'hbb33b31d),
	.w3(32'h3b6cd811),
	.w4(32'h3bad16af),
	.w5(32'hbb441994),
	.w6(32'h3be70109),
	.w7(32'h3bd36fb8),
	.w8(32'hba81263b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081122),
	.w1(32'hb99e3da8),
	.w2(32'hba8feaa0),
	.w3(32'hbb62e57e),
	.w4(32'hbaa9e356),
	.w5(32'hba978b02),
	.w6(32'hbb6b7497),
	.w7(32'hbafa66ea),
	.w8(32'hbb4f78ef),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb431f3),
	.w1(32'hbbf5a504),
	.w2(32'hbb9d3969),
	.w3(32'hbace1095),
	.w4(32'hbbabfccf),
	.w5(32'hbb7fedf4),
	.w6(32'hbb781900),
	.w7(32'hbadd9a99),
	.w8(32'hbb141e27),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee1621),
	.w1(32'hba42d851),
	.w2(32'h3a29a5ed),
	.w3(32'hba9470e2),
	.w4(32'hba5cc741),
	.w5(32'hbacc195b),
	.w6(32'h39c4ed91),
	.w7(32'h3aba686e),
	.w8(32'h3b893661),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a396422),
	.w1(32'h3a24ae9e),
	.w2(32'h3a7d3630),
	.w3(32'h3adbf349),
	.w4(32'h3b2e7d6d),
	.w5(32'h3a8a2304),
	.w6(32'h3ac68360),
	.w7(32'h3b1f5302),
	.w8(32'h3a70165b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dec067),
	.w1(32'h3a05b8f5),
	.w2(32'h3a600265),
	.w3(32'h39ec7465),
	.w4(32'h3a82134a),
	.w5(32'h398b9051),
	.w6(32'h39639b30),
	.w7(32'h3a9015af),
	.w8(32'hbb04ee44),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab722fd),
	.w1(32'h3b10d012),
	.w2(32'h3aab3be8),
	.w3(32'hba8ba647),
	.w4(32'h37f0b73b),
	.w5(32'h3b522e7e),
	.w6(32'h3a8320be),
	.w7(32'hb93b7f1d),
	.w8(32'h3b2bc0d9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4181b6),
	.w1(32'hbbaafcf4),
	.w2(32'hbb71027c),
	.w3(32'h3a8fc606),
	.w4(32'hbb283281),
	.w5(32'hba84f742),
	.w6(32'h3aba80a8),
	.w7(32'h39bbbbd6),
	.w8(32'hbb046aba),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc119d),
	.w1(32'h3b06ed42),
	.w2(32'h3b42491a),
	.w3(32'h3b459832),
	.w4(32'h3b535a34),
	.w5(32'h3b63e011),
	.w6(32'h3b393cef),
	.w7(32'h3b5d539e),
	.w8(32'h3b44a312),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18cc5a),
	.w1(32'h3c0175b9),
	.w2(32'h38e7e334),
	.w3(32'hbb030016),
	.w4(32'h3baff3f2),
	.w5(32'h3b061e70),
	.w6(32'hbb749ea5),
	.w7(32'h3a9590e0),
	.w8(32'hbba1815d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c560b),
	.w1(32'hbb5d995a),
	.w2(32'h3abc26f5),
	.w3(32'hbad97732),
	.w4(32'hbac4e6ab),
	.w5(32'h39d25a69),
	.w6(32'hbb0d40a2),
	.w7(32'hbac52363),
	.w8(32'hb8ca83dd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45694b),
	.w1(32'h39dcdf23),
	.w2(32'h3a07125e),
	.w3(32'h3ad1998d),
	.w4(32'hba5e44f3),
	.w5(32'hbaa62d93),
	.w6(32'hbb7b4c0c),
	.w7(32'h3a0414e6),
	.w8(32'h3a874835),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6639),
	.w1(32'hbb5854c2),
	.w2(32'hbb2b4fa3),
	.w3(32'hbb3afa5d),
	.w4(32'hbc19f9b7),
	.w5(32'hbb2d87d8),
	.w6(32'h3b848620),
	.w7(32'hbb4f8641),
	.w8(32'hbb197b10),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08781b),
	.w1(32'hbc0a7d9e),
	.w2(32'hbc45cccb),
	.w3(32'h3ad02aea),
	.w4(32'h3b81d4ea),
	.w5(32'hbb08471e),
	.w6(32'h3b28dc41),
	.w7(32'h3b950de2),
	.w8(32'h3c1696e7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e85e6),
	.w1(32'hba0909a6),
	.w2(32'h3a6cf324),
	.w3(32'h3b1595e1),
	.w4(32'h3ba9f880),
	.w5(32'hbb7b2e84),
	.w6(32'h3bcfd676),
	.w7(32'hbbdaafb3),
	.w8(32'hbbf9c88e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0924ba),
	.w1(32'hbaa70a9b),
	.w2(32'h3b6d4953),
	.w3(32'h3a4f8571),
	.w4(32'h3b6ab269),
	.w5(32'h3ac15a23),
	.w6(32'hbaf88827),
	.w7(32'h3b1860ce),
	.w8(32'hbc0c3581),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9add05e),
	.w1(32'hbc438777),
	.w2(32'hbc5314c5),
	.w3(32'h3b04e0df),
	.w4(32'h3aaf92af),
	.w5(32'h3b805ea7),
	.w6(32'h3b6e9d1b),
	.w7(32'h3bd4ac77),
	.w8(32'hbb556f4f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc757d59),
	.w1(32'hbcc32cc0),
	.w2(32'hbbccdee5),
	.w3(32'hbbdc1053),
	.w4(32'hbcc58449),
	.w5(32'hbb492054),
	.w6(32'h3b620ddb),
	.w7(32'hbb09161a),
	.w8(32'h3b3be485),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119b4d),
	.w1(32'hbba21e0f),
	.w2(32'h3c4a63c5),
	.w3(32'hbb287dfd),
	.w4(32'hb914dc5f),
	.w5(32'h3bb735a7),
	.w6(32'h3bf7ec5e),
	.w7(32'h3bc9f7ed),
	.w8(32'h39e5cd83),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ee6ba),
	.w1(32'hbadb3041),
	.w2(32'h3b0ecf34),
	.w3(32'h3b82ea2e),
	.w4(32'h3aca8fa2),
	.w5(32'h3bffaa0f),
	.w6(32'h3a84c803),
	.w7(32'h3c1162e7),
	.w8(32'h3c39d60e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba608fc0),
	.w1(32'hbaf12e77),
	.w2(32'h3c487cc5),
	.w3(32'h3b142834),
	.w4(32'h3abaf0b4),
	.w5(32'h3c0a52cf),
	.w6(32'h3bdeb2f7),
	.w7(32'h3bc702fe),
	.w8(32'h3b031258),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f54df),
	.w1(32'hbaa25642),
	.w2(32'hbbf41a03),
	.w3(32'h3c086870),
	.w4(32'hbc35939a),
	.w5(32'h3c29661c),
	.w6(32'h3ba074c5),
	.w7(32'hbc30c710),
	.w8(32'h3c6518eb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ac9cd),
	.w1(32'hbc602d83),
	.w2(32'h3b0283ad),
	.w3(32'h3b0e1d00),
	.w4(32'hbb99f0e0),
	.w5(32'h3bc02dcd),
	.w6(32'h3c9d92fb),
	.w7(32'h3a6d06a9),
	.w8(32'h3bd3e411),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc449a54),
	.w1(32'hbaeabcec),
	.w2(32'hbc176f99),
	.w3(32'hbc5d1c87),
	.w4(32'hbc0cf264),
	.w5(32'hbcafe07e),
	.w6(32'h3bade727),
	.w7(32'h3ad0e32a),
	.w8(32'hbcf50309),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9f878),
	.w1(32'h3c2c2c4b),
	.w2(32'h3bd6065a),
	.w3(32'hbcb7c900),
	.w4(32'h3b8926de),
	.w5(32'hb9ea24cf),
	.w6(32'hbce95e58),
	.w7(32'hbcaa53cd),
	.w8(32'h3a46d322),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44260a),
	.w1(32'h3c024c71),
	.w2(32'h3c395bab),
	.w3(32'h3aace18d),
	.w4(32'h3c06bee1),
	.w5(32'hbb3d5443),
	.w6(32'hbbb7e175),
	.w7(32'h3c245dbb),
	.w8(32'hbbcd38f1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac8d97),
	.w1(32'h3a42558e),
	.w2(32'hbbc95ee2),
	.w3(32'hbc4c7ba7),
	.w4(32'hbc4d29e4),
	.w5(32'hbb37e843),
	.w6(32'hbc0f0997),
	.w7(32'hbc28d8c2),
	.w8(32'h3bc650f9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2becc8),
	.w1(32'hbc0d6c4d),
	.w2(32'hbbfc39a0),
	.w3(32'hb9ec7926),
	.w4(32'hbb0f7a29),
	.w5(32'h3c0a8267),
	.w6(32'hbb2698bd),
	.w7(32'hba8a53bd),
	.w8(32'h3c94f17f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf9641),
	.w1(32'hbcad66f8),
	.w2(32'hbb76613f),
	.w3(32'hba5d40c8),
	.w4(32'hbc371a5b),
	.w5(32'h3bcff949),
	.w6(32'h3ca8954a),
	.w7(32'h3b7e171a),
	.w8(32'h3c3222fd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7869b),
	.w1(32'hbb426c6d),
	.w2(32'h3bb792b8),
	.w3(32'h3c146b31),
	.w4(32'h3c3131ca),
	.w5(32'h3bdc4def),
	.w6(32'h3c279d00),
	.w7(32'h3c181286),
	.w8(32'h3c50119b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fcff4),
	.w1(32'h3b97d05a),
	.w2(32'h3aac05b6),
	.w3(32'hbaee2ad1),
	.w4(32'h3b0b3900),
	.w5(32'hba29472c),
	.w6(32'h3b92c9e3),
	.w7(32'h3b1bf46d),
	.w8(32'hbb5bdc24),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca231),
	.w1(32'hbc5789e2),
	.w2(32'h3b7642b6),
	.w3(32'hbb97a465),
	.w4(32'hbc338145),
	.w5(32'h3c1667ad),
	.w6(32'hbc34f82f),
	.w7(32'hbc6d1043),
	.w8(32'h3be93ca9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ed84),
	.w1(32'hbc8bc8bd),
	.w2(32'hbb833977),
	.w3(32'h3c2d4b23),
	.w4(32'hbc3f53fc),
	.w5(32'h3b722977),
	.w6(32'hba9b97fc),
	.w7(32'h3a53c32c),
	.w8(32'h3be537e6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6a53),
	.w1(32'hbc3d224b),
	.w2(32'hbc86eaee),
	.w3(32'h3b8e66c3),
	.w4(32'hbbeaeca1),
	.w5(32'hbd02fe6c),
	.w6(32'h3c12a2ae),
	.w7(32'h37f45780),
	.w8(32'hbcc04bbb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0171db),
	.w1(32'hbcac8c31),
	.w2(32'h3b82d0cd),
	.w3(32'hbd59e095),
	.w4(32'hbcebb884),
	.w5(32'h3be6b02e),
	.w6(32'hbd3f27a2),
	.w7(32'hbd06bbb5),
	.w8(32'h3b317bd9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12ed09),
	.w1(32'h3bda8001),
	.w2(32'h3bb6103f),
	.w3(32'h3c386082),
	.w4(32'h3b24dfe4),
	.w5(32'h3c6a55ff),
	.w6(32'h3c1ed6d9),
	.w7(32'h3b8c0f62),
	.w8(32'h3c927ee0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37f55b),
	.w1(32'hbbaaa7e5),
	.w2(32'hbb209a66),
	.w3(32'hbb28a61e),
	.w4(32'hbc24ed9a),
	.w5(32'h3b2d5e9e),
	.w6(32'hbaff8547),
	.w7(32'hbb4bbe52),
	.w8(32'hb99a240c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfe743),
	.w1(32'hbb4effb9),
	.w2(32'h3bdaee3b),
	.w3(32'h3b8f035d),
	.w4(32'h3b11411c),
	.w5(32'h3c22d549),
	.w6(32'hba41263b),
	.w7(32'hb908a336),
	.w8(32'hbb110710),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8acee7b),
	.w1(32'hbc6e2dce),
	.w2(32'hbb217b5f),
	.w3(32'h3c5cf103),
	.w4(32'hb9cf966d),
	.w5(32'h3af5fc85),
	.w6(32'h3bf8b7a9),
	.w7(32'h3becf524),
	.w8(32'h3a70d3d1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f7ba),
	.w1(32'hbb7781dc),
	.w2(32'hbaffa1dc),
	.w3(32'hb9ede07e),
	.w4(32'h3b372f92),
	.w5(32'hbb9bcaf6),
	.w6(32'hbb240b2c),
	.w7(32'hbc41f58a),
	.w8(32'hbc2ca65e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1ee39),
	.w1(32'hbc026672),
	.w2(32'hbc06d314),
	.w3(32'hbbdd68e4),
	.w4(32'hbc64064b),
	.w5(32'hbc04a891),
	.w6(32'hbc26ec83),
	.w7(32'hbbe67b73),
	.w8(32'hbca28ac6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0ea2b),
	.w1(32'hbc9c6dfb),
	.w2(32'h3b37063a),
	.w3(32'hbc7ccb0e),
	.w4(32'hbca734a5),
	.w5(32'hbb8d34ab),
	.w6(32'hbbcac476),
	.w7(32'hbc1a1d27),
	.w8(32'hbc091b5f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe865da),
	.w1(32'hbbf1610a),
	.w2(32'hba30fd5e),
	.w3(32'h3b2623e7),
	.w4(32'h3c5f4603),
	.w5(32'h3b131bfd),
	.w6(32'h3aea6e79),
	.w7(32'h3cebe840),
	.w8(32'h3c9e979b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae18ccd),
	.w1(32'h3bc1faab),
	.w2(32'hbbc441c0),
	.w3(32'h3bab5136),
	.w4(32'h3c326a03),
	.w5(32'hbc8c9aa0),
	.w6(32'h3d0076dd),
	.w7(32'h3d084252),
	.w8(32'hbb443078),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc751fe3),
	.w1(32'hbb98d19d),
	.w2(32'hbc0de3b6),
	.w3(32'hbd12e834),
	.w4(32'hbca3a398),
	.w5(32'hbc579508),
	.w6(32'hbc5b7e57),
	.w7(32'hbc81fd39),
	.w8(32'hbc99736c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394eeba7),
	.w1(32'hbb0573de),
	.w2(32'hbc0bc741),
	.w3(32'hbb8e7063),
	.w4(32'h37320f33),
	.w5(32'hbbd1698b),
	.w6(32'hbd045e0b),
	.w7(32'hbc8b19c3),
	.w8(32'h3b80f60c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c071e),
	.w1(32'hbc33de8c),
	.w2(32'hbba565dd),
	.w3(32'hbbf46624),
	.w4(32'hbc3a59e4),
	.w5(32'h3ac32fa2),
	.w6(32'hbafe581c),
	.w7(32'hbb3c0394),
	.w8(32'h3a9444e3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac492f),
	.w1(32'hbb476f9a),
	.w2(32'hb89cc7c0),
	.w3(32'hbb95515e),
	.w4(32'hbbb0fc0e),
	.w5(32'hbbe1e813),
	.w6(32'hbab70ac1),
	.w7(32'hbb6270f1),
	.w8(32'hbbade160),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a71623),
	.w1(32'h3b612b63),
	.w2(32'h3b6482d2),
	.w3(32'hbc3859dd),
	.w4(32'hbc544e2e),
	.w5(32'h3ba6d588),
	.w6(32'hbb44d273),
	.w7(32'hb99e73bf),
	.w8(32'h3b089598),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491a3e),
	.w1(32'hbb058ef8),
	.w2(32'h3b6f83b3),
	.w3(32'h3b76b26c),
	.w4(32'h3c20d941),
	.w5(32'h3c1b3714),
	.w6(32'h3a4ed861),
	.w7(32'h3bd090c8),
	.w8(32'h3bc2b420),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa46b),
	.w1(32'hbbc92e55),
	.w2(32'hbc553a41),
	.w3(32'h3c42d5ec),
	.w4(32'h3b8bc9bc),
	.w5(32'hbb603582),
	.w6(32'h3c63d486),
	.w7(32'h3c342b7c),
	.w8(32'h3c080fdc),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf86e2),
	.w1(32'hbca276e0),
	.w2(32'h3b3ec5f9),
	.w3(32'hbaa9a47a),
	.w4(32'hbc710359),
	.w5(32'h38ce857c),
	.w6(32'h3c9bb77b),
	.w7(32'h3968fad1),
	.w8(32'h3c152c99),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17611f),
	.w1(32'h3ac3df34),
	.w2(32'hbb8919c7),
	.w3(32'h3c0459c4),
	.w4(32'h3c359301),
	.w5(32'hbbaa645e),
	.w6(32'h3c1f923f),
	.w7(32'h3b8a2bfc),
	.w8(32'hbbcb5379),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149684),
	.w1(32'hbb65eef6),
	.w2(32'hbb04f394),
	.w3(32'hbb544d0d),
	.w4(32'h3b8ab804),
	.w5(32'hbbc40b20),
	.w6(32'hbba1163b),
	.w7(32'hba7dcef0),
	.w8(32'hbc4e7699),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863aa10),
	.w1(32'h3c003aff),
	.w2(32'hba95b4a0),
	.w3(32'hbc0c001e),
	.w4(32'hbab037e9),
	.w5(32'h3a459fc1),
	.w6(32'hbc8b43d0),
	.w7(32'hbc6714ab),
	.w8(32'h3bfa5155),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc34e2),
	.w1(32'hba0e5ee9),
	.w2(32'hba98ac15),
	.w3(32'hbd24a595),
	.w4(32'hbc8620bc),
	.w5(32'hbb269dcf),
	.w6(32'hbd0ca405),
	.w7(32'hbce6fd13),
	.w8(32'hbbccdee0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9f45e),
	.w1(32'hbc0aae29),
	.w2(32'h3b02ef40),
	.w3(32'h3b9913e4),
	.w4(32'h3ab2e2de),
	.w5(32'h3afceea7),
	.w6(32'h3b64fe6c),
	.w7(32'h3c036f09),
	.w8(32'h3c3f592b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7809e),
	.w1(32'hbbbaf65c),
	.w2(32'hbb3406c5),
	.w3(32'h3b610fd7),
	.w4(32'h3b68f31b),
	.w5(32'h39593392),
	.w6(32'h3bdc2d6d),
	.w7(32'h3b33f894),
	.w8(32'h3bc7febd),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd878f),
	.w1(32'hbc25f63d),
	.w2(32'h394fdf28),
	.w3(32'h3bd9c329),
	.w4(32'hbb7f6788),
	.w5(32'h3afe850b),
	.w6(32'h3c782103),
	.w7(32'hbab42692),
	.w8(32'hbb1da791),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7672a3),
	.w1(32'hbc2e7230),
	.w2(32'hbc3af37d),
	.w3(32'hbb0b9314),
	.w4(32'hbc246bb4),
	.w5(32'h3a2ee978),
	.w6(32'hbb6b627b),
	.w7(32'hbc041d6a),
	.w8(32'h3ba1603f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca9a54),
	.w1(32'hbcf99eb5),
	.w2(32'hbb5ee76b),
	.w3(32'hbc2021eb),
	.w4(32'hbcaa6423),
	.w5(32'h3b116b17),
	.w6(32'h3c151a9b),
	.w7(32'h3b36950b),
	.w8(32'h3bb48dd7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1edb),
	.w1(32'hbbc70c40),
	.w2(32'hbaac4383),
	.w3(32'h3b9e90a8),
	.w4(32'h3b20e5b4),
	.w5(32'h3bfec3b8),
	.w6(32'h3aa23ffb),
	.w7(32'hbaf2c91d),
	.w8(32'h3a87e863),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4e1f4),
	.w1(32'hb75e0ea0),
	.w2(32'h3c0a9766),
	.w3(32'h3c0442d8),
	.w4(32'h3bc940d0),
	.w5(32'h3a2af95f),
	.w6(32'hb9bda2c9),
	.w7(32'h39a014e2),
	.w8(32'hbc91b9f6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7add8),
	.w1(32'hbc4ca77b),
	.w2(32'hbac8686d),
	.w3(32'hbb798c7e),
	.w4(32'hbb0bfe54),
	.w5(32'h3a40d542),
	.w6(32'hbb6d4e22),
	.w7(32'h3c303e22),
	.w8(32'h3aceec51),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf94439),
	.w1(32'hbb2335f6),
	.w2(32'hbb958787),
	.w3(32'hbb710cd8),
	.w4(32'h3bbe0c91),
	.w5(32'hbbb7ab7f),
	.w6(32'hbc144113),
	.w7(32'h3b3640b4),
	.w8(32'hbc46a37e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5feb73),
	.w1(32'hbbcbf100),
	.w2(32'h3a362451),
	.w3(32'hbc9faa48),
	.w4(32'hbc1d8f8e),
	.w5(32'h3bc08fe3),
	.w6(32'hbcab697c),
	.w7(32'hbc738745),
	.w8(32'h3c1de162),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c84c),
	.w1(32'hbb048db6),
	.w2(32'h3c3503b9),
	.w3(32'h3c1503d4),
	.w4(32'h3b9d46b9),
	.w5(32'h3b49df2b),
	.w6(32'h3c83fff5),
	.w7(32'h3c3cdcff),
	.w8(32'h3b80e937),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2a5b1),
	.w1(32'hba4a75d0),
	.w2(32'hbc756036),
	.w3(32'h3a842eeb),
	.w4(32'hbb880a46),
	.w5(32'hbbe59bcc),
	.w6(32'h3c46089c),
	.w7(32'hbb012a44),
	.w8(32'hbadee73d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5770ea),
	.w1(32'hbc997b40),
	.w2(32'h3b04cb3b),
	.w3(32'hbccb2217),
	.w4(32'hbc9da638),
	.w5(32'h3b0e5776),
	.w6(32'hbcb58bc7),
	.w7(32'hbcb0e4bc),
	.w8(32'h3b0c5d56),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0fc13),
	.w1(32'hbbc75a35),
	.w2(32'h3b2eb386),
	.w3(32'hbbe29236),
	.w4(32'hbba07a22),
	.w5(32'h3c3d4cb7),
	.w6(32'hb6d8da68),
	.w7(32'hbc103698),
	.w8(32'h3c570e20),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397b7a),
	.w1(32'hbc0b108f),
	.w2(32'hbaf55e34),
	.w3(32'h3ca4176c),
	.w4(32'h3c17a6e1),
	.w5(32'hba740219),
	.w6(32'h3cc99c0b),
	.w7(32'h3c5cfedf),
	.w8(32'hbacef7dd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd59de3),
	.w1(32'hbbc24387),
	.w2(32'hbb91d39f),
	.w3(32'h3c374ba9),
	.w4(32'h3bd04e2a),
	.w5(32'h39994f89),
	.w6(32'h3cb8d0ef),
	.w7(32'h3c58636c),
	.w8(32'h3abc3950),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc112ab4),
	.w1(32'hbbd4d634),
	.w2(32'h3add256e),
	.w3(32'hbb65267a),
	.w4(32'hbb8a1cf7),
	.w5(32'h3c6536f0),
	.w6(32'hbb1d6ec9),
	.w7(32'hbab14341),
	.w8(32'h3c1edbac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ecf9d),
	.w1(32'h3904b529),
	.w2(32'hbb3ac419),
	.w3(32'h3b8eea85),
	.w4(32'h3be43ce6),
	.w5(32'h3ad3ed50),
	.w6(32'h3a831088),
	.w7(32'h3bda10f2),
	.w8(32'h3bd75605),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28fc5b),
	.w1(32'hbcedc2c4),
	.w2(32'hbc4933e6),
	.w3(32'hbb3a3099),
	.w4(32'hbc508f2e),
	.w5(32'hbc21b579),
	.w6(32'h3b993bfb),
	.w7(32'hbc704b30),
	.w8(32'hbc6fb5a8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808d12),
	.w1(32'hbbd7ba0a),
	.w2(32'h3b5ca683),
	.w3(32'hba8ca82f),
	.w4(32'hbc467c57),
	.w5(32'hbbc47c10),
	.w6(32'h3b98cd63),
	.w7(32'hbb9c9582),
	.w8(32'hbca9bdbf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6eb13a),
	.w1(32'h3cacf736),
	.w2(32'hbb37e256),
	.w3(32'h3ba4421c),
	.w4(32'h3cab8b0f),
	.w5(32'hba0d4de8),
	.w6(32'hbca7720c),
	.w7(32'h3a865fec),
	.w8(32'h3a74aac8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff09e3),
	.w1(32'hbbd10232),
	.w2(32'hb80ef3ba),
	.w3(32'hbb8c8ff1),
	.w4(32'hbb377f28),
	.w5(32'h3a91b3ab),
	.w6(32'hbba9a01c),
	.w7(32'hbb425b59),
	.w8(32'h3876b21a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba51420),
	.w1(32'hbb8e1619),
	.w2(32'h3b83ef56),
	.w3(32'h3b3f4ff3),
	.w4(32'h3ae3d315),
	.w5(32'hbb0955ff),
	.w6(32'hba8650a1),
	.w7(32'h3a091041),
	.w8(32'hbb8935c4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e9ebc),
	.w1(32'hbbecdbab),
	.w2(32'h3aa30909),
	.w3(32'hbaaa8faf),
	.w4(32'hbbb88df1),
	.w5(32'h3c0eecca),
	.w6(32'hbb9867d1),
	.w7(32'h3ba1c054),
	.w8(32'h3be48815),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65b838),
	.w1(32'h3b61ab72),
	.w2(32'hbc8c743a),
	.w3(32'h3b875ff2),
	.w4(32'h3985752b),
	.w5(32'hbcc7a161),
	.w6(32'h3c0dff45),
	.w7(32'h3a06eeb9),
	.w8(32'hbbddf35d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1ea4b),
	.w1(32'hbcced67d),
	.w2(32'h3bd56579),
	.w3(32'hbd0575fe),
	.w4(32'hbd110d45),
	.w5(32'hba4bdd03),
	.w6(32'hbc4b1d18),
	.w7(32'hbc610608),
	.w8(32'h3c23bf11),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbae75b),
	.w1(32'hbc079055),
	.w2(32'h3ba58d0b),
	.w3(32'h3b23c336),
	.w4(32'hbb92675a),
	.w5(32'h3b7c2820),
	.w6(32'h3ad708d1),
	.w7(32'hbb26f3ed),
	.w8(32'hbbe01956),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04171a),
	.w1(32'hbc0f5a90),
	.w2(32'hbb8584c1),
	.w3(32'h3c1e66fd),
	.w4(32'h3b8ee894),
	.w5(32'h3b73a903),
	.w6(32'h391a34e8),
	.w7(32'h3bb27bb6),
	.w8(32'h3bf15442),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5b0e9),
	.w1(32'hbbe59fba),
	.w2(32'hbbb81839),
	.w3(32'hbbfb3ca7),
	.w4(32'hbc38d94a),
	.w5(32'hba8ca8f7),
	.w6(32'hbb67d093),
	.w7(32'hbcab67a6),
	.w8(32'hbaab9096),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb27d08),
	.w1(32'hbaf26640),
	.w2(32'hb9d7e002),
	.w3(32'hbad424d4),
	.w4(32'hbbb58ffe),
	.w5(32'h3be7dfea),
	.w6(32'hba4adcdc),
	.w7(32'h3ba08f9a),
	.w8(32'hbba2d797),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accf4bc),
	.w1(32'h3b06a0f8),
	.w2(32'h3c08940b),
	.w3(32'h3c202023),
	.w4(32'h3c41fc7b),
	.w5(32'h38de4437),
	.w6(32'h3b197ba3),
	.w7(32'hbb26e224),
	.w8(32'h39aa34b0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2b08f),
	.w1(32'hbc8d7b61),
	.w2(32'h3c3a70e7),
	.w3(32'h3b267fc4),
	.w4(32'hbbb1dda7),
	.w5(32'h3b8295b0),
	.w6(32'h3c1a65fd),
	.w7(32'h3bb72829),
	.w8(32'h3b710064),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85bbf8),
	.w1(32'hbbb7805e),
	.w2(32'hba90110d),
	.w3(32'hbb9cb8b9),
	.w4(32'hbc2b3f14),
	.w5(32'h3b957cfe),
	.w6(32'h3b3759a5),
	.w7(32'hbb84e0f0),
	.w8(32'h3c0dcb4b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eea144),
	.w1(32'hbb944681),
	.w2(32'hbb132f7c),
	.w3(32'h3ab57ecb),
	.w4(32'hbb8a5b21),
	.w5(32'hbb79f363),
	.w6(32'h3c1a9648),
	.w7(32'h3ad8cf97),
	.w8(32'hbbca64df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6b4f),
	.w1(32'hbc05153a),
	.w2(32'hbbb92aab),
	.w3(32'h3b31e6e0),
	.w4(32'h3c0b07ae),
	.w5(32'h3b857bf7),
	.w6(32'h3b20acf9),
	.w7(32'h3c2a8d84),
	.w8(32'h3c046a22),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22f887),
	.w1(32'hbc5c9ba1),
	.w2(32'hbb9c5bcc),
	.w3(32'hba0e0109),
	.w4(32'hba954483),
	.w5(32'hbb1d1ea8),
	.w6(32'h3b106050),
	.w7(32'h3bca5643),
	.w8(32'hbb86c40f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0abd9a),
	.w1(32'hbc13164f),
	.w2(32'hbbb8132a),
	.w3(32'hbc8b4320),
	.w4(32'hbc022d58),
	.w5(32'hbbb7fa0e),
	.w6(32'hbc29b06b),
	.w7(32'hbc1c5f05),
	.w8(32'hbbdfa131),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c221),
	.w1(32'hbb8c3d90),
	.w2(32'hbbf7dcad),
	.w3(32'hbc6371f9),
	.w4(32'hbc3c00ba),
	.w5(32'hbbe42193),
	.w6(32'hbb26bacc),
	.w7(32'hbc2c1c6a),
	.w8(32'hbc1027ec),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc484a57),
	.w1(32'hbbb3abfb),
	.w2(32'hba9a6d6d),
	.w3(32'hbc1e2e43),
	.w4(32'hbc4588bb),
	.w5(32'h3be4b02c),
	.w6(32'hbc025b63),
	.w7(32'hbbf09568),
	.w8(32'h3b32e152),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2304a3),
	.w1(32'hbbda90f1),
	.w2(32'h3b5f9990),
	.w3(32'hbbea2232),
	.w4(32'hbc343212),
	.w5(32'h3b861322),
	.w6(32'h3b715214),
	.w7(32'hbb9f5989),
	.w8(32'h3b2ab2f7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c050),
	.w1(32'hbb355e93),
	.w2(32'h3a76fc92),
	.w3(32'hbafa679c),
	.w4(32'hbbb1ffef),
	.w5(32'hbb63ce7c),
	.w6(32'hba016dc4),
	.w7(32'hbb1303dc),
	.w8(32'hbb5fb3aa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7d196),
	.w1(32'hbbe7cc57),
	.w2(32'hbc05092b),
	.w3(32'hbbffee1d),
	.w4(32'hbc2db3e0),
	.w5(32'hbbb78788),
	.w6(32'hbbe78265),
	.w7(32'hbc958056),
	.w8(32'hbc02cc14),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e6b19),
	.w1(32'hbc7a572a),
	.w2(32'hbb60603c),
	.w3(32'hbcb1e1cb),
	.w4(32'hbc8c8836),
	.w5(32'hbc683801),
	.w6(32'hbc3ca5f5),
	.w7(32'hbc8ae377),
	.w8(32'hbc5aab64),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324407),
	.w1(32'hbc3b9670),
	.w2(32'h3a45df65),
	.w3(32'hbcfaf69c),
	.w4(32'hbd03f65e),
	.w5(32'hbc0f3919),
	.w6(32'hbce03041),
	.w7(32'hbcc748fb),
	.w8(32'hbaa105e4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53147e),
	.w1(32'h3bde1057),
	.w2(32'h3c8c3248),
	.w3(32'hbcadc498),
	.w4(32'hbc117789),
	.w5(32'h3c5a9e20),
	.w6(32'hbbf43375),
	.w7(32'hbb8d18c3),
	.w8(32'hbc614e35),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbe05c),
	.w1(32'h3c2f6d3c),
	.w2(32'hbbcda2d8),
	.w3(32'h3d0bb9e4),
	.w4(32'h3cbc4855),
	.w5(32'hbca97324),
	.w6(32'hba2cd2b1),
	.w7(32'h3c029301),
	.w8(32'hbc29e6d8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60bde5),
	.w1(32'hbc343863),
	.w2(32'h3be001f4),
	.w3(32'hbd0fbe06),
	.w4(32'hbcec498d),
	.w5(32'h3c13fba1),
	.w6(32'hbc816100),
	.w7(32'hbc521de5),
	.w8(32'hb9dc0669),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d349),
	.w1(32'hbb8e8caf),
	.w2(32'hbbcea597),
	.w3(32'h3c2e55a9),
	.w4(32'h3c4f0742),
	.w5(32'hbb4629fa),
	.w6(32'h3c37f02b),
	.w7(32'h3b70ebf5),
	.w8(32'h393d5ed9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2acbca),
	.w1(32'hbbafdf57),
	.w2(32'h3b751470),
	.w3(32'h3b8ed872),
	.w4(32'h3baaab7b),
	.w5(32'hbb76aa37),
	.w6(32'h3b6e3a7f),
	.w7(32'h3bd1018e),
	.w8(32'h3b828fd6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432fcb),
	.w1(32'hba7eec85),
	.w2(32'h3b43e9a3),
	.w3(32'hbbcb911c),
	.w4(32'hbba855a2),
	.w5(32'h388f05d6),
	.w6(32'h3ac296a9),
	.w7(32'hbb257367),
	.w8(32'hbb4e3ea4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8064cc),
	.w1(32'hb9f84c26),
	.w2(32'hb88204b2),
	.w3(32'h3b382e57),
	.w4(32'h3875f2bc),
	.w5(32'hbab4324f),
	.w6(32'hb9b8c61e),
	.w7(32'h3ab78a5f),
	.w8(32'hbb34c3e1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab85e9d),
	.w1(32'h3b85bd17),
	.w2(32'hbb6f6baa),
	.w3(32'h3b68460e),
	.w4(32'h3b75b1e8),
	.w5(32'hbb31ea44),
	.w6(32'hbaf09a2b),
	.w7(32'h3b3c8e0c),
	.w8(32'hbbeb6049),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba87f6),
	.w1(32'hbca0c1c9),
	.w2(32'hbaae873e),
	.w3(32'hbc1f10c9),
	.w4(32'h3ae962a3),
	.w5(32'hbbfbb2f2),
	.w6(32'h3c0cca66),
	.w7(32'h3c8d7d44),
	.w8(32'hbb7392e0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe7e95),
	.w1(32'hbbaa4f50),
	.w2(32'h38887bbf),
	.w3(32'hbbc8b208),
	.w4(32'hba156c4c),
	.w5(32'hbbdcc4de),
	.w6(32'hbb996be2),
	.w7(32'hba2cdba9),
	.w8(32'hb9a72da4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cd69e),
	.w1(32'hbb98c280),
	.w2(32'hbb81c524),
	.w3(32'hbbdbb57e),
	.w4(32'h39e2f22e),
	.w5(32'h3b0e02db),
	.w6(32'hbb2230b8),
	.w7(32'hbba19c7f),
	.w8(32'h3c333280),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cb6c9),
	.w1(32'h3b10da17),
	.w2(32'h3c36db5e),
	.w3(32'h3bb14fba),
	.w4(32'hb9e89a95),
	.w5(32'h3b501a14),
	.w6(32'h3bbdf876),
	.w7(32'h3b3bad02),
	.w8(32'h3bf48bb1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b6e73),
	.w1(32'h3bac5a67),
	.w2(32'h3afbf946),
	.w3(32'h3c413fcc),
	.w4(32'h3b5c1646),
	.w5(32'h3b6a353e),
	.w6(32'h3c09447c),
	.w7(32'h3bbfe266),
	.w8(32'h3bf6f5a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87e09c),
	.w1(32'hbc9bc680),
	.w2(32'hbb967d25),
	.w3(32'h3c123a52),
	.w4(32'hbbeba621),
	.w5(32'hbc99114f),
	.w6(32'h3cbf7e64),
	.w7(32'h3c1e83e3),
	.w8(32'hbc6bdf08),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc737614),
	.w1(32'hbcc25f2d),
	.w2(32'h3b9d3d84),
	.w3(32'hbc8f23e5),
	.w4(32'hbc4c2151),
	.w5(32'h3a9db8b6),
	.w6(32'hbc8db6c1),
	.w7(32'hbc880fe9),
	.w8(32'h3c1876a5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc217dd),
	.w1(32'hbb871671),
	.w2(32'hbabb124a),
	.w3(32'h3c259947),
	.w4(32'h3b26b6ce),
	.w5(32'hbac4a9ac),
	.w6(32'h3c7f9beb),
	.w7(32'h3c06a9d4),
	.w8(32'h3a74cc80),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54ff34),
	.w1(32'h3ae79361),
	.w2(32'hbc1b0a1d),
	.w3(32'h3ad9758f),
	.w4(32'h3ba6765c),
	.w5(32'hbc8f3398),
	.w6(32'h3b3544a3),
	.w7(32'h3b0cd29b),
	.w8(32'hbc2af1f4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3af67d),
	.w1(32'hbc6ec0e0),
	.w2(32'hbba75b9a),
	.w3(32'hbbb00e27),
	.w4(32'hbc4e92d3),
	.w5(32'hbbc434b0),
	.w6(32'hbbee0835),
	.w7(32'hbbf995a6),
	.w8(32'hb9cf40ae),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7418a9),
	.w1(32'hbb1aa1ae),
	.w2(32'h3add6fe1),
	.w3(32'hbc87baa5),
	.w4(32'hbc0d052e),
	.w5(32'h3b6f0988),
	.w6(32'hbbc20b6e),
	.w7(32'hbb50bfdf),
	.w8(32'h3bb661e1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a505),
	.w1(32'hbc283924),
	.w2(32'hbb4b94c1),
	.w3(32'h38c7c2b9),
	.w4(32'hbbf6bb0f),
	.w5(32'hbb9aa43f),
	.w6(32'h3ad560ab),
	.w7(32'hba7eca3d),
	.w8(32'hbab4e0c3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f500),
	.w1(32'hbc42b97a),
	.w2(32'hbb977b52),
	.w3(32'hbc6a570b),
	.w4(32'hbc1be936),
	.w5(32'h3881d687),
	.w6(32'hbb628d4f),
	.w7(32'hbb6eb9c4),
	.w8(32'hbb7ed069),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdd0cc),
	.w1(32'hbcbf3cc7),
	.w2(32'h3b96ee85),
	.w3(32'hbba62f2c),
	.w4(32'hbc204370),
	.w5(32'h3bfd2e31),
	.w6(32'h3be4de5c),
	.w7(32'h390d2562),
	.w8(32'h3c2174cc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f932f),
	.w1(32'h3c8a2f37),
	.w2(32'hbb818861),
	.w3(32'h3c3b8d59),
	.w4(32'h3c9d48e0),
	.w5(32'hbbd38090),
	.w6(32'h3bef5dd7),
	.w7(32'h3c041b40),
	.w8(32'hbbd5fe27),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1091d8),
	.w1(32'h3c11c839),
	.w2(32'hbb53b966),
	.w3(32'h3a68d39b),
	.w4(32'h3c196504),
	.w5(32'hbb3dbc25),
	.w6(32'hbbb37b18),
	.w7(32'hb9413e67),
	.w8(32'h3b18c300),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b21e5),
	.w1(32'hbc12a4b7),
	.w2(32'h3bcc6ced),
	.w3(32'hbc0b7252),
	.w4(32'hbc5142f3),
	.w5(32'h3bd0a764),
	.w6(32'h3bbc9e54),
	.w7(32'h3a8e4211),
	.w8(32'h3b8e681c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b704293),
	.w1(32'h383e42b3),
	.w2(32'h3b8110a1),
	.w3(32'h3bdc1b95),
	.w4(32'h3b7fc8c0),
	.w5(32'hbaee8101),
	.w6(32'hba8a6d9c),
	.w7(32'hb9e5df05),
	.w8(32'hbb959c0c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd352f),
	.w1(32'h3aae1583),
	.w2(32'h3c840e9e),
	.w3(32'h3b38574e),
	.w4(32'h3b4ba90a),
	.w5(32'h3c78517e),
	.w6(32'hbaff5467),
	.w7(32'h3b1aa857),
	.w8(32'hbb9a3767),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17d8c),
	.w1(32'hba2876f4),
	.w2(32'hbbda6811),
	.w3(32'h3ca9c2fb),
	.w4(32'h3b14b968),
	.w5(32'hbc86cb07),
	.w6(32'hbb88852d),
	.w7(32'hbabdbec4),
	.w8(32'hbbd00899),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3496af),
	.w1(32'h3b3f56cb),
	.w2(32'h3a99f980),
	.w3(32'hbd2c4ec8),
	.w4(32'hbcee99bd),
	.w5(32'hba96ccfe),
	.w6(32'hbced72a0),
	.w7(32'hbcf3406e),
	.w8(32'hbb28e176),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2998d9),
	.w1(32'h3b95102a),
	.w2(32'h39d3efc3),
	.w3(32'h3b5946a3),
	.w4(32'h3bd11023),
	.w5(32'h3b277475),
	.w6(32'hbac867d2),
	.w7(32'h3b403121),
	.w8(32'h3bf877cb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44585c),
	.w1(32'hbbb95ae5),
	.w2(32'hba642746),
	.w3(32'h3bb4a423),
	.w4(32'h3aba4150),
	.w5(32'h3b31fe5f),
	.w6(32'h3c3820b0),
	.w7(32'h3ae6a94a),
	.w8(32'hbb589f0f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959a763),
	.w1(32'hb7eccdf2),
	.w2(32'h3b992b5d),
	.w3(32'hba71a7b1),
	.w4(32'h3a997b35),
	.w5(32'h3c94a6d3),
	.w6(32'hbb8bc56c),
	.w7(32'hbbaf18a0),
	.w8(32'h3be64c34),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd04682),
	.w1(32'hb950fa08),
	.w2(32'h3c1d6c60),
	.w3(32'h3ce57291),
	.w4(32'h3cca6dbe),
	.w5(32'h3bc54a0c),
	.w6(32'h3c7ed4cb),
	.w7(32'h3c98f77c),
	.w8(32'h3c103127),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52de69),
	.w1(32'hbb012b4e),
	.w2(32'h3ba6e823),
	.w3(32'hb88f708f),
	.w4(32'hbc1c6ada),
	.w5(32'h3bf48687),
	.w6(32'h3b39a0f7),
	.w7(32'hbbc1d805),
	.w8(32'h3bef74a3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d2124),
	.w1(32'h3b1b7d7a),
	.w2(32'hbc0a6eb9),
	.w3(32'h3ae04628),
	.w4(32'h3b3d94b2),
	.w5(32'hbb9215aa),
	.w6(32'h382a2d79),
	.w7(32'hbb1434b7),
	.w8(32'h3c860f77),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b0186),
	.w1(32'hbbb6c573),
	.w2(32'h3b651cca),
	.w3(32'h3c0532fb),
	.w4(32'hbb403577),
	.w5(32'h3bae3146),
	.w6(32'h3c35385a),
	.w7(32'h3b85e8bc),
	.w8(32'h3b168e33),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9018bf),
	.w1(32'hbb9b0d66),
	.w2(32'hba9a5537),
	.w3(32'h3c28294f),
	.w4(32'h3b8df4bd),
	.w5(32'hba4eb099),
	.w6(32'h3b13018f),
	.w7(32'h3b9b6a77),
	.w8(32'hbb8d1000),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c2285d),
	.w1(32'hb9601803),
	.w2(32'hbb5bcf50),
	.w3(32'hbb47e50b),
	.w4(32'hbb0da03b),
	.w5(32'h3b0616bc),
	.w6(32'hbbf8073c),
	.w7(32'hba6607a9),
	.w8(32'h3a283492),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ab40f),
	.w1(32'hbc11361b),
	.w2(32'h3a0ef05f),
	.w3(32'hb9bfed83),
	.w4(32'hbbf73b5b),
	.w5(32'hbaa553b0),
	.w6(32'h3b84053d),
	.w7(32'h3a67a128),
	.w8(32'h3a82961d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c126307),
	.w1(32'h3b134819),
	.w2(32'h39c5b031),
	.w3(32'h3c452e1a),
	.w4(32'h3bd0c4b7),
	.w5(32'h3983b721),
	.w6(32'h3be59f27),
	.w7(32'h3b9a85ba),
	.w8(32'h3a9baad1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f0c82),
	.w1(32'h3a5c0c1e),
	.w2(32'h3b4b7321),
	.w3(32'h3a00a798),
	.w4(32'hb93228a3),
	.w5(32'h3b383160),
	.w6(32'h3a4cc003),
	.w7(32'hba4e0f9a),
	.w8(32'h3974b966),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf74c9),
	.w1(32'h3be24182),
	.w2(32'h3bda66b6),
	.w3(32'h3a8016c1),
	.w4(32'h3b58ed23),
	.w5(32'hbb0f10d9),
	.w6(32'h3b16852e),
	.w7(32'h3baa8812),
	.w8(32'hbbda80c1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48c6f2),
	.w1(32'h3ac49d4e),
	.w2(32'h3ad93a77),
	.w3(32'h3c842740),
	.w4(32'h3cc4d2a9),
	.w5(32'hba164f5e),
	.w6(32'hbc1991d4),
	.w7(32'hbbb942c4),
	.w8(32'h3af0000d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8229d1),
	.w1(32'hbb0aab74),
	.w2(32'hba4a3c23),
	.w3(32'hb9a73b20),
	.w4(32'hbb4ec623),
	.w5(32'h3b549474),
	.w6(32'h3b6ac201),
	.w7(32'h3b0c9e94),
	.w8(32'hbc1240ec),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675002),
	.w1(32'h3c1cbd9d),
	.w2(32'hbc08a2ce),
	.w3(32'h3c29a0bb),
	.w4(32'h3c60d443),
	.w5(32'h3bb026d5),
	.w6(32'hbbaf2cb1),
	.w7(32'hbb201971),
	.w8(32'hb84ccf4a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0185),
	.w1(32'hbab173fa),
	.w2(32'hbb27a3b1),
	.w3(32'h3c0a4bb3),
	.w4(32'h3ac89252),
	.w5(32'hbb2a3173),
	.w6(32'h3b0d4329),
	.w7(32'h3c00dc7e),
	.w8(32'hba517a1f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08d5b8),
	.w1(32'hbae8fd94),
	.w2(32'hba382a15),
	.w3(32'hbaa28039),
	.w4(32'hba802321),
	.w5(32'h3b092555),
	.w6(32'hb98ce7bf),
	.w7(32'h3a5ee2a0),
	.w8(32'h3c3fa9a2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b19e0),
	.w1(32'hbba0f3e8),
	.w2(32'h39ac4720),
	.w3(32'h3b7e3209),
	.w4(32'hbbffb68d),
	.w5(32'h3aa19b15),
	.w6(32'h3c327aaa),
	.w7(32'hba3b4935),
	.w8(32'hba5de5b6),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab21b79),
	.w1(32'h3b17312f),
	.w2(32'hbc5cc4f6),
	.w3(32'h3add5b20),
	.w4(32'h3b9fe8e2),
	.w5(32'hbc1c025a),
	.w6(32'h38aa75fd),
	.w7(32'h3aef88cb),
	.w8(32'h3b02e2ce),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2f58d),
	.w1(32'hbbdfa5de),
	.w2(32'h3b3b8a9f),
	.w3(32'h3b933227),
	.w4(32'h3b5d5239),
	.w5(32'hbb258513),
	.w6(32'h3b93d0ae),
	.w7(32'hbc0f0729),
	.w8(32'hbb15d237),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009bd6),
	.w1(32'h3b609b86),
	.w2(32'h3ba0c9fe),
	.w3(32'h3aecedaa),
	.w4(32'h3b57c7b6),
	.w5(32'hbbeda570),
	.w6(32'h3ba86b3e),
	.w7(32'h3bab38b2),
	.w8(32'hbc04572b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d723),
	.w1(32'h3bdd29f4),
	.w2(32'h3aed5490),
	.w3(32'hbc30f5fc),
	.w4(32'hbbe20fec),
	.w5(32'h3989fb17),
	.w6(32'hbb8adf57),
	.w7(32'hbbc8343b),
	.w8(32'h39eb2a31),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa47fce),
	.w1(32'h3b4e076f),
	.w2(32'h3a5c12da),
	.w3(32'h3b6dac71),
	.w4(32'h3bde90a4),
	.w5(32'h3a310b84),
	.w6(32'h3bb920c0),
	.w7(32'h3c783685),
	.w8(32'h38ed52fd),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba35f9f),
	.w1(32'h39beb39b),
	.w2(32'h3c3f282e),
	.w3(32'h3bca2675),
	.w4(32'hba5847ed),
	.w5(32'h3b60a794),
	.w6(32'hbb4537c7),
	.w7(32'hba10db2d),
	.w8(32'h3b5ef34f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8acad),
	.w1(32'h39f30dda),
	.w2(32'hbb39ae9a),
	.w3(32'h3953d4ee),
	.w4(32'hbb9bc625),
	.w5(32'hbc57d88b),
	.w6(32'h3b9b13d6),
	.w7(32'h3ba1de0c),
	.w8(32'hbc6e7823),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03054d),
	.w1(32'h3bc5c6d0),
	.w2(32'h3a93cda8),
	.w3(32'hbab556c7),
	.w4(32'h3bdc42f0),
	.w5(32'h3abe75a5),
	.w6(32'hbca520ef),
	.w7(32'hbc15f1f6),
	.w8(32'hbb010a74),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a95d9),
	.w1(32'h3b53dafc),
	.w2(32'h3b90e45e),
	.w3(32'h3b3ff2bd),
	.w4(32'hb9d04e18),
	.w5(32'hbb85c690),
	.w6(32'h39002200),
	.w7(32'hba58458a),
	.w8(32'hbba49ded),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e99c),
	.w1(32'hbc109cc0),
	.w2(32'hbc3513ad),
	.w3(32'h3afcd156),
	.w4(32'hb9688b75),
	.w5(32'hba0aede5),
	.w6(32'hbb9e308b),
	.w7(32'hbb902b8b),
	.w8(32'hba8273af),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba534f3),
	.w1(32'hbc6ca994),
	.w2(32'hbb6257ed),
	.w3(32'h3b9c14aa),
	.w4(32'h3c0b2c82),
	.w5(32'hbc173a9a),
	.w6(32'h3c14e827),
	.w7(32'h3c82a98f),
	.w8(32'hbbe218d7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0e514),
	.w1(32'hbc1f3498),
	.w2(32'hba29cbee),
	.w3(32'hbc66a1dd),
	.w4(32'hbc40f7d1),
	.w5(32'hbb85f025),
	.w6(32'hbc31e7ac),
	.w7(32'hbb2c95a0),
	.w8(32'hbb938f06),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15e326),
	.w1(32'hbba7fcfe),
	.w2(32'h3b442cb7),
	.w3(32'hbbbd3c68),
	.w4(32'hbba2856e),
	.w5(32'h3b6d056a),
	.w6(32'hbb7f291d),
	.w7(32'hbb52d73a),
	.w8(32'h3a40ef1d),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b688bd1),
	.w1(32'h3b93ed60),
	.w2(32'h3868ebd0),
	.w3(32'h3bd8eacd),
	.w4(32'h3ba61b09),
	.w5(32'hba8c11e2),
	.w6(32'h3bb4adc5),
	.w7(32'h3bb86abe),
	.w8(32'hbc39c4d5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedbb9c),
	.w1(32'h3c11d243),
	.w2(32'hbbb06995),
	.w3(32'hbb2eacce),
	.w4(32'hbb31f75d),
	.w5(32'h3af3b981),
	.w6(32'hbc462680),
	.w7(32'hbbfc5487),
	.w8(32'h3be4c0b2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30fcd8),
	.w1(32'hbc555641),
	.w2(32'hbae0c41f),
	.w3(32'h3b45128c),
	.w4(32'h3a96fbcb),
	.w5(32'h3c2227b0),
	.w6(32'h3befb702),
	.w7(32'h3bf2d087),
	.w8(32'h3bc83d89),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7fed2),
	.w1(32'hbc3712bf),
	.w2(32'hbc008bb9),
	.w3(32'h3bf05005),
	.w4(32'h38fdbfad),
	.w5(32'h3bb13757),
	.w6(32'h3a06cfb2),
	.w7(32'h3b232f73),
	.w8(32'h3c1dfe94),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bd7d7),
	.w1(32'hbca5cb23),
	.w2(32'h3b6b9986),
	.w3(32'h3c136a17),
	.w4(32'hbb814ad0),
	.w5(32'hba54eeef),
	.w6(32'h3bc59804),
	.w7(32'h3bd21a78),
	.w8(32'hbbac6cbf),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ed260),
	.w1(32'hbb344d41),
	.w2(32'h3c36284e),
	.w3(32'hbac700e4),
	.w4(32'hba390e8b),
	.w5(32'hbba9430b),
	.w6(32'hbc3bf30f),
	.w7(32'hbc60627d),
	.w8(32'h3bc4e098),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d3e2a),
	.w1(32'h3c4143e3),
	.w2(32'hbc2ebf98),
	.w3(32'hbb6b908c),
	.w4(32'h3b25dc3c),
	.w5(32'h3be214ef),
	.w6(32'h3a9f9290),
	.w7(32'h3b3b3562),
	.w8(32'h3c11173a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11fd8a),
	.w1(32'hbbe5d29d),
	.w2(32'hbb221658),
	.w3(32'h3b6926ca),
	.w4(32'h3ab42a54),
	.w5(32'h3b94465d),
	.w6(32'h3bd02eff),
	.w7(32'h3b80099f),
	.w8(32'hbbff4971),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3304),
	.w1(32'hbc05fbd4),
	.w2(32'hba02ca46),
	.w3(32'h3c407d51),
	.w4(32'h3c14b914),
	.w5(32'hbb88022c),
	.w6(32'h3a37e1c3),
	.w7(32'h3bf9b26f),
	.w8(32'hbbd6537e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c2db),
	.w1(32'h3bb853a0),
	.w2(32'hb9d21054),
	.w3(32'hbb6a62c4),
	.w4(32'hbaa3c21f),
	.w5(32'h3a3ea078),
	.w6(32'hbb4373d6),
	.w7(32'h3ab16bd2),
	.w8(32'hbb75ae41),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe5609),
	.w1(32'h3be6993d),
	.w2(32'h3c328f77),
	.w3(32'hba41277c),
	.w4(32'h3bb0056b),
	.w5(32'hbb80305a),
	.w6(32'hbbced22e),
	.w7(32'hba3d483e),
	.w8(32'hbb4db378),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce4f6),
	.w1(32'h3b1afa97),
	.w2(32'hba11efcf),
	.w3(32'hbb04a9c8),
	.w4(32'hba66dec7),
	.w5(32'hbc022c68),
	.w6(32'hb9b30965),
	.w7(32'hbb99c1f5),
	.w8(32'hbbea566c),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41b40c),
	.w1(32'h3bde4ccf),
	.w2(32'hbab569b1),
	.w3(32'h3b0d52a8),
	.w4(32'hbbcda7a4),
	.w5(32'hbb4d3b00),
	.w6(32'h3b654674),
	.w7(32'hbb101524),
	.w8(32'hbb9631a2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44e216),
	.w1(32'hbbb2155e),
	.w2(32'h3a507ada),
	.w3(32'h3ac56278),
	.w4(32'h3a84eebb),
	.w5(32'hb7987500),
	.w6(32'h3a038977),
	.w7(32'h3b135a98),
	.w8(32'hbb0eeeb2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b306085),
	.w1(32'h3b9ac3bf),
	.w2(32'hba709350),
	.w3(32'hbb931103),
	.w4(32'hbb38fb40),
	.w5(32'hbbc56bf4),
	.w6(32'hbbebe16f),
	.w7(32'hbb25ce8f),
	.w8(32'hba6eea6f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7ebe),
	.w1(32'h3aac1c2b),
	.w2(32'hbbda0219),
	.w3(32'hbb856ae8),
	.w4(32'hbb50040e),
	.w5(32'h3ac69bab),
	.w6(32'hba1fdd50),
	.w7(32'h3b104116),
	.w8(32'h3c0ec63d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefc1a8),
	.w1(32'h3acbbf36),
	.w2(32'hbbd534a5),
	.w3(32'hb9d675e6),
	.w4(32'hba0fd609),
	.w5(32'hbae51daf),
	.w6(32'h3c0359e4),
	.w7(32'h3c1f4f81),
	.w8(32'h3a866fa1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67369c),
	.w1(32'hbc046431),
	.w2(32'h3add0424),
	.w3(32'hbacec4e6),
	.w4(32'hba673c48),
	.w5(32'h3ad79774),
	.w6(32'h39c0d948),
	.w7(32'h3a4679ff),
	.w8(32'hba006652),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec7540),
	.w1(32'h39a9b073),
	.w2(32'hbbd10a32),
	.w3(32'h3ac3b818),
	.w4(32'h393417b0),
	.w5(32'hbb568fe9),
	.w6(32'h3b0a4fc0),
	.w7(32'h3a3b0546),
	.w8(32'hbc43582d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5ab11),
	.w1(32'hbb723413),
	.w2(32'hbac23e4f),
	.w3(32'hbacdeee8),
	.w4(32'h3a345438),
	.w5(32'h3b540615),
	.w6(32'hbbc937e5),
	.w7(32'hbba07dfb),
	.w8(32'h3c07b14c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf410fa),
	.w1(32'hbbd4a4be),
	.w2(32'h3aebe0a6),
	.w3(32'h3b7e4ecc),
	.w4(32'h382f3883),
	.w5(32'hba364622),
	.w6(32'h3bbe5518),
	.w7(32'h3b46d71b),
	.w8(32'hba89007d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf0626),
	.w1(32'hba4be175),
	.w2(32'h39b5b9e5),
	.w3(32'h3aae2776),
	.w4(32'hbacf3647),
	.w5(32'hbba02cc0),
	.w6(32'h3a13c9d9),
	.w7(32'hbabfed4c),
	.w8(32'hbaf81218),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2af5a),
	.w1(32'hbad60d53),
	.w2(32'hbb9d018d),
	.w3(32'hbb9a493b),
	.w4(32'hbbb6fb05),
	.w5(32'hbba32c4e),
	.w6(32'h39623669),
	.w7(32'h3b31b014),
	.w8(32'hbbc38cc1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabad1cf),
	.w1(32'h37de618f),
	.w2(32'hbb4651b4),
	.w3(32'hbbae2a79),
	.w4(32'h3a9e3696),
	.w5(32'hbb584530),
	.w6(32'hbc035e05),
	.w7(32'hbbb1cddc),
	.w8(32'hbc3be80a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059ad0),
	.w1(32'h38f816f7),
	.w2(32'hbbbf9f63),
	.w3(32'hbc038ea5),
	.w4(32'hbc0524d2),
	.w5(32'hb93c5dcd),
	.w6(32'hbc3fe35c),
	.w7(32'hbbcacd84),
	.w8(32'h3c682e2a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41ea0d),
	.w1(32'hbc03f029),
	.w2(32'hbb19415c),
	.w3(32'h3a98ea98),
	.w4(32'hbafbe19b),
	.w5(32'hbb0868b8),
	.w6(32'h3c936754),
	.w7(32'h3c6a9b7f),
	.w8(32'hbb81afb0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d6380),
	.w1(32'hbab4a317),
	.w2(32'hb9daf68b),
	.w3(32'h3ae9299c),
	.w4(32'h3ad10e42),
	.w5(32'hbb18a71e),
	.w6(32'hba81037b),
	.w7(32'h3ac03352),
	.w8(32'hbbdeb802),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7dac0),
	.w1(32'h3bebfc3e),
	.w2(32'hbaa83aae),
	.w3(32'hb88dd3de),
	.w4(32'hbb1945c6),
	.w5(32'h3c630a28),
	.w6(32'hbbc8bc74),
	.w7(32'hbb57d79c),
	.w8(32'h3c392e21),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2d013),
	.w1(32'hbc5075c8),
	.w2(32'hb90781e5),
	.w3(32'h3c152655),
	.w4(32'hbbc40ce0),
	.w5(32'h3c2f5d78),
	.w6(32'h3be31347),
	.w7(32'h3be7dac3),
	.w8(32'h3bd05b9c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a91c1),
	.w1(32'hbc351e67),
	.w2(32'hbab8a773),
	.w3(32'h3ae0cef5),
	.w4(32'h3af83357),
	.w5(32'hbbeb4d89),
	.w6(32'hbaefaaf9),
	.w7(32'h3bd472cb),
	.w8(32'hbc4eaad0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9b98a),
	.w1(32'hbb90b043),
	.w2(32'h3b463f58),
	.w3(32'hbb78e1b8),
	.w4(32'h3b175525),
	.w5(32'h3a036571),
	.w6(32'hbb89ffac),
	.w7(32'hbbaf33c5),
	.w8(32'h3b0d9c57),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8112ed),
	.w1(32'hba8d8e0a),
	.w2(32'hba6fbee4),
	.w3(32'hb8391fdd),
	.w4(32'hb9f2afed),
	.w5(32'h399eaaf6),
	.w6(32'hba3756bb),
	.w7(32'hba1ae029),
	.w8(32'h3adee082),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1e64f),
	.w1(32'hbbd82131),
	.w2(32'h38fab290),
	.w3(32'h3a30d68b),
	.w4(32'hbb3c36dc),
	.w5(32'hba807711),
	.w6(32'h3bd195cc),
	.w7(32'h3bad60d4),
	.w8(32'h3ae6c4a7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab729),
	.w1(32'hb756fd8d),
	.w2(32'hbb6d10a5),
	.w3(32'h394ee492),
	.w4(32'hbb449efa),
	.w5(32'hbbd42923),
	.w6(32'h3b64a31f),
	.w7(32'h3ab4155d),
	.w8(32'hbb9dc8b2),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dc99),
	.w1(32'hbaf8e7da),
	.w2(32'hbb9bcdff),
	.w3(32'hbc0d71a1),
	.w4(32'hbb2ceede),
	.w5(32'hbc079272),
	.w6(32'h3b2dc024),
	.w7(32'hbaf44afd),
	.w8(32'hbbc2f927),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b802d78),
	.w1(32'hbb1f5af7),
	.w2(32'hba09fbdd),
	.w3(32'hbc31cb5c),
	.w4(32'hbb4a7e4d),
	.w5(32'h3aa22c2c),
	.w6(32'hbc325be8),
	.w7(32'hbb59f419),
	.w8(32'hbb640f53),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86effe),
	.w1(32'hbbaf2f0a),
	.w2(32'hbc1273ff),
	.w3(32'hbb7ffc1c),
	.w4(32'hbba30d1a),
	.w5(32'h3aa9b97b),
	.w6(32'hbbc7d4d2),
	.w7(32'hbb97f9c4),
	.w8(32'h3a0dec6e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331fc6),
	.w1(32'hbbf5364c),
	.w2(32'hba170aa6),
	.w3(32'hbbc79633),
	.w4(32'hbb19c987),
	.w5(32'h3b14d044),
	.w6(32'h39f58836),
	.w7(32'hba329526),
	.w8(32'hbaa80d1c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1075b2),
	.w1(32'hbbb4637f),
	.w2(32'h3bb232e6),
	.w3(32'h3bb19970),
	.w4(32'hba644f5b),
	.w5(32'h3b4fbb48),
	.w6(32'h3b26e1f8),
	.w7(32'h3b64eb88),
	.w8(32'h3b944ef4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a0106),
	.w1(32'h3aacd56a),
	.w2(32'hbbf84052),
	.w3(32'h3b7f611e),
	.w4(32'h3b4f90ef),
	.w5(32'hbb36a083),
	.w6(32'h3b87c361),
	.w7(32'h3ba63314),
	.w8(32'h3ba9903d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc525907),
	.w1(32'hbc74a2ed),
	.w2(32'hbb8d96ee),
	.w3(32'h39ea4aae),
	.w4(32'hb9db88ff),
	.w5(32'hbb01c2e5),
	.w6(32'h3b8ba322),
	.w7(32'h3b0c2a77),
	.w8(32'hbb1bdbf7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d3ec6),
	.w1(32'hbb829283),
	.w2(32'hbb8147e6),
	.w3(32'h39ae279d),
	.w4(32'h3b0a1359),
	.w5(32'hba3fe0b4),
	.w6(32'hbc12a81c),
	.w7(32'hbc07f808),
	.w8(32'hbabc73fe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cbee5),
	.w1(32'hbb310e04),
	.w2(32'h3ad9ad19),
	.w3(32'h3b17b7da),
	.w4(32'h3b1a091d),
	.w5(32'hbbeec1d8),
	.w6(32'h3950bc70),
	.w7(32'hb8a721a7),
	.w8(32'hba3bf7a3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3925d3),
	.w1(32'h3c11ab20),
	.w2(32'h3b9f76ce),
	.w3(32'hba5f6b8f),
	.w4(32'h3ae1884e),
	.w5(32'h3b39a8e7),
	.w6(32'h3b0a7647),
	.w7(32'h39cf077f),
	.w8(32'h3b85dd4b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc19dfa),
	.w1(32'h3c096ce7),
	.w2(32'h3bdff273),
	.w3(32'h3bab5907),
	.w4(32'h3bd0e6d8),
	.w5(32'h3a38d821),
	.w6(32'h3b27c302),
	.w7(32'h3b291ba7),
	.w8(32'h3b113237),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc21fe),
	.w1(32'h3bdffcf4),
	.w2(32'h3b14b014),
	.w3(32'hbb26baf8),
	.w4(32'hbb0934e6),
	.w5(32'h3c06ff4b),
	.w6(32'h3aab1795),
	.w7(32'hbaf16869),
	.w8(32'h3c0e1a1d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e843f),
	.w1(32'hbbe72246),
	.w2(32'h3bd4b368),
	.w3(32'hbb1f63be),
	.w4(32'hbba79abc),
	.w5(32'h3bd17dd6),
	.w6(32'h3b80c647),
	.w7(32'h3b16fa93),
	.w8(32'hbb205097),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b4612),
	.w1(32'h3b38b7f0),
	.w2(32'h3a38667c),
	.w3(32'h3c47c28c),
	.w4(32'hbc5071c4),
	.w5(32'h3baaec57),
	.w6(32'hbbd409b5),
	.w7(32'hbc21fa5e),
	.w8(32'hbb4137e7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae85360),
	.w1(32'hbbbea28b),
	.w2(32'hbbce0209),
	.w3(32'h3c035c2b),
	.w4(32'h3c14fea4),
	.w5(32'hbbe77339),
	.w6(32'hbb0b0247),
	.w7(32'hbba6a034),
	.w8(32'hbc0f71cd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22bac6),
	.w1(32'hbbfc9650),
	.w2(32'h3bd2fe51),
	.w3(32'hbb6f6965),
	.w4(32'hbbcfa000),
	.w5(32'h3c65ed2a),
	.w6(32'hbc12d5c0),
	.w7(32'hbbac0ac4),
	.w8(32'h3c5b628d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfde5c1),
	.w1(32'hbbfe64a4),
	.w2(32'h3b3e539d),
	.w3(32'h3c40f951),
	.w4(32'hb906400c),
	.w5(32'hba9cf87f),
	.w6(32'h3c1086f9),
	.w7(32'h3add4b8c),
	.w8(32'hb9d0941d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6549a),
	.w1(32'h3aa8a95f),
	.w2(32'hba663c50),
	.w3(32'h3b406ee8),
	.w4(32'h3bb2eb8b),
	.w5(32'hbc183710),
	.w6(32'h3b997365),
	.w7(32'h3b931dcc),
	.w8(32'hbc51a25a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50a5f8),
	.w1(32'h3baeb858),
	.w2(32'h3b45d94d),
	.w3(32'hbaa688c4),
	.w4(32'h3c3ed450),
	.w5(32'h3b9b00c2),
	.w6(32'hbbefa6fc),
	.w7(32'hbbc0b43c),
	.w8(32'hbbcf7b71),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e674b),
	.w1(32'h3b7ff1b2),
	.w2(32'hbb22ab22),
	.w3(32'h3be23e98),
	.w4(32'h3ba287b7),
	.w5(32'hbaaa9ae8),
	.w6(32'hbbd9223a),
	.w7(32'hbc1bc5f1),
	.w8(32'h39bfb4f9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b631b38),
	.w1(32'hbc6aa521),
	.w2(32'hbb380b9c),
	.w3(32'h3c0606a5),
	.w4(32'hbb94cc4e),
	.w5(32'h3acd8619),
	.w6(32'h3a722d6d),
	.w7(32'h38e8d25a),
	.w8(32'h3aa39454),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807ed2),
	.w1(32'hbbfb0e9c),
	.w2(32'hbc40cd11),
	.w3(32'h39dade10),
	.w4(32'hbba59606),
	.w5(32'hbb92b527),
	.w6(32'hbb20992b),
	.w7(32'hbb020244),
	.w8(32'h3a25c637),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b3138),
	.w1(32'hbc1487eb),
	.w2(32'hbb9ae134),
	.w3(32'hbb91638d),
	.w4(32'hbb83f6ac),
	.w5(32'hba6cca95),
	.w6(32'h3b871c4b),
	.w7(32'hbb785959),
	.w8(32'hbaf39338),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5cf8b),
	.w1(32'hbc5299d6),
	.w2(32'hbb8e1b9c),
	.w3(32'hbb0d702f),
	.w4(32'hbc1ddf81),
	.w5(32'h3a3be84d),
	.w6(32'hbb2ba786),
	.w7(32'hbb133518),
	.w8(32'h3b039bb5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5953b0),
	.w1(32'hbb4c9b9b),
	.w2(32'h3bafdcea),
	.w3(32'hba4d855f),
	.w4(32'h3a9ad77e),
	.w5(32'h3a82bed5),
	.w6(32'h3ab367d4),
	.w7(32'h3b524dd8),
	.w8(32'hbb431b9f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e31e),
	.w1(32'h3a389c92),
	.w2(32'hbb6412cc),
	.w3(32'h3ab65407),
	.w4(32'h3bcc1b8d),
	.w5(32'hbbb78c35),
	.w6(32'hbb9f5f3c),
	.w7(32'hbbcc87c8),
	.w8(32'hbc06fdea),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e0b2),
	.w1(32'hb9f48774),
	.w2(32'h3c26bbee),
	.w3(32'hbb9db5c3),
	.w4(32'hbbd8b916),
	.w5(32'h3bcdabfe),
	.w6(32'hbbd02c13),
	.w7(32'hbb2d43a3),
	.w8(32'hbc9198ba),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c3bb5),
	.w1(32'h3c1d85e5),
	.w2(32'h3a83eeba),
	.w3(32'h3c03038f),
	.w4(32'h3c25cd9b),
	.w5(32'hbbb49d05),
	.w6(32'hbc7f7515),
	.w7(32'hbc4ca0cc),
	.w8(32'hbbeb1b6c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012fb5),
	.w1(32'hbb77acb6),
	.w2(32'hba8cc897),
	.w3(32'hbbb0f8de),
	.w4(32'h3b8e0e54),
	.w5(32'h3b511c50),
	.w6(32'hbb9a8f5d),
	.w7(32'hbb37d279),
	.w8(32'hba849e09),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29fe68),
	.w1(32'hbbb61aeb),
	.w2(32'hbbf761e8),
	.w3(32'h3b0de5f4),
	.w4(32'hbbb74654),
	.w5(32'hbb0e2720),
	.w6(32'h3bb06600),
	.w7(32'h3c052d4d),
	.w8(32'h3c11b8f8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab08c20),
	.w1(32'hbbb9f446),
	.w2(32'h3c24a519),
	.w3(32'h3bb833c2),
	.w4(32'hba01cda2),
	.w5(32'hbbe529b3),
	.w6(32'h3c372fae),
	.w7(32'h3bb096a8),
	.w8(32'hbc50ada4),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafc07a),
	.w1(32'h3c3a394d),
	.w2(32'hb926e4f7),
	.w3(32'h3b5d716d),
	.w4(32'h3c42bf38),
	.w5(32'hbab20702),
	.w6(32'hbc2101fc),
	.w7(32'hbbcdaf75),
	.w8(32'h3bfb24e5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0a755),
	.w1(32'hbc296e07),
	.w2(32'h3b21abab),
	.w3(32'h3a739e99),
	.w4(32'hbbf5407d),
	.w5(32'h3ad5609a),
	.w6(32'h3c08c4f8),
	.w7(32'h3b20eb7a),
	.w8(32'h3b0b02c9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba616c),
	.w1(32'h3a3c5264),
	.w2(32'hb8c7f38c),
	.w3(32'h3a0de0b0),
	.w4(32'h3b07817b),
	.w5(32'h3b111452),
	.w6(32'hb87a5bef),
	.w7(32'h3a316fa1),
	.w8(32'hbb06d582),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f608f),
	.w1(32'h3b35ce99),
	.w2(32'h39c2a66f),
	.w3(32'h3bce8210),
	.w4(32'h3c5e9e99),
	.w5(32'hbb33fcd2),
	.w6(32'hbb48905f),
	.w7(32'hbb9392f1),
	.w8(32'hbb1712e2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38532a4d),
	.w1(32'hbb022f50),
	.w2(32'h3b0b9ce9),
	.w3(32'hbb05b121),
	.w4(32'hba16e23d),
	.w5(32'h3b7e83e0),
	.w6(32'hbb767b64),
	.w7(32'hbb96d7e9),
	.w8(32'hbc05ea70),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87eb30),
	.w1(32'hbbc457df),
	.w2(32'hbbe68150),
	.w3(32'h3c530784),
	.w4(32'h3b2b45f6),
	.w5(32'hbb9217cb),
	.w6(32'hbb7848b8),
	.w7(32'hbac9e871),
	.w8(32'hbc180b6e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09ee9e),
	.w1(32'h3c37f269),
	.w2(32'hbb83c3fd),
	.w3(32'h3b05a13f),
	.w4(32'h3bff7fcf),
	.w5(32'hbbb5533c),
	.w6(32'hbb16f50c),
	.w7(32'h3ab6206c),
	.w8(32'hbb80ae5d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44331b),
	.w1(32'h3b326b31),
	.w2(32'hb987f9ef),
	.w3(32'h3b78221d),
	.w4(32'hba006c01),
	.w5(32'h3a415588),
	.w6(32'hbb359733),
	.w7(32'hba9e5ba7),
	.w8(32'h3a6f33f7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c903c),
	.w1(32'hbb4864ff),
	.w2(32'hbb5b7f82),
	.w3(32'h39917415),
	.w4(32'h3a0c0765),
	.w5(32'h375315e1),
	.w6(32'h3b89100c),
	.w7(32'h3b4e3d3d),
	.w8(32'h3b28ce23),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b02d2),
	.w1(32'hbb2c2842),
	.w2(32'hbc2d6e30),
	.w3(32'h3ad891ee),
	.w4(32'hb965e094),
	.w5(32'h3b64cbaa),
	.w6(32'h3aa52f2c),
	.w7(32'h3b00ae20),
	.w8(32'h3b851346),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ffbe3),
	.w1(32'hbc480641),
	.w2(32'hba4026bf),
	.w3(32'h3bcd878b),
	.w4(32'h3b9a2ef7),
	.w5(32'hbad6bfaa),
	.w6(32'hba5a6e36),
	.w7(32'h3acf9776),
	.w8(32'hbb983090),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba737ebb),
	.w1(32'hb9148f72),
	.w2(32'hbc1ff3f0),
	.w3(32'hbb11d760),
	.w4(32'hbb034623),
	.w5(32'h3bb02353),
	.w6(32'hbba2fb20),
	.w7(32'hbb81f39a),
	.w8(32'h3c23f42f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf8930f),
	.w1(32'hbcaa295a),
	.w2(32'hbb940137),
	.w3(32'h3ada2d1e),
	.w4(32'hbb4cf2c2),
	.w5(32'hbb4eecc5),
	.w6(32'h3bf834fa),
	.w7(32'h3b1ac818),
	.w8(32'hbc088142),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc022c8),
	.w1(32'hbbdb610c),
	.w2(32'hbb4e7f67),
	.w3(32'hbb00b8d0),
	.w4(32'hbba35713),
	.w5(32'hbb9ed5b2),
	.w6(32'hbb83b6d4),
	.w7(32'hbba6bf68),
	.w8(32'hbbe4cd8c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3f363),
	.w1(32'hbbaf9a6c),
	.w2(32'h3ad5543e),
	.w3(32'hbb4f2637),
	.w4(32'hbad090a2),
	.w5(32'h3b9d27a6),
	.w6(32'hbc8e7d32),
	.w7(32'hbb33bc23),
	.w8(32'h395fb546),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule