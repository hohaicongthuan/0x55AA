module layer_10_featuremap_117(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeba16),
	.w1(32'hbb683f4d),
	.w2(32'hbbca46af),
	.w3(32'hb88b454a),
	.w4(32'hba665614),
	.w5(32'hba96b004),
	.w6(32'hb9823188),
	.w7(32'hbadd7575),
	.w8(32'hba443d9a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3ea22),
	.w1(32'h3995425c),
	.w2(32'h3aa2f981),
	.w3(32'hbabd3d43),
	.w4(32'hba0117be),
	.w5(32'h3a43ebea),
	.w6(32'hba944cf3),
	.w7(32'h398f6cac),
	.w8(32'h37114f36),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2d2f0),
	.w1(32'h3a59f81d),
	.w2(32'h3a77cfd7),
	.w3(32'h3aab410f),
	.w4(32'h3a8e5aef),
	.w5(32'h3aa90114),
	.w6(32'hba41aad3),
	.w7(32'hbacd253c),
	.w8(32'hbae10a6b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16b457),
	.w1(32'h3b61ccd6),
	.w2(32'h3b612316),
	.w3(32'h3a9b85ef),
	.w4(32'hba5f33fe),
	.w5(32'hba195abd),
	.w6(32'h3a3bae84),
	.w7(32'hba3a8246),
	.w8(32'h3afe346f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2aa5),
	.w1(32'hbb2fdcf6),
	.w2(32'h3ab8e779),
	.w3(32'h3b3ed212),
	.w4(32'hbb67d0a7),
	.w5(32'hb9dd6aed),
	.w6(32'h3a6107ed),
	.w7(32'h3acb544e),
	.w8(32'h3af6bfc6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe49ea),
	.w1(32'hb8125ea0),
	.w2(32'h3aa382ab),
	.w3(32'h3a557366),
	.w4(32'hbaf584df),
	.w5(32'hb8dc2291),
	.w6(32'h3a786210),
	.w7(32'h3a6eb379),
	.w8(32'h3a4f4f86),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a485799),
	.w1(32'h3b1cc042),
	.w2(32'h3b53d4ec),
	.w3(32'hb98ca9a1),
	.w4(32'h3a3d8b59),
	.w5(32'h3b25c075),
	.w6(32'hb9e780b5),
	.w7(32'h3a880d9e),
	.w8(32'h3a996c13),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb8fa8),
	.w1(32'hba0aafd7),
	.w2(32'h38ab364a),
	.w3(32'h3ac857c5),
	.w4(32'hbaea2211),
	.w5(32'hba49a4b2),
	.w6(32'h3a0583ad),
	.w7(32'h3a5a5679),
	.w8(32'h3a8b6952),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a034f30),
	.w1(32'hb9de7bf9),
	.w2(32'h3a8e3d48),
	.w3(32'hba51faec),
	.w4(32'hba0a84a7),
	.w5(32'h3aca0cb2),
	.w6(32'hb8944de9),
	.w7(32'h3a2d13f5),
	.w8(32'hba278253),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4298dd),
	.w1(32'h3a24a38d),
	.w2(32'h3a9bf39a),
	.w3(32'hba03e79b),
	.w4(32'hb99666d0),
	.w5(32'h3abba1da),
	.w6(32'hbb179aed),
	.w7(32'hb99bf69c),
	.w8(32'hba9ad322),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbb20),
	.w1(32'hba5b04d6),
	.w2(32'h39d9823b),
	.w3(32'hba55f8d9),
	.w4(32'hbaf93f43),
	.w5(32'hba977e2d),
	.w6(32'hbab14bb8),
	.w7(32'hbb05be29),
	.w8(32'hbaf1eb49),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1ab73),
	.w1(32'hb9d4fed3),
	.w2(32'hb9f382f0),
	.w3(32'hba863ee7),
	.w4(32'hbadb5261),
	.w5(32'hbb0cd183),
	.w6(32'h3b57194e),
	.w7(32'h3b0c4f68),
	.w8(32'h3bcd0765),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c8d20),
	.w1(32'hb96ac4ab),
	.w2(32'hbaad1550),
	.w3(32'h3a6fcb32),
	.w4(32'hbac44844),
	.w5(32'hbad264c2),
	.w6(32'h3a91cce6),
	.w7(32'h39776fb2),
	.w8(32'h3a170542),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6d4a),
	.w1(32'hbb30d433),
	.w2(32'hb9c6c7ea),
	.w3(32'hbad55ecd),
	.w4(32'hbb566722),
	.w5(32'hbaa315f7),
	.w6(32'hba292bef),
	.w7(32'h3ae66048),
	.w8(32'h3b0f3fa2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d78a),
	.w1(32'hbac60884),
	.w2(32'h39864ec1),
	.w3(32'h39e356fc),
	.w4(32'hbba73119),
	.w5(32'hbbac2fae),
	.w6(32'h3bd0a961),
	.w7(32'h3bdf461a),
	.w8(32'h3c18c701),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bfe8a),
	.w1(32'hb9dcb7fd),
	.w2(32'h3aa63b98),
	.w3(32'hbb047fa6),
	.w4(32'hbb04ddfc),
	.w5(32'hb9cb2433),
	.w6(32'h39078a8f),
	.w7(32'h399c508a),
	.w8(32'h3aa38444),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d4bc0d),
	.w1(32'hbb0ae05a),
	.w2(32'h3b17e097),
	.w3(32'hba878aba),
	.w4(32'h3bb0618b),
	.w5(32'h3c2bec26),
	.w6(32'hbb5cdc46),
	.w7(32'h3ad8b932),
	.w8(32'hbb89be76),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac45514),
	.w1(32'h3a1c9877),
	.w2(32'h3b05daf4),
	.w3(32'h3c117c11),
	.w4(32'hba95d067),
	.w5(32'h3ad51171),
	.w6(32'hbadfcc3d),
	.w7(32'hb967e839),
	.w8(32'h37fd8eb2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a3d5c),
	.w1(32'h3a92244f),
	.w2(32'h3aac2a8f),
	.w3(32'h39d8a05f),
	.w4(32'hba0746b5),
	.w5(32'h3a7a0765),
	.w6(32'h39e36932),
	.w7(32'hb871ddbe),
	.w8(32'hbab59abe),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba947677),
	.w1(32'h38cd0515),
	.w2(32'h3ab58916),
	.w3(32'hbaac8fbd),
	.w4(32'hba145743),
	.w5(32'h3a84e25d),
	.w6(32'h3aabfdf3),
	.w7(32'h3aceff8b),
	.w8(32'hb8a267f2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b124e1),
	.w1(32'h3ad84a06),
	.w2(32'hbb501621),
	.w3(32'hba82a72c),
	.w4(32'h3ab2e011),
	.w5(32'hbb54f117),
	.w6(32'h3af2e2a2),
	.w7(32'hba5d6b63),
	.w8(32'h3a79eaa7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9728f8),
	.w1(32'hbb246b37),
	.w2(32'h3b68ace3),
	.w3(32'hbaaf1d9d),
	.w4(32'hbb229c12),
	.w5(32'h3a0c70c0),
	.w6(32'h3a81e664),
	.w7(32'h3aeab5a9),
	.w8(32'hb887a39f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e7385),
	.w1(32'h3c9b5425),
	.w2(32'h3c18df5a),
	.w3(32'h3b213a72),
	.w4(32'h3b661afe),
	.w5(32'hbb29475f),
	.w6(32'h3b97e103),
	.w7(32'hbbb29788),
	.w8(32'h38ce3d3b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b823d),
	.w1(32'hb9ca92f5),
	.w2(32'h3a6cb812),
	.w3(32'hbaf1ea2e),
	.w4(32'hbac3dbf7),
	.w5(32'hba1daec3),
	.w6(32'h3a1e20d3),
	.w7(32'h3ab6e276),
	.w8(32'h3b29f08e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b9f5f),
	.w1(32'h3aa8866f),
	.w2(32'h3ad97942),
	.w3(32'hba1ef6e2),
	.w4(32'hba29f609),
	.w5(32'h3a990f76),
	.w6(32'hbab97205),
	.w7(32'hbb629cbc),
	.w8(32'hbb18c42c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7ef47),
	.w1(32'hba00f829),
	.w2(32'h3aefcdba),
	.w3(32'h3abcced6),
	.w4(32'h3b491509),
	.w5(32'h3bc972f2),
	.w6(32'hbbd39b0d),
	.w7(32'h39bf7127),
	.w8(32'hba9e4292),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8ff35),
	.w1(32'hb9711045),
	.w2(32'hb9a41d6d),
	.w3(32'h3b6a3a74),
	.w4(32'hba8fa1f4),
	.w5(32'hba979ad7),
	.w6(32'h3a9aec3e),
	.w7(32'h39aaf30d),
	.w8(32'h39da26c0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9828fbd),
	.w1(32'h391c81bb),
	.w2(32'h3a44d947),
	.w3(32'hbb0b26d5),
	.w4(32'hbb42cba1),
	.w5(32'hbaeba35d),
	.w6(32'hbad3853e),
	.w7(32'hbacc00ab),
	.w8(32'h3a2fe7d6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93419d),
	.w1(32'h3b2dcd3e),
	.w2(32'h3c0f61e7),
	.w3(32'hba39b7d2),
	.w4(32'h3bd1f24e),
	.w5(32'h3c5ad679),
	.w6(32'h3a888625),
	.w7(32'h3bd6d531),
	.w8(32'hbbbfbb9b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22cb1c),
	.w1(32'h3addd20c),
	.w2(32'h3a9f09a4),
	.w3(32'hbb246d5e),
	.w4(32'h3c8da738),
	.w5(32'h3c6f86f7),
	.w6(32'h3ba9c53f),
	.w7(32'h3bcdb3e0),
	.w8(32'h3b5e525c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196fd1),
	.w1(32'h39e61f91),
	.w2(32'hbb118c67),
	.w3(32'h3c50e787),
	.w4(32'hb87005d6),
	.w5(32'hbb1d09f4),
	.w6(32'h3acadf6f),
	.w7(32'hba3d443b),
	.w8(32'h3a1756ea),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5df14),
	.w1(32'hb98638b2),
	.w2(32'hba8d300e),
	.w3(32'hbab8232d),
	.w4(32'hbab52f8c),
	.w5(32'hbb0c29ec),
	.w6(32'h3a2d107d),
	.w7(32'hb9ed0cc8),
	.w8(32'h398f6f54),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b6aac),
	.w1(32'hbb51e6db),
	.w2(32'h3a4e1254),
	.w3(32'hbaf139f8),
	.w4(32'hbb3498a6),
	.w5(32'h3ad37d8a),
	.w6(32'hbadb6e1e),
	.w7(32'h3a71345e),
	.w8(32'hbb5be783),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305bf1),
	.w1(32'h3b5faf11),
	.w2(32'h3aefeaea),
	.w3(32'hb980371b),
	.w4(32'h3bd6c509),
	.w5(32'h3b69a1ac),
	.w6(32'h3bd8a8d1),
	.w7(32'h3b64579d),
	.w8(32'hbbf52989),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0633eb),
	.w1(32'h3aa816be),
	.w2(32'h3a7729a1),
	.w3(32'hbbfbaa44),
	.w4(32'hbaddb8b6),
	.w5(32'hba2d90fe),
	.w6(32'hbaf33195),
	.w7(32'hbac50dec),
	.w8(32'hbb82edfc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb011517),
	.w1(32'h3937f26c),
	.w2(32'hbaa83d6d),
	.w3(32'hbb2e6f08),
	.w4(32'hbacc6def),
	.w5(32'hbafa2509),
	.w6(32'hb86f7f6c),
	.w7(32'hbaf9befb),
	.w8(32'h3a1d4508),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab55362),
	.w1(32'hb98f2337),
	.w2(32'h3b239d54),
	.w3(32'h3997ac90),
	.w4(32'hbb2a520c),
	.w5(32'h3a99cd8b),
	.w6(32'h39424228),
	.w7(32'h3af295fb),
	.w8(32'h3ac0d503),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ae8f2),
	.w1(32'h3b07e55b),
	.w2(32'h3b534892),
	.w3(32'h3a999d98),
	.w4(32'h3a8b50a4),
	.w5(32'h3b0ed0bb),
	.w6(32'h399a9b6f),
	.w7(32'h3a4f2966),
	.w8(32'h3ac06f7e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec0fe1),
	.w1(32'h3a5da41a),
	.w2(32'h3ad89ebd),
	.w3(32'h3a9161de),
	.w4(32'hb9e1eac8),
	.w5(32'h3926967b),
	.w6(32'h3ac066ea),
	.w7(32'h3b299172),
	.w8(32'h3b665575),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3acb5),
	.w1(32'h3aa5f59a),
	.w2(32'h3ad25afc),
	.w3(32'h39a4e89b),
	.w4(32'h3a411684),
	.w5(32'h3a8b00cc),
	.w6(32'h3a290d14),
	.w7(32'h3a91616c),
	.w8(32'h39b1c2eb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ed4b2),
	.w1(32'h3b88bb5b),
	.w2(32'hbbfefd65),
	.w3(32'h3a0e3d10),
	.w4(32'h3c9c8e76),
	.w5(32'h3bc4c7cf),
	.w6(32'h3c214a18),
	.w7(32'h3a81e4f1),
	.w8(32'h3b97269d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73a6c7),
	.w1(32'h3b0898e0),
	.w2(32'h3b09804a),
	.w3(32'h3c1006eb),
	.w4(32'h3a1571dc),
	.w5(32'hb944267b),
	.w6(32'h385760ad),
	.w7(32'hbaa8fa2c),
	.w8(32'hba9699c8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39555f9b),
	.w1(32'h390fd634),
	.w2(32'hbaf924ad),
	.w3(32'hba0c5ff2),
	.w4(32'h3995848c),
	.w5(32'hbaff5218),
	.w6(32'h3ae0c082),
	.w7(32'hba749589),
	.w8(32'hbaacbed7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a03e8),
	.w1(32'hbb0c796b),
	.w2(32'h3b72db23),
	.w3(32'hbae846f5),
	.w4(32'hbae7f6c7),
	.w5(32'h3b95e062),
	.w6(32'hbb84004e),
	.w7(32'h3aeeb02a),
	.w8(32'h3ab5c0aa),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99945d1),
	.w1(32'hbaabf180),
	.w2(32'h3b6ec1d5),
	.w3(32'h3a8b2e6e),
	.w4(32'hbb404b14),
	.w5(32'hbac5ba38),
	.w6(32'hba60e5f8),
	.w7(32'h3a4ebe9d),
	.w8(32'hb9b52e45),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55c45e),
	.w1(32'h3a9c144a),
	.w2(32'h3b0ff292),
	.w3(32'hb8f4082d),
	.w4(32'hbab83165),
	.w5(32'hba0262d1),
	.w6(32'h392880b4),
	.w7(32'h385ae1e7),
	.w8(32'h3a2185cf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a769d4),
	.w1(32'h396f9bc5),
	.w2(32'h38f03f1e),
	.w3(32'hba9992c3),
	.w4(32'hbb5f292d),
	.w5(32'hbb1d0c67),
	.w6(32'h3ba84a4d),
	.w7(32'h3b957218),
	.w8(32'h3ba48562),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19bbe8),
	.w1(32'h3c030c47),
	.w2(32'h3ca0568e),
	.w3(32'hb8a502f4),
	.w4(32'h3bf07aff),
	.w5(32'h3cb0805a),
	.w6(32'h3add7d89),
	.w7(32'h3c3e19bf),
	.w8(32'hbc02b35c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b813aee),
	.w1(32'hb711bb4c),
	.w2(32'hbaafe86c),
	.w3(32'h3a4c6151),
	.w4(32'hb9f846b0),
	.w5(32'hbaba4f84),
	.w6(32'h3a90483a),
	.w7(32'hbab4c54a),
	.w8(32'hba9aa290),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28af79),
	.w1(32'hba60651c),
	.w2(32'h39424166),
	.w3(32'hba9b153d),
	.w4(32'hbac005c7),
	.w5(32'hba3b2f6b),
	.w6(32'h39e1a315),
	.w7(32'h3ad6845b),
	.w8(32'h3b2baded),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae915d1),
	.w1(32'h3ad2ce9b),
	.w2(32'h39986134),
	.w3(32'h3a40a842),
	.w4(32'h3a900154),
	.w5(32'h3b323c32),
	.w6(32'h3a133554),
	.w7(32'h3a77aa16),
	.w8(32'h3a991f0d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73a571),
	.w1(32'h3af8bb3f),
	.w2(32'h3b6245d8),
	.w3(32'h3a98962b),
	.w4(32'hbb15443d),
	.w5(32'hbaf98f61),
	.w6(32'h3a0bb4c1),
	.w7(32'hba0723d3),
	.w8(32'h3b8e18c6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b621494),
	.w1(32'h3b007f82),
	.w2(32'h3a9b73c0),
	.w3(32'h3a91e576),
	.w4(32'h3a6e5c75),
	.w5(32'h3a093c13),
	.w6(32'h3b17b82b),
	.w7(32'h399c7460),
	.w8(32'h3b2da0b7),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60aacf),
	.w1(32'hbafa29bf),
	.w2(32'h3b2a763c),
	.w3(32'h3ace6db5),
	.w4(32'hbb687132),
	.w5(32'h3a1ce935),
	.w6(32'hb8f9bc70),
	.w7(32'h3a63a9f4),
	.w8(32'h3a517468),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b6f3c),
	.w1(32'hbb550e52),
	.w2(32'hbb026902),
	.w3(32'h3a2243dc),
	.w4(32'hbb06fd60),
	.w5(32'hba39d81c),
	.w6(32'hbb002f53),
	.w7(32'hba4d2cb5),
	.w8(32'hbb4c4f11),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb404e0f),
	.w1(32'hbb98c4c7),
	.w2(32'hbc696c8c),
	.w3(32'hbb131f19),
	.w4(32'h3ac6b6b2),
	.w5(32'hbc11b88c),
	.w6(32'h3b8192c7),
	.w7(32'hbb71a756),
	.w8(32'h3bfdb944),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4951c),
	.w1(32'hb9a253eb),
	.w2(32'hbb1e1f78),
	.w3(32'hba892f11),
	.w4(32'h3b00169a),
	.w5(32'hba571729),
	.w6(32'h3a128c45),
	.w7(32'hbb099dd8),
	.w8(32'hbab1330c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf2e4c),
	.w1(32'hbb651fff),
	.w2(32'hbb7edc56),
	.w3(32'hbb0b0ad0),
	.w4(32'hbb5474c2),
	.w5(32'hbae24853),
	.w6(32'hb89081a7),
	.w7(32'hba8808ac),
	.w8(32'h3b0eb157),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05740e),
	.w1(32'h3b0e677c),
	.w2(32'h3ad838de),
	.w3(32'hbadf13cc),
	.w4(32'h3a7e8570),
	.w5(32'h3a729088),
	.w6(32'h3a421190),
	.w7(32'h39b22716),
	.w8(32'h399ead1b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9edec),
	.w1(32'hba9e7bc5),
	.w2(32'hb90e2e41),
	.w3(32'h3ad8ac39),
	.w4(32'hbb0b6d22),
	.w5(32'hba919b06),
	.w6(32'hb85185fd),
	.w7(32'h3a81b60e),
	.w8(32'h3af41073),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac25659),
	.w1(32'hba06acd3),
	.w2(32'hb8456d5b),
	.w3(32'hb821fa3e),
	.w4(32'hba80e14a),
	.w5(32'hba50c34f),
	.w6(32'hba4e0303),
	.w7(32'hbaadc824),
	.w8(32'hbaf1c43c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b88fa1),
	.w1(32'hba8f2c16),
	.w2(32'h3b0d396f),
	.w3(32'hba7eb929),
	.w4(32'hba89f9fa),
	.w5(32'h3a3f533b),
	.w6(32'h39f31bd4),
	.w7(32'h3b14d9f4),
	.w8(32'h3b09f1ab),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af633d2),
	.w1(32'hbac4b722),
	.w2(32'h3b244722),
	.w3(32'h3a5f2243),
	.w4(32'h39c9946f),
	.w5(32'h3b26b1fb),
	.w6(32'h3a37ddad),
	.w7(32'hba7e832b),
	.w8(32'hbb88db4d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39809610),
	.w1(32'hbb003b86),
	.w2(32'h3abcf063),
	.w3(32'h3a03b389),
	.w4(32'hbae72f72),
	.w5(32'h3b245275),
	.w6(32'hbb4b0268),
	.w7(32'h3a2f915b),
	.w8(32'hb98a6544),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03ce78),
	.w1(32'hba5d14d0),
	.w2(32'hba42053a),
	.w3(32'h3a28d812),
	.w4(32'hbad08555),
	.w5(32'hba28bc54),
	.w6(32'hba8ebd09),
	.w7(32'hbadce6ec),
	.w8(32'hbb13a9e3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbb9b6),
	.w1(32'hbb58764c),
	.w2(32'hbb67a2b4),
	.w3(32'hbaa4d9fa),
	.w4(32'hbaa0ac73),
	.w5(32'h3a37ca1c),
	.w6(32'hbb063ddf),
	.w7(32'hbb298b8f),
	.w8(32'hba57f46a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8f88a),
	.w1(32'hba46a317),
	.w2(32'hbbbcfb4a),
	.w3(32'hbad8ee18),
	.w4(32'h3bffd5a5),
	.w5(32'hb80c5d6a),
	.w6(32'h3ba37114),
	.w7(32'hba77731d),
	.w8(32'h3be03152),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3618e3),
	.w1(32'h3c8dbd39),
	.w2(32'h3bb26fd6),
	.w3(32'h3b88b285),
	.w4(32'h3cb6f2a5),
	.w5(32'h3c50eac4),
	.w6(32'h3c34fda2),
	.w7(32'h39b586ff),
	.w8(32'h3adbbd4b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c352073),
	.w1(32'hb903070c),
	.w2(32'h39b7a697),
	.w3(32'h3c3b8199),
	.w4(32'hbaaa250e),
	.w5(32'hbabde396),
	.w6(32'h3a899bb3),
	.w7(32'h39973b09),
	.w8(32'h3b37b1da),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949dfa4),
	.w1(32'hba5ec2ec),
	.w2(32'hbafe26ea),
	.w3(32'hba291921),
	.w4(32'hba4d8297),
	.w5(32'h3a4aa163),
	.w6(32'hbafa29b2),
	.w7(32'hba92766d),
	.w8(32'h3aba8fd2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812288),
	.w1(32'h3a7018e0),
	.w2(32'h3a73e841),
	.w3(32'hbb041390),
	.w4(32'hb9876b32),
	.w5(32'h39a9cac2),
	.w6(32'hba92cff0),
	.w7(32'hba8a7e83),
	.w8(32'hba822c8d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a072e39),
	.w1(32'hba0ca565),
	.w2(32'hb9a99a35),
	.w3(32'h395cf106),
	.w4(32'hbad4bfa4),
	.w5(32'hba7dc249),
	.w6(32'h3aa3c0a5),
	.w7(32'h3a5e77df),
	.w8(32'h3b23b616),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33b6d8),
	.w1(32'hba36411f),
	.w2(32'hb8b8cf32),
	.w3(32'hb7565cd1),
	.w4(32'hbadd15cf),
	.w5(32'hba4ad916),
	.w6(32'h39dce98d),
	.w7(32'h3a4584c3),
	.w8(32'h3b105bc1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cef4f),
	.w1(32'h3a821702),
	.w2(32'hba9505a9),
	.w3(32'h3986c2f4),
	.w4(32'hba412f4c),
	.w5(32'hbb2ca4ce),
	.w6(32'h3a32413e),
	.w7(32'hbae97317),
	.w8(32'hb982eb20),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11cb8a),
	.w1(32'h3b13a695),
	.w2(32'h3b3253c3),
	.w3(32'hbaab29ce),
	.w4(32'h39a340f0),
	.w5(32'h3ab39917),
	.w6(32'h3ae0020f),
	.w7(32'h399d0aa3),
	.w8(32'hb9cabc85),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01d107),
	.w1(32'hbb379e18),
	.w2(32'hba4ee44e),
	.w3(32'h3a89403c),
	.w4(32'hbb85396e),
	.w5(32'hbb834a8a),
	.w6(32'hb95d845f),
	.w7(32'h3add42a4),
	.w8(32'h3bf61dac),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cc402),
	.w1(32'hbb18f026),
	.w2(32'hb99083c7),
	.w3(32'hba7f08ef),
	.w4(32'hbb6a4761),
	.w5(32'hb9f03da6),
	.w6(32'hba48c499),
	.w7(32'h3a74f105),
	.w8(32'h3ae44865),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964394c),
	.w1(32'h3a1724f3),
	.w2(32'h3a991d57),
	.w3(32'hba535221),
	.w4(32'h381565e2),
	.w5(32'h3978a355),
	.w6(32'hb9b16f46),
	.w7(32'hbb1c57f4),
	.w8(32'hbb057296),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985c482),
	.w1(32'hbb1b33d3),
	.w2(32'h3a66233d),
	.w3(32'h395a5d5f),
	.w4(32'hb970d474),
	.w5(32'h3bab4f2e),
	.w6(32'hbbb439a4),
	.w7(32'hbb2c720a),
	.w8(32'hbbb0986c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7abf),
	.w1(32'h3afff6ed),
	.w2(32'hbb0fc2b0),
	.w3(32'h3a88da0c),
	.w4(32'h3a897f80),
	.w5(32'hbb333fe9),
	.w6(32'h3b3d2879),
	.w7(32'hba87ad71),
	.w8(32'h396899ce),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d57cb9),
	.w1(32'h3c43f8ea),
	.w2(32'hbba0ec36),
	.w3(32'hba6a73a8),
	.w4(32'h3c91abd2),
	.w5(32'hba87e3b9),
	.w6(32'h3c68b8f6),
	.w7(32'hbb6dda24),
	.w8(32'h3b059be2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f62fd),
	.w1(32'h3abd7440),
	.w2(32'h3b31db15),
	.w3(32'h39d9c4e0),
	.w4(32'h394ff885),
	.w5(32'h3a663ce2),
	.w6(32'h392a2f98),
	.w7(32'h3a79b256),
	.w8(32'hb985f98b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76205f),
	.w1(32'h3b027c1f),
	.w2(32'h3b3133ab),
	.w3(32'h3a0de048),
	.w4(32'h3b32715a),
	.w5(32'h3b8063d6),
	.w6(32'h3877295e),
	.w7(32'hba59aeb3),
	.w8(32'hba73e776),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace1ba3),
	.w1(32'h3a31f59f),
	.w2(32'h39e80193),
	.w3(32'h3b155163),
	.w4(32'h394eb06a),
	.w5(32'hb9b648a1),
	.w6(32'h39879e24),
	.w7(32'hb9ea5853),
	.w8(32'hba2bc2af),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d720e1),
	.w1(32'h3c1d14b9),
	.w2(32'h3c5d6d39),
	.w3(32'h3913c0f9),
	.w4(32'h3a7cee3e),
	.w5(32'h3ba8e9ab),
	.w6(32'h3bf2d8e8),
	.w7(32'h3bcfb5a3),
	.w8(32'hbbaf62aa),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf99c9e),
	.w1(32'h392bf967),
	.w2(32'hb81dffc0),
	.w3(32'hbbddd22b),
	.w4(32'h3b2db6b4),
	.w5(32'h3ac33962),
	.w6(32'h3a7e238b),
	.w7(32'h3a5e8185),
	.w8(32'h3b1a61b5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc9357),
	.w1(32'hbb1cc5e6),
	.w2(32'hba90cde4),
	.w3(32'h3b6e17f4),
	.w4(32'hba8ca9da),
	.w5(32'h3a85f9ca),
	.w6(32'hbb27f649),
	.w7(32'hba221f26),
	.w8(32'h39896039),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb052df4),
	.w1(32'h378e545e),
	.w2(32'hbb0241f2),
	.w3(32'h3928fe5b),
	.w4(32'h397712d2),
	.w5(32'hbb089804),
	.w6(32'h3a69768b),
	.w7(32'hba5f681f),
	.w8(32'h39511235),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf167d),
	.w1(32'hbaed230e),
	.w2(32'hbb169930),
	.w3(32'hba769748),
	.w4(32'hba9f6080),
	.w5(32'hbab14ace),
	.w6(32'hba317a1a),
	.w7(32'hba55865c),
	.w8(32'hbb1d5e9d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21b56b),
	.w1(32'h3a4e8f7e),
	.w2(32'hbb1132bb),
	.w3(32'hbb17a754),
	.w4(32'h397883a5),
	.w5(32'hbb3c355a),
	.w6(32'h3aa2187d),
	.w7(32'hba911d71),
	.w8(32'h3a1f9c8a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39273d8d),
	.w1(32'h3b2bf8f8),
	.w2(32'h3adc057e),
	.w3(32'hba9e1a1a),
	.w4(32'h38bfe1c7),
	.w5(32'hba6b7533),
	.w6(32'h3a5e3e3a),
	.w7(32'h39a2e2e2),
	.w8(32'h3a37517c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e314f),
	.w1(32'h3acb5007),
	.w2(32'h3b0dbdfd),
	.w3(32'hba6c6a1c),
	.w4(32'h3a03c275),
	.w5(32'h3aee0cc2),
	.w6(32'hb8cdd097),
	.w7(32'h38a899a2),
	.w8(32'h38d03b19),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb31a9),
	.w1(32'h3b15524b),
	.w2(32'h3a64d58f),
	.w3(32'h3a91b0dd),
	.w4(32'h3823f1e3),
	.w5(32'hba0e93dd),
	.w6(32'hb74b498e),
	.w7(32'hba016811),
	.w8(32'hbabfda13),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf7a45),
	.w1(32'h3c2288b2),
	.w2(32'hbbceca84),
	.w3(32'hba25ebc1),
	.w4(32'h3c5f53ff),
	.w5(32'hbb88cb55),
	.w6(32'h3c45a11f),
	.w7(32'hbb510a26),
	.w8(32'h3b124fbc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eeaadf),
	.w1(32'h3b07f1d7),
	.w2(32'h3ae823bd),
	.w3(32'hba2f55f0),
	.w4(32'hba34f4d6),
	.w5(32'hba586122),
	.w6(32'hba6eb009),
	.w7(32'hbaceb372),
	.w8(32'hbab466dc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b146c6e),
	.w1(32'hba967fc7),
	.w2(32'hba16140f),
	.w3(32'hba5e550c),
	.w4(32'hbae187b8),
	.w5(32'hba67a104),
	.w6(32'h39e2b513),
	.w7(32'h39d4147a),
	.w8(32'h3a8d7da5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e027d),
	.w1(32'h3c4dd068),
	.w2(32'h3b895485),
	.w3(32'hba126278),
	.w4(32'h3bc3551f),
	.w5(32'hbaaf8653),
	.w6(32'h3ba5a573),
	.w7(32'hbb9f275c),
	.w8(32'hbb195e03),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02e4be),
	.w1(32'h3a82adc6),
	.w2(32'hbabdde0c),
	.w3(32'hbb1b5743),
	.w4(32'h3a815940),
	.w5(32'h3b71e9c8),
	.w6(32'h3a9b8a88),
	.w7(32'hba49735c),
	.w8(32'hb9ed6b52),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b209c3),
	.w1(32'h3b39cf69),
	.w2(32'h3b58fae9),
	.w3(32'h3a1c7c8b),
	.w4(32'h392aed7e),
	.w5(32'h3a7ec7dd),
	.w6(32'hb9fa2589),
	.w7(32'h39697b67),
	.w8(32'hbb04b4f6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33b06f),
	.w1(32'h3af4a592),
	.w2(32'h38e903dc),
	.w3(32'h3ad4882e),
	.w4(32'h3ad84843),
	.w5(32'h3b2e7289),
	.w6(32'h3b10b760),
	.w7(32'hbaaf4f64),
	.w8(32'hba83a125),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e71528),
	.w1(32'hbb48821a),
	.w2(32'hbbe382af),
	.w3(32'h3b02358f),
	.w4(32'hbacf04cb),
	.w5(32'hba91b83b),
	.w6(32'hbaa893b8),
	.w7(32'hbb9523fd),
	.w8(32'hb980bfed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76833c),
	.w1(32'hbacbada2),
	.w2(32'hbb02627b),
	.w3(32'hbb4703f0),
	.w4(32'hbb35286e),
	.w5(32'hbb8d30c7),
	.w6(32'h3ad5522d),
	.w7(32'hbaded10a),
	.w8(32'h3b8bce26),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a698d1f),
	.w1(32'hbb7fba53),
	.w2(32'hba02bb8a),
	.w3(32'hbaaf73b1),
	.w4(32'hbba65e02),
	.w5(32'hba839574),
	.w6(32'hbac31a6e),
	.w7(32'h3aaeb026),
	.w8(32'h3b467816),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30463f),
	.w1(32'hba5b4010),
	.w2(32'hba39c8c3),
	.w3(32'hbaea3bf3),
	.w4(32'hbb3445c4),
	.w5(32'hbb0208df),
	.w6(32'h39ce8652),
	.w7(32'h39bfdeae),
	.w8(32'h3b18bc13),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35fb18),
	.w1(32'hbaa3691b),
	.w2(32'h39f95926),
	.w3(32'h3a51886a),
	.w4(32'hbb2b01c9),
	.w5(32'h3938a9c8),
	.w6(32'h39bf903e),
	.w7(32'h3a3fad64),
	.w8(32'h3ac222b4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c15ec),
	.w1(32'h3a33b6d4),
	.w2(32'h3a643b58),
	.w3(32'hb9b31b78),
	.w4(32'h39786c47),
	.w5(32'h3a5aedb8),
	.w6(32'h3a8f41f4),
	.w7(32'h3a2064ec),
	.w8(32'h3613169d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cc0bd),
	.w1(32'h3ad4bac4),
	.w2(32'h3b233da5),
	.w3(32'hbabd4d08),
	.w4(32'hba7d8b34),
	.w5(32'hbabe519a),
	.w6(32'hb9c0492f),
	.w7(32'hbabbff87),
	.w8(32'hbb173c89),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284d8a),
	.w1(32'h3b4878a1),
	.w2(32'h3903c89f),
	.w3(32'hba2e2cb9),
	.w4(32'h39d05a82),
	.w5(32'hbb102d51),
	.w6(32'h3ad19daf),
	.w7(32'hba00f9fa),
	.w8(32'h3a7bfecd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f287),
	.w1(32'hbab30f21),
	.w2(32'h3914a749),
	.w3(32'hba54add3),
	.w4(32'hbb0f6023),
	.w5(32'hb9decefd),
	.w6(32'hba0f6b2e),
	.w7(32'h3a7272a1),
	.w8(32'h3ad18e0e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a803630),
	.w1(32'h3a72d3b3),
	.w2(32'h3b1515f6),
	.w3(32'h3916d02a),
	.w4(32'hba43b46f),
	.w5(32'hb97433e6),
	.w6(32'h3ab7b1fb),
	.w7(32'h3a2044b8),
	.w8(32'h3a06b3d0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff7cfe),
	.w1(32'h3a995483),
	.w2(32'h3b0d1c88),
	.w3(32'h3ab36649),
	.w4(32'hbabf3628),
	.w5(32'hb9ec8ea3),
	.w6(32'h39ed8690),
	.w7(32'h3a793800),
	.w8(32'h3b326e9a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05a732),
	.w1(32'hbbd92647),
	.w2(32'h3aa1cd9a),
	.w3(32'hb9b9fe20),
	.w4(32'hbb9952b5),
	.w5(32'hbb197a15),
	.w6(32'hbb3cbf32),
	.w7(32'h39622b9c),
	.w8(32'h3a50c52f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809a30),
	.w1(32'hb7fb5335),
	.w2(32'h3afffdb5),
	.w3(32'h3ab91c7a),
	.w4(32'hbb3141e4),
	.w5(32'hb9122615),
	.w6(32'h3a266b53),
	.w7(32'h3a8eba6b),
	.w8(32'h3b1f208f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1089e4),
	.w1(32'h3b3990f1),
	.w2(32'h3a5ac25a),
	.w3(32'h39d28134),
	.w4(32'hba90f607),
	.w5(32'hbb172f0a),
	.w6(32'h3b2f60ea),
	.w7(32'h3b1e812c),
	.w8(32'h3af59f5f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a637eaf),
	.w1(32'hbb75ccaa),
	.w2(32'hbb1c9892),
	.w3(32'hbaeacff3),
	.w4(32'hbb8b3a48),
	.w5(32'hbb2745a3),
	.w6(32'hbb0e0795),
	.w7(32'hb94511eb),
	.w8(32'hbb2a5484),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fd6c4),
	.w1(32'hbb6027b0),
	.w2(32'hba4875f4),
	.w3(32'hbb387dc8),
	.w4(32'hbb736bc3),
	.w5(32'hba48068d),
	.w6(32'hbaba7d1c),
	.w7(32'h3a991733),
	.w8(32'h3ae29076),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e83d86),
	.w1(32'hbaa55bcd),
	.w2(32'hba14c595),
	.w3(32'hba64430d),
	.w4(32'hbaec064a),
	.w5(32'hba762a7e),
	.w6(32'h39bca3e0),
	.w7(32'h3a1f80ab),
	.w8(32'h3a8cae50),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d62cb),
	.w1(32'hbae1dbf2),
	.w2(32'hb91cc707),
	.w3(32'hba86c72e),
	.w4(32'hbb2c00ac),
	.w5(32'hba40439d),
	.w6(32'hb958ba3e),
	.w7(32'h3a8ff7b0),
	.w8(32'h3a967db8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9811a09),
	.w1(32'hba80fd47),
	.w2(32'h39e9607b),
	.w3(32'hba6a1d5a),
	.w4(32'hbad95e11),
	.w5(32'hbb473665),
	.w6(32'h3b1e222c),
	.w7(32'h3b4b5788),
	.w8(32'h3b29232d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b5992),
	.w1(32'hb9e89445),
	.w2(32'hba8cd203),
	.w3(32'hbaf0d62f),
	.w4(32'hbad67450),
	.w5(32'h3a892cfa),
	.w6(32'hb9d7658e),
	.w7(32'hbab1167e),
	.w8(32'hba58e5e6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7445e),
	.w1(32'h39917adb),
	.w2(32'h39f63f97),
	.w3(32'hbace6684),
	.w4(32'hbb816a1c),
	.w5(32'hbb626545),
	.w6(32'h39ff0555),
	.w7(32'hba412e6c),
	.w8(32'h3a771eaa),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb735),
	.w1(32'h3b26424b),
	.w2(32'h3aafc7a2),
	.w3(32'hbad64706),
	.w4(32'hba89eab4),
	.w5(32'hb98a92f6),
	.w6(32'h3b0248ff),
	.w7(32'h3aa7e7f7),
	.w8(32'h39092ca8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a081685),
	.w1(32'hbaa7fda7),
	.w2(32'h3a02ce0d),
	.w3(32'hbb081903),
	.w4(32'hbb05f042),
	.w5(32'hba483dba),
	.w6(32'h39c79e6d),
	.w7(32'h3aadacfe),
	.w8(32'h3b1b3ba7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e181),
	.w1(32'hbad64761),
	.w2(32'h3ad53ec1),
	.w3(32'hb8808ff5),
	.w4(32'hbabfae5e),
	.w5(32'hbb15102d),
	.w6(32'h3a9bddee),
	.w7(32'h3b0cd874),
	.w8(32'h3aafbffb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb622e64),
	.w1(32'h3a6b71d2),
	.w2(32'h3a784f41),
	.w3(32'hbba3e78e),
	.w4(32'h359be1a2),
	.w5(32'h3a76e3a5),
	.w6(32'h3a8efd31),
	.w7(32'h3a4a0778),
	.w8(32'h3ab45ce3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac90b74),
	.w1(32'h3add2cff),
	.w2(32'hba9260f1),
	.w3(32'h3ab7ab66),
	.w4(32'h3a903231),
	.w5(32'hbac581c2),
	.w6(32'h3b1d1388),
	.w7(32'hb881376b),
	.w8(32'h3a12bbd3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0baa3),
	.w1(32'h38373018),
	.w2(32'h37225ac8),
	.w3(32'hba9c144f),
	.w4(32'h38105fd9),
	.w5(32'hb7de0291),
	.w6(32'h37570a0f),
	.w7(32'h37e1cc9a),
	.w8(32'hb79bdc7c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d56dfc),
	.w1(32'hb8ca8d8d),
	.w2(32'h388ee058),
	.w3(32'hb9dd3871),
	.w4(32'hba4eb92d),
	.w5(32'hb9dbfb8e),
	.w6(32'hb88d98f5),
	.w7(32'hb935a377),
	.w8(32'hb897ccf0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3685e9),
	.w1(32'h3a27f862),
	.w2(32'h3a448e47),
	.w3(32'h3912257b),
	.w4(32'h3917c5e8),
	.w5(32'h395174c7),
	.w6(32'h398e0d46),
	.w7(32'h3983321f),
	.w8(32'h39bce26c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901daa4),
	.w1(32'h38ae887f),
	.w2(32'h38d63b15),
	.w3(32'hb740a668),
	.w4(32'hb835233e),
	.w5(32'hb801b4a6),
	.w6(32'h37c8038c),
	.w7(32'hb71710b9),
	.w8(32'h38390e7a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad2697),
	.w1(32'hb8587b4a),
	.w2(32'hb8eaf40e),
	.w3(32'hb9502f33),
	.w4(32'hb963b188),
	.w5(32'hb94328bd),
	.w6(32'hb8f5b854),
	.w7(32'hb88c6e32),
	.w8(32'hb8bf1e7f),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b5d401),
	.w1(32'h38a4908c),
	.w2(32'h396ae876),
	.w3(32'hb7c5be1d),
	.w4(32'hb78b1900),
	.w5(32'h388d0d86),
	.w6(32'h38f38af6),
	.w7(32'h38dc320e),
	.w8(32'h39430d33),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391eaea1),
	.w1(32'h38b5fbc5),
	.w2(32'h39301a57),
	.w3(32'hb91d9791),
	.w4(32'hb802e5b3),
	.w5(32'hb7cfd479),
	.w6(32'h382606c4),
	.w7(32'h38a122b9),
	.w8(32'h391e64ce),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995862c),
	.w1(32'h39975155),
	.w2(32'h3a1b0c88),
	.w3(32'hb9047002),
	.w4(32'h38129bda),
	.w5(32'hb51ce966),
	.w6(32'h390c9d46),
	.w7(32'h39894565),
	.w8(32'h39be3d8a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7919ee),
	.w1(32'h3a6eff23),
	.w2(32'h3a857dea),
	.w3(32'h37df1b44),
	.w4(32'h394cd742),
	.w5(32'h393918b4),
	.w6(32'h3996dac7),
	.w7(32'h39836ff0),
	.w8(32'h39e5aa84),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810b6e6),
	.w1(32'h39247622),
	.w2(32'h3999aaad),
	.w3(32'h35ffd82a),
	.w4(32'h385d4f1b),
	.w5(32'h384628a7),
	.w6(32'h39ab2a18),
	.w7(32'h399018c5),
	.w8(32'h39960746),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebccf8),
	.w1(32'h39833661),
	.w2(32'h39a19ae5),
	.w3(32'h37c9e678),
	.w4(32'hb8bb6c7d),
	.w5(32'hb8e955b3),
	.w6(32'h38f352ed),
	.w7(32'h3838c013),
	.w8(32'h391828dd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a657d49),
	.w1(32'h3a3addf5),
	.w2(32'h3a4221e8),
	.w3(32'h39cf0d8c),
	.w4(32'h393401ca),
	.w5(32'h396a7d70),
	.w6(32'h39eba6ef),
	.w7(32'h399ccad9),
	.w8(32'h39c6c57f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8d207),
	.w1(32'hb8312e3e),
	.w2(32'h396593ba),
	.w3(32'hb924414a),
	.w4(32'hb9826a13),
	.w5(32'h3745e31e),
	.w6(32'h390c915b),
	.w7(32'h396172a9),
	.w8(32'h39968512),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a303b5),
	.w1(32'h39c87f50),
	.w2(32'h397ecd96),
	.w3(32'h37324b1f),
	.w4(32'h37fb8841),
	.w5(32'hb8891e44),
	.w6(32'h391069a0),
	.w7(32'h39015bb2),
	.w8(32'h39942bd9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380d32ac),
	.w1(32'h39083fda),
	.w2(32'h391c90d6),
	.w3(32'hb7f5ab14),
	.w4(32'h386f6be2),
	.w5(32'h38475562),
	.w6(32'h385f899d),
	.w7(32'h38e0ffbe),
	.w8(32'h391d92b8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4315a),
	.w1(32'h39810651),
	.w2(32'h3a92a064),
	.w3(32'hb9c5a62e),
	.w4(32'h399d04b9),
	.w5(32'h3a4a7ec7),
	.w6(32'h3a7fc3c3),
	.w7(32'h3ab45f00),
	.w8(32'h3aafb953),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4a975),
	.w1(32'h39e6a73e),
	.w2(32'h39df6dcf),
	.w3(32'h3998cd6e),
	.w4(32'h39b40125),
	.w5(32'h39b60dc4),
	.w6(32'h39e680da),
	.w7(32'h39dc00ba),
	.w8(32'h3a0c58e4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ca55ce),
	.w1(32'h37d0195d),
	.w2(32'h37c1a0e1),
	.w3(32'h38343592),
	.w4(32'h37e1053e),
	.w5(32'h38343ee5),
	.w6(32'h37b1bc35),
	.w7(32'h37edaa74),
	.w8(32'h3757cf81),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb593b160),
	.w1(32'h35a15be1),
	.w2(32'h3779223a),
	.w3(32'h37114721),
	.w4(32'h368ee36b),
	.w5(32'h35e0305e),
	.w6(32'h37ae97c2),
	.w7(32'h3787ff3b),
	.w8(32'h37bf3823),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936399c),
	.w1(32'h39563113),
	.w2(32'h3991176a),
	.w3(32'h39078797),
	.w4(32'h384ade71),
	.w5(32'h38eb4e4f),
	.w6(32'h39357be7),
	.w7(32'h389a66e0),
	.w8(32'h39370f27),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00e02c),
	.w1(32'h3a350198),
	.w2(32'h3a2afcf7),
	.w3(32'h39c3fe17),
	.w4(32'h39cb7817),
	.w5(32'h3a065c1b),
	.w6(32'h3a1a900e),
	.w7(32'h3a266a7a),
	.w8(32'h3a3d95e7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d01b66),
	.w1(32'h39ec19dd),
	.w2(32'h3a1ddd50),
	.w3(32'hb7a88184),
	.w4(32'hb8a87977),
	.w5(32'h390f7eb4),
	.w6(32'h39b0262a),
	.w7(32'h39969e0c),
	.w8(32'h3a157f32),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361f1a37),
	.w1(32'hb695c175),
	.w2(32'hb682c1ec),
	.w3(32'h368b1e50),
	.w4(32'hb69d252f),
	.w5(32'h33830b36),
	.w6(32'hb5a13963),
	.w7(32'hb596301b),
	.w8(32'hb6982586),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f576),
	.w1(32'h3a32f028),
	.w2(32'h3a2b5fa6),
	.w3(32'h385bee9d),
	.w4(32'h396283ae),
	.w5(32'h390c70f0),
	.w6(32'h39a78815),
	.w7(32'h39c41493),
	.w8(32'h3a176da5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40fd91),
	.w1(32'h39db8090),
	.w2(32'h3a36d824),
	.w3(32'h393c7714),
	.w4(32'h3985fa50),
	.w5(32'h3951bddf),
	.w6(32'h39709320),
	.w7(32'h39cbc1ce),
	.w8(32'h398e0cbe),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e45d0),
	.w1(32'h3a1d9fbb),
	.w2(32'h39dfb816),
	.w3(32'h3996e6cc),
	.w4(32'h36d8248c),
	.w5(32'hb8dfa015),
	.w6(32'h39a0b79e),
	.w7(32'h38d67089),
	.w8(32'h39770d1a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37de0044),
	.w1(32'h3a716607),
	.w2(32'h3ab32f87),
	.w3(32'hb79c7e3f),
	.w4(32'h3a814f2a),
	.w5(32'h3a8d04ec),
	.w6(32'h39e96e81),
	.w7(32'h3a812218),
	.w8(32'h3a48c55d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39225444),
	.w1(32'h393cfac8),
	.w2(32'h395c8fe6),
	.w3(32'h392acca3),
	.w4(32'h38708fdf),
	.w5(32'h38ed1d03),
	.w6(32'h39664c2f),
	.w7(32'h3936f1d2),
	.w8(32'h39167176),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923b6a5),
	.w1(32'h37bac812),
	.w2(32'hb95f2f3a),
	.w3(32'hb93589f1),
	.w4(32'h38385800),
	.w5(32'hb9200d97),
	.w6(32'hb937fb36),
	.w7(32'h38596c7e),
	.w8(32'hb98d93d4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dca2f),
	.w1(32'h3967b968),
	.w2(32'h385af346),
	.w3(32'h383d1eb6),
	.w4(32'h39ae66f8),
	.w5(32'hb6e0233e),
	.w6(32'h39d394b0),
	.w7(32'h39eb873e),
	.w8(32'h39e70c73),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d501d),
	.w1(32'h39a61938),
	.w2(32'h3a2beca6),
	.w3(32'hb909de4f),
	.w4(32'hb8550106),
	.w5(32'h399e5525),
	.w6(32'h396aec1b),
	.w7(32'h399f8398),
	.w8(32'h3a0d06ea),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fb9bf2),
	.w1(32'h352e2c61),
	.w2(32'h396419a4),
	.w3(32'hb92afd62),
	.w4(32'hb8d09476),
	.w5(32'h387e0c6f),
	.w6(32'h38c6cae8),
	.w7(32'h38f49d7c),
	.w8(32'h395f0534),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39970816),
	.w1(32'h394a8b94),
	.w2(32'h3942b2ef),
	.w3(32'h3900e158),
	.w4(32'h37d7c147),
	.w5(32'h38b3c5d3),
	.w6(32'h38db078f),
	.w7(32'h386a3630),
	.w8(32'h39015ec2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3702b5d9),
	.w1(32'hb7f12c6e),
	.w2(32'hb7558c72),
	.w3(32'h365801b1),
	.w4(32'hb6bcea7b),
	.w5(32'hb4112ba6),
	.w6(32'h378710c1),
	.w7(32'h37885189),
	.w8(32'h37b063f9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a052b7a),
	.w1(32'h39ec59ef),
	.w2(32'h3a0a814f),
	.w3(32'h3886236c),
	.w4(32'h36c06d31),
	.w5(32'h3892f5d1),
	.w6(32'h3985d6b0),
	.w7(32'h39219a30),
	.w8(32'h3926ea4d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986e580),
	.w1(32'h39942b77),
	.w2(32'h39a163d1),
	.w3(32'h38e25554),
	.w4(32'h38b57478),
	.w5(32'h395287df),
	.w6(32'h387b1aa9),
	.w7(32'h38817b6e),
	.w8(32'h3962c1b8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f201ec),
	.w1(32'h3877a0a0),
	.w2(32'h3984e43f),
	.w3(32'hb9214dcd),
	.w4(32'h39714872),
	.w5(32'h39a1565b),
	.w6(32'h394e12a7),
	.w7(32'h39b2142b),
	.w8(32'h39d30b14),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7bd44),
	.w1(32'h388d4a95),
	.w2(32'h384bec10),
	.w3(32'h38bb14d8),
	.w4(32'h388a2697),
	.w5(32'h37c6bac2),
	.w6(32'h38c01111),
	.w7(32'h39158c76),
	.w8(32'h37e395fd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de1663),
	.w1(32'hb73a68b1),
	.w2(32'hb916d91d),
	.w3(32'hb9acd2bf),
	.w4(32'hb9587a5d),
	.w5(32'hb9351d12),
	.w6(32'hb986a3da),
	.w7(32'hb97503ee),
	.w8(32'hb96fd319),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9102e9e),
	.w1(32'hb8647637),
	.w2(32'hb847b234),
	.w3(32'hb929dfed),
	.w4(32'hb89903fa),
	.w5(32'hb83e1bec),
	.w6(32'hb90adf79),
	.w7(32'hb885b168),
	.w8(32'hb86a496f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390615b5),
	.w1(32'h38b98f63),
	.w2(32'hb6645369),
	.w3(32'h38e20220),
	.w4(32'h38eb36ff),
	.w5(32'h382282db),
	.w6(32'h38621acc),
	.w7(32'h38efaae1),
	.w8(32'hb7e50304),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846f94f),
	.w1(32'h399cc954),
	.w2(32'h399c5d2c),
	.w3(32'h38f148b7),
	.w4(32'h39b37cfa),
	.w5(32'h38baf3f6),
	.w6(32'h398f274b),
	.w7(32'h39a85f51),
	.w8(32'h39b370d0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0912c0),
	.w1(32'h3a37308e),
	.w2(32'h3a2daa58),
	.w3(32'h39b86432),
	.w4(32'h386eb1ea),
	.w5(32'h39927d80),
	.w6(32'h3a43ab7f),
	.w7(32'h39deb0be),
	.w8(32'h3a335cbb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f286d),
	.w1(32'h3900602a),
	.w2(32'hb7a14f07),
	.w3(32'h38490531),
	.w4(32'h3816b4f1),
	.w5(32'hb7bef120),
	.w6(32'h381a10cb),
	.w7(32'h38d4af96),
	.w8(32'hb85bfdaf),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f0f3c),
	.w1(32'h39ae8660),
	.w2(32'h39e20c98),
	.w3(32'h369e328c),
	.w4(32'h399beb0c),
	.w5(32'h388f385b),
	.w6(32'h3994ae5a),
	.w7(32'h3a02e1f7),
	.w8(32'h39ab90a7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cbcd1),
	.w1(32'h382376b5),
	.w2(32'h39055907),
	.w3(32'hb9da38ee),
	.w4(32'hb9279775),
	.w5(32'hb8f1556a),
	.w6(32'hb98f690c),
	.w7(32'hb8d06b23),
	.w8(32'hb8a96ac3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20dca6),
	.w1(32'h3a10b92c),
	.w2(32'h3a66d950),
	.w3(32'hb940545e),
	.w4(32'h38bde907),
	.w5(32'h38c207f5),
	.w6(32'hb80fa9fb),
	.w7(32'h39641e09),
	.w8(32'h3a2dcbc7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b067f4),
	.w1(32'h39dc7e95),
	.w2(32'h3a034ba2),
	.w3(32'hb9cf2eda),
	.w4(32'hb9985c9b),
	.w5(32'hb95d7078),
	.w6(32'hb95a5b9a),
	.w7(32'hb9236e7a),
	.w8(32'hb7265058),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256277),
	.w1(32'h3a666467),
	.w2(32'h3a1676b7),
	.w3(32'h391dd1c7),
	.w4(32'h39cf553e),
	.w5(32'h384cbcbd),
	.w6(32'h38ab5e8c),
	.w7(32'h3982d2bd),
	.w8(32'h396dd18f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8ffe3),
	.w1(32'hb79f373b),
	.w2(32'hb6ca4724),
	.w3(32'hb7dc6ef7),
	.w4(32'hb7fed39d),
	.w5(32'h382d7b87),
	.w6(32'hb820dbf2),
	.w7(32'hb6f058b3),
	.w8(32'h381b5701),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39036b48),
	.w1(32'h38ba5891),
	.w2(32'h38c1948c),
	.w3(32'hb7cc1017),
	.w4(32'hb80adee6),
	.w5(32'hb98cc8b0),
	.w6(32'h392a1d98),
	.w7(32'h393136d0),
	.w8(32'h38ebde1a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360a2867),
	.w1(32'hb6a240ed),
	.w2(32'hb5dc4264),
	.w3(32'h36ea7cb0),
	.w4(32'h362968eb),
	.w5(32'h3660f3db),
	.w6(32'h365df473),
	.w7(32'h35e27107),
	.w8(32'h3601abd0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e96a3c),
	.w1(32'h390c148d),
	.w2(32'h39157e50),
	.w3(32'hb7622ba2),
	.w4(32'h3581c770),
	.w5(32'hb689c24d),
	.w6(32'h378de304),
	.w7(32'h36822a23),
	.w8(32'hb79d6d31),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a8b24a),
	.w1(32'hb846ac54),
	.w2(32'hb71e24e3),
	.w3(32'hb7f8bc9b),
	.w4(32'hb7c9b654),
	.w5(32'hb798bc30),
	.w6(32'h37e1a3c0),
	.w7(32'h388c53a5),
	.w8(32'h37f119e7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d0e6a),
	.w1(32'h382693f3),
	.w2(32'h397b02cc),
	.w3(32'hb9a35c03),
	.w4(32'hb9a6750c),
	.w5(32'hb9ad4e1c),
	.w6(32'hb93f693c),
	.w7(32'hb8458a23),
	.w8(32'h38a714e6),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb609287a),
	.w1(32'hb5ae080c),
	.w2(32'hb529eb26),
	.w3(32'h3580614e),
	.w4(32'hb5f1ec9e),
	.w5(32'hb5567812),
	.w6(32'h36c8a301),
	.w7(32'h361f70d4),
	.w8(32'hb68ac015),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d719a),
	.w1(32'h389602a4),
	.w2(32'h37b0150f),
	.w3(32'h38482034),
	.w4(32'h3889bae3),
	.w5(32'h3720a7e7),
	.w6(32'h37de23c3),
	.w7(32'h384b8365),
	.w8(32'h3748f2ea),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a93786),
	.w1(32'h378094a5),
	.w2(32'h39557b36),
	.w3(32'hb98ffeb7),
	.w4(32'hb8f54a3b),
	.w5(32'h37c100ca),
	.w6(32'hb8b29eb0),
	.w7(32'h3889b018),
	.w8(32'h390fe827),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ab1b0),
	.w1(32'h396ebcaf),
	.w2(32'h39f9b9b8),
	.w3(32'h39436133),
	.w4(32'hb85b4460),
	.w5(32'h365403c4),
	.w6(32'h38e03115),
	.w7(32'h392cc6fd),
	.w8(32'h3993171e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087db4),
	.w1(32'h39bf25ca),
	.w2(32'h397b8961),
	.w3(32'h39cba777),
	.w4(32'hb94982b0),
	.w5(32'h3948b35a),
	.w6(32'h3a15f5fd),
	.w7(32'hb9169297),
	.w8(32'h3832e9cd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3852f33a),
	.w1(32'h36736522),
	.w2(32'hb6753a73),
	.w3(32'hb6dc254c),
	.w4(32'hb840aa65),
	.w5(32'hb7af9938),
	.w6(32'hb81c4c07),
	.w7(32'hb8471444),
	.w8(32'hb8092224),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb723),
	.w1(32'h3a6c6b68),
	.w2(32'h3a6d9e77),
	.w3(32'h3a3226b2),
	.w4(32'h397da0e3),
	.w5(32'h39669e6f),
	.w6(32'h39d80274),
	.w7(32'h397d83ed),
	.w8(32'h3a3f7ca7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c16836),
	.w1(32'h3a8ebefc),
	.w2(32'h3ab6a372),
	.w3(32'hba3c5c99),
	.w4(32'h39a385c2),
	.w5(32'h39b798a5),
	.w6(32'h39c5ba34),
	.w7(32'h3a1d9cae),
	.w8(32'h3a547655),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c5434),
	.w1(32'h396ba9ab),
	.w2(32'h38af5fed),
	.w3(32'h37f93a6b),
	.w4(32'h38c3290f),
	.w5(32'h390385e9),
	.w6(32'h37b923fe),
	.w7(32'h38826e65),
	.w8(32'h387a9503),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61954d5),
	.w1(32'hb783d27a),
	.w2(32'hb6db20f1),
	.w3(32'hb66e3ec2),
	.w4(32'hb729d1ba),
	.w5(32'hb71345ae),
	.w6(32'hb75f164d),
	.w7(32'hb6e4ddbf),
	.w8(32'hb70f9940),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908e84a),
	.w1(32'h3931647f),
	.w2(32'h384e20bb),
	.w3(32'h393a3350),
	.w4(32'h3936966e),
	.w5(32'h36af8a06),
	.w6(32'h38aededd),
	.w7(32'h38c4bc93),
	.w8(32'hb6e63ba6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368ab6db),
	.w1(32'h36385ecf),
	.w2(32'h35b9b864),
	.w3(32'h37382365),
	.w4(32'h36238604),
	.w5(32'hb48596a9),
	.w6(32'h36c277a5),
	.w7(32'hb6a01194),
	.w8(32'hb7344532),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d8ea),
	.w1(32'h398e3ef0),
	.w2(32'h39390bce),
	.w3(32'h3951c510),
	.w4(32'h390a2ac6),
	.w5(32'h3901ec90),
	.w6(32'h3953b974),
	.w7(32'h38c76334),
	.w8(32'h38f0b21e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995306d),
	.w1(32'h39f5164b),
	.w2(32'h39f7020c),
	.w3(32'hb859b25c),
	.w4(32'h39304732),
	.w5(32'h39adf79a),
	.w6(32'h38fdc845),
	.w7(32'h39724347),
	.w8(32'h39e82a56),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b35aa0),
	.w1(32'h3976d652),
	.w2(32'h39d63769),
	.w3(32'h399c8039),
	.w4(32'h381a7f80),
	.w5(32'h38d877cd),
	.w6(32'h39d73a07),
	.w7(32'h39aa0c73),
	.w8(32'h39ddbca2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1a7ca),
	.w1(32'h37defbbb),
	.w2(32'h37f7c360),
	.w3(32'hb84653b0),
	.w4(32'h36c8a01f),
	.w5(32'h369ab8f8),
	.w6(32'hb7b62f1f),
	.w7(32'h384dad00),
	.w8(32'h37dd480e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a510d8f),
	.w1(32'h3a48ae7a),
	.w2(32'h3a61ec40),
	.w3(32'h39508e18),
	.w4(32'h39644596),
	.w5(32'h39af3917),
	.w6(32'h39ca66de),
	.w7(32'h399019b8),
	.w8(32'h3a0eb0ef),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390edb78),
	.w1(32'h397dbcc1),
	.w2(32'h3969a290),
	.w3(32'h3981f537),
	.w4(32'h39a17089),
	.w5(32'h39c0a7be),
	.w6(32'h38ea28de),
	.w7(32'h399ee3fd),
	.w8(32'h39bf2f39),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb33ad222),
	.w1(32'hb70ffbaa),
	.w2(32'hb50bafc0),
	.w3(32'h36b00c4b),
	.w4(32'hb5e0269b),
	.w5(32'h36d62311),
	.w6(32'h369e98ff),
	.w7(32'h35a238fa),
	.w8(32'h36c9c072),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390548e1),
	.w1(32'h388f425e),
	.w2(32'hb81deac4),
	.w3(32'h38508577),
	.w4(32'h375dedd6),
	.w5(32'hb9165156),
	.w6(32'h388f2bff),
	.w7(32'h374535fd),
	.w8(32'h37946f11),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362c3130),
	.w1(32'hb78c7783),
	.w2(32'hb6a1749d),
	.w3(32'h37a5b466),
	.w4(32'h36113986),
	.w5(32'h375eb519),
	.w6(32'h3750176c),
	.w7(32'h3634671c),
	.w8(32'h36ea3c7e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8ad82),
	.w1(32'h39e0e77f),
	.w2(32'h3a0b9eed),
	.w3(32'h381acd08),
	.w4(32'h390c4cd0),
	.w5(32'h39959468),
	.w6(32'h395dcdac),
	.w7(32'h3987e519),
	.w8(32'h39ec878e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a26074),
	.w1(32'h39def9a3),
	.w2(32'h3a12c5ef),
	.w3(32'h3882c4f2),
	.w4(32'h3904f2b4),
	.w5(32'h394be4ce),
	.w6(32'h391b5774),
	.w7(32'h3997e2d8),
	.w8(32'h3959653d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6a1bb),
	.w1(32'h39988566),
	.w2(32'h39e11e0f),
	.w3(32'hb939a751),
	.w4(32'h3860c9ae),
	.w5(32'h389ce618),
	.w6(32'h38cc2384),
	.w7(32'h399f8100),
	.w8(32'h39a8c1f7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83d962c),
	.w1(32'hb8f0309d),
	.w2(32'hb87e7402),
	.w3(32'hb8c6399f),
	.w4(32'hb8c7dbc4),
	.w5(32'hb8818ce6),
	.w6(32'hb89977ec),
	.w7(32'hb8662dba),
	.w8(32'hb8455cdb),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38918b32),
	.w1(32'h39a78bd2),
	.w2(32'h3a30a1f4),
	.w3(32'hb9ae13d5),
	.w4(32'h372f1290),
	.w5(32'h39568923),
	.w6(32'h3907362d),
	.w7(32'h39b27e5e),
	.w8(32'h3a150000),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10ad0f),
	.w1(32'h39a3709a),
	.w2(32'h399d960b),
	.w3(32'h398a2997),
	.w4(32'h39964469),
	.w5(32'hb816372f),
	.w6(32'h39b1fae1),
	.w7(32'h395353ec),
	.w8(32'h396d275e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b71d8),
	.w1(32'h38e5ad01),
	.w2(32'h39d6f71b),
	.w3(32'hb977f242),
	.w4(32'hb98be27c),
	.w5(32'hb895b711),
	.w6(32'h39139570),
	.w7(32'h397174f2),
	.w8(32'h3a059ce8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37220e14),
	.w1(32'hb599ef09),
	.w2(32'hb6defd00),
	.w3(32'h37af8ebf),
	.w4(32'h36e4e1ab),
	.w5(32'h350f9401),
	.w6(32'h362fec75),
	.w7(32'hb699c6d7),
	.w8(32'hb7228a16),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb667c030),
	.w1(32'hb703a426),
	.w2(32'hb69a3c37),
	.w3(32'hb5ca39e2),
	.w4(32'hb527c01e),
	.w5(32'hb5c7f66b),
	.w6(32'hb6a76c9e),
	.w7(32'hb6aff5e4),
	.w8(32'hb68f382f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8fd0b),
	.w1(32'h39c10b1b),
	.w2(32'h39bafd9b),
	.w3(32'hb94a4358),
	.w4(32'hb8cd0a82),
	.w5(32'h383a061c),
	.w6(32'hb88e6b77),
	.w7(32'hb7f5b76b),
	.w8(32'h390eccf9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfe9a4),
	.w1(32'h3a2a5d48),
	.w2(32'h3a148f65),
	.w3(32'h382d02c7),
	.w4(32'h398dbe65),
	.w5(32'h3984e493),
	.w6(32'h39818665),
	.w7(32'h39f5db34),
	.w8(32'h3a32d79f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1d6dd),
	.w1(32'h39a1f66f),
	.w2(32'h39b02330),
	.w3(32'h3943280f),
	.w4(32'h3889814f),
	.w5(32'hb8a4a1cd),
	.w6(32'h39edb1a9),
	.w7(32'h39fcfe1f),
	.w8(32'h3a076578),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e0821),
	.w1(32'h39cc9f48),
	.w2(32'h39834394),
	.w3(32'hb94ce88a),
	.w4(32'hb92e3c2a),
	.w5(32'hb9a4ad89),
	.w6(32'hb8cbbfec),
	.w7(32'hb99a94fb),
	.w8(32'hb94472f4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aa379f),
	.w1(32'h312971c2),
	.w2(32'h3729646a),
	.w3(32'h38080c31),
	.w4(32'hb82296c3),
	.w5(32'hb7b13d98),
	.w6(32'hb85f2f06),
	.w7(32'hb7141feb),
	.w8(32'hb69b1b83),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a1c0d),
	.w1(32'h35c50f3c),
	.w2(32'h37c70039),
	.w3(32'hb8839411),
	.w4(32'hb8f61681),
	.w5(32'hb8a75291),
	.w6(32'h37332f52),
	.w7(32'hb71fddfc),
	.w8(32'hb6e0eb26),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6927f7),
	.w1(32'h3a3f4276),
	.w2(32'h3a4bfa8c),
	.w3(32'h3a805e0d),
	.w4(32'h3a163ac9),
	.w5(32'h3a77b0c1),
	.w6(32'h3a103d2e),
	.w7(32'h39236f60),
	.w8(32'h3a0080f0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4364af),
	.w1(32'h3a170d76),
	.w2(32'h3a24d77c),
	.w3(32'h38ab3900),
	.w4(32'hb8940c96),
	.w5(32'h3987bcd1),
	.w6(32'h38df0586),
	.w7(32'h3909c44c),
	.w8(32'h39ee1800),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d28ee),
	.w1(32'h39dcde74),
	.w2(32'h39d351d2),
	.w3(32'h3a07fd08),
	.w4(32'hb966a73d),
	.w5(32'h3894dc0c),
	.w6(32'h39e9328c),
	.w7(32'hb893e071),
	.w8(32'h39707404),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cb361c),
	.w1(32'h39056601),
	.w2(32'h39de7468),
	.w3(32'hb9492ae4),
	.w4(32'h37a7c5cc),
	.w5(32'h39b22110),
	.w6(32'h38a2ffec),
	.w7(32'h39724c7f),
	.w8(32'h39ad93e6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391876e9),
	.w1(32'h398e3ee3),
	.w2(32'h3a2629f6),
	.w3(32'hb90a2955),
	.w4(32'h38db7486),
	.w5(32'h396922e5),
	.w6(32'h39113650),
	.w7(32'h39b71d81),
	.w8(32'h39e4f5f9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e20020),
	.w1(32'hb632f1e6),
	.w2(32'hb5d87a03),
	.w3(32'h371e40a7),
	.w4(32'hb5959a46),
	.w5(32'h35076f60),
	.w6(32'h358e5bdd),
	.w7(32'hb59d70f5),
	.w8(32'h357c59ff),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6aeb4a0),
	.w1(32'hb6d4fbd9),
	.w2(32'hb6a8eb9b),
	.w3(32'hb65eebd0),
	.w4(32'hb62c6d7b),
	.w5(32'h34082911),
	.w6(32'hb64aae0c),
	.w7(32'hb6c37400),
	.w8(32'hb6873953),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d77aaa),
	.w1(32'hb92e549b),
	.w2(32'hb8ae90a1),
	.w3(32'hb94cd919),
	.w4(32'hb8feb6b4),
	.w5(32'hb85c8312),
	.w6(32'hb7aeb309),
	.w7(32'hb6c358c7),
	.w8(32'hb67028cd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36160302),
	.w1(32'hb6b249a0),
	.w2(32'hb6879abc),
	.w3(32'h36bc32a6),
	.w4(32'hb5a502d1),
	.w5(32'h36499ed2),
	.w6(32'hb67a7f8c),
	.w7(32'hb63a6074),
	.w8(32'h36dd8cf6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963f439),
	.w1(32'h39734b5a),
	.w2(32'h390f861b),
	.w3(32'h38755959),
	.w4(32'h38d4813d),
	.w5(32'h3912e476),
	.w6(32'h38a2dbf4),
	.w7(32'h38aae423),
	.w8(32'h38390532),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6f403),
	.w1(32'hb84984cc),
	.w2(32'h390a08cf),
	.w3(32'hb82c0e80),
	.w4(32'hb95c77f8),
	.w5(32'hb875999b),
	.w6(32'h391b7c66),
	.w7(32'h39a028fe),
	.w8(32'h3a06de93),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925bf6c),
	.w1(32'h39543e64),
	.w2(32'h3998b16b),
	.w3(32'h36eae77b),
	.w4(32'h38162008),
	.w5(32'h38e0fef4),
	.w6(32'h3969fd50),
	.w7(32'h39630aaa),
	.w8(32'h39aca104),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a0aff2),
	.w1(32'hb70b5ba7),
	.w2(32'hb6c01643),
	.w3(32'hb797918c),
	.w4(32'hb6a5b118),
	.w5(32'hb684af8d),
	.w6(32'hb7a4ce30),
	.w7(32'hb747388a),
	.w8(32'hb7192f8c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47b5bf),
	.w1(32'h3a0b75c2),
	.w2(32'h3a518ea7),
	.w3(32'h3a23583d),
	.w4(32'hb9a71d85),
	.w5(32'hb8178fef),
	.w6(32'h3a2db2a2),
	.w7(32'hb8ca898b),
	.w8(32'h39a20518),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9dfaa),
	.w1(32'h39c8b032),
	.w2(32'h39c56917),
	.w3(32'h38f1e2b2),
	.w4(32'h39023e78),
	.w5(32'h391815c3),
	.w6(32'h387b82f7),
	.w7(32'h390eff66),
	.w8(32'h3958e6c1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb551254d),
	.w1(32'hb72a4fda),
	.w2(32'hb751a088),
	.w3(32'h36d98567),
	.w4(32'hb652d091),
	.w5(32'hb5a47660),
	.w6(32'hb58afd46),
	.w7(32'hb5c0a2b4),
	.w8(32'hb651820a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2e477),
	.w1(32'h39a11598),
	.w2(32'h398f6924),
	.w3(32'hb7340f64),
	.w4(32'hb88dcb2b),
	.w5(32'h383772eb),
	.w6(32'h390fcfaa),
	.w7(32'hb70686c9),
	.w8(32'h384c269b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3f5e2f9),
	.w1(32'h382658e4),
	.w2(32'hb5a98417),
	.w3(32'h356395ae),
	.w4(32'h386edc18),
	.w5(32'hb65f1025),
	.w6(32'hb6aa1c8f),
	.w7(32'h383296c3),
	.w8(32'h35407717),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868693c),
	.w1(32'hb6f64e0f),
	.w2(32'hb81fc248),
	.w3(32'hb8f0b646),
	.w4(32'hb8e158e6),
	.w5(32'hb8eeae4c),
	.w6(32'hb8c93ff4),
	.w7(32'hb8dff71e),
	.w8(32'hb89c0cde),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f9450),
	.w1(32'hb721f10b),
	.w2(32'hb64e5757),
	.w3(32'hb64b5390),
	.w4(32'hb6a69e94),
	.w5(32'h35df3816),
	.w6(32'hb60d45eb),
	.w7(32'hb5a12a71),
	.w8(32'h360d258e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb755ec1d),
	.w1(32'hb6c45af1),
	.w2(32'hb6fc4ba9),
	.w3(32'hb71c2466),
	.w4(32'hb656ff3c),
	.w5(32'hb6d12c0a),
	.w6(32'hb713baf7),
	.w7(32'hb60ae844),
	.w8(32'hb6a7f427),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38984c4e),
	.w1(32'h38d36252),
	.w2(32'h39484026),
	.w3(32'h3766d4ee),
	.w4(32'h388a3c06),
	.w5(32'h39341ea7),
	.w6(32'h3927bae0),
	.w7(32'h39158fa3),
	.w8(32'h39445193),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6636e2),
	.w1(32'h3a23c460),
	.w2(32'h3a253790),
	.w3(32'h391fee96),
	.w4(32'h39750338),
	.w5(32'hb94e4423),
	.w6(32'h3988c511),
	.w7(32'h39946e7a),
	.w8(32'h3a10b6a9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08193e),
	.w1(32'h3a019c78),
	.w2(32'h3a179ad9),
	.w3(32'h3940af58),
	.w4(32'h391a03d8),
	.w5(32'h3905b423),
	.w6(32'h39820af8),
	.w7(32'h38f7b8f5),
	.w8(32'h398e952a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14cbf5),
	.w1(32'h3a4261a6),
	.w2(32'h3a1c2467),
	.w3(32'hb6c4e06f),
	.w4(32'h398a2285),
	.w5(32'h38837f52),
	.w6(32'h3972fbdd),
	.w7(32'h3976d5aa),
	.w8(32'h39c8c567),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a6d706),
	.w1(32'h3607dd70),
	.w2(32'hb6736655),
	.w3(32'h371046b2),
	.w4(32'hb6264e2f),
	.w5(32'hb761c5d7),
	.w6(32'hb6156c01),
	.w7(32'hb4ea5fdb),
	.w8(32'hb728f20c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ed3f59),
	.w1(32'hb7adc59b),
	.w2(32'hb7be2b3b),
	.w3(32'hb8a1aaa1),
	.w4(32'hb88e4ee1),
	.w5(32'hb8584d01),
	.w6(32'hb7dfcc5a),
	.w7(32'h366cdefc),
	.w8(32'h3709e1eb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ac5d21),
	.w1(32'hb66b501b),
	.w2(32'hb60c5d3c),
	.w3(32'h372aa141),
	.w4(32'h36853d56),
	.w5(32'h36e05cf5),
	.w6(32'hb5862904),
	.w7(32'h35eaeb8c),
	.w8(32'h35ac17fd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60c87dc),
	.w1(32'hb648255a),
	.w2(32'hb6680c0e),
	.w3(32'h343f12a9),
	.w4(32'hb48589d1),
	.w5(32'hb56fe40b),
	.w6(32'hb5d824db),
	.w7(32'h3519044b),
	.w8(32'hb64c1e4b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab3b54),
	.w1(32'h390053df),
	.w2(32'h39d03509),
	.w3(32'hb8871039),
	.w4(32'hb7a74fef),
	.w5(32'hb702c1b6),
	.w6(32'h382f744f),
	.w7(32'h38c14e64),
	.w8(32'h399e4a1d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb749d3a6),
	.w1(32'hb845e7f2),
	.w2(32'hb8f7794b),
	.w3(32'h386ab247),
	.w4(32'hb72a5d29),
	.w5(32'hb8be702a),
	.w6(32'hb789aba7),
	.w7(32'hb8815fb2),
	.w8(32'hb8c019f3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390bdcc7),
	.w1(32'h38ad1f51),
	.w2(32'h38c0f5ed),
	.w3(32'h38376b73),
	.w4(32'hb6fd4a0f),
	.w5(32'h37d25bbf),
	.w6(32'hb75edff8),
	.w7(32'h3817aed7),
	.w8(32'hb5db9b67),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890a1e2),
	.w1(32'h3912e6d5),
	.w2(32'h393f43e1),
	.w3(32'h3681c5da),
	.w4(32'hb6413d16),
	.w5(32'h37ad9b37),
	.w6(32'hb710d8b8),
	.w7(32'h3839ccf7),
	.w8(32'h389c2cc1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38053389),
	.w1(32'h379c2fb4),
	.w2(32'h36a907de),
	.w3(32'h3826d1c1),
	.w4(32'h372bc768),
	.w5(32'hb66b6677),
	.w6(32'h37cdde89),
	.w7(32'h377a8e0e),
	.w8(32'hb4eb6711),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39169bf3),
	.w1(32'h38e2900a),
	.w2(32'h392af50b),
	.w3(32'hb744f6a6),
	.w4(32'hb792a7a6),
	.w5(32'h3822829d),
	.w6(32'h37e409b8),
	.w7(32'h382c88cb),
	.w8(32'h38f5e520),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373b62ec),
	.w1(32'hb66f7b5e),
	.w2(32'hb7db6537),
	.w3(32'hb7f53f8f),
	.w4(32'hb78cde93),
	.w5(32'hb7adaff2),
	.w6(32'hb7bea36d),
	.w7(32'h37b1c515),
	.w8(32'h378ba530),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965aa84),
	.w1(32'h36b0c940),
	.w2(32'h3a325447),
	.w3(32'hba4b36fe),
	.w4(32'hba058cee),
	.w5(32'hba11796d),
	.w6(32'hb9b3158a),
	.w7(32'hb93229b3),
	.w8(32'h38ada7eb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ecc4e2),
	.w1(32'hb9d2db21),
	.w2(32'hb9e3bece),
	.w3(32'hb7f923a5),
	.w4(32'hba0bbd7e),
	.w5(32'hb97b1c8f),
	.w6(32'hb99a7640),
	.w7(32'hb9f86741),
	.w8(32'hb9078fe8),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95529ae),
	.w1(32'hb8ceec79),
	.w2(32'hb6ce6192),
	.w3(32'hb9624a83),
	.w4(32'hb9751a95),
	.w5(32'hb853b5a2),
	.w6(32'h37adaa15),
	.w7(32'h39059244),
	.w8(32'h395609a1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule