module layer_8_featuremap_176(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0e119),
	.w1(32'hbbe6f6b7),
	.w2(32'hbbff821c),
	.w3(32'hbbd89d88),
	.w4(32'h3a84176e),
	.w5(32'hba73546a),
	.w6(32'h3b0d8c7f),
	.w7(32'h3ae93bc0),
	.w8(32'h3a98b4ce),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85360f),
	.w1(32'hbcf33018),
	.w2(32'hbd096c7c),
	.w3(32'hbc0e0be0),
	.w4(32'hbc760806),
	.w5(32'hbcaac70b),
	.w6(32'hbc5d3e06),
	.w7(32'hbc373648),
	.w8(32'h3c330387),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadea26),
	.w1(32'hb9163999),
	.w2(32'h3977a87f),
	.w3(32'h3b73dc19),
	.w4(32'hb81fab57),
	.w5(32'h3a64de96),
	.w6(32'hb991c95e),
	.w7(32'hbb859fbb),
	.w8(32'hbb4381f6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0739fa),
	.w1(32'hbb8f409f),
	.w2(32'hba4d9f8f),
	.w3(32'hbaa41a1c),
	.w4(32'hbb8ebd4c),
	.w5(32'hbbdde1a7),
	.w6(32'hbb29e8d3),
	.w7(32'hb91a9b94),
	.w8(32'hbb3486aa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d1056),
	.w1(32'hbcb4d26d),
	.w2(32'hbcb8a953),
	.w3(32'hbbbdd624),
	.w4(32'hbb2b5630),
	.w5(32'hbbb7974d),
	.w6(32'hbc3ad416),
	.w7(32'hbc7b454d),
	.w8(32'hbb91bbc6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc457309),
	.w1(32'hbc12a91f),
	.w2(32'h3be409a0),
	.w3(32'hba76303a),
	.w4(32'hbb1e8b86),
	.w5(32'hba6a109b),
	.w6(32'h3a434070),
	.w7(32'h3c0362e3),
	.w8(32'hbb606055),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2883),
	.w1(32'h3cdd7ce0),
	.w2(32'h3d0ef4f0),
	.w3(32'h3ac2b320),
	.w4(32'h3c9818a8),
	.w5(32'h3cd829df),
	.w6(32'h3bf14c2a),
	.w7(32'h3c15fc29),
	.w8(32'hbc36a294),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ca79a),
	.w1(32'hba7ea28c),
	.w2(32'h3aaf5e7d),
	.w3(32'hbb40a6eb),
	.w4(32'hbb11d81f),
	.w5(32'hbbafe8f0),
	.w6(32'h3b7a1d0a),
	.w7(32'h3b0215a2),
	.w8(32'hba94dde9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0467d7),
	.w1(32'h3b1f698b),
	.w2(32'h3c156d45),
	.w3(32'h3b4c3941),
	.w4(32'h3c76f9d8),
	.w5(32'h3cb7a722),
	.w6(32'hbb971e54),
	.w7(32'hbae7455f),
	.w8(32'h3b5dc98f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b411384),
	.w1(32'hbaddda33),
	.w2(32'hbc175a8b),
	.w3(32'h3c84cb6b),
	.w4(32'hbb4b5364),
	.w5(32'hbabaaee6),
	.w6(32'h3a8c836a),
	.w7(32'h3a24dd6c),
	.w8(32'hbbc4ac9f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecb4ee),
	.w1(32'hbc1de843),
	.w2(32'hbc36e32f),
	.w3(32'hbae57da6),
	.w4(32'hbb51e805),
	.w5(32'hbbca1f0b),
	.w6(32'hba7eb8ec),
	.w7(32'hbbbc4583),
	.w8(32'hb928a3be),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992f27),
	.w1(32'hbb445e93),
	.w2(32'hbb57f055),
	.w3(32'hbae0184e),
	.w4(32'h3b607ce4),
	.w5(32'hbb4bd9a8),
	.w6(32'h3a1a4801),
	.w7(32'h3b28346c),
	.w8(32'hbaae4c10),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc404e07),
	.w1(32'h3ae70d5e),
	.w2(32'hba1cba98),
	.w3(32'hbc3665c2),
	.w4(32'hbad50c38),
	.w5(32'h39ab08c2),
	.w6(32'hbac2b450),
	.w7(32'hbb3e9623),
	.w8(32'hbb8cf6f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c739f),
	.w1(32'hbbe4d7b9),
	.w2(32'hb98c0646),
	.w3(32'hbbb06c7f),
	.w4(32'hbba2fe1d),
	.w5(32'hbaba5dc4),
	.w6(32'hbbd06603),
	.w7(32'hbb4d6258),
	.w8(32'hbb84e307),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d4f52),
	.w1(32'hbc93a2da),
	.w2(32'hbca27094),
	.w3(32'h3bc27b14),
	.w4(32'hbcc1288b),
	.w5(32'hbcd89f1c),
	.w6(32'hbc69fd94),
	.w7(32'hbc04a081),
	.w8(32'hbaae48ac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7dfa5),
	.w1(32'hba73c61f),
	.w2(32'hba04a3d4),
	.w3(32'hbc61f260),
	.w4(32'hbaa1d5be),
	.w5(32'hba3780da),
	.w6(32'hb9aa87e4),
	.w7(32'h38b8309f),
	.w8(32'hbb9b8923),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba118a44),
	.w1(32'h3acc07c0),
	.w2(32'h3b590c3f),
	.w3(32'hba87c648),
	.w4(32'hb8a06f41),
	.w5(32'hbb8af478),
	.w6(32'h3a83dbe9),
	.w7(32'h3bc07c16),
	.w8(32'h394fb423),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6879),
	.w1(32'hbc17e23e),
	.w2(32'hbbaefdb0),
	.w3(32'hbbdfed39),
	.w4(32'hbb434886),
	.w5(32'hbba453ed),
	.w6(32'hbb5fbf63),
	.w7(32'h3ab1f1f2),
	.w8(32'hbab05093),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba989c4),
	.w1(32'h38b6e6e9),
	.w2(32'hbb7fe96c),
	.w3(32'h3b236821),
	.w4(32'h3bc1c536),
	.w5(32'hbb857d13),
	.w6(32'h3cbe4f21),
	.w7(32'h3c87a101),
	.w8(32'h3c0e0854),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139c8c),
	.w1(32'h3d0f887e),
	.w2(32'h3d39c0ee),
	.w3(32'hbb9e72d0),
	.w4(32'h3c911177),
	.w5(32'h3d07ffa1),
	.w6(32'h3c30d345),
	.w7(32'h3c6c5270),
	.w8(32'hbca64718),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbde60),
	.w1(32'h3a4e1290),
	.w2(32'hbb0fb48b),
	.w3(32'hbb2b35de),
	.w4(32'hbae20231),
	.w5(32'hbbd0c246),
	.w6(32'hb9f9f3f3),
	.w7(32'hbbcb6b9d),
	.w8(32'hbbd4261d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf290a5),
	.w1(32'hb83865fd),
	.w2(32'h39c27c39),
	.w3(32'hbaec7dd9),
	.w4(32'hb9204a86),
	.w5(32'h3b42b82c),
	.w6(32'hbbc290b6),
	.w7(32'hbb212ca3),
	.w8(32'hb902cb2c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4464e),
	.w1(32'hbb911731),
	.w2(32'hbc56d0dd),
	.w3(32'h3c341730),
	.w4(32'h3a1ad9ad),
	.w5(32'hbbc59e89),
	.w6(32'h3c2d819b),
	.w7(32'h3ba38e8c),
	.w8(32'h3bf1ac26),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5f66f),
	.w1(32'h37813a33),
	.w2(32'hb9e6fd0a),
	.w3(32'h3ade9006),
	.w4(32'hbb4adb8f),
	.w5(32'hba675197),
	.w6(32'hbc18042c),
	.w7(32'hbbe592bb),
	.w8(32'hbc21b12e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44a8a6),
	.w1(32'h3beebfcf),
	.w2(32'hb6ee109c),
	.w3(32'hbb29cdc2),
	.w4(32'hb8813e57),
	.w5(32'hbae57cfc),
	.w6(32'h3b31780e),
	.w7(32'h39a65454),
	.w8(32'hba98e8ae),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa306c5),
	.w1(32'hbc03d53d),
	.w2(32'hbbe428eb),
	.w3(32'hbac0e30f),
	.w4(32'h3ab5770b),
	.w5(32'hbad5fd41),
	.w6(32'h3c2bcad1),
	.w7(32'h3990ef98),
	.w8(32'hba8cd96b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ccd39),
	.w1(32'h3aada976),
	.w2(32'hbb47e8d2),
	.w3(32'hbbbc5bf8),
	.w4(32'h3b1f1969),
	.w5(32'hba00cdd8),
	.w6(32'hba4a607d),
	.w7(32'h3ac78af7),
	.w8(32'hbb79569a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37ac17),
	.w1(32'hbb8af99c),
	.w2(32'hbc858265),
	.w3(32'h3cb11b5a),
	.w4(32'h3c3fad5a),
	.w5(32'hbc469ae1),
	.w6(32'h3d388af8),
	.w7(32'h3c22411d),
	.w8(32'h3b979b57),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ae269),
	.w1(32'hbab34f69),
	.w2(32'h3c1f2c43),
	.w3(32'hbbbdb07f),
	.w4(32'h3b7734a6),
	.w5(32'h3c6677fb),
	.w6(32'h3b2c2118),
	.w7(32'h3c3bc8ac),
	.w8(32'h3c66f0ee),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d5ee5),
	.w1(32'h3ab16f5f),
	.w2(32'hbaf223e1),
	.w3(32'h3c8248c9),
	.w4(32'h3a01dad8),
	.w5(32'hbb8213b4),
	.w6(32'hb91703be),
	.w7(32'h3b1ce100),
	.w8(32'hbc2bb243),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc974cb6),
	.w1(32'h3bd3f588),
	.w2(32'h3c007d46),
	.w3(32'hbcc30469),
	.w4(32'h3bae07d1),
	.w5(32'h3b8eca43),
	.w6(32'h39ab3b47),
	.w7(32'hbb2dea37),
	.w8(32'hbb587a3c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a9fd4),
	.w1(32'hbb99efb2),
	.w2(32'hb97eb153),
	.w3(32'h3b6e7d07),
	.w4(32'hbb3dde7f),
	.w5(32'hbb4d079a),
	.w6(32'hbc0263ca),
	.w7(32'hbbf0fd97),
	.w8(32'hbb817266),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b521206),
	.w1(32'h3ba2b060),
	.w2(32'hb97f9f80),
	.w3(32'h3b1ead13),
	.w4(32'h3b7bebf5),
	.w5(32'h3b433fb9),
	.w6(32'h3bbdf1da),
	.w7(32'h3b94dd2d),
	.w8(32'hbb118595),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbfad8),
	.w1(32'h3b59473f),
	.w2(32'h3a0b788a),
	.w3(32'hbbb0df8d),
	.w4(32'h3b67d409),
	.w5(32'h3b0b94f3),
	.w6(32'h3b9ee1bb),
	.w7(32'h3b0444ff),
	.w8(32'hbb862fdd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b699a5b),
	.w1(32'h3b5a5f24),
	.w2(32'h3bee04b2),
	.w3(32'hbaf82310),
	.w4(32'h3aa92f59),
	.w5(32'h39f3dde7),
	.w6(32'hbbe9f7a9),
	.w7(32'hbac3a5ea),
	.w8(32'hbb1dd60d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4721df),
	.w1(32'hbbb50058),
	.w2(32'hbaf77ffb),
	.w3(32'hbb2f98dd),
	.w4(32'hba3fc30d),
	.w5(32'hbae0e14c),
	.w6(32'h3b2fa16b),
	.w7(32'h3b21669d),
	.w8(32'h3b871119),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20606d),
	.w1(32'hbbd3e6db),
	.w2(32'hbbad5691),
	.w3(32'hba812803),
	.w4(32'hbaf09237),
	.w5(32'hbb1a64d1),
	.w6(32'hbc1c3fc6),
	.w7(32'hbc0877df),
	.w8(32'hbc399f7d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc9b0d),
	.w1(32'hbd64cab2),
	.w2(32'hbd94b9c3),
	.w3(32'hbba439fe),
	.w4(32'hbd302977),
	.w5(32'hbd7bf047),
	.w6(32'hbcb3526f),
	.w7(32'hbcb2b9d3),
	.w8(32'h3c8b64b3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc317b97),
	.w1(32'hbb4fa92d),
	.w2(32'hbb47544e),
	.w3(32'hbc29bd83),
	.w4(32'h3be4e732),
	.w5(32'h3b42c681),
	.w6(32'hbba68158),
	.w7(32'h3a7d1338),
	.w8(32'hbb8b46ac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e5701),
	.w1(32'h3b0ba1af),
	.w2(32'hba912df3),
	.w3(32'h3b9efc0b),
	.w4(32'hbb42c335),
	.w5(32'hbb7b1ace),
	.w6(32'h399880bb),
	.w7(32'hbaafcb24),
	.w8(32'hbad406d2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a81d5),
	.w1(32'hbc6510f1),
	.w2(32'hbc926bf4),
	.w3(32'hbca1f8a7),
	.w4(32'hbc0348f6),
	.w5(32'hbc794532),
	.w6(32'h3b261ad5),
	.w7(32'h3b923b40),
	.w8(32'hba950dce),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00046b),
	.w1(32'h3c5ca866),
	.w2(32'h3a4dfc50),
	.w3(32'hbab4354c),
	.w4(32'h3be4a351),
	.w5(32'hbb29bcef),
	.w6(32'h3c080d9c),
	.w7(32'h3ab20453),
	.w8(32'hbbf24059),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b5e10),
	.w1(32'h39997f72),
	.w2(32'hbad667bc),
	.w3(32'hbb9de70d),
	.w4(32'h39ec1d37),
	.w5(32'hba9cdce8),
	.w6(32'hbafb62aa),
	.w7(32'hbb48ea13),
	.w8(32'hbaabf14b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7713b),
	.w1(32'hbb787a63),
	.w2(32'hbb55e00d),
	.w3(32'hbb5e8317),
	.w4(32'hbbff756d),
	.w5(32'hbba43e15),
	.w6(32'hbc02af28),
	.w7(32'hbba64899),
	.w8(32'hbbd1b380),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978a12),
	.w1(32'hbba7f2f2),
	.w2(32'hbba17cc6),
	.w3(32'hb9e9be07),
	.w4(32'hbb5ed36d),
	.w5(32'hbc24309a),
	.w6(32'h3bf6b330),
	.w7(32'h3ae60141),
	.w8(32'h3b2eb2b7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a6e51),
	.w1(32'hbc2f32e0),
	.w2(32'h3c0f3ce6),
	.w3(32'hbb8bfdf0),
	.w4(32'hbc95ee6c),
	.w5(32'hba4548a2),
	.w6(32'hbcc5e1fc),
	.w7(32'hbbff059b),
	.w8(32'hbc8e00ab),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fe49b),
	.w1(32'h39fc3d68),
	.w2(32'h3ae4d781),
	.w3(32'hbbd985d1),
	.w4(32'hb9026095),
	.w5(32'hb994a6ef),
	.w6(32'hbb1c617b),
	.w7(32'hbb6a96d3),
	.w8(32'hbbb2fec4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e4f87),
	.w1(32'hbb592a55),
	.w2(32'hbbb43215),
	.w3(32'h3aa28e99),
	.w4(32'hba8bfa84),
	.w5(32'hbc134317),
	.w6(32'h3aa08312),
	.w7(32'h3b084254),
	.w8(32'h3b52b8f1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2a7e),
	.w1(32'hbaf34470),
	.w2(32'hbba98f4f),
	.w3(32'hba9bdceb),
	.w4(32'h3acac583),
	.w5(32'hba22801f),
	.w6(32'hbadae3e1),
	.w7(32'h3b0d11cb),
	.w8(32'h3b72dbab),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6418b2),
	.w1(32'hbbb06cbe),
	.w2(32'h3b097f69),
	.w3(32'h3a100b56),
	.w4(32'hbaec1060),
	.w5(32'hbb30943e),
	.w6(32'h3a34aca5),
	.w7(32'hbaac5900),
	.w8(32'h3b9fd2b8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba20310),
	.w1(32'hbc71cb3d),
	.w2(32'hbd028b79),
	.w3(32'hbc22085d),
	.w4(32'hbc85e0de),
	.w5(32'hbcaa9161),
	.w6(32'hbc1d1a11),
	.w7(32'hbc0560c5),
	.w8(32'h3bba1a29),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987b7d),
	.w1(32'hb98418d0),
	.w2(32'h3b890666),
	.w3(32'hbb9440c3),
	.w4(32'hbc012c74),
	.w5(32'hbc227571),
	.w6(32'h3c80a8b9),
	.w7(32'h3c860538),
	.w8(32'h3c177670),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d71d),
	.w1(32'hbda56473),
	.w2(32'hbdd050ef),
	.w3(32'h3a5e4da4),
	.w4(32'hbd83996f),
	.w5(32'hbdb1f1e9),
	.w6(32'hbd131f46),
	.w7(32'hbd20f02e),
	.w8(32'h3bd1daa9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b8ad3),
	.w1(32'hbacdf2ac),
	.w2(32'hbc0e54e2),
	.w3(32'hbcc8c430),
	.w4(32'h3b5945c0),
	.w5(32'hba4b9272),
	.w6(32'h3ae83d30),
	.w7(32'hbb7eba6b),
	.w8(32'h39fb2ad1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ee3a2),
	.w1(32'hbb1e2e79),
	.w2(32'h3b831e19),
	.w3(32'h3b60d6c5),
	.w4(32'hba846ab0),
	.w5(32'hb91a8bac),
	.w6(32'hb94b13e4),
	.w7(32'hb9a636e9),
	.w8(32'hbb017e6e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13e461),
	.w1(32'hbc3fb878),
	.w2(32'hbc6caf1a),
	.w3(32'hba184cd7),
	.w4(32'hbbefaca4),
	.w5(32'hbc1f1019),
	.w6(32'h3b42b667),
	.w7(32'hbbaee16f),
	.w8(32'h3af5bf62),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecbf23),
	.w1(32'h3b9918ec),
	.w2(32'hbc064d76),
	.w3(32'hbb4c008d),
	.w4(32'h3b0f2547),
	.w5(32'hbb8636b6),
	.w6(32'h3bcafe98),
	.w7(32'hbc03e343),
	.w8(32'hbb47e1f3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd985e5),
	.w1(32'hbbfbf907),
	.w2(32'h3aec79d9),
	.w3(32'hbc4b03da),
	.w4(32'hbba5d683),
	.w5(32'hbb06c381),
	.w6(32'hbbccb5b1),
	.w7(32'hba64c90b),
	.w8(32'hbb71da86),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724831),
	.w1(32'hbc3803bc),
	.w2(32'hbc46dd0e),
	.w3(32'hbb984426),
	.w4(32'hbc103e22),
	.w5(32'hbc62cebe),
	.w6(32'hb9a3a134),
	.w7(32'hbb0f18ed),
	.w8(32'h3bca3eea),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49740f),
	.w1(32'hbb84dce0),
	.w2(32'hbbfdbefe),
	.w3(32'hbb341cb2),
	.w4(32'hbbc79c5e),
	.w5(32'hbbcdf1a5),
	.w6(32'hbb916a9c),
	.w7(32'hbc05d879),
	.w8(32'hbbef5034),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98a18a),
	.w1(32'h3b96b82d),
	.w2(32'h3af31040),
	.w3(32'h3a0bd916),
	.w4(32'hbaaf8b62),
	.w5(32'hbbbbcdef),
	.w6(32'hbb2f345f),
	.w7(32'hbb66ad19),
	.w8(32'hbc16e7ec),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba742bd3),
	.w1(32'h3bc374bb),
	.w2(32'h3be707c6),
	.w3(32'hbbf845c0),
	.w4(32'h3c5e75de),
	.w5(32'h3c640203),
	.w6(32'hbb2c78d0),
	.w7(32'hbb0da29f),
	.w8(32'hbbc63104),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0b44),
	.w1(32'hbc8d375c),
	.w2(32'hbc47d150),
	.w3(32'h3c0e928e),
	.w4(32'hbc5638f1),
	.w5(32'hbc404765),
	.w6(32'hbbb29d48),
	.w7(32'hbbb05324),
	.w8(32'hbc58e781),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc175d89),
	.w1(32'h3c3eef07),
	.w2(32'h3c268b11),
	.w3(32'hbc22ff0c),
	.w4(32'h3c1e5ba8),
	.w5(32'h3bf8750c),
	.w6(32'h3c5c0d2b),
	.w7(32'h3c191933),
	.w8(32'h3c0cef71),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9af31),
	.w1(32'hbcbf7091),
	.w2(32'hbcfb826f),
	.w3(32'h3bc7fb5a),
	.w4(32'hbca8e1fc),
	.w5(32'hbcf68fc9),
	.w6(32'hbb8f5231),
	.w7(32'hb9b76d9b),
	.w8(32'h3ca5cdad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92d426),
	.w1(32'h3a144e99),
	.w2(32'h381cc7e1),
	.w3(32'h3b537953),
	.w4(32'hb9bd7ca3),
	.w5(32'h3b519b29),
	.w6(32'h3a8419c2),
	.w7(32'h3b089575),
	.w8(32'hb915f619),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae82074),
	.w1(32'h38b6c031),
	.w2(32'hbab07826),
	.w3(32'h3a9bd509),
	.w4(32'hbb061ca6),
	.w5(32'hbb5f03b1),
	.w6(32'h3a440050),
	.w7(32'hb90abd80),
	.w8(32'hba35efc0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913929),
	.w1(32'hbb8338b0),
	.w2(32'hbc1a3a2f),
	.w3(32'hbb10103e),
	.w4(32'hba6a9908),
	.w5(32'hbb320e19),
	.w6(32'h3b016ee3),
	.w7(32'hbb4e2aaa),
	.w8(32'hbc15783d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27917e),
	.w1(32'hbb9c1e80),
	.w2(32'h3af4bc7d),
	.w3(32'hbbcbf950),
	.w4(32'hbb7a8a60),
	.w5(32'h3b8e6f5a),
	.w6(32'hbbd7f693),
	.w7(32'hbb018e42),
	.w8(32'hbb34204f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef4a3),
	.w1(32'h3b3904e8),
	.w2(32'hba462ff9),
	.w3(32'h3b7e4eb1),
	.w4(32'h3ae430ec),
	.w5(32'hbb737a21),
	.w6(32'h3c5c7ad5),
	.w7(32'h3b83e6f8),
	.w8(32'h3be1ab38),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bd37a),
	.w1(32'h3c941179),
	.w2(32'h3c84ad22),
	.w3(32'h3a4e945d),
	.w4(32'h3c474749),
	.w5(32'h3c1ab940),
	.w6(32'h3c991bec),
	.w7(32'h3c8cd911),
	.w8(32'h3cb54314),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4d0ff),
	.w1(32'hbbec8cb8),
	.w2(32'hbba82de6),
	.w3(32'h3c97613c),
	.w4(32'hb9982512),
	.w5(32'hbb810589),
	.w6(32'hbab2f2a0),
	.w7(32'hbaac0ce1),
	.w8(32'hbaa646d0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4988b0),
	.w1(32'h3b36639f),
	.w2(32'hb95bda8e),
	.w3(32'hba8bbee4),
	.w4(32'hbb3335b1),
	.w5(32'hbb2d46e4),
	.w6(32'h3a6ad5ff),
	.w7(32'h39f59f03),
	.w8(32'hbaea7a3d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c619a),
	.w1(32'hbc11b8cb),
	.w2(32'hbbfaca47),
	.w3(32'hba443dc2),
	.w4(32'hbbc43dfe),
	.w5(32'hbc02f7c8),
	.w6(32'hbb4db5fa),
	.w7(32'hbb41a9e3),
	.w8(32'hbb67f0b4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ecc0),
	.w1(32'h3be744b2),
	.w2(32'h3c00ac54),
	.w3(32'hbbafbca4),
	.w4(32'h3c09b89c),
	.w5(32'h3b8d1c79),
	.w6(32'h39ab63eb),
	.w7(32'h3ab45ce3),
	.w8(32'h3b166475),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec1123),
	.w1(32'hbb4f3c1b),
	.w2(32'hbb7d8d5c),
	.w3(32'h3c050b52),
	.w4(32'hbb8f408e),
	.w5(32'hbbdb72d5),
	.w6(32'h3c2230c2),
	.w7(32'h3b70a767),
	.w8(32'h3b49cf36),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4eaa72),
	.w1(32'hba83fee1),
	.w2(32'h3acc9675),
	.w3(32'h3a1758b8),
	.w4(32'h3b1dfda4),
	.w5(32'hbb9873a7),
	.w6(32'h3aff3d75),
	.w7(32'hbb22088d),
	.w8(32'h39c18d82),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1ec22),
	.w1(32'h3a18aab6),
	.w2(32'hbbe5e8c1),
	.w3(32'h3b39594b),
	.w4(32'h3be36248),
	.w5(32'hbbd91d3a),
	.w6(32'h3c4d1c79),
	.w7(32'h39257f18),
	.w8(32'hba638448),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f3bee),
	.w1(32'h3b9ea1b4),
	.w2(32'h3acde723),
	.w3(32'hbbbead22),
	.w4(32'hbb7d2f98),
	.w5(32'hbba74627),
	.w6(32'h3b3a6a49),
	.w7(32'h3b6ee82c),
	.w8(32'h3992c2d9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54cb19),
	.w1(32'hb94e7afe),
	.w2(32'hbb8f3233),
	.w3(32'hb9ee640d),
	.w4(32'hba8b8c1c),
	.w5(32'hb9b75541),
	.w6(32'hbbccc6a0),
	.w7(32'hbae2b20c),
	.w8(32'hbb27f7c0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb469c33),
	.w1(32'h3b8337ff),
	.w2(32'h3bb5e072),
	.w3(32'h3b5cc35c),
	.w4(32'h3bc966ec),
	.w5(32'h3bb34c2c),
	.w6(32'h3b3ac961),
	.w7(32'h3b9a3ec7),
	.w8(32'h3b859f71),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29faa),
	.w1(32'hbbf18261),
	.w2(32'hbb0b9b87),
	.w3(32'h39582f1c),
	.w4(32'hbc02bd71),
	.w5(32'hba416a9f),
	.w6(32'hbbf56562),
	.w7(32'hbc2007f8),
	.w8(32'hbc03a19a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dfacd9),
	.w1(32'hbba5262e),
	.w2(32'hbc032b9f),
	.w3(32'hbac9f1e7),
	.w4(32'h3808b025),
	.w5(32'hbc271544),
	.w6(32'h3c183266),
	.w7(32'h3bb61ad6),
	.w8(32'h3bb69e14),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6d480),
	.w1(32'hbc8dcdf3),
	.w2(32'hbc754044),
	.w3(32'hbc96aa45),
	.w4(32'hbc3abee9),
	.w5(32'hbc9bbd51),
	.w6(32'hbb438fb9),
	.w7(32'h3b1f0ac6),
	.w8(32'hbc1f6e91),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0f3b6),
	.w1(32'hbc232a33),
	.w2(32'hbc258d33),
	.w3(32'hbbb9f55d),
	.w4(32'hbbb3ce80),
	.w5(32'hbc258c45),
	.w6(32'h3b1f5a27),
	.w7(32'h3bc8d07a),
	.w8(32'hba794762),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a652c52),
	.w1(32'hbb5bc613),
	.w2(32'hb9d77d59),
	.w3(32'h3bb07fc3),
	.w4(32'hbbc411bb),
	.w5(32'hbba27ca3),
	.w6(32'h3bc922b2),
	.w7(32'h3addcd5f),
	.w8(32'h3b9b0cf4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f20ad),
	.w1(32'h3b6e1cdd),
	.w2(32'h3b7ef3fb),
	.w3(32'hbab0aebe),
	.w4(32'hbb792239),
	.w5(32'hba693c1e),
	.w6(32'h3bf62719),
	.w7(32'h3bbd9d70),
	.w8(32'h3bb7684c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac39526),
	.w1(32'h3bce1edf),
	.w2(32'h3bccef3b),
	.w3(32'hbb3e4ac4),
	.w4(32'hb9d9978e),
	.w5(32'hbaaed584),
	.w6(32'h3b9dffbc),
	.w7(32'h3c21bcc2),
	.w8(32'h3b17d608),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5746),
	.w1(32'h3a4eb964),
	.w2(32'h3a4007ce),
	.w3(32'hbaa29ea7),
	.w4(32'hbb8c500f),
	.w5(32'hbb920c23),
	.w6(32'hbaa46d8b),
	.w7(32'hba8aab86),
	.w8(32'hb9b2ebfc),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba1fa6),
	.w1(32'hba94c4f0),
	.w2(32'h3b0382c3),
	.w3(32'hbb8c860e),
	.w4(32'hba05c18e),
	.w5(32'hbb5e1398),
	.w6(32'h3ac5b197),
	.w7(32'h3b59ce83),
	.w8(32'h3b8fc2ce),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ccd5b),
	.w1(32'hbbaf5156),
	.w2(32'hbbb296cb),
	.w3(32'hbb6bfcf4),
	.w4(32'hbb458b08),
	.w5(32'hbbd3908d),
	.w6(32'hba4be924),
	.w7(32'hbbf836a0),
	.w8(32'hbbf96a70),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc64128),
	.w1(32'hbaa7ebca),
	.w2(32'h3af1aec9),
	.w3(32'hbaa27bc1),
	.w4(32'h3b50c257),
	.w5(32'h3addf225),
	.w6(32'hbba10aca),
	.w7(32'hbaca8343),
	.w8(32'h39dcb371),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910b94),
	.w1(32'h3c337afc),
	.w2(32'h3c98368b),
	.w3(32'h3b472877),
	.w4(32'h3c1b1993),
	.w5(32'h3cb00801),
	.w6(32'h39a95f33),
	.w7(32'h3b5afda4),
	.w8(32'hbb326ae7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155746),
	.w1(32'hba97e2f5),
	.w2(32'hba1d72a0),
	.w3(32'h3c41646d),
	.w4(32'h3b7f2fad),
	.w5(32'h3b8ef8ee),
	.w6(32'h3b4dfc2d),
	.w7(32'h3bb76211),
	.w8(32'h3bf97a37),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c059),
	.w1(32'h38e7b420),
	.w2(32'h3b0aa0c9),
	.w3(32'h3c2807d6),
	.w4(32'h3b916691),
	.w5(32'h3b5ad123),
	.w6(32'hbaedcc4a),
	.w7(32'hba958309),
	.w8(32'hbb0efe2a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5261),
	.w1(32'hbc083e30),
	.w2(32'hbc1428fc),
	.w3(32'h3aabef69),
	.w4(32'hbc2d665e),
	.w5(32'hbc4465f8),
	.w6(32'hbb8662a7),
	.w7(32'hbb51af11),
	.w8(32'hbbe763d4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809453),
	.w1(32'hba8cf447),
	.w2(32'hbc305892),
	.w3(32'hbb89f5bd),
	.w4(32'hba5bde23),
	.w5(32'hbc0284ea),
	.w6(32'h3c2eb334),
	.w7(32'h3b8f921c),
	.w8(32'h3b8c55fd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b50c7),
	.w1(32'h3900d27c),
	.w2(32'hbb35b0c4),
	.w3(32'hbb8f25d2),
	.w4(32'hb993d86a),
	.w5(32'hbad26dba),
	.w6(32'hbb63e3bb),
	.w7(32'hbab7fece),
	.w8(32'hba707747),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9810d72),
	.w1(32'h3b27d9de),
	.w2(32'h3a1dc5da),
	.w3(32'h3a1259b1),
	.w4(32'hba62450c),
	.w5(32'hbb938f31),
	.w6(32'h3aaf16a9),
	.w7(32'hb8c6bb2f),
	.w8(32'hba3a5096),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdc0b1),
	.w1(32'hb7f5e820),
	.w2(32'h3af44130),
	.w3(32'hbb11b458),
	.w4(32'h3a73a922),
	.w5(32'hbb860b7b),
	.w6(32'h3b2ac251),
	.w7(32'hbb29097a),
	.w8(32'h3abee2bb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2aea6),
	.w1(32'h3be44bbe),
	.w2(32'h3b374a72),
	.w3(32'hbb87818c),
	.w4(32'h3a3da18e),
	.w5(32'hbabd8563),
	.w6(32'h3b496480),
	.w7(32'h3a48f417),
	.w8(32'h3b7a6f27),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92a695),
	.w1(32'h3b4a3f41),
	.w2(32'h3b96f23c),
	.w3(32'h3a64a906),
	.w4(32'h3b247e1d),
	.w5(32'h3b184e87),
	.w6(32'h3c078cb8),
	.w7(32'h3a8f9ded),
	.w8(32'h3a7343ed),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80c9a8),
	.w1(32'hbc038b93),
	.w2(32'hb8230030),
	.w3(32'h3a138c5b),
	.w4(32'h3b0cda41),
	.w5(32'h39ce1887),
	.w6(32'hbadd0197),
	.w7(32'hbbdf561e),
	.w8(32'hbbadebe3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68755b),
	.w1(32'hba9b20d4),
	.w2(32'hbb108b0b),
	.w3(32'hbb070f7b),
	.w4(32'h376af388),
	.w5(32'hbb974941),
	.w6(32'hba5d15ee),
	.w7(32'hba926809),
	.w8(32'hba3bbe6c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb4653),
	.w1(32'h3b123e74),
	.w2(32'h3b3649df),
	.w3(32'hbbc3f8ba),
	.w4(32'hba83cc70),
	.w5(32'hbb0c0e31),
	.w6(32'hbabd2b59),
	.w7(32'hbb856a8a),
	.w8(32'hbb692872),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab4609),
	.w1(32'hbcb2a39a),
	.w2(32'hbc43cdc3),
	.w3(32'h3b10caeb),
	.w4(32'hbceb3e3b),
	.w5(32'hbccd340b),
	.w6(32'hbc36e336),
	.w7(32'h3b6053dc),
	.w8(32'h3c58b70e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2da470),
	.w1(32'h3b6cc4ff),
	.w2(32'h3b4c96b3),
	.w3(32'h3a8c24a2),
	.w4(32'hbbe21bff),
	.w5(32'hbc008a1f),
	.w6(32'h3bd261c9),
	.w7(32'h3bd6a5a9),
	.w8(32'h3b2b04b6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ebbb9),
	.w1(32'h3a5b99cf),
	.w2(32'hbb84fb2e),
	.w3(32'hbbebac4a),
	.w4(32'hba98890a),
	.w5(32'hbb86a20e),
	.w6(32'hbb736c68),
	.w7(32'hbc07f642),
	.w8(32'hbb23a69c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58530),
	.w1(32'h3b05d2ed),
	.w2(32'h3b00fe7d),
	.w3(32'hbc000717),
	.w4(32'hb94b17a2),
	.w5(32'h3b403b07),
	.w6(32'h3afa7bee),
	.w7(32'h3a995e42),
	.w8(32'h3b1307c2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a3392),
	.w1(32'hbcf0b56c),
	.w2(32'hbd15a346),
	.w3(32'h3ba2acbc),
	.w4(32'hbc8d4985),
	.w5(32'hbccdb6f7),
	.w6(32'hbc1cbb15),
	.w7(32'hbc19d7f1),
	.w8(32'h3c48e455),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3d80),
	.w1(32'hbb1242a5),
	.w2(32'hbb875907),
	.w3(32'h3b2209b0),
	.w4(32'hbb83286f),
	.w5(32'h39c4c562),
	.w6(32'hbb930b1c),
	.w7(32'hbb0292d5),
	.w8(32'h3af263b7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc288523),
	.w1(32'h3cb1b931),
	.w2(32'h3ceb4518),
	.w3(32'hbba0184c),
	.w4(32'h3c887d30),
	.w5(32'h3ccae408),
	.w6(32'h3c3be5f9),
	.w7(32'h3c87bd31),
	.w8(32'h3b198cb9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76dbda),
	.w1(32'hbc567d09),
	.w2(32'hb9dbe83d),
	.w3(32'h3c3ca898),
	.w4(32'hbbf4c7e5),
	.w5(32'hbb29f79e),
	.w6(32'hbc58c9a6),
	.w7(32'hbc0f6c0d),
	.w8(32'hbb1aefdc),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b030a8b),
	.w1(32'h3abc5210),
	.w2(32'h3af24425),
	.w3(32'h38d2396e),
	.w4(32'hba4b1952),
	.w5(32'hb995609b),
	.w6(32'hba81d9c8),
	.w7(32'hba8e87f3),
	.w8(32'hbb1b2eab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a3564),
	.w1(32'h3adc2a2e),
	.w2(32'h3b8432ca),
	.w3(32'hbb58f28f),
	.w4(32'hba07cbe0),
	.w5(32'hbaa35969),
	.w6(32'hba5935cd),
	.w7(32'hbbb64317),
	.w8(32'hbb304c0c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af53c8),
	.w1(32'hbd2ce5cd),
	.w2(32'hbd559b32),
	.w3(32'hbacf813a),
	.w4(32'hbd00e0b8),
	.w5(32'hbd32d2fe),
	.w6(32'hbc99691b),
	.w7(32'hbc9906b4),
	.w8(32'h3be574b2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc557aab),
	.w1(32'h3b65a794),
	.w2(32'h3af0a9eb),
	.w3(32'hbc0b0942),
	.w4(32'h3b49daa9),
	.w5(32'hba034b86),
	.w6(32'hba99f6a8),
	.w7(32'h3a969fdb),
	.w8(32'hbba2e6ef),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2d416),
	.w1(32'hbbb25a61),
	.w2(32'hbbf8e5e5),
	.w3(32'hbb0fe78c),
	.w4(32'hbbe65d24),
	.w5(32'hbba8970c),
	.w6(32'hbae36fb4),
	.w7(32'hb8fa4729),
	.w8(32'h39e0e81b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12613f),
	.w1(32'h3bd7ed4c),
	.w2(32'hbac0648b),
	.w3(32'h3b8bcd76),
	.w4(32'h3b8fb06d),
	.w5(32'h3b3dfee9),
	.w6(32'hbaea17a3),
	.w7(32'hbb933d01),
	.w8(32'h3aea2b51),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3efe24),
	.w1(32'h3b3fafaf),
	.w2(32'hba210af6),
	.w3(32'h3af71bb1),
	.w4(32'h3a918d85),
	.w5(32'hbabee5e2),
	.w6(32'hbaa99ffc),
	.w7(32'hbb49ad18),
	.w8(32'hbb8833b8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb263aef),
	.w1(32'hbb87a8ae),
	.w2(32'hba56899a),
	.w3(32'hbb329edf),
	.w4(32'hbbca1a65),
	.w5(32'hbc06e31a),
	.w6(32'hbbd2fedb),
	.w7(32'hbbfc49cd),
	.w8(32'hbbaf35a3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba816e22),
	.w1(32'h3b89202b),
	.w2(32'h3b92ed2f),
	.w3(32'h3ba15f17),
	.w4(32'h3bd31b2b),
	.w5(32'h3ba1334d),
	.w6(32'hba5e7027),
	.w7(32'h3bf78dc8),
	.w8(32'h38245686),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb52737),
	.w1(32'h3c72ddbd),
	.w2(32'h3ca95599),
	.w3(32'h3b5628a4),
	.w4(32'h3c9f67a0),
	.w5(32'h3cc2665e),
	.w6(32'h3c46ce2c),
	.w7(32'h3c54ed66),
	.w8(32'h3c1a7f8e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c3a35),
	.w1(32'hbbd81780),
	.w2(32'hbb6d2a7e),
	.w3(32'h3ca0f18d),
	.w4(32'hbc0c82d6),
	.w5(32'h3a32448b),
	.w6(32'hbc263b0f),
	.w7(32'hbaaf389d),
	.w8(32'h39295d28),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf0ecc),
	.w1(32'hbacfcf24),
	.w2(32'h3b11f68f),
	.w3(32'h3b46e18d),
	.w4(32'hbb6911fa),
	.w5(32'hbaaf4260),
	.w6(32'h39c2cc5e),
	.w7(32'h3a909f5d),
	.w8(32'hbabc6f47),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb965e86),
	.w1(32'hbb0dd93a),
	.w2(32'hba7c5be3),
	.w3(32'h3aa4e854),
	.w4(32'hb71a98c6),
	.w5(32'hbb212c8e),
	.w6(32'hbb47a26d),
	.w7(32'hbbce0ef0),
	.w8(32'h3a80d3b9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a087),
	.w1(32'hbad18929),
	.w2(32'hbae00080),
	.w3(32'h3a557428),
	.w4(32'h3aaca59d),
	.w5(32'hbaf2ea30),
	.w6(32'h3abb042a),
	.w7(32'h39dfd65d),
	.w8(32'h3a970bf0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a817591),
	.w1(32'h3bd435ac),
	.w2(32'hbb314251),
	.w3(32'hb9be6352),
	.w4(32'h3bae3124),
	.w5(32'h3af78a66),
	.w6(32'h3ae3391a),
	.w7(32'hbb6c571e),
	.w8(32'hbb7585be),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule