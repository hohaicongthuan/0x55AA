module layer_10_featuremap_225(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4805f),
	.w1(32'h3a87ce3b),
	.w2(32'hbb8f7267),
	.w3(32'h3b669add),
	.w4(32'h3ba3db2c),
	.w5(32'h3cb8d066),
	.w6(32'hbb918286),
	.w7(32'h3b83e410),
	.w8(32'h3b70ee95),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c864d1a),
	.w1(32'h3caae832),
	.w2(32'h3c397281),
	.w3(32'hbc240faf),
	.w4(32'hbc09b87e),
	.w5(32'hbb294828),
	.w6(32'h3c2eef06),
	.w7(32'h3c346d4d),
	.w8(32'hbae082dc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92b413),
	.w1(32'h3a62da92),
	.w2(32'h3c90d92f),
	.w3(32'hbc82de5f),
	.w4(32'h3dbb8c35),
	.w5(32'h3bbb4538),
	.w6(32'hbba5428e),
	.w7(32'hbbcffbdc),
	.w8(32'hbb870dac),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00fcfd),
	.w1(32'hbb345706),
	.w2(32'h3a2c1270),
	.w3(32'h3ccb7535),
	.w4(32'h3b8103ba),
	.w5(32'hbb87487c),
	.w6(32'h3b8d43f6),
	.w7(32'hbbd972f5),
	.w8(32'hbc34f3f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70faba),
	.w1(32'hbb10b972),
	.w2(32'hbb6e3c33),
	.w3(32'hbba9420e),
	.w4(32'h3cf133b4),
	.w5(32'h3a2315dc),
	.w6(32'h3b1751ff),
	.w7(32'h3b78cbec),
	.w8(32'h3bf8c424),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf21de),
	.w1(32'h3bd72099),
	.w2(32'hbb2b9666),
	.w3(32'hbc735593),
	.w4(32'hbb072c0b),
	.w5(32'h3aadb78f),
	.w6(32'hba84dd30),
	.w7(32'hbb7508fb),
	.w8(32'hbc903bc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ad0f0),
	.w1(32'hb95d83bc),
	.w2(32'hbb873416),
	.w3(32'h3b92b050),
	.w4(32'h3c177835),
	.w5(32'h3c2e07eb),
	.w6(32'h3b7bf3a2),
	.w7(32'h3b60404d),
	.w8(32'hb964eea3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ca9e3),
	.w1(32'h3b154a6f),
	.w2(32'h3ab50b1f),
	.w3(32'hbbff388c),
	.w4(32'hbb2ec2b0),
	.w5(32'hbb691e76),
	.w6(32'h397e8a2c),
	.w7(32'hbc212a2b),
	.w8(32'h3a72c850),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c707f62),
	.w1(32'hbc2e0800),
	.w2(32'h3b86f4ea),
	.w3(32'h3c6df6b4),
	.w4(32'hbb326ab6),
	.w5(32'h3a969356),
	.w6(32'h3b55113b),
	.w7(32'hbbfd2353),
	.w8(32'hb9d52f0a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8980f3),
	.w1(32'hb90b8a55),
	.w2(32'h3bec2bfc),
	.w3(32'hbc0934dd),
	.w4(32'hbb174f8a),
	.w5(32'hbc0e3dea),
	.w6(32'h3cb9d508),
	.w7(32'h3c6a4f66),
	.w8(32'hb8fe008f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35c57),
	.w1(32'h3b87f779),
	.w2(32'hbc1fc9b3),
	.w3(32'h3c503c95),
	.w4(32'hbbdb31bc),
	.w5(32'h39ba6330),
	.w6(32'h3b9e963f),
	.w7(32'hbc067672),
	.w8(32'h3b8e1b4c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6b5ab),
	.w1(32'hbc2fd524),
	.w2(32'h3b400b71),
	.w3(32'h3c4652bb),
	.w4(32'h3c8235fa),
	.w5(32'hbb0027e2),
	.w6(32'hb922732b),
	.w7(32'hb7b4b458),
	.w8(32'hbb324ca4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c014),
	.w1(32'h3b4108a3),
	.w2(32'hbc3b1423),
	.w3(32'hbbfbf38e),
	.w4(32'hbba46bab),
	.w5(32'h3b9a4da8),
	.w6(32'hbb83e3f0),
	.w7(32'h3c65991b),
	.w8(32'hbc3445ae),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf546a8),
	.w1(32'h3c5b05b2),
	.w2(32'h3a53007b),
	.w3(32'h3c1062f6),
	.w4(32'h3c97ceef),
	.w5(32'hbbba2614),
	.w6(32'hbc3a84fb),
	.w7(32'hbab2c0b7),
	.w8(32'h3bd47acd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4a55ac),
	.w1(32'hbc04ee93),
	.w2(32'hbbbef4b8),
	.w3(32'h3bb3ae5a),
	.w4(32'hb9244bbe),
	.w5(32'h3c4439af),
	.w6(32'hbcb21585),
	.w7(32'h3be8d907),
	.w8(32'hbacdb22f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1db14),
	.w1(32'hbbb2b55d),
	.w2(32'h3aa6e5b1),
	.w3(32'hbb0c4184),
	.w4(32'hbbe468e4),
	.w5(32'h3ac29351),
	.w6(32'hbc2e447e),
	.w7(32'h3c122d73),
	.w8(32'h3c1e7715),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273acf),
	.w1(32'h3b504ee4),
	.w2(32'h3c45a34d),
	.w3(32'hbbd14b4d),
	.w4(32'hb762aff9),
	.w5(32'hb9ac0cf3),
	.w6(32'h389a983a),
	.w7(32'hbc091436),
	.w8(32'h3b9020a2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd821),
	.w1(32'h3b2f677b),
	.w2(32'h3bdbbf22),
	.w3(32'hbc3c7f48),
	.w4(32'hbb937a6f),
	.w5(32'hb97d7285),
	.w6(32'h3c713bdf),
	.w7(32'h3c3b574c),
	.w8(32'h3afc4203),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbacf9),
	.w1(32'hbbbbeb50),
	.w2(32'hbbc27bbd),
	.w3(32'h3c07e92f),
	.w4(32'h39186923),
	.w5(32'h3d30400d),
	.w6(32'h3aff882a),
	.w7(32'h3c038005),
	.w8(32'h3b9fed39),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c2e2b),
	.w1(32'hbc229fee),
	.w2(32'h3c06320f),
	.w3(32'hbb37aede),
	.w4(32'h3c9225d6),
	.w5(32'hbb18b7e2),
	.w6(32'hbb62fa27),
	.w7(32'h3ba26242),
	.w8(32'h38dc9643),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c160d85),
	.w1(32'h396edc33),
	.w2(32'h3c198a89),
	.w3(32'h3c814d15),
	.w4(32'hbab4374a),
	.w5(32'hbc5631e0),
	.w6(32'hbbd7fdaf),
	.w7(32'h3bbf2098),
	.w8(32'h3a745794),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb11176),
	.w1(32'h3c0dabdc),
	.w2(32'hbb8d1b31),
	.w3(32'h3b0b8656),
	.w4(32'h3b26216f),
	.w5(32'hbb88e4cf),
	.w6(32'h3c24dc59),
	.w7(32'h38319f8c),
	.w8(32'h3c087222),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aded858),
	.w1(32'hba4beda4),
	.w2(32'h3be2ab7e),
	.w3(32'hbbd790a1),
	.w4(32'hbc163b07),
	.w5(32'h3cc3b5d0),
	.w6(32'hbb719d99),
	.w7(32'hbc269a64),
	.w8(32'h3beb6287),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a8981),
	.w1(32'hbc43d7c3),
	.w2(32'h3ad99b0d),
	.w3(32'hbc8f297d),
	.w4(32'hbba07f7f),
	.w5(32'hbc54441b),
	.w6(32'hbc92d6f3),
	.w7(32'h3d0f2557),
	.w8(32'hbc01faa9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97e6fb),
	.w1(32'h3b002bdf),
	.w2(32'hbc86bb75),
	.w3(32'hbad3dc88),
	.w4(32'hbb9f486d),
	.w5(32'h3bd78fb6),
	.w6(32'hbbdb4f24),
	.w7(32'hbc49f8d7),
	.w8(32'h3ca5ec65),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b73d4),
	.w1(32'hbc680a34),
	.w2(32'hbc69a87d),
	.w3(32'h3bd72020),
	.w4(32'hbc1e2e40),
	.w5(32'h3c0329a4),
	.w6(32'hb9f695e6),
	.w7(32'hbc41b047),
	.w8(32'hb999ede3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc107cea),
	.w1(32'h3c812937),
	.w2(32'h3bf0fe55),
	.w3(32'hb9cc5994),
	.w4(32'hba0280e4),
	.w5(32'h3b5dd865),
	.w6(32'h3c1518bc),
	.w7(32'h3b3181b3),
	.w8(32'h3c16f7bc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39abd5),
	.w1(32'h3c7f3b97),
	.w2(32'hb8829684),
	.w3(32'h3c2bf1e7),
	.w4(32'h3ba7e641),
	.w5(32'hbb91c6e9),
	.w6(32'hb8e91417),
	.w7(32'hba7b0a84),
	.w8(32'h3bd492a8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb120d98),
	.w1(32'hbbd3fa9f),
	.w2(32'h3c177433),
	.w3(32'h3c568f11),
	.w4(32'h3b579a13),
	.w5(32'hbb7232e7),
	.w6(32'hbc3d4fba),
	.w7(32'h3be48128),
	.w8(32'hbb4afb8b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002e04),
	.w1(32'hbac9cfd8),
	.w2(32'h3abb2dcc),
	.w3(32'h3c0dbd0b),
	.w4(32'hbb87739a),
	.w5(32'h3c59dfca),
	.w6(32'h3c2aa475),
	.w7(32'hbc97106a),
	.w8(32'h3c6a2e89),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10901f),
	.w1(32'h3a9ed3e4),
	.w2(32'hbc07ec49),
	.w3(32'h3bb87674),
	.w4(32'h3c3d9f7b),
	.w5(32'hbc05ca1f),
	.w6(32'hbb74863b),
	.w7(32'h3b2710fe),
	.w8(32'hbbe3c99d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1d67d),
	.w1(32'hbb835ac0),
	.w2(32'hbb488010),
	.w3(32'hbb9bff9f),
	.w4(32'hbb72026a),
	.w5(32'hbae3200c),
	.w6(32'hbbd3b8bd),
	.w7(32'h3c0d6a41),
	.w8(32'hbbfef8b8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e1817),
	.w1(32'h3c78443f),
	.w2(32'hbba68c1d),
	.w3(32'h3bc74a5b),
	.w4(32'h3c57a7b5),
	.w5(32'hbaa0dc3a),
	.w6(32'hbb7c4966),
	.w7(32'h3c10a976),
	.w8(32'hbbaed340),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa656a5),
	.w1(32'h3a30d9c1),
	.w2(32'hbb921b7b),
	.w3(32'hbb3ae599),
	.w4(32'h3c2c1d9d),
	.w5(32'h3bd3a04f),
	.w6(32'h3b35e629),
	.w7(32'hbba83dfd),
	.w8(32'h39ff61c0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bb8c0),
	.w1(32'h3bf6aa00),
	.w2(32'h3c8c853b),
	.w3(32'h3b47c249),
	.w4(32'h3bcac828),
	.w5(32'hbc7a04fc),
	.w6(32'hbb224b14),
	.w7(32'hbbdf11ea),
	.w8(32'h3b276368),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba903ed),
	.w1(32'h3beac11c),
	.w2(32'hbbc4caf4),
	.w3(32'hbafbea71),
	.w4(32'h3cb6b29e),
	.w5(32'h3c57ddd0),
	.w6(32'h3bbbe466),
	.w7(32'hbbb742df),
	.w8(32'h3ba657d3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ebc9),
	.w1(32'hbb825cfa),
	.w2(32'h3b1cc7ba),
	.w3(32'h3aa4e85f),
	.w4(32'hbb35be26),
	.w5(32'h3b37c781),
	.w6(32'h3b25e26e),
	.w7(32'h3c1f9361),
	.w8(32'h39f89963),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b9d0d),
	.w1(32'hba175183),
	.w2(32'h3c70b5bb),
	.w3(32'hbbd64bd6),
	.w4(32'hbbb6f183),
	.w5(32'h3931cd06),
	.w6(32'h3c3ee68e),
	.w7(32'hbb282694),
	.w8(32'h3c891ca9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcbf9d),
	.w1(32'h3bb991c7),
	.w2(32'hbc5c319d),
	.w3(32'hbc87b0e8),
	.w4(32'hbb541968),
	.w5(32'h3afc7192),
	.w6(32'h3be06905),
	.w7(32'h3c4cd151),
	.w8(32'h3c2f754c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce4e7b),
	.w1(32'hbb2d9fbd),
	.w2(32'h3c0abfb6),
	.w3(32'h3b066154),
	.w4(32'h3a846778),
	.w5(32'h3c1cca69),
	.w6(32'hbb79b230),
	.w7(32'hbbcb3f66),
	.w8(32'h3c0eb5ab),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3654eee0),
	.w1(32'hbce14f24),
	.w2(32'h3bd3a1b3),
	.w3(32'hbb5c8bbe),
	.w4(32'hbc4140ac),
	.w5(32'h3b0cb842),
	.w6(32'h39fbd4f4),
	.w7(32'h3b8c49bc),
	.w8(32'h3a29f7be),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae5bbb),
	.w1(32'h3b66dbf1),
	.w2(32'hbbb917f4),
	.w3(32'hbcbccfc1),
	.w4(32'h39944206),
	.w5(32'h3ae7387b),
	.w6(32'hbc44af9b),
	.w7(32'h3b597813),
	.w8(32'hbaea9e42),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2afcdf),
	.w1(32'h3ac2bc10),
	.w2(32'h3ba0d048),
	.w3(32'hbba479e5),
	.w4(32'h3bb6504e),
	.w5(32'hbc61c911),
	.w6(32'h3b0fd956),
	.w7(32'h3b3134d5),
	.w8(32'hbbb9e505),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba507f),
	.w1(32'h3b25e642),
	.w2(32'h3887bcf7),
	.w3(32'hbc1f714a),
	.w4(32'hbc3ed623),
	.w5(32'h3b0a4039),
	.w6(32'hbbb6b473),
	.w7(32'h3b27cbca),
	.w8(32'hba1e9496),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5a115),
	.w1(32'h3b8b2711),
	.w2(32'hbc1a41cd),
	.w3(32'hbbc6b2b1),
	.w4(32'hbb39ef91),
	.w5(32'h3c3f04ef),
	.w6(32'h39d77f25),
	.w7(32'hbb48ce0f),
	.w8(32'hb78083bc),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba497),
	.w1(32'h3b9303a6),
	.w2(32'hbc49c3a8),
	.w3(32'h3c31a15d),
	.w4(32'h3bb85086),
	.w5(32'h3bba9d70),
	.w6(32'hbb8392a3),
	.w7(32'hbbf37521),
	.w8(32'h3c1d1b49),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7ee7),
	.w1(32'h39a0b709),
	.w2(32'h3c91a7ef),
	.w3(32'h3aec24c1),
	.w4(32'h3ae4560a),
	.w5(32'h3bacf01f),
	.w6(32'hba1fcbaa),
	.w7(32'hbbaf1322),
	.w8(32'h3bdaef6d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50417f),
	.w1(32'hbb947899),
	.w2(32'hbb8eaa1f),
	.w3(32'hbc4ea32d),
	.w4(32'hba1b57b6),
	.w5(32'h3a22ee1b),
	.w6(32'h3bb22379),
	.w7(32'hbb359ea0),
	.w8(32'hbbffcf7a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a905d2e),
	.w1(32'h3afc35f0),
	.w2(32'h3bcab505),
	.w3(32'h3c8800a5),
	.w4(32'hbc145473),
	.w5(32'hbb73cc52),
	.w6(32'hbb5f81d6),
	.w7(32'h3b29c4c5),
	.w8(32'h3a15f07c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876ecba),
	.w1(32'h3a67a35f),
	.w2(32'h3b97305e),
	.w3(32'hbb966822),
	.w4(32'h3c0f2d8c),
	.w5(32'hbbdb8f76),
	.w6(32'hbb618144),
	.w7(32'hbb54b1a1),
	.w8(32'h39ada4ca),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d253f9),
	.w1(32'hb9754f29),
	.w2(32'hb988b94b),
	.w3(32'h3c0869d5),
	.w4(32'hbba6258d),
	.w5(32'h38d267a6),
	.w6(32'h3a98588c),
	.w7(32'h39965f5f),
	.w8(32'h3a6e44c8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6be9f),
	.w1(32'h3c8f4482),
	.w2(32'hbb21feec),
	.w3(32'hbb11c2af),
	.w4(32'h3b520fa3),
	.w5(32'h3c8e47ba),
	.w6(32'hbc3348c6),
	.w7(32'h3ac2e415),
	.w8(32'h3b19fe48),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18f1fa),
	.w1(32'h3b01f435),
	.w2(32'h3c27de0a),
	.w3(32'h3c4dccfe),
	.w4(32'h3b94dcb8),
	.w5(32'hbb3fc339),
	.w6(32'hbb1f4b34),
	.w7(32'h3c2f7758),
	.w8(32'h3c0d50ab),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ec514),
	.w1(32'h3bc61fcd),
	.w2(32'h3be13e4b),
	.w3(32'h3bd2ec61),
	.w4(32'h3b3891fa),
	.w5(32'hbc013f78),
	.w6(32'hbbe46ef4),
	.w7(32'hbb512c91),
	.w8(32'hbc8d636d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b998a),
	.w1(32'hbbaab608),
	.w2(32'h3c7fc47a),
	.w3(32'hbb95b42a),
	.w4(32'h3babe93f),
	.w5(32'h3bd1c7da),
	.w6(32'h3c45f679),
	.w7(32'hbbd88ec5),
	.w8(32'h3c3926e5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafa4a2),
	.w1(32'hbbc172f6),
	.w2(32'h3b5d165d),
	.w3(32'h3b12d937),
	.w4(32'hbba275a7),
	.w5(32'h3b5b92f8),
	.w6(32'hbb7d4712),
	.w7(32'h3b01509d),
	.w8(32'h3b04dac4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fec36),
	.w1(32'h3b88eeae),
	.w2(32'h3b22355e),
	.w3(32'h3a712cff),
	.w4(32'h3c46bee8),
	.w5(32'h3c20d075),
	.w6(32'hbac70e6f),
	.w7(32'h3a73d9ce),
	.w8(32'h3af44105),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc5526),
	.w1(32'hbaa013b6),
	.w2(32'h3cc77a52),
	.w3(32'hbbaa90e3),
	.w4(32'h3c52f1ca),
	.w5(32'h3bf7b382),
	.w6(32'hb9da6053),
	.w7(32'hbbd2b9cd),
	.w8(32'hbbcb86e8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096af7),
	.w1(32'h3c8e1558),
	.w2(32'h3b0b175f),
	.w3(32'hbc3e689b),
	.w4(32'h3ae88575),
	.w5(32'h3b47a22d),
	.w6(32'hbbb5ec4c),
	.w7(32'hbb13d6f5),
	.w8(32'hbb46a083),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eaf95),
	.w1(32'hba7baf34),
	.w2(32'h3c107950),
	.w3(32'h3b9fd5b7),
	.w4(32'hbb35ad00),
	.w5(32'h3b7e69b2),
	.w6(32'h3c2fa6c6),
	.w7(32'hbb99b02a),
	.w8(32'hbb5bdd59),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ed8ff),
	.w1(32'hb8b8dc3e),
	.w2(32'h3afa2a3b),
	.w3(32'hbbdb57f1),
	.w4(32'hbbe7baff),
	.w5(32'h3c3f4ddb),
	.w6(32'h3bc652a6),
	.w7(32'h3b10ceb8),
	.w8(32'hbadd2f34),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad82a93),
	.w1(32'hbaad7877),
	.w2(32'h3b168d4a),
	.w3(32'hbb2b3563),
	.w4(32'hbb4bf8d0),
	.w5(32'hbb0d5a09),
	.w6(32'h3b6698ff),
	.w7(32'h3b65e092),
	.w8(32'h3c4d91d7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c697cd5),
	.w1(32'hbaa88b03),
	.w2(32'h39787d1b),
	.w3(32'h3b48e861),
	.w4(32'h3b785449),
	.w5(32'hbc30dd7e),
	.w6(32'hbb7b01eb),
	.w7(32'h3b9372be),
	.w8(32'h38ad2fc7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd48c71),
	.w1(32'h3bf536ac),
	.w2(32'hb9ae0a6c),
	.w3(32'hbb669c7c),
	.w4(32'h3c0941da),
	.w5(32'h3b8cc8c2),
	.w6(32'hbcf91a41),
	.w7(32'hbc5e2e6a),
	.w8(32'hbc02af95),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b453866),
	.w1(32'h3c60620c),
	.w2(32'h3a245be9),
	.w3(32'hba7aef0e),
	.w4(32'hbbda27e4),
	.w5(32'h3be4dc07),
	.w6(32'h3c4ed6ac),
	.w7(32'hbc0a0c19),
	.w8(32'hbc291024),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc479a),
	.w1(32'hbc7d5dd2),
	.w2(32'h3a46d2a4),
	.w3(32'hbbb27a75),
	.w4(32'h3b105cd0),
	.w5(32'hbb0e0c16),
	.w6(32'h3c365c52),
	.w7(32'h3b3a3d2b),
	.w8(32'h393376cf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5aa1ea),
	.w1(32'h3c1f30cc),
	.w2(32'hbb7b98b1),
	.w3(32'h3c96c3b7),
	.w4(32'hbb4d5758),
	.w5(32'h3b914d14),
	.w6(32'hb8a57de1),
	.w7(32'hbc8286da),
	.w8(32'h3bada2d5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6ab96),
	.w1(32'h3a2b6c41),
	.w2(32'hbb56315d),
	.w3(32'h3b6b4dbf),
	.w4(32'h3aa2cb72),
	.w5(32'hbb8bc39d),
	.w6(32'hbaf88398),
	.w7(32'h3b4c577b),
	.w8(32'h3b9cfdf5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d23b7),
	.w1(32'h3bca4fbb),
	.w2(32'hbb0d346e),
	.w3(32'h3acb24e8),
	.w4(32'h37a81218),
	.w5(32'h3c12afee),
	.w6(32'hbc57bcfb),
	.w7(32'hbb8e7405),
	.w8(32'hbc311048),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f9c02),
	.w1(32'hba185ccf),
	.w2(32'h39855965),
	.w3(32'hbb2c00d7),
	.w4(32'hbb50f097),
	.w5(32'h3b9f9908),
	.w6(32'hbb86659f),
	.w7(32'hbb4f03ba),
	.w8(32'hbac09d7c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f304e1),
	.w1(32'hb9629935),
	.w2(32'h3ba6e2bc),
	.w3(32'hbc3e0404),
	.w4(32'h37d5cb1c),
	.w5(32'h3bc4349d),
	.w6(32'h3c1112ed),
	.w7(32'hbb46ff49),
	.w8(32'h3ba3bb4c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc531eea),
	.w1(32'h3b5667ce),
	.w2(32'h3c534b02),
	.w3(32'hbaa7f68c),
	.w4(32'h3c4fbd02),
	.w5(32'h3ba1ffcc),
	.w6(32'hbc533b27),
	.w7(32'hbad7ac83),
	.w8(32'h3a89f7c4),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c22448),
	.w1(32'h3aaff992),
	.w2(32'h3a156e83),
	.w3(32'hbb22df5b),
	.w4(32'h3be72fe6),
	.w5(32'hbc1de885),
	.w6(32'h3aa0ffc0),
	.w7(32'hbb5606a3),
	.w8(32'hbb4b4df8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba956e12),
	.w1(32'h36c2f85a),
	.w2(32'hbbfabdb6),
	.w3(32'h3bc3bcbd),
	.w4(32'h3aaf636e),
	.w5(32'hbbbef22e),
	.w6(32'h3badfb8e),
	.w7(32'h3b9906c9),
	.w8(32'hbb47d5bf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f042b),
	.w1(32'h3add1c15),
	.w2(32'h381e8bc3),
	.w3(32'h3b84761f),
	.w4(32'hbb472332),
	.w5(32'h3ac2e660),
	.w6(32'hbbda2840),
	.w7(32'hbbd9c5c3),
	.w8(32'hbb5ffdb6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef6c2),
	.w1(32'hbc1df769),
	.w2(32'h3b63052e),
	.w3(32'h3b104de6),
	.w4(32'h3c5dafac),
	.w5(32'h3c5d07f1),
	.w6(32'hbb0f459b),
	.w7(32'h39a3c1ab),
	.w8(32'hbb840ad6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78861c),
	.w1(32'h3b94e3c8),
	.w2(32'hbb2b4602),
	.w3(32'h3b767fb2),
	.w4(32'hbad0c163),
	.w5(32'hb7a34135),
	.w6(32'h3b8c7b7f),
	.w7(32'h3b509397),
	.w8(32'h3ab8e737),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b1fd1),
	.w1(32'hbb9e7a65),
	.w2(32'hbc5e4b28),
	.w3(32'h38a4c74a),
	.w4(32'h3be33fda),
	.w5(32'hba8ae4a3),
	.w6(32'h3ba847e5),
	.w7(32'hbc423897),
	.w8(32'h3bc929e2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cfaeed),
	.w1(32'h3b12ea2a),
	.w2(32'h3a66c251),
	.w3(32'hbbca566b),
	.w4(32'hb8f0bed7),
	.w5(32'hbbbdfc7a),
	.w6(32'h3b54331c),
	.w7(32'h3b4a7d96),
	.w8(32'hb9fae68d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f0574),
	.w1(32'hb90dbbce),
	.w2(32'hbc8899d1),
	.w3(32'hbb1b99bc),
	.w4(32'hbb1d8288),
	.w5(32'h3c187982),
	.w6(32'h39834468),
	.w7(32'hbc0af246),
	.w8(32'hba7760e8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b877ebb),
	.w1(32'hbbe37e83),
	.w2(32'hbb338ddb),
	.w3(32'hbb9e9b2a),
	.w4(32'h3b8298b2),
	.w5(32'h3b59a58a),
	.w6(32'h3cccdc1e),
	.w7(32'hbb98675f),
	.w8(32'hbb73dd13),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75bd2f),
	.w1(32'h3bb043b7),
	.w2(32'hba8a3189),
	.w3(32'hbc28d76d),
	.w4(32'h3af989c6),
	.w5(32'h3c86ab49),
	.w6(32'hb84df301),
	.w7(32'hbb1a89b0),
	.w8(32'h3b310d92),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb999e6c),
	.w1(32'hbb6f827d),
	.w2(32'h3acfbff7),
	.w3(32'hbb090083),
	.w4(32'hbb273507),
	.w5(32'h3c20d94a),
	.w6(32'h3cafb91c),
	.w7(32'hbad9d998),
	.w8(32'h3c6e3300),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14502a),
	.w1(32'hbba87b69),
	.w2(32'hba2b040e),
	.w3(32'h3cb74b09),
	.w4(32'h3b29cf38),
	.w5(32'hbc3bf5ba),
	.w6(32'hbbdcbbb8),
	.w7(32'hbc5b8570),
	.w8(32'h3c40f854),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcdcbd),
	.w1(32'h399015d6),
	.w2(32'hbbb88257),
	.w3(32'hbcb409df),
	.w4(32'h3bea865b),
	.w5(32'hbc0455de),
	.w6(32'h3c955ec4),
	.w7(32'h3c9259d3),
	.w8(32'hbccf67c0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34f381),
	.w1(32'h3b0eb7c5),
	.w2(32'h3ac2bdba),
	.w3(32'hbc1eff6e),
	.w4(32'h3c8201bf),
	.w5(32'h3c859bf1),
	.w6(32'h3d0939a5),
	.w7(32'h3ba99e64),
	.w8(32'hbccb138b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccef933),
	.w1(32'h3b63c059),
	.w2(32'hbce3dc5b),
	.w3(32'h3caf7ccc),
	.w4(32'h3bb7c891),
	.w5(32'h3cc0dbab),
	.w6(32'h399e5d71),
	.w7(32'h3be13a8e),
	.w8(32'h3b877d90),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9b01),
	.w1(32'hbce64fbd),
	.w2(32'hbc87867a),
	.w3(32'hbc48f159),
	.w4(32'h3c1b5f7c),
	.w5(32'h3c8e03b2),
	.w6(32'hbb65eea4),
	.w7(32'h3bd433cf),
	.w8(32'hbcbad5da),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e9c6a),
	.w1(32'hbc451336),
	.w2(32'h3b971572),
	.w3(32'h3a8f4195),
	.w4(32'h392ffad8),
	.w5(32'hbc5025f0),
	.w6(32'hbc1dae57),
	.w7(32'hbc18d71a),
	.w8(32'h3c8c59b3),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bef2a),
	.w1(32'hbd2c15a6),
	.w2(32'hbc07aee5),
	.w3(32'h3c515835),
	.w4(32'h3b23305e),
	.w5(32'hba9a2b85),
	.w6(32'h3c15adf0),
	.w7(32'h3c3c4f82),
	.w8(32'hbb0ecba3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ab747),
	.w1(32'h3bb24e9b),
	.w2(32'h3c6d7f18),
	.w3(32'h3bbc840b),
	.w4(32'hbc76a7bb),
	.w5(32'h3b33a8b4),
	.w6(32'hbb540bae),
	.w7(32'h3b3b9065),
	.w8(32'h3b0f72a0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c4971),
	.w1(32'hbb148a44),
	.w2(32'hbcbe8dec),
	.w3(32'h3c145cb5),
	.w4(32'h3be424fc),
	.w5(32'h3b0b41b3),
	.w6(32'h3a864b35),
	.w7(32'hbc01bb60),
	.w8(32'h3c08513c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6aee),
	.w1(32'h3c05beb3),
	.w2(32'h3c509920),
	.w3(32'h3b333444),
	.w4(32'hbb0e6622),
	.w5(32'h3c106a28),
	.w6(32'h3c23dd74),
	.w7(32'hbd001831),
	.w8(32'hbc07ab8b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0542a5),
	.w1(32'h3ba9279e),
	.w2(32'h3c299fb0),
	.w3(32'hbb297ccf),
	.w4(32'hbc2c1636),
	.w5(32'hbc29924e),
	.w6(32'hbc323ade),
	.w7(32'hba5f62ff),
	.w8(32'h3a1d9316),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c188600),
	.w1(32'h3be3263b),
	.w2(32'h38a4f974),
	.w3(32'hbc17323d),
	.w4(32'h3c363319),
	.w5(32'h3c835ddd),
	.w6(32'h3ae608ce),
	.w7(32'h3b1d4577),
	.w8(32'hb9a2663a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75ad46),
	.w1(32'hbcabcb16),
	.w2(32'hbc1a7ac2),
	.w3(32'hbc452cd2),
	.w4(32'h3c13253c),
	.w5(32'hbb0630cc),
	.w6(32'hbbd371a8),
	.w7(32'h3c3562cf),
	.w8(32'h3b182734),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc882d6),
	.w1(32'h3c19bd60),
	.w2(32'h3b3fd00e),
	.w3(32'h3bc6c813),
	.w4(32'h3cde9f50),
	.w5(32'h3bdbfc86),
	.w6(32'hbc138337),
	.w7(32'h3b82c134),
	.w8(32'hb81d59c8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7fe06),
	.w1(32'hbbe05b9f),
	.w2(32'hbc39442a),
	.w3(32'h3ad52a8f),
	.w4(32'hbb750310),
	.w5(32'hbb65c67c),
	.w6(32'hbc4262c3),
	.w7(32'h3c1e9e88),
	.w8(32'hbcaacf14),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1324a8),
	.w1(32'h3b643da5),
	.w2(32'h3ac326b3),
	.w3(32'h3b1fe095),
	.w4(32'hbbaf36dc),
	.w5(32'hbaef8bd0),
	.w6(32'hb98e9509),
	.w7(32'h3b762f0b),
	.w8(32'h3a9aa240),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f363f),
	.w1(32'h3b9d7215),
	.w2(32'h3a773505),
	.w3(32'h3c6c0d80),
	.w4(32'h3c3b527a),
	.w5(32'hbb13e1fc),
	.w6(32'hbb858e2b),
	.w7(32'h3c92dd76),
	.w8(32'h3a5a6fd4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb813cc2),
	.w1(32'hbc3fcb0f),
	.w2(32'hbc27c7c2),
	.w3(32'h3a5eccf1),
	.w4(32'h3baf4907),
	.w5(32'hba812b8f),
	.w6(32'hba8b1d48),
	.w7(32'hbc577666),
	.w8(32'hbd04c480),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2931ce),
	.w1(32'h3afd585f),
	.w2(32'h39bdd870),
	.w3(32'h3b0552d7),
	.w4(32'h3b874216),
	.w5(32'hb8d7dcbc),
	.w6(32'h3b07f591),
	.w7(32'hbc74f8da),
	.w8(32'hbbd6c52e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83e95b),
	.w1(32'hbacc77d0),
	.w2(32'h3bd71c85),
	.w3(32'hbae878e5),
	.w4(32'hbc426a6f),
	.w5(32'hbaa5e341),
	.w6(32'hbc17ad21),
	.w7(32'h3baa55b9),
	.w8(32'hbbbb2650),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7028b),
	.w1(32'h3bd64ab1),
	.w2(32'h3c0f14d2),
	.w3(32'h3a100375),
	.w4(32'hbc1184b2),
	.w5(32'hbc03a444),
	.w6(32'hbad20a59),
	.w7(32'hba10ce69),
	.w8(32'hbc3bc9fa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b8775),
	.w1(32'h3a37e2e1),
	.w2(32'hbc1b54db),
	.w3(32'h3b1b9575),
	.w4(32'hbca1b83c),
	.w5(32'hbc51bd14),
	.w6(32'hbc43381e),
	.w7(32'hbc059be2),
	.w8(32'h3c08386f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aded429),
	.w1(32'h39caaf15),
	.w2(32'hbcadc2ab),
	.w3(32'h3c403f46),
	.w4(32'hbcc0ef45),
	.w5(32'h3b908024),
	.w6(32'h3b7ec9f3),
	.w7(32'h3b73645a),
	.w8(32'hbcabd52b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5a1a1),
	.w1(32'h3c64a322),
	.w2(32'h3b542387),
	.w3(32'hbc09bdd6),
	.w4(32'hba8f4898),
	.w5(32'h3ada6cdc),
	.w6(32'h3b3bd15f),
	.w7(32'h3c1be48f),
	.w8(32'h385d1237),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc225891),
	.w1(32'hbb5b8502),
	.w2(32'h366746ca),
	.w3(32'hbb7cc970),
	.w4(32'hbc80e538),
	.w5(32'hbbf7b097),
	.w6(32'h3aab3732),
	.w7(32'h3b9378ed),
	.w8(32'hbc3f4c01),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc28fca),
	.w1(32'hbb987613),
	.w2(32'h3c369c8f),
	.w3(32'hbb678f67),
	.w4(32'hbc105b2a),
	.w5(32'h3c1199a0),
	.w6(32'h3c5319b5),
	.w7(32'h3bcd0a54),
	.w8(32'h3c4eef89),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16a8a6),
	.w1(32'h3b3ad793),
	.w2(32'h3c3833e3),
	.w3(32'hb7950b9c),
	.w4(32'hbbb0ebee),
	.w5(32'h390e6b94),
	.w6(32'hbc62933f),
	.w7(32'h3c2fa188),
	.w8(32'h389cd9f5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a8b13),
	.w1(32'hbc19d336),
	.w2(32'h3cd97077),
	.w3(32'hbc298baf),
	.w4(32'h3af7c842),
	.w5(32'h3d2e197e),
	.w6(32'h3b9985b4),
	.w7(32'h3aef4e24),
	.w8(32'hbb0269a2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e1629),
	.w1(32'hbc85c60e),
	.w2(32'h3bc8b470),
	.w3(32'h39961bc8),
	.w4(32'hbca11eeb),
	.w5(32'hbc6d4720),
	.w6(32'hbc8b31c8),
	.w7(32'h3bf60d6a),
	.w8(32'h3c8c7e3e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805bd4),
	.w1(32'hbaa709bb),
	.w2(32'h3b885be6),
	.w3(32'hbb28abd0),
	.w4(32'h3b0895f2),
	.w5(32'h3c3efef8),
	.w6(32'hbb43d6f2),
	.w7(32'hbc139556),
	.w8(32'h3c27476b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aafb7),
	.w1(32'hbc17292e),
	.w2(32'h3c07892e),
	.w3(32'hbba19bc6),
	.w4(32'h3ac8be4f),
	.w5(32'h37f7527e),
	.w6(32'h3b9db4cc),
	.w7(32'hbc4a20cd),
	.w8(32'h3ab1ecd4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e96df),
	.w1(32'h3978b806),
	.w2(32'hbbc0f20d),
	.w3(32'h3ac09c2b),
	.w4(32'h3b6fa0e6),
	.w5(32'hbb7c08b0),
	.w6(32'hba13f05a),
	.w7(32'hb9ebd6ee),
	.w8(32'hbbdad71d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c01b8),
	.w1(32'hbb86d43e),
	.w2(32'h39b7ecb2),
	.w3(32'hba6245f5),
	.w4(32'h3a9f8b0f),
	.w5(32'h3b6568fe),
	.w6(32'h3c8c9d9e),
	.w7(32'hbb1addd3),
	.w8(32'h3a678055),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27119c),
	.w1(32'hbc66193d),
	.w2(32'hbbc696b9),
	.w3(32'hbc2cd525),
	.w4(32'hbb00803e),
	.w5(32'hbbff58e7),
	.w6(32'h3cc1e774),
	.w7(32'h3b5acd43),
	.w8(32'hbbd2e60c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1722aa),
	.w1(32'hbb26246e),
	.w2(32'h3c0f793e),
	.w3(32'h3b431529),
	.w4(32'h3b877271),
	.w5(32'h3b1732da),
	.w6(32'hbab5d665),
	.w7(32'hbc08184d),
	.w8(32'h3a73c007),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e2574),
	.w1(32'hbc4e0929),
	.w2(32'hbb9ddf8c),
	.w3(32'hbb83debd),
	.w4(32'hba80f8b0),
	.w5(32'hbc26849b),
	.w6(32'hbbc9cb86),
	.w7(32'h3b033908),
	.w8(32'hbc6a096a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebfa5f),
	.w1(32'h3b861d75),
	.w2(32'h3ab1092a),
	.w3(32'h3b43fbea),
	.w4(32'hbbc6c5c3),
	.w5(32'h3a106f8e),
	.w6(32'h3af76f91),
	.w7(32'h3ced30d8),
	.w8(32'hbc172598),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c367cb8),
	.w1(32'h39a57522),
	.w2(32'h3c18c2b6),
	.w3(32'hbd21324f),
	.w4(32'hbc862146),
	.w5(32'h3c412973),
	.w6(32'h3aa4d099),
	.w7(32'h3c08dda2),
	.w8(32'hbb0bd038),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4226f8),
	.w1(32'hbc395421),
	.w2(32'h3a1a628d),
	.w3(32'h3bc9eef6),
	.w4(32'hb9b7ad6f),
	.w5(32'h3be054b3),
	.w6(32'h3bbbda78),
	.w7(32'hbb5845d5),
	.w8(32'hbbb74f4b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b992),
	.w1(32'hbb0bec70),
	.w2(32'hba334984),
	.w3(32'hbb8e83a1),
	.w4(32'hbb9124f1),
	.w5(32'hbb247ccb),
	.w6(32'hbc940efc),
	.w7(32'h3a65745d),
	.w8(32'hba8486ac),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5be439),
	.w1(32'h3b470ca4),
	.w2(32'hbb993d40),
	.w3(32'h392455ce),
	.w4(32'hbc553c61),
	.w5(32'hbbc97087),
	.w6(32'h3b5cabce),
	.w7(32'hbc2ad86f),
	.w8(32'h3c078164),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7ed86),
	.w1(32'hbc022223),
	.w2(32'hbc0d2304),
	.w3(32'hbb0ac7d3),
	.w4(32'hbbbf9c8d),
	.w5(32'h3b9a6c6c),
	.w6(32'h3ab39beb),
	.w7(32'hbb88b8a3),
	.w8(32'hba27db80),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce181),
	.w1(32'h3521cb89),
	.w2(32'h3c3afcbb),
	.w3(32'hbb502274),
	.w4(32'h3b04791e),
	.w5(32'hbc834bfc),
	.w6(32'h3b9d74c3),
	.w7(32'hbabe4a0c),
	.w8(32'h3acf8b88),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc127393),
	.w1(32'hb99da7c0),
	.w2(32'hbb229cbd),
	.w3(32'hbc0d6725),
	.w4(32'hbc8b294a),
	.w5(32'h3acafd80),
	.w6(32'hbb67c95e),
	.w7(32'h3c91088e),
	.w8(32'hbc29cda6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4202ab),
	.w1(32'h3b345079),
	.w2(32'h39d37a0e),
	.w3(32'hbb8124f0),
	.w4(32'hba64c32a),
	.w5(32'hbb67bd9a),
	.w6(32'h3bfc1a08),
	.w7(32'h3bdfb222),
	.w8(32'hbae8fead),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5130a0),
	.w1(32'h3be40c2b),
	.w2(32'hba1c81e5),
	.w3(32'hbcb18f1d),
	.w4(32'hbc27fbce),
	.w5(32'hbc673c91),
	.w6(32'hbc31c539),
	.w7(32'h3c1185a8),
	.w8(32'h3a5bc248),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2955f8),
	.w1(32'hbb9e7369),
	.w2(32'h3b88aaac),
	.w3(32'hbba1460a),
	.w4(32'hbbdeef3f),
	.w5(32'hbbe347ec),
	.w6(32'h38abd316),
	.w7(32'hbb28433b),
	.w8(32'hbb5816a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d31a4),
	.w1(32'hbb2100fd),
	.w2(32'hbbe447a8),
	.w3(32'h3c0a1810),
	.w4(32'hbc0b508c),
	.w5(32'h3c21fa57),
	.w6(32'hb6c70c72),
	.w7(32'hbbc48552),
	.w8(32'hbc1e0260),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658f58),
	.w1(32'h3bc9dae8),
	.w2(32'hbba73099),
	.w3(32'h3b67f4b8),
	.w4(32'h3b8879f5),
	.w5(32'hba6a7526),
	.w6(32'h3bab9b7a),
	.w7(32'hb987d15d),
	.w8(32'hbc7a8507),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdee30),
	.w1(32'h3c7f0714),
	.w2(32'hbc121039),
	.w3(32'h3beb4044),
	.w4(32'hbc0011b0),
	.w5(32'h3b136e5e),
	.w6(32'hbc07b1a0),
	.w7(32'hbc35e957),
	.w8(32'hbc0f5eb6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63502d),
	.w1(32'hba969151),
	.w2(32'hbba60132),
	.w3(32'hbc5db541),
	.w4(32'h3b102540),
	.w5(32'h3be42d6f),
	.w6(32'hbb79d4f3),
	.w7(32'hbab7da7e),
	.w8(32'hbb86f5ec),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51a191),
	.w1(32'hbc110ce9),
	.w2(32'h3a573fbb),
	.w3(32'hbb8d834f),
	.w4(32'hbacd7f98),
	.w5(32'h3c8075d0),
	.w6(32'h3adfe788),
	.w7(32'hbb50a0d1),
	.w8(32'hbb4a991f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952ce86),
	.w1(32'hb9ae9cac),
	.w2(32'hba8eaa6b),
	.w3(32'h3b88c42d),
	.w4(32'h3ab5c445),
	.w5(32'hbc318033),
	.w6(32'h3a0bd13e),
	.w7(32'hb96f699a),
	.w8(32'hbb5ec7f6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa47d32),
	.w1(32'hbc297574),
	.w2(32'hbb876081),
	.w3(32'h39fe4d92),
	.w4(32'hbc182817),
	.w5(32'h3b7829d2),
	.w6(32'hbb243450),
	.w7(32'hbbfa7482),
	.w8(32'hba5b7f6c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8fb1e),
	.w1(32'h3a4d1a21),
	.w2(32'hbb03341a),
	.w3(32'h3c3b1a37),
	.w4(32'h3b503a7c),
	.w5(32'hba377752),
	.w6(32'hbabd24a7),
	.w7(32'h3b07a347),
	.w8(32'h3c3a8b9f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ccc67),
	.w1(32'hbae9d759),
	.w2(32'h3c4347ce),
	.w3(32'hbba322d2),
	.w4(32'h3b5e4293),
	.w5(32'h3a8ec7d7),
	.w6(32'h3b951c26),
	.w7(32'hba458ab7),
	.w8(32'h393c4ae8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372fd8c6),
	.w1(32'hbabb577e),
	.w2(32'hbbc2b493),
	.w3(32'h3c5c9da6),
	.w4(32'hbc71e407),
	.w5(32'h3cf0fa14),
	.w6(32'h3c617d43),
	.w7(32'hbaff0d10),
	.w8(32'hbb6282a3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4377dc),
	.w1(32'hbbeb4a93),
	.w2(32'h3c20332d),
	.w3(32'h3a67729e),
	.w4(32'h3b962b73),
	.w5(32'h3b7e963e),
	.w6(32'hbb9d1dd5),
	.w7(32'h3b8006d2),
	.w8(32'h3bbe24bb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae03491),
	.w1(32'hbb543013),
	.w2(32'h3c0cde57),
	.w3(32'h3c4d0313),
	.w4(32'h3bedbedc),
	.w5(32'hbbb36cb1),
	.w6(32'h3b639c5e),
	.w7(32'hbbe4370b),
	.w8(32'h3c98db54),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2c21),
	.w1(32'h3b59de09),
	.w2(32'h3b330a87),
	.w3(32'hbc363a0a),
	.w4(32'h3be812ff),
	.w5(32'h3c34deec),
	.w6(32'h3bb4de8f),
	.w7(32'hb8d94951),
	.w8(32'h3c1db98b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f2458),
	.w1(32'hbc8433cd),
	.w2(32'h3bdae427),
	.w3(32'hba912e42),
	.w4(32'hba680b81),
	.w5(32'h39ae10e0),
	.w6(32'h3aba34c9),
	.w7(32'h3ca2cd97),
	.w8(32'h3bed9d85),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98832ac),
	.w1(32'h3be1ab34),
	.w2(32'hbc278a04),
	.w3(32'hbafd2bf7),
	.w4(32'hbc32a791),
	.w5(32'hbb1963f7),
	.w6(32'h3c514add),
	.w7(32'hbbca9e6c),
	.w8(32'hbbc2044c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeb77a),
	.w1(32'hba9378a4),
	.w2(32'hbac870b5),
	.w3(32'hbb41ca43),
	.w4(32'hbb01e63d),
	.w5(32'hba241cc0),
	.w6(32'hbbaf0503),
	.w7(32'hbb8b573b),
	.w8(32'h3b4d813a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedc3b0),
	.w1(32'h3c08c444),
	.w2(32'hbbf91122),
	.w3(32'hbc01f20c),
	.w4(32'h3b5cd4c9),
	.w5(32'hbaa7327f),
	.w6(32'h3cb582bb),
	.w7(32'hba5bc508),
	.w8(32'hbb24b68a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65868c),
	.w1(32'hbbab547b),
	.w2(32'h3a3c3270),
	.w3(32'hbb825784),
	.w4(32'hbb86f1f6),
	.w5(32'hbba8959e),
	.w6(32'h3c3a7247),
	.w7(32'h3c61fc12),
	.w8(32'hba872b83),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eec9a),
	.w1(32'hbbb3ef78),
	.w2(32'h3a82b8d1),
	.w3(32'h3bbea66b),
	.w4(32'h3c50c033),
	.w5(32'hbb72470d),
	.w6(32'h3b8f0bda),
	.w7(32'hbc35f2e4),
	.w8(32'h3a5eceb3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c125a95),
	.w1(32'hbba10bc3),
	.w2(32'h3b7671cc),
	.w3(32'h39cdbd65),
	.w4(32'hbb460d56),
	.w5(32'h3a8c3e79),
	.w6(32'h3ce8d34d),
	.w7(32'h3c6fd889),
	.w8(32'h3b04bace),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073995),
	.w1(32'h3c371ecb),
	.w2(32'h3a2be496),
	.w3(32'hbbe3b00b),
	.w4(32'h3c1bc053),
	.w5(32'hb9316f91),
	.w6(32'hba39ec4d),
	.w7(32'hb90760f4),
	.w8(32'hbbc37f29),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30bbed),
	.w1(32'h3af56e80),
	.w2(32'h3c832f0b),
	.w3(32'hb9e31618),
	.w4(32'h3c9de777),
	.w5(32'hba4c73f4),
	.w6(32'hbbc87568),
	.w7(32'hb9601b2a),
	.w8(32'hbc005aa3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1368b6),
	.w1(32'h3bce8039),
	.w2(32'h3b83cfaa),
	.w3(32'h39680c21),
	.w4(32'hbc4adfb3),
	.w5(32'hbabd14e3),
	.w6(32'h3c1d5ac7),
	.w7(32'h3b127415),
	.w8(32'h3b19d8de),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c8938),
	.w1(32'hba838ffe),
	.w2(32'hba896f20),
	.w3(32'hbaa0627e),
	.w4(32'h3bcc27dd),
	.w5(32'hb708afdb),
	.w6(32'hb8a4cb32),
	.w7(32'h3bda67c7),
	.w8(32'hbab72079),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2295b),
	.w1(32'h3b20472b),
	.w2(32'hbac2db24),
	.w3(32'hbcbb2beb),
	.w4(32'h3c839e9c),
	.w5(32'h3b7f73c2),
	.w6(32'hbb302622),
	.w7(32'h3bd42e2b),
	.w8(32'hbc830ca4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb16f41),
	.w1(32'h3bc36c9c),
	.w2(32'hbb41216b),
	.w3(32'hbb4f1e31),
	.w4(32'hbbb3b320),
	.w5(32'h3be890e7),
	.w6(32'h3af22a1a),
	.w7(32'h3b999972),
	.w8(32'hbbdc74b8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab249cc),
	.w1(32'h3b60d92d),
	.w2(32'hbbf53e4d),
	.w3(32'hb9ce88ad),
	.w4(32'hbb556e50),
	.w5(32'hba9a50b3),
	.w6(32'h3b04bf81),
	.w7(32'hbc238231),
	.w8(32'hbc1b22eb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e4f3),
	.w1(32'h3bf2a784),
	.w2(32'hbb14d4a3),
	.w3(32'h3b181c4d),
	.w4(32'h3b192967),
	.w5(32'h3bfa675a),
	.w6(32'hbc01acfa),
	.w7(32'hb8719e71),
	.w8(32'hbbd8f931),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376479),
	.w1(32'hb846d01d),
	.w2(32'hb6658ee2),
	.w3(32'hbb871482),
	.w4(32'hbc1a1967),
	.w5(32'h3b1ac942),
	.w6(32'h398cc428),
	.w7(32'h3c1bed41),
	.w8(32'h3b90124b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13652c),
	.w1(32'hbbcf50dc),
	.w2(32'h3ba04b07),
	.w3(32'h3bfbdbe4),
	.w4(32'hbc01c6c4),
	.w5(32'h39b899ab),
	.w6(32'h3b707775),
	.w7(32'h3c0d6949),
	.w8(32'hbb200e9b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba509c7e),
	.w1(32'hba95c329),
	.w2(32'h3c0d4c90),
	.w3(32'h3b431cef),
	.w4(32'h3c88ddd9),
	.w5(32'h3c6c28cf),
	.w6(32'h3bf6ac22),
	.w7(32'h3b8135d0),
	.w8(32'hbc1d38bf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21def5),
	.w1(32'hbb7afcd3),
	.w2(32'hbc2160a5),
	.w3(32'hbb3d3584),
	.w4(32'hbbd2529c),
	.w5(32'h38650ccb),
	.w6(32'hba0975c7),
	.w7(32'h3986b10b),
	.w8(32'h3cdbf70c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c3788),
	.w1(32'h3bf17cb2),
	.w2(32'hbb689206),
	.w3(32'hbacb22fe),
	.w4(32'h3b987c2c),
	.w5(32'h3b20401b),
	.w6(32'hbc3eb092),
	.w7(32'hbb8ff76a),
	.w8(32'h3c0a617e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c2e1),
	.w1(32'hbb895a50),
	.w2(32'hbb3f0adb),
	.w3(32'h3bb02c62),
	.w4(32'h3bd09724),
	.w5(32'h384f8591),
	.w6(32'h3b1b57f1),
	.w7(32'hbbd12144),
	.w8(32'h3bba588d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86c26b),
	.w1(32'h3b8514f2),
	.w2(32'h3b338d13),
	.w3(32'hbb345c5d),
	.w4(32'h3ab8539e),
	.w5(32'hbbd16dc1),
	.w6(32'hbb811383),
	.w7(32'hb9896925),
	.w8(32'hba728474),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1616f5),
	.w1(32'hbab2532a),
	.w2(32'h3a94a7c1),
	.w3(32'h3c68fe65),
	.w4(32'h39ad80cf),
	.w5(32'h3c42d918),
	.w6(32'h3ba352bf),
	.w7(32'h3bde747e),
	.w8(32'h3cb4b3a1),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db33d),
	.w1(32'h3bdd67d9),
	.w2(32'h3b190e56),
	.w3(32'hbb736ced),
	.w4(32'h3c12f591),
	.w5(32'h3b97be7d),
	.w6(32'h38e705f3),
	.w7(32'hbbdead60),
	.w8(32'h3c16eb98),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31f64c),
	.w1(32'h3b8ee1b8),
	.w2(32'hbcc2ae1a),
	.w3(32'h3ba5b717),
	.w4(32'h3bbf0d9f),
	.w5(32'h3c993415),
	.w6(32'hbc135323),
	.w7(32'hbcdd6ac6),
	.w8(32'h3b207eb0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac002c),
	.w1(32'hbbb01265),
	.w2(32'h3c3e4e26),
	.w3(32'hbb4f6dd1),
	.w4(32'h3c918445),
	.w5(32'hba2d5294),
	.w6(32'hbc8f78af),
	.w7(32'h3bdb434a),
	.w8(32'h3c210308),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f0efb),
	.w1(32'h3bbb6788),
	.w2(32'hbbf35be5),
	.w3(32'h3c805257),
	.w4(32'h3b84abb4),
	.w5(32'h3b27d5ef),
	.w6(32'hba5d24ff),
	.w7(32'h3c9d256f),
	.w8(32'hb9c64bf0),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6459c0),
	.w1(32'h392d4687),
	.w2(32'hb9d7735a),
	.w3(32'h3ba8bb23),
	.w4(32'h3b8a4453),
	.w5(32'h3bfd5711),
	.w6(32'h3b0ddea4),
	.w7(32'h3c2e7580),
	.w8(32'h3b938b26),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1d5e5),
	.w1(32'h3b7a300e),
	.w2(32'h3c1b393d),
	.w3(32'h3a91faab),
	.w4(32'h3c517eff),
	.w5(32'hbc3add52),
	.w6(32'h3c264b4c),
	.w7(32'h39d6b566),
	.w8(32'hbb1c2997),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c086e24),
	.w1(32'h3b96511d),
	.w2(32'h3c033127),
	.w3(32'h3a5778b2),
	.w4(32'h3adf1ba2),
	.w5(32'hbb92ec9e),
	.w6(32'h3c04d6bb),
	.w7(32'h3b040ef9),
	.w8(32'h3bd74115),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92cbb2),
	.w1(32'hbc1a522a),
	.w2(32'hbb9a5dd2),
	.w3(32'hbc1f9893),
	.w4(32'hbba775af),
	.w5(32'h3c508a5c),
	.w6(32'hbba5641e),
	.w7(32'h38c21ad0),
	.w8(32'hbba4064a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ec11c),
	.w1(32'h3b8290a2),
	.w2(32'h3c0bf3d2),
	.w3(32'h3b62682d),
	.w4(32'hbbdda86b),
	.w5(32'h3c81555a),
	.w6(32'hbbbef491),
	.w7(32'hb901d7ae),
	.w8(32'hbbee68ef),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5166),
	.w1(32'hbba3d509),
	.w2(32'h3c59e018),
	.w3(32'hbb25fd3d),
	.w4(32'hba50a04c),
	.w5(32'h3972ea3a),
	.w6(32'hbbc52060),
	.w7(32'h3bf02dea),
	.w8(32'hbb0b5318),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c250418),
	.w1(32'h3b7ecf35),
	.w2(32'h3b8f473b),
	.w3(32'hb90b6a8b),
	.w4(32'h3a0a9a28),
	.w5(32'hbac2926d),
	.w6(32'h3a0c18ae),
	.w7(32'hbbbeebeb),
	.w8(32'h3bc8afd7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc908eef),
	.w1(32'hbc26965e),
	.w2(32'hbbc8e785),
	.w3(32'h3b94fd96),
	.w4(32'h3c9bb64a),
	.w5(32'h3b8ad8a8),
	.w6(32'hbb8e4069),
	.w7(32'h3c680a9c),
	.w8(32'hba94d05d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb32708),
	.w1(32'hb99d444c),
	.w2(32'h3afbc3a9),
	.w3(32'h3c1b7a9d),
	.w4(32'h3bb7994c),
	.w5(32'h3c60a8bc),
	.w6(32'h3a1393b2),
	.w7(32'h3be23967),
	.w8(32'h3b758676),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a400815),
	.w1(32'h3ba0783f),
	.w2(32'h3c19c726),
	.w3(32'hbc08ef8d),
	.w4(32'h3b810e2a),
	.w5(32'hbb7a56a1),
	.w6(32'h3bd2f9b2),
	.w7(32'hbb1475d0),
	.w8(32'h3cb92f78),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb880b77a),
	.w1(32'hbbd3da01),
	.w2(32'hbbad549f),
	.w3(32'h3c5cb2f4),
	.w4(32'hbb1a6f4d),
	.w5(32'h3c43ba8a),
	.w6(32'h3b7c2f62),
	.w7(32'h3c1a8bae),
	.w8(32'hbb18de5a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c191e),
	.w1(32'h3bab48fc),
	.w2(32'h3ba2c7f4),
	.w3(32'h3c202f64),
	.w4(32'hbb8825e2),
	.w5(32'h3aa9dabd),
	.w6(32'h3bc26b21),
	.w7(32'hbb5ed37c),
	.w8(32'hb982582e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a7736),
	.w1(32'h3b9cce51),
	.w2(32'hbb1c0d16),
	.w3(32'h3c09537b),
	.w4(32'hbb2e7202),
	.w5(32'hbb34088b),
	.w6(32'hb712032f),
	.w7(32'hbbe2630c),
	.w8(32'hba3a5ecd),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f1fa7),
	.w1(32'hbbbc1058),
	.w2(32'h3c06c1ae),
	.w3(32'hba6d8033),
	.w4(32'hbb8635e7),
	.w5(32'h3b936150),
	.w6(32'h3b887139),
	.w7(32'h3c5dca00),
	.w8(32'hba27022a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa0f82),
	.w1(32'hbb7b1d18),
	.w2(32'hbbc95ac6),
	.w3(32'h3b2f2010),
	.w4(32'h3c99cd16),
	.w5(32'h3abe8bdf),
	.w6(32'h3a999e32),
	.w7(32'h3bf7d107),
	.w8(32'h36a989f8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc685084),
	.w1(32'hbc3617de),
	.w2(32'hbc030ddb),
	.w3(32'h3ba42b8f),
	.w4(32'h3bdec964),
	.w5(32'h39dd6209),
	.w6(32'h3c004860),
	.w7(32'h3aec5387),
	.w8(32'hbb27c7cd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fe75a),
	.w1(32'hb9998c67),
	.w2(32'h3a9c50ca),
	.w3(32'hba86ea6a),
	.w4(32'h3c10994f),
	.w5(32'hba9dbfb5),
	.w6(32'h3c23021f),
	.w7(32'h3bf2b1ba),
	.w8(32'hbb328861),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa65e7),
	.w1(32'h3c39f20e),
	.w2(32'hba00a155),
	.w3(32'hb81ebb9d),
	.w4(32'hbaa8db00),
	.w5(32'h3aa07b4d),
	.w6(32'h3a9a74b2),
	.w7(32'h3b72b78f),
	.w8(32'h3bd456f0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2edc4f),
	.w1(32'h3c02858a),
	.w2(32'hbb063805),
	.w3(32'h3c101e6a),
	.w4(32'h39d633e3),
	.w5(32'h39fd2a1b),
	.w6(32'h3c85860e),
	.w7(32'h3b12676b),
	.w8(32'h3c9c1e8f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1332dc),
	.w1(32'hbc1b6074),
	.w2(32'h3b4b22d4),
	.w3(32'hb921af95),
	.w4(32'hbbbded43),
	.w5(32'h3b1634ff),
	.w6(32'h3c24243e),
	.w7(32'h3b84f6ad),
	.w8(32'hbb0f2501),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aa236),
	.w1(32'h3c5d2ab8),
	.w2(32'hbc009d87),
	.w3(32'h3b5a3b4a),
	.w4(32'hba5de0a5),
	.w5(32'hbb144a98),
	.w6(32'hba8ecac6),
	.w7(32'h3b8f13cc),
	.w8(32'h3b989240),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39615702),
	.w1(32'h3cc23e3c),
	.w2(32'h3c06e6d4),
	.w3(32'hbbb29238),
	.w4(32'hbc12a0f1),
	.w5(32'hbb41990b),
	.w6(32'h3ba68764),
	.w7(32'h3b98d3c4),
	.w8(32'h3bc03071),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0228cb),
	.w1(32'h3c02cf5f),
	.w2(32'h3a2ce670),
	.w3(32'hb92bc12b),
	.w4(32'h3891d6ae),
	.w5(32'h3aa2f8d4),
	.w6(32'h38389f33),
	.w7(32'hbbd33b5e),
	.w8(32'h3b092b80),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ada213),
	.w1(32'hbb6e3547),
	.w2(32'h3bf010ea),
	.w3(32'h3adc327e),
	.w4(32'hbc58cfcc),
	.w5(32'hb9dce973),
	.w6(32'h3b863ec1),
	.w7(32'h3ce8e3af),
	.w8(32'h3ac07ede),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2bd0f),
	.w1(32'h3c767647),
	.w2(32'h3a7e0126),
	.w3(32'h3ba71951),
	.w4(32'hba11f2f1),
	.w5(32'h3bb068fe),
	.w6(32'h3be8362c),
	.w7(32'h3afb0b49),
	.w8(32'h398f62cb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19951),
	.w1(32'hbbf15c53),
	.w2(32'hbc1bad8f),
	.w3(32'h3cba3b54),
	.w4(32'h3b12a1c4),
	.w5(32'h3bbb659a),
	.w6(32'h3c0d02b0),
	.w7(32'h3be72fe2),
	.w8(32'h3b8d66ad),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b437055),
	.w1(32'hbc0ba5d0),
	.w2(32'hbbaf63e7),
	.w3(32'hbca57172),
	.w4(32'h3c2f6f0b),
	.w5(32'hbc23ff3f),
	.w6(32'h3b4c05d0),
	.w7(32'hb9d6d7d1),
	.w8(32'h3c878304),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb022),
	.w1(32'hbaa56cfb),
	.w2(32'hbc103f68),
	.w3(32'h3bf3677f),
	.w4(32'hbb2d6ce2),
	.w5(32'hbbd7ed56),
	.w6(32'h3b3c345b),
	.w7(32'hb992d255),
	.w8(32'h3b66b571),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb2ecc),
	.w1(32'hbc5bbe51),
	.w2(32'h3c3854d7),
	.w3(32'hbc3df4cb),
	.w4(32'hbb1f633c),
	.w5(32'h3ba24fc3),
	.w6(32'hbb0a5db2),
	.w7(32'hbb84f92c),
	.w8(32'h3a9b605e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f67db),
	.w1(32'hbaf0314e),
	.w2(32'h3c182e76),
	.w3(32'hbbcd40d3),
	.w4(32'hbb93e0f6),
	.w5(32'h3bef0da0),
	.w6(32'h3ac090d1),
	.w7(32'hbb9984f8),
	.w8(32'h3c39d16c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ccf08),
	.w1(32'hbb76f331),
	.w2(32'h3ce47942),
	.w3(32'h3bc6c20a),
	.w4(32'hbc409a92),
	.w5(32'h3bf83993),
	.w6(32'hbb32dbb8),
	.w7(32'hbba2743f),
	.w8(32'hbbcc2a53),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a59c6),
	.w1(32'hbc61889b),
	.w2(32'h3b0fe785),
	.w3(32'hbc3adc43),
	.w4(32'h3bb4d889),
	.w5(32'hbcc71434),
	.w6(32'h3c1ad623),
	.w7(32'h3b704722),
	.w8(32'hbba38938),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67c5c0),
	.w1(32'h3b736c21),
	.w2(32'h3c9e14d5),
	.w3(32'h3b83462f),
	.w4(32'hbbbc0fa2),
	.w5(32'hbbf0ade4),
	.w6(32'hbbe30512),
	.w7(32'hbad5ab45),
	.w8(32'hbbf92345),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9951fae),
	.w1(32'hb9ead256),
	.w2(32'hbb5667d8),
	.w3(32'h3b0d3214),
	.w4(32'hbb1da56e),
	.w5(32'hbb0a6f0e),
	.w6(32'hbb8747be),
	.w7(32'hbabb2a20),
	.w8(32'h3a8cc8df),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2303b8),
	.w1(32'hbb85e2c9),
	.w2(32'hbc275c6d),
	.w3(32'h3c20e218),
	.w4(32'hbc3225f5),
	.w5(32'h3c69a076),
	.w6(32'hbb7507e5),
	.w7(32'hbaa6e84b),
	.w8(32'hb9f8233d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18670f),
	.w1(32'h3bafee1b),
	.w2(32'hbb8b94ef),
	.w3(32'hbae6f611),
	.w4(32'h3b0d9182),
	.w5(32'hba5863d4),
	.w6(32'h3c01c773),
	.w7(32'hbc39f0fc),
	.w8(32'h3a75aee8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7681c8),
	.w1(32'hbbe97bf1),
	.w2(32'hbb9262bd),
	.w3(32'hbb5e4759),
	.w4(32'h3c1c6148),
	.w5(32'h3c15131f),
	.w6(32'hbb520e87),
	.w7(32'h3b9ba00c),
	.w8(32'h3b4c02f6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c633f62),
	.w1(32'hbc0a6fbe),
	.w2(32'hbb295e49),
	.w3(32'h3a6b89dd),
	.w4(32'hbc9b1d10),
	.w5(32'hbae78d6b),
	.w6(32'hbbd18b7b),
	.w7(32'hbb47e708),
	.w8(32'hbbceb5a2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad05fd2),
	.w1(32'hbc2c06d8),
	.w2(32'hb8e97992),
	.w3(32'h3c942979),
	.w4(32'h3847df9e),
	.w5(32'h3b87fe1d),
	.w6(32'h3cb202f3),
	.w7(32'h3c6fa440),
	.w8(32'h3c88c0c6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa082a),
	.w1(32'hbc012bad),
	.w2(32'hbafd1a92),
	.w3(32'hbb91c574),
	.w4(32'hbb8c278e),
	.w5(32'h3aea71c7),
	.w6(32'hbb385c77),
	.w7(32'h3b639b51),
	.w8(32'hbc616e0d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4386ac),
	.w1(32'h3bd00920),
	.w2(32'h35d90872),
	.w3(32'h3b94dbd8),
	.w4(32'hb9db47e6),
	.w5(32'h3b991153),
	.w6(32'hbc11fe0a),
	.w7(32'h3ca01dac),
	.w8(32'h398c17b9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd80c91),
	.w1(32'hbb0dc25d),
	.w2(32'hbc066641),
	.w3(32'h3cd4236c),
	.w4(32'hbb6480ff),
	.w5(32'hbb88766a),
	.w6(32'hba3cb66b),
	.w7(32'h3ba52aa8),
	.w8(32'hb845a517),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15a96e),
	.w1(32'hbc66995c),
	.w2(32'h3b8635a5),
	.w3(32'hbb16d37a),
	.w4(32'h3a894703),
	.w5(32'h3babaaab),
	.w6(32'hbc9bd03a),
	.w7(32'hbc9db13d),
	.w8(32'h3c7a049c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7adbc),
	.w1(32'h3c5abc0b),
	.w2(32'h3b2a5f1e),
	.w3(32'hbc2bd1ce),
	.w4(32'h3c0f1f05),
	.w5(32'h3c2d2919),
	.w6(32'hbc0ddc28),
	.w7(32'hbc44cf4a),
	.w8(32'hbc4f5c4d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afffd),
	.w1(32'h3b09cf61),
	.w2(32'hbb8e00a5),
	.w3(32'hbbafdbb4),
	.w4(32'hbae8a4da),
	.w5(32'h3b925951),
	.w6(32'hbbd2bf41),
	.w7(32'h389b094e),
	.w8(32'hbb495ccb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd39de5),
	.w1(32'h3be1621e),
	.w2(32'h3a95b9df),
	.w3(32'h3c01aa10),
	.w4(32'h3b8b02c8),
	.w5(32'h38af7bba),
	.w6(32'hbb1fd0ec),
	.w7(32'hb726ce91),
	.w8(32'hbc412669),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef7ed6),
	.w1(32'hbcc3d9e8),
	.w2(32'h3c34e0cb),
	.w3(32'hbaf0ce32),
	.w4(32'hbc2f6674),
	.w5(32'h3b334182),
	.w6(32'h3b8c7329),
	.w7(32'hb992ba84),
	.w8(32'hb917be25),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb569d12),
	.w1(32'hbb4ec6ab),
	.w2(32'hbc139e5f),
	.w3(32'h3bd763cf),
	.w4(32'hb98b0380),
	.w5(32'h3c2500d6),
	.w6(32'hbbfcb867),
	.w7(32'hbc02a78b),
	.w8(32'hbc1d2c31),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b5b54),
	.w1(32'hbca94408),
	.w2(32'hbb0a09eb),
	.w3(32'h39bf8a0e),
	.w4(32'h3bccdb46),
	.w5(32'hbc60785f),
	.w6(32'hbb12cc66),
	.w7(32'hba2bbee9),
	.w8(32'hb9d99014),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f601c),
	.w1(32'h3b58999d),
	.w2(32'hbb29b5b5),
	.w3(32'hbc536de9),
	.w4(32'h3c0b2989),
	.w5(32'hbc8f677c),
	.w6(32'hbbeb1a51),
	.w7(32'h3a50e4b5),
	.w8(32'h3b945650),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c93dc),
	.w1(32'hbbc654f4),
	.w2(32'h38a4a07a),
	.w3(32'h3c6e2fb1),
	.w4(32'hbc07291e),
	.w5(32'hba9be847),
	.w6(32'h3a976687),
	.w7(32'h3aa50803),
	.w8(32'hbb070235),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc99feb),
	.w1(32'h3b0ceb5d),
	.w2(32'hbb971436),
	.w3(32'hbac49b3e),
	.w4(32'hb9828631),
	.w5(32'hbc6509d6),
	.w6(32'h39e66806),
	.w7(32'hbb5d3f9f),
	.w8(32'h3ba87f45),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93b3e7),
	.w1(32'h3c20f391),
	.w2(32'hbc369a93),
	.w3(32'hbb33112f),
	.w4(32'hbc156657),
	.w5(32'hbbd2652b),
	.w6(32'h3c1122ad),
	.w7(32'hbb45b411),
	.w8(32'h3bd2aab8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a101f28),
	.w1(32'hbbe8efc2),
	.w2(32'h3b7bf922),
	.w3(32'h3af5e453),
	.w4(32'h3c84a48f),
	.w5(32'h3b8a2f6c),
	.w6(32'hba0f850d),
	.w7(32'hbbdf3e33),
	.w8(32'hbbbd5450),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a8758),
	.w1(32'hba0d7aa6),
	.w2(32'h3c117435),
	.w3(32'hbc2595d8),
	.w4(32'h3c177ec1),
	.w5(32'h3ca64209),
	.w6(32'h3c3e2a89),
	.w7(32'hbb6e1b08),
	.w8(32'hbbf51549),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca0d95),
	.w1(32'hb8333e37),
	.w2(32'h3c4eb1a0),
	.w3(32'hb9e674de),
	.w4(32'hbc031cce),
	.w5(32'hbc4f848e),
	.w6(32'h394a4f6b),
	.w7(32'h3a28e19d),
	.w8(32'hba9f9a5f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc596010),
	.w1(32'hbc2fcaa7),
	.w2(32'hbbcd6f41),
	.w3(32'h3cb1abe2),
	.w4(32'hbbe2ecb5),
	.w5(32'hbb4e20fb),
	.w6(32'hb9bd485c),
	.w7(32'hbc99d509),
	.w8(32'hbb4bb624),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39883f6c),
	.w1(32'hbc281b58),
	.w2(32'hba248680),
	.w3(32'hbc380dad),
	.w4(32'hbbb24c62),
	.w5(32'hbbd0822c),
	.w6(32'hbb86968b),
	.w7(32'hb831fbd1),
	.w8(32'h3c4eba21),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb53373),
	.w1(32'hbd4b5593),
	.w2(32'h3c598a8b),
	.w3(32'hbbe4731a),
	.w4(32'h3b7f27eb),
	.w5(32'h3a39c2a9),
	.w6(32'h3b2fb481),
	.w7(32'hbb8ec4ea),
	.w8(32'h3b6ed658),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc883bac),
	.w1(32'h3bca0f7f),
	.w2(32'hbaf953a1),
	.w3(32'h3c355d52),
	.w4(32'hbc27566e),
	.w5(32'h3c3b02de),
	.w6(32'hbb3ff9ca),
	.w7(32'hbb52fb0a),
	.w8(32'hbc780625),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6c5a94),
	.w1(32'h3b990be6),
	.w2(32'hba71dd4e),
	.w3(32'hbc3f9753),
	.w4(32'h3abefcce),
	.w5(32'hba820b87),
	.w6(32'hbc4b489b),
	.w7(32'hba5617a5),
	.w8(32'h3bc70632),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ee802),
	.w1(32'h3b8928e2),
	.w2(32'h3aaee858),
	.w3(32'h3aadd0ff),
	.w4(32'h3cfd32e6),
	.w5(32'hbc63eaf7),
	.w6(32'hba0a851b),
	.w7(32'h3b18f1ee),
	.w8(32'hbb9ddf5a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ed6f2),
	.w1(32'hbb2b8571),
	.w2(32'hbc45886b),
	.w3(32'hbb2b8fd6),
	.w4(32'hbba57dd1),
	.w5(32'h39c626df),
	.w6(32'h3c4ef987),
	.w7(32'h3ad896c1),
	.w8(32'hbc174246),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba847505),
	.w1(32'h3bcaaa00),
	.w2(32'hba8d1433),
	.w3(32'h3bafeff6),
	.w4(32'h3b4b5cce),
	.w5(32'hbaf67868),
	.w6(32'hb76b7ee5),
	.w7(32'hbb6eaff8),
	.w8(32'hbbf902a7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5267),
	.w1(32'hbc459c2e),
	.w2(32'hbc0b25bf),
	.w3(32'hbc1c4810),
	.w4(32'hbcaf6296),
	.w5(32'h3cbb8f69),
	.w6(32'hbc5f3d90),
	.w7(32'hbbdbdb6f),
	.w8(32'hbba59a48),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f186),
	.w1(32'hbbed7d75),
	.w2(32'hbc6554d5),
	.w3(32'h3bba29ca),
	.w4(32'h3c0389e5),
	.w5(32'h3bd0caac),
	.w6(32'h3bd1e9f7),
	.w7(32'h3c05e7ea),
	.w8(32'hbc61b443),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60548f),
	.w1(32'h3c2883a3),
	.w2(32'h3b259fb7),
	.w3(32'hbc92aa86),
	.w4(32'hba7dc13c),
	.w5(32'hbb99cf42),
	.w6(32'hbad02b09),
	.w7(32'hbaa41b43),
	.w8(32'h39d1b074),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb13ee),
	.w1(32'hbbd68be2),
	.w2(32'hbc4ec581),
	.w3(32'h3b242399),
	.w4(32'h3ba059f2),
	.w5(32'h3c451891),
	.w6(32'h3c6a1951),
	.w7(32'h3942a0ee),
	.w8(32'hb8886205),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07bcae),
	.w1(32'hbb2e358d),
	.w2(32'hbbf0d5f4),
	.w3(32'h3b0ad95c),
	.w4(32'hbaa70954),
	.w5(32'hbb366eaa),
	.w6(32'hbc0b4d19),
	.w7(32'hbc5ce1ae),
	.w8(32'hbbc96f5f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d3c52),
	.w1(32'hbb017794),
	.w2(32'h3bedd6fb),
	.w3(32'h38085edc),
	.w4(32'h3b182254),
	.w5(32'h3a31187b),
	.w6(32'hbb992ea4),
	.w7(32'h3cfd9d98),
	.w8(32'hba4744d0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842ecb),
	.w1(32'h3bcc6422),
	.w2(32'h3b6e36f9),
	.w3(32'h3c55f41d),
	.w4(32'h39f722e0),
	.w5(32'h3c214218),
	.w6(32'h3ccea9c1),
	.w7(32'hbb10daa4),
	.w8(32'hbb14a347),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85efc9),
	.w1(32'hbb64bef6),
	.w2(32'h3c5991f5),
	.w3(32'h3ae85a4b),
	.w4(32'hbc1b9d17),
	.w5(32'h3c893332),
	.w6(32'hbc10556d),
	.w7(32'hbb6b3966),
	.w8(32'h3c71e0b0),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af301),
	.w1(32'hbaf12253),
	.w2(32'hbc26580a),
	.w3(32'hbc0747df),
	.w4(32'h3a782e0b),
	.w5(32'hbc012655),
	.w6(32'hbab847da),
	.w7(32'h3ba2c87b),
	.w8(32'h39b3cadd),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81839e),
	.w1(32'hbb81c17a),
	.w2(32'hb8064ffc),
	.w3(32'hbc08ba4c),
	.w4(32'h3b496390),
	.w5(32'hbca79690),
	.w6(32'hbaae9dff),
	.w7(32'hbc400023),
	.w8(32'hbb6373ab),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb492ff24),
	.w1(32'h3adfe6f3),
	.w2(32'hbb4efc50),
	.w3(32'hbc5620b5),
	.w4(32'hbabfe868),
	.w5(32'h3c37632e),
	.w6(32'h3c0c5f20),
	.w7(32'h3c3471d1),
	.w8(32'hbc017ade),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9246a1),
	.w1(32'hb9ba5271),
	.w2(32'h3b41f8d7),
	.w3(32'hbc015453),
	.w4(32'hbba63f9c),
	.w5(32'h3ab5b8d9),
	.w6(32'hbc37ccde),
	.w7(32'hbb5b4b4d),
	.w8(32'hbbf808f0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886565),
	.w1(32'h3c14609f),
	.w2(32'h3bb82db3),
	.w3(32'hbb028ade),
	.w4(32'hbc190112),
	.w5(32'h3b8ec532),
	.w6(32'hbc87068e),
	.w7(32'hbc71c9d6),
	.w8(32'hbc0559e8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81d11b),
	.w1(32'h3c08c421),
	.w2(32'h3c3ef8ab),
	.w3(32'hbb419faf),
	.w4(32'h3c0cc11b),
	.w5(32'hbaa1b374),
	.w6(32'hbc3e7994),
	.w7(32'h3b650f55),
	.w8(32'hbbcdd953),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5fec5),
	.w1(32'h3d07d127),
	.w2(32'h3a50404e),
	.w3(32'hbbd0a98b),
	.w4(32'hbbb18ae7),
	.w5(32'h39a65dd9),
	.w6(32'h3b93ec3f),
	.w7(32'hbb8a1756),
	.w8(32'hbb3722be),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359786),
	.w1(32'h3b909c2a),
	.w2(32'hba27e16e),
	.w3(32'hba239189),
	.w4(32'h3b29eeb0),
	.w5(32'hbb64af75),
	.w6(32'hbbceb4f5),
	.w7(32'h3b417c20),
	.w8(32'h3a35c006),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64c4e8),
	.w1(32'h3d20aacb),
	.w2(32'hbc6dad94),
	.w3(32'h3bd33d38),
	.w4(32'h39460dae),
	.w5(32'hbbab55a0),
	.w6(32'hbb25ec42),
	.w7(32'hb9df11c0),
	.w8(32'hbce780d5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57b269),
	.w1(32'h3c120782),
	.w2(32'h3b4a3d46),
	.w3(32'h3b0c2fd3),
	.w4(32'hbc21caa3),
	.w5(32'h3bd64400),
	.w6(32'hbc542174),
	.w7(32'h3be6c529),
	.w8(32'h3b486b58),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e0c2),
	.w1(32'hbbcb1c58),
	.w2(32'h3c93b5b6),
	.w3(32'h3bfa7c3c),
	.w4(32'hbb32c504),
	.w5(32'hbbad9471),
	.w6(32'hbc03e9b8),
	.w7(32'h3bf400b1),
	.w8(32'h3c562adb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bf9c0),
	.w1(32'hbc44bb68),
	.w2(32'hbb69e692),
	.w3(32'hbbd5f798),
	.w4(32'hbc29d90c),
	.w5(32'hbc392bad),
	.w6(32'hbcf59719),
	.w7(32'h3ca4170a),
	.w8(32'hbbe4ab1e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fc75a),
	.w1(32'hbb421634),
	.w2(32'h3b91494d),
	.w3(32'hbc14136b),
	.w4(32'h3b8a0ac9),
	.w5(32'hbb8ba9cd),
	.w6(32'hbb89982e),
	.w7(32'hbbc7e4ed),
	.w8(32'hbb48f4c3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcc340),
	.w1(32'h3d41f89c),
	.w2(32'hbb307abf),
	.w3(32'hbcc9e699),
	.w4(32'hbafa416f),
	.w5(32'hbb849544),
	.w6(32'hbb85acaf),
	.w7(32'h3b73311c),
	.w8(32'h3c1ed3fa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule