module layer_10_featuremap_145(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bbeb4),
	.w1(32'h39acd858),
	.w2(32'hbb2567fe),
	.w3(32'hbaa94de3),
	.w4(32'hb93c1e5e),
	.w5(32'hbb688353),
	.w6(32'h3b0ddd0c),
	.w7(32'hba2d8def),
	.w8(32'h3b682e18),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81cf45),
	.w1(32'h3b163d88),
	.w2(32'h3b1f6b5c),
	.w3(32'hba9473ec),
	.w4(32'h3b07f10d),
	.w5(32'h3a744101),
	.w6(32'h3ae31779),
	.w7(32'h392ae571),
	.w8(32'h3a1d2788),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5c439),
	.w1(32'hbacb8413),
	.w2(32'hb94c9209),
	.w3(32'h39e4c531),
	.w4(32'hba035528),
	.w5(32'hba8c3e99),
	.w6(32'hba9808b8),
	.w7(32'hbaf3fe15),
	.w8(32'hbb1e0c1b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ebf33d),
	.w1(32'h3b4d4c52),
	.w2(32'h3ac0dc35),
	.w3(32'hbabf3784),
	.w4(32'hbb7c5104),
	.w5(32'hbbeaed24),
	.w6(32'hb9b0db66),
	.w7(32'h399f9041),
	.w8(32'hb95fb9c7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeae99f),
	.w1(32'hbb07a7ba),
	.w2(32'hbb4ee8c5),
	.w3(32'hbbd0c219),
	.w4(32'h3a0c16c9),
	.w5(32'hba11fc63),
	.w6(32'hbac7bbe0),
	.w7(32'hbace7c02),
	.w8(32'hbad02c5e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860d8e),
	.w1(32'h3a4990cb),
	.w2(32'hba9b0e6d),
	.w3(32'hbb04393d),
	.w4(32'hb63910cd),
	.w5(32'hbaf14eee),
	.w6(32'h3a971f55),
	.w7(32'hba5f1642),
	.w8(32'h3a2add0a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e96183),
	.w1(32'h3b6cbb86),
	.w2(32'h3b7cc019),
	.w3(32'h394b619c),
	.w4(32'h3b4fd7b7),
	.w5(32'h3aaa160f),
	.w6(32'h3a2f1e22),
	.w7(32'h3b350ce7),
	.w8(32'h3b139465),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d9715),
	.w1(32'h3b31e5c5),
	.w2(32'h3abdb5ec),
	.w3(32'h3ad9ff59),
	.w4(32'h3b72d00e),
	.w5(32'h3acae11b),
	.w6(32'h3ba57279),
	.w7(32'h3b708bc3),
	.w8(32'h3b21bb52),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71695d),
	.w1(32'hbb299d70),
	.w2(32'h3954b51c),
	.w3(32'hba6469c5),
	.w4(32'hbafbdc85),
	.w5(32'h3a932fc6),
	.w6(32'hbb178a63),
	.w7(32'hba24b5f6),
	.w8(32'h3a3fa43f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c8f2),
	.w1(32'h3b611731),
	.w2(32'h3b868f38),
	.w3(32'h3b66fdc9),
	.w4(32'h395ff7df),
	.w5(32'h3a05d879),
	.w6(32'h3b784bdb),
	.w7(32'h3a57af5c),
	.w8(32'h3ad681f0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80746a),
	.w1(32'hba79565b),
	.w2(32'hbad40146),
	.w3(32'hbb0219e6),
	.w4(32'h3a39b64d),
	.w5(32'hbae4cbe5),
	.w6(32'h3b6bc327),
	.w7(32'h3a91ca45),
	.w8(32'hbb265894),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb338b6),
	.w1(32'h3a8c8fe7),
	.w2(32'h3b1488d2),
	.w3(32'hbb9af85c),
	.w4(32'h3ab1febf),
	.w5(32'h3a32bb9f),
	.w6(32'h3b64b46b),
	.w7(32'h3afa650b),
	.w8(32'h3b573c01),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc0e9e),
	.w1(32'hb9bb3552),
	.w2(32'h3b6fb68a),
	.w3(32'h3ae58f41),
	.w4(32'h3ab7df13),
	.w5(32'h3b29082a),
	.w6(32'h3a2a42e8),
	.w7(32'h398b6c8a),
	.w8(32'h3af8b095),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e5dfa),
	.w1(32'h3b48131f),
	.w2(32'h39888a74),
	.w3(32'hb81ab5d5),
	.w4(32'h3b19f843),
	.w5(32'h39461fd0),
	.w6(32'h3b8c8ebf),
	.w7(32'h3b1857bc),
	.w8(32'h3ace8145),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65cf43),
	.w1(32'h3a46e1f6),
	.w2(32'hb9e60008),
	.w3(32'hbaa5ec76),
	.w4(32'h3bd39609),
	.w5(32'h3b27c2f1),
	.w6(32'h3b10332c),
	.w7(32'h3b20c349),
	.w8(32'h3afb4900),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cf7ef),
	.w1(32'h3abc9b4c),
	.w2(32'h3b447083),
	.w3(32'h3a94ab14),
	.w4(32'h3915aca5),
	.w5(32'h3afdeca9),
	.w6(32'h3a50d9f4),
	.w7(32'h39b3f5da),
	.w8(32'h3b3e94e0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce7d03),
	.w1(32'hbad09260),
	.w2(32'h3c2c0209),
	.w3(32'h399e0f21),
	.w4(32'hba42c5be),
	.w5(32'h3c756f7d),
	.w6(32'hbbd02cb3),
	.w7(32'h3bcc0ed1),
	.w8(32'hba5c1fd8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fd0d8),
	.w1(32'h3b513ae0),
	.w2(32'h3bab8e65),
	.w3(32'h3ca3658d),
	.w4(32'h3b5892ce),
	.w5(32'h3b57ba7e),
	.w6(32'h3b869e7d),
	.w7(32'h3b9017e9),
	.w8(32'h3b6d0d4b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c25d5),
	.w1(32'h39f5d673),
	.w2(32'h3a8c1e99),
	.w3(32'h3a97ae0d),
	.w4(32'h3a33e64a),
	.w5(32'h3a861dcf),
	.w6(32'hb9965812),
	.w7(32'h39178d36),
	.w8(32'h3b2f43ec),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d9106),
	.w1(32'hbad62238),
	.w2(32'h3a217624),
	.w3(32'h3a151908),
	.w4(32'hbaa12d65),
	.w5(32'h3a6319a9),
	.w6(32'hbaba1ca7),
	.w7(32'h38be7678),
	.w8(32'h3a3069c1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06aa33),
	.w1(32'hbad78400),
	.w2(32'hbade278e),
	.w3(32'h3958e6d1),
	.w4(32'hb9c29968),
	.w5(32'hba936e9f),
	.w6(32'hbada1caf),
	.w7(32'hbaef89c5),
	.w8(32'h399a043a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865794a),
	.w1(32'hbb2183d0),
	.w2(32'h3c2ca98c),
	.w3(32'hba72f261),
	.w4(32'h39bb90a0),
	.w5(32'hbb61d169),
	.w6(32'hbaa716a3),
	.w7(32'hba4367ba),
	.w8(32'h3b8b9c8f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8669d),
	.w1(32'h3b79bb6c),
	.w2(32'h3c806769),
	.w3(32'hbb191a9e),
	.w4(32'hbbc32563),
	.w5(32'h3c7fc44c),
	.w6(32'h39bc9b24),
	.w7(32'h3ba019fd),
	.w8(32'h3ad1f43f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3589),
	.w1(32'h3aa77673),
	.w2(32'h3b478a32),
	.w3(32'hbb6748e3),
	.w4(32'hb8e6d495),
	.w5(32'h3ae206a5),
	.w6(32'h3aaf5e1a),
	.w7(32'hba6fced4),
	.w8(32'h3ab430ce),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa85adb),
	.w1(32'hba8e63db),
	.w2(32'h3b4c3b51),
	.w3(32'h3b02c1fa),
	.w4(32'hba4cbbaf),
	.w5(32'h3b81982f),
	.w6(32'h3ac24732),
	.w7(32'hbacdeb8d),
	.w8(32'h3a759a91),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b406d6b),
	.w1(32'h3baafdbc),
	.w2(32'h3be52bed),
	.w3(32'h3b716c5c),
	.w4(32'hba8f8988),
	.w5(32'h3ab28471),
	.w6(32'hbb071078),
	.w7(32'hb9126e67),
	.w8(32'hbbdb0c7d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435b02),
	.w1(32'hb965f350),
	.w2(32'h3a44c9e2),
	.w3(32'h3ad4063f),
	.w4(32'h3a4ece89),
	.w5(32'h3a864c5c),
	.w6(32'hb9086d69),
	.w7(32'h398b4ec2),
	.w8(32'h39195ebc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae56d03),
	.w1(32'hb9e5ec4e),
	.w2(32'h3b0ec82d),
	.w3(32'hba81a230),
	.w4(32'hbb56ff5a),
	.w5(32'h37e3a2d6),
	.w6(32'h3af7b38e),
	.w7(32'hba4f2ab2),
	.w8(32'h3a853a68),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990d62d),
	.w1(32'hbb900724),
	.w2(32'h3ae5d48d),
	.w3(32'hba39aff2),
	.w4(32'hbb4d0d59),
	.w5(32'h3b8cc948),
	.w6(32'hbbcddc2f),
	.w7(32'hb9bb5e74),
	.w8(32'h3b90ae9f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0294e9),
	.w1(32'hbb9830d5),
	.w2(32'h3b8557eb),
	.w3(32'h3c0f860d),
	.w4(32'h3b8bd092),
	.w5(32'h3c6f46b7),
	.w6(32'hbc0184bc),
	.w7(32'hbad92ffb),
	.w8(32'h3c065f74),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c880268),
	.w1(32'hba87eb78),
	.w2(32'hba93cff6),
	.w3(32'h3cd5b13c),
	.w4(32'h39e4b288),
	.w5(32'h39ce6867),
	.w6(32'hba86b92c),
	.w7(32'hbae7a079),
	.w8(32'hba179a92),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24c6ec),
	.w1(32'h3a46f51b),
	.w2(32'h3a481b2a),
	.w3(32'h39d42505),
	.w4(32'h3a52e0e3),
	.w5(32'hb94dce7e),
	.w6(32'hb9c732fd),
	.w7(32'hb998acac),
	.w8(32'hb9ea40f3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9597297),
	.w1(32'hbaf102f5),
	.w2(32'h3a6ecf53),
	.w3(32'hba909d03),
	.w4(32'hbba7e90b),
	.w5(32'hbaa00f83),
	.w6(32'hbaff117c),
	.w7(32'hb98b9b40),
	.w8(32'h3b92fbb8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcedd05),
	.w1(32'hbaeefe93),
	.w2(32'hbb9ab24e),
	.w3(32'h3b6d010c),
	.w4(32'hba1967a5),
	.w5(32'hbb48eb78),
	.w6(32'hbb192089),
	.w7(32'hbb8c95af),
	.w8(32'hbaf4df5d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc137ba1),
	.w1(32'h3b07c9d7),
	.w2(32'h3af93dc9),
	.w3(32'hbc11d3e1),
	.w4(32'h39cd46ed),
	.w5(32'hb9b1e5db),
	.w6(32'h3a21fee7),
	.w7(32'hba45ec55),
	.w8(32'hb89fedf5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b7b01),
	.w1(32'h39de61a7),
	.w2(32'hba69fd05),
	.w3(32'hb91acb8d),
	.w4(32'h3af986de),
	.w5(32'h39f1c767),
	.w6(32'hb9b2eb2f),
	.w7(32'hba8651a9),
	.w8(32'h3a67d83a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3f9c4),
	.w1(32'h398e1164),
	.w2(32'h3ae917ea),
	.w3(32'hb5070780),
	.w4(32'h3ac654e4),
	.w5(32'h3b2b5dfc),
	.w6(32'hba1abb8b),
	.w7(32'hbb1e1068),
	.w8(32'h3ac55350),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bdc67),
	.w1(32'hbb81b91f),
	.w2(32'h3acba25c),
	.w3(32'h3ad17135),
	.w4(32'hbb8381cd),
	.w5(32'h3ac81dd0),
	.w6(32'h389f4932),
	.w7(32'hbbc2c802),
	.w8(32'hba4193be),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9028b),
	.w1(32'hbbdb3555),
	.w2(32'hb92e1560),
	.w3(32'hbabadf0b),
	.w4(32'hbbdfaa14),
	.w5(32'h3a1530db),
	.w6(32'h3ae58ba2),
	.w7(32'hbbb53132),
	.w8(32'hb9226000),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0ef17),
	.w1(32'h3a8c372a),
	.w2(32'h3a6a381a),
	.w3(32'h394a9c08),
	.w4(32'h3ac622c4),
	.w5(32'h3ab2ef57),
	.w6(32'h3a9a905d),
	.w7(32'h39e263f7),
	.w8(32'h3a0436e2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0b4f5),
	.w1(32'hbbcb64e9),
	.w2(32'hbb73c355),
	.w3(32'h394012cb),
	.w4(32'h3c0a70ab),
	.w5(32'h3c381644),
	.w6(32'hbc189d61),
	.w7(32'hbafbb13f),
	.w8(32'h3bc6df5d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c242db2),
	.w1(32'hba0cb716),
	.w2(32'hba0132f6),
	.w3(32'h3cbc9b2f),
	.w4(32'h3b11ed8d),
	.w5(32'hb995e2b0),
	.w6(32'hba1876cc),
	.w7(32'hba321667),
	.w8(32'h3a530d4d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f821f),
	.w1(32'hba7267c8),
	.w2(32'h3b140d88),
	.w3(32'h3a03727c),
	.w4(32'hba7accb0),
	.w5(32'h3ae69a1f),
	.w6(32'hbb27d536),
	.w7(32'h39514a4f),
	.w8(32'h389f094f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236479),
	.w1(32'h3bd07492),
	.w2(32'h3b8a6cab),
	.w3(32'h3b325c55),
	.w4(32'h3b388136),
	.w5(32'hba8358c7),
	.w6(32'h3c1b2748),
	.w7(32'h3ba0a47a),
	.w8(32'h3ace369b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68cc03),
	.w1(32'hbad2ee6b),
	.w2(32'h3b237084),
	.w3(32'hbbd29e63),
	.w4(32'hba1ab72e),
	.w5(32'h3b291a91),
	.w6(32'h3a6c7ba5),
	.w7(32'hbb0e1d0f),
	.w8(32'hba808152),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb026ad8),
	.w1(32'hba724d28),
	.w2(32'h3bbcc8ae),
	.w3(32'hb88bffa0),
	.w4(32'hba3f766d),
	.w5(32'h3aa87e17),
	.w6(32'hba8aaaea),
	.w7(32'hbb300d6f),
	.w8(32'h3aecd806),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb751e373),
	.w1(32'hbb02aa04),
	.w2(32'h3b396376),
	.w3(32'hbb103535),
	.w4(32'hbb0133c6),
	.w5(32'h3b1712de),
	.w6(32'hbad4616c),
	.w7(32'h3a7aaea8),
	.w8(32'h3b15ccb6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a4ba),
	.w1(32'h3b5c1b9c),
	.w2(32'h3c3cf284),
	.w3(32'h3bc1fd58),
	.w4(32'h3b7c28f9),
	.w5(32'h3c5016e1),
	.w6(32'h39a83eec),
	.w7(32'h3c35546d),
	.w8(32'h3bf43f0a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2616ad),
	.w1(32'hb98f343e),
	.w2(32'h3abe4601),
	.w3(32'h3beae7fb),
	.w4(32'hb952ed39),
	.w5(32'h3a1d3467),
	.w6(32'hbace1b4c),
	.w7(32'hb93a605a),
	.w8(32'h3a132443),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8875dc3),
	.w1(32'h3ac81494),
	.w2(32'hba1439b4),
	.w3(32'hb99dfa8e),
	.w4(32'h3ad5fd84),
	.w5(32'hb9c4a5fa),
	.w6(32'h3b2db120),
	.w7(32'h3a298245),
	.w8(32'hb965d321),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac7b34),
	.w1(32'h39da7c41),
	.w2(32'hba015645),
	.w3(32'hba193966),
	.w4(32'h39c5c438),
	.w5(32'hb9cb3879),
	.w6(32'h3a883435),
	.w7(32'h3a972ed6),
	.w8(32'h38eb5dd6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4894ad),
	.w1(32'h3b0ad0e3),
	.w2(32'h3a8f710b),
	.w3(32'hb9a0d074),
	.w4(32'hbb35e221),
	.w5(32'h3a4021f7),
	.w6(32'h3b55891a),
	.w7(32'hba5f110a),
	.w8(32'h39f53fdb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b046970),
	.w1(32'h39d4a945),
	.w2(32'h39d4f2f4),
	.w3(32'h3ab5b713),
	.w4(32'h39e6bd73),
	.w5(32'hb9ac8ab5),
	.w6(32'hba749bcc),
	.w7(32'hba8f0efc),
	.w8(32'h3a178670),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a30ad),
	.w1(32'h3b1cdbad),
	.w2(32'h3b5325f4),
	.w3(32'h3b3e3093),
	.w4(32'h3b5c1c77),
	.w5(32'h3b1a4bb0),
	.w6(32'h3b900e98),
	.w7(32'h3b679129),
	.w8(32'h3b8a54a6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba075c65),
	.w1(32'hba5bfca3),
	.w2(32'h3bf98524),
	.w3(32'hbb089eee),
	.w4(32'hbba6d439),
	.w5(32'h3b8f2671),
	.w6(32'hbadcbab1),
	.w7(32'h3bb4dcd5),
	.w8(32'hbb168f58),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b589741),
	.w1(32'hbc6bb380),
	.w2(32'hbc77b614),
	.w3(32'h390b5d23),
	.w4(32'h3bd7a35a),
	.w5(32'h3bb2339e),
	.w6(32'hbc3e4179),
	.w7(32'hbc3796bf),
	.w8(32'h3ba006f6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d25e2),
	.w1(32'hba23cfd7),
	.w2(32'h3b02f99a),
	.w3(32'h3caac7d1),
	.w4(32'h3b3042ff),
	.w5(32'h3ae9dd15),
	.w6(32'h3a3f5c46),
	.w7(32'h3b290e55),
	.w8(32'h3b17a899),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073435),
	.w1(32'h3b03451e),
	.w2(32'hbad565d1),
	.w3(32'h3b1489ad),
	.w4(32'h3b8f91ae),
	.w5(32'hb9fbecb0),
	.w6(32'h3b8559fb),
	.w7(32'hb9ce5e03),
	.w8(32'h3b2efcad),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d6abb),
	.w1(32'h3b01b21f),
	.w2(32'h389822fb),
	.w3(32'hbb1194af),
	.w4(32'h3a080a04),
	.w5(32'hbab6aaa5),
	.w6(32'h3af3f0c7),
	.w7(32'h376d807c),
	.w8(32'hb8f97093),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6beca0),
	.w1(32'h3a2391a2),
	.w2(32'h3980934a),
	.w3(32'hba8daff5),
	.w4(32'h3a16b089),
	.w5(32'h399f5c9e),
	.w6(32'h3a3dcb51),
	.w7(32'h39b68ca0),
	.w8(32'h393adc9e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39111bb5),
	.w1(32'h3a38ef5a),
	.w2(32'h3b06ed18),
	.w3(32'h39b5a0e6),
	.w4(32'h3a15216d),
	.w5(32'h3af855d2),
	.w6(32'hb985c5ee),
	.w7(32'hba36dc16),
	.w8(32'h3a4145e4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2421c),
	.w1(32'hbaddcf92),
	.w2(32'hb9553247),
	.w3(32'h3ab2558b),
	.w4(32'h3b0de77c),
	.w5(32'h3b04930b),
	.w6(32'h39bf2f2d),
	.w7(32'h3a3c5ce1),
	.w8(32'h39bd5b79),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1a63a),
	.w1(32'h3b0ed78c),
	.w2(32'h3a976f9d),
	.w3(32'h3ac382d6),
	.w4(32'h395f3aba),
	.w5(32'h3b148de9),
	.w6(32'h3afa7d96),
	.w7(32'hb8bcedd9),
	.w8(32'h3b688fdc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8f718),
	.w1(32'h3b1dd929),
	.w2(32'hba09dd3a),
	.w3(32'h3b8a1be0),
	.w4(32'h3a210654),
	.w5(32'hbb44a762),
	.w6(32'h3b8a413c),
	.w7(32'h3ac0cc7b),
	.w8(32'hbab32cbd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514ec4),
	.w1(32'hba86f6d7),
	.w2(32'hb9493cd3),
	.w3(32'hbb95b9b5),
	.w4(32'hbae61efe),
	.w5(32'hba0aa5e4),
	.w6(32'hba952bba),
	.w7(32'h3884c56d),
	.w8(32'h3a92d28c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa57a86),
	.w1(32'hb9d75804),
	.w2(32'h3afdff2d),
	.w3(32'h3a4a2cd0),
	.w4(32'hba370401),
	.w5(32'hbb0966e3),
	.w6(32'h3ad7745b),
	.w7(32'hba217fe2),
	.w8(32'h3b0cdcd8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb913c),
	.w1(32'hbb381f0d),
	.w2(32'h3a3e1079),
	.w3(32'hbb2935d1),
	.w4(32'h3c08d2aa),
	.w5(32'h3bf8d616),
	.w6(32'hbc1d22af),
	.w7(32'hbbe5d62f),
	.w8(32'h3b6b8f96),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbd479),
	.w1(32'h3b238fbb),
	.w2(32'h3c27866e),
	.w3(32'h3c985f12),
	.w4(32'h392c05bf),
	.w5(32'h3c38a012),
	.w6(32'hbb599f89),
	.w7(32'h3bae7285),
	.w8(32'h3b90ed49),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c60b7),
	.w1(32'hba09b4df),
	.w2(32'h3b18e302),
	.w3(32'h3b16b726),
	.w4(32'hbaa116ed),
	.w5(32'h3a98df52),
	.w6(32'hba19b5f1),
	.w7(32'hbb191c2a),
	.w8(32'h3a94ad8c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b04a),
	.w1(32'hbbb887e2),
	.w2(32'h3af942a9),
	.w3(32'h3aa5154d),
	.w4(32'hbb5b5942),
	.w5(32'h3b519efd),
	.w6(32'h3a428a39),
	.w7(32'hbbc8a5df),
	.w8(32'h3b255a67),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0c59e),
	.w1(32'h3ab59366),
	.w2(32'h3ab7e847),
	.w3(32'hbae6f3b3),
	.w4(32'h3ac0ac5f),
	.w5(32'h3837e0a5),
	.w6(32'h3a1a94aa),
	.w7(32'h3a583fe9),
	.w8(32'hb9767e3b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dec861),
	.w1(32'h39a4793a),
	.w2(32'h3a443a06),
	.w3(32'hb98df91b),
	.w4(32'h3a73fd88),
	.w5(32'h39fd4ea6),
	.w6(32'h3a9820e7),
	.w7(32'h396cd3bf),
	.w8(32'hb9a6e7ca),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903473e),
	.w1(32'h39986c04),
	.w2(32'h3902926d),
	.w3(32'hba76f3bb),
	.w4(32'h3984409b),
	.w5(32'h387a71a5),
	.w6(32'h39ca4e77),
	.w7(32'h392e94c5),
	.w8(32'hb90892b5),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c6001),
	.w1(32'h3a2d4cf9),
	.w2(32'h39bab72b),
	.w3(32'hba43ce19),
	.w4(32'h3a722c51),
	.w5(32'h398a50c8),
	.w6(32'hba8062ed),
	.w7(32'hba49281f),
	.w8(32'hba37e5b5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b4517),
	.w1(32'h3b047b57),
	.w2(32'h3929a63d),
	.w3(32'hba3b3ab2),
	.w4(32'h3abca8ab),
	.w5(32'hb9edc0fe),
	.w6(32'h3b4255ca),
	.w7(32'h3a7648d0),
	.w8(32'h3a5047af),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac65071),
	.w1(32'h3bcfbfc7),
	.w2(32'h3bb734b3),
	.w3(32'h3ad8c3b0),
	.w4(32'h3af15273),
	.w5(32'h3b1c5b37),
	.w6(32'h3bd0da6b),
	.w7(32'h3bf5ed5d),
	.w8(32'h3b0e0314),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f79ea),
	.w1(32'h3afec8e4),
	.w2(32'h3b2c5786),
	.w3(32'h3b8bbf94),
	.w4(32'h3a5d04b6),
	.w5(32'h3ae3f398),
	.w6(32'h3b7a6a1c),
	.w7(32'h3aeab0a9),
	.w8(32'h3b078b22),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0626b),
	.w1(32'h3a375415),
	.w2(32'h3b3864c0),
	.w3(32'h3b6228a3),
	.w4(32'h3afc14dd),
	.w5(32'h3b6e09fd),
	.w6(32'h3b554f45),
	.w7(32'hba759ef7),
	.w8(32'h3b1c7911),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f022),
	.w1(32'h3bb03f6d),
	.w2(32'h3ca71adf),
	.w3(32'h3b137d6b),
	.w4(32'hbba329b2),
	.w5(32'h3c4877b8),
	.w6(32'h3aff1319),
	.w7(32'h3c485cd7),
	.w8(32'hbb20ca7a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c411938),
	.w1(32'hbac9915e),
	.w2(32'hb9e79aaa),
	.w3(32'h3b6bc264),
	.w4(32'h38f0c7ed),
	.w5(32'h39df8e95),
	.w6(32'hbad6675d),
	.w7(32'hbb05c137),
	.w8(32'h38b90dc4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5226c3),
	.w1(32'hbb8d1e84),
	.w2(32'hbbd1a9e8),
	.w3(32'h3a60ac3d),
	.w4(32'h3c034711),
	.w5(32'h3bd293a2),
	.w6(32'hbb9cd437),
	.w7(32'hbb6b56e3),
	.w8(32'h3b887632),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3d8b3),
	.w1(32'h3a9802c0),
	.w2(32'h3b4f05e5),
	.w3(32'h3c36e800),
	.w4(32'h3b2b6c57),
	.w5(32'h3b53ec6b),
	.w6(32'h3aae51d4),
	.w7(32'h3aea34f0),
	.w8(32'h3b134496),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ceaf4),
	.w1(32'hbb136561),
	.w2(32'hbac4bf54),
	.w3(32'h3ab96981),
	.w4(32'h3a982f0a),
	.w5(32'h3b62b49a),
	.w6(32'hbb83e38b),
	.w7(32'hbb047428),
	.w8(32'hba75539d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25d103),
	.w1(32'h3b0dc612),
	.w2(32'h3acc098d),
	.w3(32'h3bccad5b),
	.w4(32'h3ac8b7a4),
	.w5(32'h37220bb0),
	.w6(32'h3a34db6a),
	.w7(32'h397a5497),
	.w8(32'h3aa81b07),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5893d8),
	.w1(32'h3b0cc320),
	.w2(32'h3a22721a),
	.w3(32'hb8832b40),
	.w4(32'h3b0439c0),
	.w5(32'h3ab090e8),
	.w6(32'hbb247497),
	.w7(32'h39f93664),
	.w8(32'hbb389f0d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a360),
	.w1(32'hb97f6382),
	.w2(32'h3a81f037),
	.w3(32'hbb308e28),
	.w4(32'h3b94c594),
	.w5(32'h3bab492d),
	.w6(32'hbb0630c2),
	.w7(32'hbad204f9),
	.w8(32'h392509f6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9675f2),
	.w1(32'hb8081d76),
	.w2(32'h3a9501a9),
	.w3(32'h3c12e9a0),
	.w4(32'hbb8f02a7),
	.w5(32'hba54b4a7),
	.w6(32'h3b255373),
	.w7(32'hba81dbbe),
	.w8(32'hb9ce6bc5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27525),
	.w1(32'hbb05afce),
	.w2(32'hbaa1287e),
	.w3(32'hbb21c170),
	.w4(32'hb9a1b5d6),
	.w5(32'h392a483b),
	.w6(32'hbae9600c),
	.w7(32'hbb1cf5cc),
	.w8(32'hba1427c0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f36179),
	.w1(32'hb9ede7c8),
	.w2(32'h3ba382d5),
	.w3(32'h3aa80d78),
	.w4(32'hbb7981eb),
	.w5(32'h3a778134),
	.w6(32'hbacdc17e),
	.w7(32'h3b1c796f),
	.w8(32'hbabb0019),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6ff0),
	.w1(32'h38727e5b),
	.w2(32'h3aedf908),
	.w3(32'h3b21a7da),
	.w4(32'h3b16e737),
	.w5(32'h3b5ddb8d),
	.w6(32'h391d0f5a),
	.w7(32'h39959b7b),
	.w8(32'h3a8496f9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b04ee),
	.w1(32'hbb1848c0),
	.w2(32'hb927663d),
	.w3(32'hb9befdab),
	.w4(32'hbb180596),
	.w5(32'h39e56577),
	.w6(32'hbab922d7),
	.w7(32'hbb74d4cf),
	.w8(32'hbab3bb43),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a136f11),
	.w1(32'h3a890d99),
	.w2(32'h3b6fd57f),
	.w3(32'h3934753f),
	.w4(32'h39d399e0),
	.w5(32'h3afb2402),
	.w6(32'h3819ec18),
	.w7(32'h3acf1980),
	.w8(32'h3ab03f38),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfac5f),
	.w1(32'h39c07ae9),
	.w2(32'h3b1d70a7),
	.w3(32'h3aba9bc7),
	.w4(32'hb9e5f896),
	.w5(32'h3af40bce),
	.w6(32'h3908d5d6),
	.w7(32'hba139b3e),
	.w8(32'h3a7e8018),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b5104),
	.w1(32'hbbd1d7c6),
	.w2(32'hbb8ea6d9),
	.w3(32'h3b641265),
	.w4(32'h3ba55fc8),
	.w5(32'h3be055d1),
	.w6(32'hbbb4c370),
	.w7(32'hbb294790),
	.w8(32'h3bae96d8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b602bae),
	.w1(32'h3960d72e),
	.w2(32'h3acfb145),
	.w3(32'h3c163272),
	.w4(32'hbaaa2443),
	.w5(32'hbadb8b07),
	.w6(32'hba9c0c77),
	.w7(32'hbb3af659),
	.w8(32'hbaa7e5e4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ed153),
	.w1(32'h39d85704),
	.w2(32'h3b9557aa),
	.w3(32'h3a472284),
	.w4(32'hba8cac4a),
	.w5(32'hba89c7fe),
	.w6(32'h3b9e5196),
	.w7(32'hb6c701aa),
	.w8(32'h3b8e8679),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6813d),
	.w1(32'h3b4dbc5e),
	.w2(32'h3c5af729),
	.w3(32'hbadd0c67),
	.w4(32'hbb5beeb9),
	.w5(32'h3c30d411),
	.w6(32'hba7ae5df),
	.w7(32'h3bd23c2e),
	.w8(32'hbb44318e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6abb61),
	.w1(32'hbaf58b7b),
	.w2(32'h39ab9c7a),
	.w3(32'hbbc988f6),
	.w4(32'hbb694c88),
	.w5(32'h38d82826),
	.w6(32'hbb174d14),
	.w7(32'hba5d8fb6),
	.w8(32'h3a51741b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef6397),
	.w1(32'h3a97da15),
	.w2(32'h3b8b5c42),
	.w3(32'hbb8eabd8),
	.w4(32'hba0194b6),
	.w5(32'h3b1e584b),
	.w6(32'h39026d0b),
	.w7(32'hb8456386),
	.w8(32'h3b2c56ee),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9719d2),
	.w1(32'hbb1bc200),
	.w2(32'h3af8888f),
	.w3(32'h3b95fac0),
	.w4(32'h3a9ad171),
	.w5(32'h3ba95e9b),
	.w6(32'hb8b3ac84),
	.w7(32'hbb1065a7),
	.w8(32'h3b9be92f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ec598),
	.w1(32'hbba21a1b),
	.w2(32'hba7f6131),
	.w3(32'h3b5587aa),
	.w4(32'hbbc0dec6),
	.w5(32'hbb56bb87),
	.w6(32'hbac019ac),
	.w7(32'hbc0de898),
	.w8(32'hbab57fc5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99c94f),
	.w1(32'h3a5d3562),
	.w2(32'h3c0cbbca),
	.w3(32'h3a32d0ec),
	.w4(32'h3b640293),
	.w5(32'h3aa22654),
	.w6(32'h3b3ed8d1),
	.w7(32'h39802f95),
	.w8(32'h3b087343),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7e572),
	.w1(32'h3a9a0008),
	.w2(32'h3aeae111),
	.w3(32'h3ad647ec),
	.w4(32'hb97a4e0e),
	.w5(32'h3a1a00cc),
	.w6(32'h3b98852b),
	.w7(32'h3acb301e),
	.w8(32'h3aee0d6c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa1e58),
	.w1(32'h39263cba),
	.w2(32'h3a0266aa),
	.w3(32'hbb0fb69b),
	.w4(32'h3a39878d),
	.w5(32'h39037eae),
	.w6(32'h3aa63d33),
	.w7(32'h3a14efb5),
	.w8(32'hb8efd833),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c8b43),
	.w1(32'h3a9d54bf),
	.w2(32'h3b178778),
	.w3(32'h3b31ca0d),
	.w4(32'h3a808ce2),
	.w5(32'h3b13c2f2),
	.w6(32'h3b942300),
	.w7(32'h3a8ff41e),
	.w8(32'h3b051621),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08f60a),
	.w1(32'hb9642e21),
	.w2(32'h3b7b04cd),
	.w3(32'h3a34f041),
	.w4(32'h3a92254e),
	.w5(32'h3ba9896e),
	.w6(32'hb954276c),
	.w7(32'h3ac59330),
	.w8(32'h3b40fe50),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821f2a),
	.w1(32'hba659e8a),
	.w2(32'h391e6b9c),
	.w3(32'h3a692c7f),
	.w4(32'hb867db62),
	.w5(32'hba49eaab),
	.w6(32'hb990bc06),
	.w7(32'hbae2db07),
	.w8(32'hbb123dd9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b3990),
	.w1(32'hbad02b35),
	.w2(32'hbae3e924),
	.w3(32'hb9fbec67),
	.w4(32'hb9a4d38f),
	.w5(32'h37c41b33),
	.w6(32'hbaa5e31b),
	.w7(32'hbae657fa),
	.w8(32'hba842a2a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a502327),
	.w1(32'h3b313190),
	.w2(32'h3b6fbdd0),
	.w3(32'h3b66fc5b),
	.w4(32'h3b3c4446),
	.w5(32'h3b1d8296),
	.w6(32'h3bae2705),
	.w7(32'h3b809a92),
	.w8(32'h3b4bca2c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391bd93e),
	.w1(32'h3af817e0),
	.w2(32'h3ac8fab4),
	.w3(32'h39fdb562),
	.w4(32'h3ab6efbe),
	.w5(32'h3ae4b26f),
	.w6(32'h3b589f25),
	.w7(32'hba016589),
	.w8(32'h3ab856d0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a258534),
	.w1(32'h3aae7984),
	.w2(32'h3a653825),
	.w3(32'h3a1ba3bb),
	.w4(32'h39b4daa5),
	.w5(32'h3ab4d58a),
	.w6(32'h3ae8692e),
	.w7(32'hb9790fa1),
	.w8(32'h3b32221a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7807df7),
	.w1(32'hb9dcaf32),
	.w2(32'hbaa79bf4),
	.w3(32'hb91d3581),
	.w4(32'hbb035954),
	.w5(32'h3a7b922a),
	.w6(32'h3b065ecb),
	.w7(32'hbb072be0),
	.w8(32'h39fe46aa),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134d39),
	.w1(32'hbad0f343),
	.w2(32'hbac95f9f),
	.w3(32'h39efd59a),
	.w4(32'hbaa89acc),
	.w5(32'hba67e99a),
	.w6(32'h3a3d3a9f),
	.w7(32'hbaa3f0d7),
	.w8(32'h3a634d56),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7dd8a),
	.w1(32'h3b0724b9),
	.w2(32'h3b1ffda1),
	.w3(32'h39399d6d),
	.w4(32'h3a557fd0),
	.w5(32'hbb056616),
	.w6(32'h3b02ec5b),
	.w7(32'h39b4c0ca),
	.w8(32'h3a715c37),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6045fc),
	.w1(32'h3a13da1a),
	.w2(32'h3a6d8954),
	.w3(32'hb8c6237d),
	.w4(32'hb94feb95),
	.w5(32'h3a18f9e2),
	.w6(32'h3982e105),
	.w7(32'h3b19ffd6),
	.w8(32'h3b38ae92),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73874e),
	.w1(32'h3a55643c),
	.w2(32'h3952fdc6),
	.w3(32'hbac9f081),
	.w4(32'h398f6354),
	.w5(32'hb9a93ce8),
	.w6(32'h3b724ba6),
	.w7(32'h3b0e4ece),
	.w8(32'hb78a219e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96a8e1),
	.w1(32'hb9988858),
	.w2(32'h3986b0ed),
	.w3(32'hbac2485b),
	.w4(32'h39f49d71),
	.w5(32'h3a3224ad),
	.w6(32'h3aa79c66),
	.w7(32'h3a7c9a63),
	.w8(32'h398c9f43),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f00ca1),
	.w1(32'h37ea00f9),
	.w2(32'hb981e255),
	.w3(32'h38da11ae),
	.w4(32'h390f5f09),
	.w5(32'hb8b034e6),
	.w6(32'h3b086608),
	.w7(32'h3a4f51b6),
	.w8(32'h398f1fb5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ddcdf2),
	.w1(32'hba25603c),
	.w2(32'h3b98c40b),
	.w3(32'hb9367e00),
	.w4(32'h3b53c4f0),
	.w5(32'h3aae89c9),
	.w6(32'h3af663a5),
	.w7(32'hb911a0df),
	.w8(32'h3a24ee46),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb613341),
	.w1(32'hbb0f8471),
	.w2(32'h3b407cdc),
	.w3(32'h399733f7),
	.w4(32'hbb20713b),
	.w5(32'h3a5d934c),
	.w6(32'hbb19f663),
	.w7(32'hbaa3b543),
	.w8(32'h3a44e6bd),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d31fd),
	.w1(32'h3a2904e6),
	.w2(32'hba4c5ea8),
	.w3(32'hba816dc8),
	.w4(32'h3a34afae),
	.w5(32'h398e2d69),
	.w6(32'hba747b91),
	.w7(32'hbb5569e3),
	.w8(32'hbaecfbd6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4b4ae),
	.w1(32'hb9bdf18f),
	.w2(32'h3a531eac),
	.w3(32'h3ac17bb5),
	.w4(32'hba844358),
	.w5(32'h39edbeca),
	.w6(32'hbaaa92e1),
	.w7(32'hbaad343c),
	.w8(32'h399caf77),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54b523),
	.w1(32'h39a462c6),
	.w2(32'h3a632128),
	.w3(32'h3a909805),
	.w4(32'h3a92a4e3),
	.w5(32'h3ae03803),
	.w6(32'h3b690949),
	.w7(32'h39802b62),
	.w8(32'h3b031dbe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67ef54),
	.w1(32'h3b96b6ab),
	.w2(32'h3c5e6f2e),
	.w3(32'hba09dc33),
	.w4(32'h3af4f6f8),
	.w5(32'h3846aab0),
	.w6(32'hb8c75c9a),
	.w7(32'h3b4a711d),
	.w8(32'h3b811682),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8be1),
	.w1(32'hbad3f1e5),
	.w2(32'hbb1dabe7),
	.w3(32'hba6a160d),
	.w4(32'hba6106d8),
	.w5(32'hbb465c3d),
	.w6(32'hbaca5036),
	.w7(32'hbb41fbfb),
	.w8(32'hb7e85ac8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70046d),
	.w1(32'hbb0bb165),
	.w2(32'hbaabcfe8),
	.w3(32'h39a68227),
	.w4(32'hb9ea7f45),
	.w5(32'hb998674b),
	.w6(32'hbb36354b),
	.w7(32'hbb1c2012),
	.w8(32'hba9cbd03),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d3e16),
	.w1(32'h394e6af5),
	.w2(32'h395bfabe),
	.w3(32'h3a188724),
	.w4(32'h3a0999d7),
	.w5(32'h397c271d),
	.w6(32'h3a5688e0),
	.w7(32'h39fcdbf9),
	.w8(32'h39da6c64),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319501),
	.w1(32'h3a38ca11),
	.w2(32'h3abde51c),
	.w3(32'hb98f2585),
	.w4(32'h3a539b08),
	.w5(32'h3a85ec22),
	.w6(32'hba6bf109),
	.w7(32'h398057a1),
	.w8(32'h3a86cf73),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a327ebd),
	.w1(32'h3a92041f),
	.w2(32'h3b16ac0f),
	.w3(32'h39da44b2),
	.w4(32'h39dc6220),
	.w5(32'h3ab69b19),
	.w6(32'h39d4742c),
	.w7(32'h3a167572),
	.w8(32'h3aef5143),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947479b),
	.w1(32'h3907d9e8),
	.w2(32'h395a4823),
	.w3(32'h380dead7),
	.w4(32'hb7bd001d),
	.w5(32'h3875c196),
	.w6(32'hb8c035ef),
	.w7(32'hb8b519ad),
	.w8(32'hb595b16e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f012b9),
	.w1(32'h38a2330b),
	.w2(32'h39c272db),
	.w3(32'h39db009a),
	.w4(32'h3894f09e),
	.w5(32'h39c78202),
	.w6(32'h39ecf3cf),
	.w7(32'h3942930a),
	.w8(32'h3a22727a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a98f01),
	.w1(32'hb763fe7b),
	.w2(32'h39f1aa72),
	.w3(32'h3a451edc),
	.w4(32'h389c854c),
	.w5(32'h39dbd212),
	.w6(32'h3a0855b3),
	.w7(32'hb5c900a6),
	.w8(32'h3a06c2a1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e755a4),
	.w1(32'h3991c60a),
	.w2(32'h3a61d954),
	.w3(32'h3983351e),
	.w4(32'hb7f6b061),
	.w5(32'h39e229b5),
	.w6(32'h390e405a),
	.w7(32'hb88641c2),
	.w8(32'h3a0015df),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81611),
	.w1(32'h3aad9989),
	.w2(32'h3ab4ccf1),
	.w3(32'h3ab86ac9),
	.w4(32'h39b850f3),
	.w5(32'h3a1202a6),
	.w6(32'h3aa4f8ab),
	.w7(32'h39c1415e),
	.w8(32'h3a155526),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a156bd8),
	.w1(32'h3abf9082),
	.w2(32'h3b3fe087),
	.w3(32'h3a9cfe22),
	.w4(32'h3a94bf86),
	.w5(32'h3b04fcdb),
	.w6(32'h3aa7bc08),
	.w7(32'h3a9a463b),
	.w8(32'h3b07980a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57d35e),
	.w1(32'hba41d98e),
	.w2(32'h39dc4d2b),
	.w3(32'h3a2ff035),
	.w4(32'hba2aceaf),
	.w5(32'h3a2ac813),
	.w6(32'h39c7d94f),
	.w7(32'hba5850e3),
	.w8(32'h3a72f319),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95438a),
	.w1(32'h38a1c395),
	.w2(32'h3a11378a),
	.w3(32'h3a499720),
	.w4(32'hba83356d),
	.w5(32'hb9781e2c),
	.w6(32'h3964d1f6),
	.w7(32'hba2e53f8),
	.w8(32'h3a2c5586),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a934707),
	.w1(32'h39fab773),
	.w2(32'h3a6fe017),
	.w3(32'h39ff3447),
	.w4(32'h37248f72),
	.w5(32'h39c80711),
	.w6(32'hb94f2f5e),
	.w7(32'hb9bd8532),
	.w8(32'h3a3a041e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a942ebd),
	.w1(32'hb924b69b),
	.w2(32'h394e5f0a),
	.w3(32'h3a482ba9),
	.w4(32'hba010e1b),
	.w5(32'h39a082ba),
	.w6(32'h3a1df984),
	.w7(32'hba13960a),
	.w8(32'h39c4f65a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32f615),
	.w1(32'h3a27535f),
	.w2(32'h3ac67f06),
	.w3(32'hb873a457),
	.w4(32'hb9d33a44),
	.w5(32'h39bee8c8),
	.w6(32'hb9dc754c),
	.w7(32'hb9c9da87),
	.w8(32'h3a44c423),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b376a8),
	.w1(32'h38504ca8),
	.w2(32'h39eb7ffa),
	.w3(32'h39d456d1),
	.w4(32'hb6baf305),
	.w5(32'h398d5c96),
	.w6(32'h39d40b44),
	.w7(32'h3843e573),
	.w8(32'h39dc0878),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3f03b),
	.w1(32'hbb412a41),
	.w2(32'hb9a864db),
	.w3(32'h3b31927c),
	.w4(32'hbaebfdfd),
	.w5(32'h3a97b2f4),
	.w6(32'h3b4be48e),
	.w7(32'hbadd1059),
	.w8(32'h3a9a27aa),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae27830),
	.w1(32'hb9b7c0d3),
	.w2(32'hb9c24bce),
	.w3(32'h3acefb47),
	.w4(32'hb8f7e44a),
	.w5(32'h3887d7a9),
	.w6(32'h3add2353),
	.w7(32'h3926bede),
	.w8(32'h3a2bec22),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7620b34),
	.w1(32'h380ee31a),
	.w2(32'hb68c7d04),
	.w3(32'h35d0a0c4),
	.w4(32'h384de132),
	.w5(32'h381b4b8b),
	.w6(32'h37c27b70),
	.w7(32'h37d78b0c),
	.w8(32'h379a5fdc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6851772),
	.w1(32'hb797fad8),
	.w2(32'h35ca843f),
	.w3(32'h358a90d3),
	.w4(32'hb721fd22),
	.w5(32'hb7e02a55),
	.w6(32'h37932e6d),
	.w7(32'hb755dab1),
	.w8(32'hb8e04986),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d03e7d),
	.w1(32'hb8f45b04),
	.w2(32'h394ba618),
	.w3(32'h3a02f697),
	.w4(32'hb98794c8),
	.w5(32'hb8cf5492),
	.w6(32'h39d8e0b5),
	.w7(32'hb91ab554),
	.w8(32'h392ee7fc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238f1e),
	.w1(32'hb8a9448d),
	.w2(32'h39eeffe2),
	.w3(32'h3af1cec5),
	.w4(32'hba30eaa2),
	.w5(32'h3a66803c),
	.w6(32'h3aa862b5),
	.w7(32'hba76f2f8),
	.w8(32'h3a956505),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf6f56),
	.w1(32'hb915dc94),
	.w2(32'h3afd11db),
	.w3(32'h3babba8b),
	.w4(32'h3aafe7a8),
	.w5(32'h3ad550a7),
	.w6(32'h3b4dad9a),
	.w7(32'h3acbd219),
	.w8(32'h3b266dd8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7257244),
	.w1(32'h37939c44),
	.w2(32'hb79924ff),
	.w3(32'hb713b6b9),
	.w4(32'h37704d1c),
	.w5(32'hb80372ff),
	.w6(32'h37753986),
	.w7(32'hb747d892),
	.w8(32'hb6dc3bff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaede91),
	.w1(32'h3a9b7dd0),
	.w2(32'h3b3106b3),
	.w3(32'h3ab4bbd4),
	.w4(32'h3a1619d3),
	.w5(32'h3aca8f56),
	.w6(32'h3acd3e6d),
	.w7(32'h3a0a61c9),
	.w8(32'h3aebee76),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4062d9),
	.w1(32'h39fb2f6e),
	.w2(32'h3a944145),
	.w3(32'h3aabcc7c),
	.w4(32'h39b0f202),
	.w5(32'h3a130e66),
	.w6(32'h3ab5ee2f),
	.w7(32'h39bd4c4e),
	.w8(32'h3a5e93ed),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a732ab4),
	.w1(32'h3af9dabb),
	.w2(32'h3b4fd878),
	.w3(32'h3aba6732),
	.w4(32'h3a9c5777),
	.w5(32'h3afdbae7),
	.w6(32'h3a23d5de),
	.w7(32'h39a249f9),
	.w8(32'h3a8d9ead),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76c65ac),
	.w1(32'hbb05dc62),
	.w2(32'h3aafc50e),
	.w3(32'h39ecaa50),
	.w4(32'hbb1c752f),
	.w5(32'h3a8d854a),
	.w6(32'h3a7a7f32),
	.w7(32'hbb35d640),
	.w8(32'hb8260526),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d5b24),
	.w1(32'hba255148),
	.w2(32'hb9904bee),
	.w3(32'h3a258496),
	.w4(32'hba160572),
	.w5(32'h38f7ee37),
	.w6(32'h3a4b1a31),
	.w7(32'hba1f3e18),
	.w8(32'h3821736c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d2b3a),
	.w1(32'hb95836fa),
	.w2(32'hb984645f),
	.w3(32'hb99c5d43),
	.w4(32'hb95ac570),
	.w5(32'hb970f45e),
	.w6(32'hb926f73b),
	.w7(32'hb95cb724),
	.w8(32'hb951a18f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b794c),
	.w1(32'hbb033342),
	.w2(32'hb990b892),
	.w3(32'hba9a8557),
	.w4(32'hbb28f05f),
	.w5(32'hb9df9152),
	.w6(32'hba9b0e2e),
	.w7(32'hbb4ab276),
	.w8(32'hbab7ee64),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a30b5),
	.w1(32'hbacd8865),
	.w2(32'h39660a7c),
	.w3(32'h3a9ef129),
	.w4(32'hbaf76c41),
	.w5(32'h3a28ec87),
	.w6(32'h3a0be550),
	.w7(32'hbb1c9b25),
	.w8(32'h39199086),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba493cbb),
	.w1(32'hbae7ac9a),
	.w2(32'h389ca3d1),
	.w3(32'hba29afeb),
	.w4(32'hbae6d38d),
	.w5(32'h3731dc90),
	.w6(32'h385fdd58),
	.w7(32'hbac9ab9c),
	.w8(32'hb941a34c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39609c16),
	.w1(32'h3973080a),
	.w2(32'h39d724a0),
	.w3(32'h399c5b7a),
	.w4(32'h397af3ec),
	.w5(32'h39abea9e),
	.w6(32'h396beb59),
	.w7(32'h37480a5c),
	.w8(32'h393a1c93),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372b6691),
	.w1(32'h383df079),
	.w2(32'h38612004),
	.w3(32'h3909dcb4),
	.w4(32'h38dfb547),
	.w5(32'h389b6646),
	.w6(32'h39273d04),
	.w7(32'h38acaf31),
	.w8(32'h38d11514),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dbddd),
	.w1(32'h3a4e2d4e),
	.w2(32'h3ac4a9c6),
	.w3(32'h39378a92),
	.w4(32'h399b34c4),
	.w5(32'h3a540471),
	.w6(32'hb90e8aa6),
	.w7(32'h38f23538),
	.w8(32'h3a7d89f2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a1fdf7),
	.w1(32'h38325272),
	.w2(32'h39baa760),
	.w3(32'hb8ff216b),
	.w4(32'hb7a6e30d),
	.w5(32'h3970a8b9),
	.w6(32'hb885575b),
	.w7(32'hb86b2fc4),
	.w8(32'hb58c97a8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982c98b),
	.w1(32'hba90f61d),
	.w2(32'hb83d1e17),
	.w3(32'hba36ced1),
	.w4(32'hbac4a763),
	.w5(32'hb9848a2f),
	.w6(32'hba5e9030),
	.w7(32'hbae2f694),
	.w8(32'hba6ea9ba),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91af461),
	.w1(32'hb8c7bc72),
	.w2(32'hb847478d),
	.w3(32'hb922acc8),
	.w4(32'hb8d67e0c),
	.w5(32'hb899f302),
	.w6(32'hb8ebcb04),
	.w7(32'hb8b61661),
	.w8(32'hb816dcea),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a11186),
	.w1(32'h3a1fdf94),
	.w2(32'h3b432531),
	.w3(32'h3a1d943f),
	.w4(32'h3aa217fc),
	.w5(32'h3b633b58),
	.w6(32'hba434fe9),
	.w7(32'h39f8395f),
	.w8(32'h3b4d0b58),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75e7cd6),
	.w1(32'hb64c0f6d),
	.w2(32'hb78c6522),
	.w3(32'hb7c7001a),
	.w4(32'h35148fed),
	.w5(32'hb7158ca2),
	.w6(32'h36cef1dd),
	.w7(32'h37d44fdb),
	.w8(32'hb7f0cdcd),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd74e0),
	.w1(32'hb87b18c1),
	.w2(32'hb8cf3a3e),
	.w3(32'hb86dbf78),
	.w4(32'hb863f35b),
	.w5(32'hb89b55dd),
	.w6(32'hb838e9bd),
	.w7(32'hb85f3a29),
	.w8(32'hb7caea8a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0474dd),
	.w1(32'hb9aa297f),
	.w2(32'h399b337f),
	.w3(32'hb7d62797),
	.w4(32'hba505beb),
	.w5(32'h397ada7d),
	.w6(32'hb95abd75),
	.w7(32'hba82c1e9),
	.w8(32'h3903338e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4fa54),
	.w1(32'h3910c40e),
	.w2(32'h3b5accdc),
	.w3(32'h3871bb18),
	.w4(32'hba4c70de),
	.w5(32'h3b274529),
	.w6(32'hb99181dc),
	.w7(32'hbaa51155),
	.w8(32'h3b1022dc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d6201),
	.w1(32'hba8adc15),
	.w2(32'h39ea5a0d),
	.w3(32'hba93ff03),
	.w4(32'hba7f01b5),
	.w5(32'h3994db1e),
	.w6(32'hb966e0e3),
	.w7(32'hba3651a3),
	.w8(32'h39ab77c7),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eacf0),
	.w1(32'h395ec332),
	.w2(32'h3adf5129),
	.w3(32'h3adc2c08),
	.w4(32'h3920bd2a),
	.w5(32'h3ab7f044),
	.w6(32'h3abfc7a6),
	.w7(32'hb876755b),
	.w8(32'h3aca3602),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac4626),
	.w1(32'h39235b04),
	.w2(32'h3a23cdb2),
	.w3(32'h3a1414dd),
	.w4(32'h37697509),
	.w5(32'h39a6e3f9),
	.w6(32'h3a1b7201),
	.w7(32'h38d3d732),
	.w8(32'h37d86ffb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3512af),
	.w1(32'h3a2845e5),
	.w2(32'h3b34ee11),
	.w3(32'h3b2548c1),
	.w4(32'hba511a4e),
	.w5(32'h3af971b6),
	.w6(32'h3abf9f0f),
	.w7(32'hb74bfaa5),
	.w8(32'h3b1de7e3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9342ee),
	.w1(32'h38d7e63b),
	.w2(32'h3b0c502f),
	.w3(32'h39fb7291),
	.w4(32'hba81bbf7),
	.w5(32'h3a8be560),
	.w6(32'h39a4d04a),
	.w7(32'hba6eb1e9),
	.w8(32'h3a84ced9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa24a16),
	.w1(32'h3ab6ffae),
	.w2(32'h3b3de02d),
	.w3(32'h3a84a591),
	.w4(32'h3a2e2f3a),
	.w5(32'h3aef78b7),
	.w6(32'h3a1dd55f),
	.w7(32'h39fa2c2c),
	.w8(32'h3aeb5ba5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376426f1),
	.w1(32'h38be6bc3),
	.w2(32'h375a8337),
	.w3(32'h37cac81d),
	.w4(32'h38b40327),
	.w5(32'hb44c7ea6),
	.w6(32'h38cb1e27),
	.w7(32'h38843656),
	.w8(32'hb8a8c169),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94d946),
	.w1(32'h3a273366),
	.w2(32'h3a22a89b),
	.w3(32'h3a3adf75),
	.w4(32'h35945948),
	.w5(32'h3831a361),
	.w6(32'h3a33a89c),
	.w7(32'h38402dce),
	.w8(32'h39c53287),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb760c388),
	.w1(32'hb7398a3b),
	.w2(32'hb884713c),
	.w3(32'h3662d47b),
	.w4(32'h37117b8c),
	.w5(32'hb83c626b),
	.w6(32'hb6e2107a),
	.w7(32'hb74b4793),
	.w8(32'hb8172064),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a239480),
	.w1(32'h3a02adaf),
	.w2(32'h3a911410),
	.w3(32'h39eb0103),
	.w4(32'h39ce02b5),
	.w5(32'h3a5d2ec3),
	.w6(32'h39a928cc),
	.w7(32'h3a090bab),
	.w8(32'h3a61b0d9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb2d99),
	.w1(32'hb939a958),
	.w2(32'hb903de11),
	.w3(32'h398970db),
	.w4(32'hb8fa581c),
	.w5(32'hb7bff06b),
	.w6(32'h398ec12e),
	.w7(32'hb948a8f3),
	.w8(32'h38acabc9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adea89e),
	.w1(32'h3a8ab9da),
	.w2(32'h3b0d3ac0),
	.w3(32'h3b4f56bb),
	.w4(32'h3a4ee145),
	.w5(32'h3aa4c94f),
	.w6(32'h3b3e5b99),
	.w7(32'h3a3c57f0),
	.w8(32'h3ac0ba44),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b4032b),
	.w1(32'hb7c0df90),
	.w2(32'h36818c91),
	.w3(32'hb7fc4736),
	.w4(32'hb5041fb0),
	.w5(32'h37c1e4e9),
	.w6(32'hb750b66e),
	.w7(32'h37227f77),
	.w8(32'hb6e94f9b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7de4fad),
	.w1(32'h37fb6b69),
	.w2(32'h37633f40),
	.w3(32'hb7a04dec),
	.w4(32'h37f4984e),
	.w5(32'h365f5ff6),
	.w6(32'h37b6a588),
	.w7(32'h380351dc),
	.w8(32'hb7ec5620),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e9820),
	.w1(32'hb8c37eba),
	.w2(32'h3912e1c4),
	.w3(32'h37cb8bea),
	.w4(32'hb9a9d257),
	.w5(32'h38356768),
	.w6(32'h395804b5),
	.w7(32'hba082ae2),
	.w8(32'h385a7966),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6bec5),
	.w1(32'h3a1ba829),
	.w2(32'h3a94f6dd),
	.w3(32'hba2275a1),
	.w4(32'hba240b29),
	.w5(32'h3a0c24c5),
	.w6(32'hba3f5780),
	.w7(32'hba129489),
	.w8(32'h3a6b8279),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3883),
	.w1(32'h389d2a1f),
	.w2(32'h3a62e64f),
	.w3(32'h3a1bee10),
	.w4(32'hb9bf78e5),
	.w5(32'h3a2a4717),
	.w6(32'h38f81e20),
	.w7(32'hba0d013f),
	.w8(32'h3a4780b3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b2971),
	.w1(32'hb881c70a),
	.w2(32'h38b4a74a),
	.w3(32'h386b6ed5),
	.w4(32'hb88789eb),
	.w5(32'h37e1e59d),
	.w6(32'h393d4f8f),
	.w7(32'hb81fa976),
	.w8(32'hb8a1ca10),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a087523),
	.w1(32'hba71cf18),
	.w2(32'h3b88f338),
	.w3(32'hbab4f8d3),
	.w4(32'hbb458a28),
	.w5(32'h3ac0767e),
	.w6(32'hbbbaa670),
	.w7(32'hbb6cf92b),
	.w8(32'hba955256),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40489f),
	.w1(32'hb942b0cd),
	.w2(32'h3b1bb31b),
	.w3(32'h3ad2e34d),
	.w4(32'hbb0fe6ac),
	.w5(32'h3a9009f2),
	.w6(32'h3ab6493b),
	.w7(32'hbb2cfb46),
	.w8(32'h3937e758),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38155364),
	.w1(32'h3950f0c7),
	.w2(32'h39d371a7),
	.w3(32'hb934bee4),
	.w4(32'h3921097a),
	.w5(32'h39954e92),
	.w6(32'h3728389b),
	.w7(32'h39ac45f0),
	.w8(32'h39c31377),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c38e0c),
	.w1(32'h3714136e),
	.w2(32'hb8a8733c),
	.w3(32'h38332c31),
	.w4(32'h381f9b0b),
	.w5(32'hb881b4a1),
	.w6(32'h37cafc8b),
	.w7(32'hb6e5eb0c),
	.w8(32'h37e05281),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ada82b),
	.w1(32'hb60f6dba),
	.w2(32'hb7b66466),
	.w3(32'h3796ec53),
	.w4(32'hb7890357),
	.w5(32'hb8117aed),
	.w6(32'h36d7dc32),
	.w7(32'h375866da),
	.w8(32'hb80b39f8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8130d97),
	.w1(32'h371cd0cc),
	.w2(32'hb7d03dc9),
	.w3(32'hb808630f),
	.w4(32'h379b7cba),
	.w5(32'hb7a52c28),
	.w6(32'h35c9e4e9),
	.w7(32'h372d8517),
	.w8(32'hb78d5c98),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ec061),
	.w1(32'h396d6560),
	.w2(32'h3a3d00bf),
	.w3(32'hb8812bc4),
	.w4(32'h398f723b),
	.w5(32'h3a0f0e45),
	.w6(32'hb9722dd8),
	.w7(32'h39dabe9e),
	.w8(32'h3a26e469),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0763fe),
	.w1(32'h3a94ac0d),
	.w2(32'h3aa41d98),
	.w3(32'h3adbae62),
	.w4(32'h39b8998c),
	.w5(32'h3ac7fda0),
	.w6(32'h3a0a3537),
	.w7(32'hb86509a8),
	.w8(32'h3af33cc8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a67a1),
	.w1(32'h3a5eddb6),
	.w2(32'h3afd586e),
	.w3(32'h3b6266b9),
	.w4(32'h3a3c00ac),
	.w5(32'h3ad64463),
	.w6(32'h3b46dde8),
	.w7(32'h3a98de2c),
	.w8(32'h3b1b448b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983dcd7),
	.w1(32'h37c137c7),
	.w2(32'h388c02cb),
	.w3(32'h397df638),
	.w4(32'hb915ea88),
	.w5(32'h37cd2c8c),
	.w6(32'h380a8b16),
	.w7(32'hb893aaef),
	.w8(32'h395edd27),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff2bbf),
	.w1(32'h3abf2548),
	.w2(32'h3b47e6cf),
	.w3(32'h3add7fb6),
	.w4(32'h3a91504d),
	.w5(32'h3b11ba80),
	.w6(32'h3a8d2706),
	.w7(32'h39abffb5),
	.w8(32'h3add9f8c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b22301),
	.w1(32'hb80179a6),
	.w2(32'h3a235d78),
	.w3(32'h3a882f01),
	.w4(32'h3a0399a3),
	.w5(32'h3a4f4d55),
	.w6(32'h3a5f398e),
	.w7(32'h3a093a5c),
	.w8(32'h3a465ba0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c9c794),
	.w1(32'hb70478ee),
	.w2(32'hb84d9c82),
	.w3(32'hb7bb9090),
	.w4(32'h36c9af02),
	.w5(32'hb8078769),
	.w6(32'hb7a82444),
	.w7(32'hb6f13b5f),
	.w8(32'hb812b78f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12439),
	.w1(32'h3a90d5f7),
	.w2(32'h3a1c1070),
	.w3(32'h3a1d60e3),
	.w4(32'h3a10813a),
	.w5(32'h38526345),
	.w6(32'h3a52ea4a),
	.w7(32'h39c67589),
	.w8(32'h3985a976),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb884db82),
	.w1(32'hb78aff89),
	.w2(32'hb905b92a),
	.w3(32'hb85943a6),
	.w4(32'hb69c7cac),
	.w5(32'hb8dd9a4c),
	.w6(32'hb800cc5b),
	.w7(32'hb7a81828),
	.w8(32'hb8cc5161),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32278c),
	.w1(32'h39825bd0),
	.w2(32'h3ae7eb05),
	.w3(32'h3a13f118),
	.w4(32'h394d55d7),
	.w5(32'h3ab4c371),
	.w6(32'h39fa0076),
	.w7(32'h394a5459),
	.w8(32'h3abfde08),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeccdf),
	.w1(32'hbaf5c6f5),
	.w2(32'h3a1a33ab),
	.w3(32'h3980c350),
	.w4(32'hbb3676ad),
	.w5(32'h3a3c24f1),
	.w6(32'h39ee090c),
	.w7(32'hbb52f736),
	.w8(32'h38fec10c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67855c),
	.w1(32'hb93446e4),
	.w2(32'h3abe44bf),
	.w3(32'h39f22f39),
	.w4(32'hba39fb9c),
	.w5(32'h3a94119f),
	.w6(32'h39a09451),
	.w7(32'hba774272),
	.w8(32'h3a89f594),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc83d7),
	.w1(32'hba495ee1),
	.w2(32'h3867be63),
	.w3(32'hba10745a),
	.w4(32'hba47f24c),
	.w5(32'h3888daf6),
	.w6(32'hb988209d),
	.w7(32'hba4affa8),
	.w8(32'hb8c0b5c5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ad937),
	.w1(32'hb947951d),
	.w2(32'h3acd4377),
	.w3(32'h3a92c821),
	.w4(32'hba4fc2bf),
	.w5(32'h3a9472b6),
	.w6(32'h3ab2c851),
	.w7(32'hba0586fa),
	.w8(32'h3ade71c0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a6144),
	.w1(32'h3a4e1225),
	.w2(32'h3aaed0df),
	.w3(32'h3ab1394e),
	.w4(32'h39f31c4b),
	.w5(32'h3a3d368e),
	.w6(32'h3aa7f3b0),
	.w7(32'h3a1a5610),
	.w8(32'h3a8247e1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39b141),
	.w1(32'h3a0ee5b7),
	.w2(32'h3b344a8c),
	.w3(32'h3bd8367d),
	.w4(32'h3b1fc77c),
	.w5(32'h3b3bef39),
	.w6(32'h3b85881d),
	.w7(32'h3b08df4c),
	.w8(32'h3b4be5a9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90116bf),
	.w1(32'hb79311d8),
	.w2(32'hb7d1eca5),
	.w3(32'hb920ea9f),
	.w4(32'hb6e7df0f),
	.w5(32'hb77d63ee),
	.w6(32'hb8437f76),
	.w7(32'hb7dd31d7),
	.w8(32'hb7e6e9ef),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a9725),
	.w1(32'h3790207d),
	.w2(32'h3488054e),
	.w3(32'h378426d9),
	.w4(32'h387072b6),
	.w5(32'h37e6f7a9),
	.w6(32'h384ebdc0),
	.w7(32'hb70c3a72),
	.w8(32'hb668823e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43a87b),
	.w1(32'hba0c9e94),
	.w2(32'h3ae56c21),
	.w3(32'h3a5374bb),
	.w4(32'hba656d18),
	.w5(32'h3ad62bbd),
	.w6(32'hb6fd605c),
	.w7(32'hba820c89),
	.w8(32'h3aeeb869),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b647c),
	.w1(32'hb9659deb),
	.w2(32'h3b244472),
	.w3(32'hb9c1da77),
	.w4(32'hbab66f4a),
	.w5(32'h3acaed48),
	.w6(32'hba5c7cfb),
	.w7(32'hbac35ec7),
	.w8(32'h3a7b077d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95ec61),
	.w1(32'hb9b2c0cf),
	.w2(32'h3accb716),
	.w3(32'h3a5e9c83),
	.w4(32'hba88ba9d),
	.w5(32'h3a54d8c7),
	.w6(32'h3a190ae8),
	.w7(32'hba947c7b),
	.w8(32'h3a8e2652),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a838b1),
	.w1(32'h3a88f7fd),
	.w2(32'h3a885795),
	.w3(32'h3999dbcc),
	.w4(32'h3a003a7e),
	.w5(32'h39de0001),
	.w6(32'h39850050),
	.w7(32'h3a75d270),
	.w8(32'h3a31ff1b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ec391),
	.w1(32'h38f8c9b2),
	.w2(32'hb7da00aa),
	.w3(32'h3743932e),
	.w4(32'h37f0f55f),
	.w5(32'hb82ad3d7),
	.w6(32'h38711a47),
	.w7(32'h38a4be6c),
	.w8(32'hb7f428e4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984bb9e),
	.w1(32'h39b1fccc),
	.w2(32'h39300b27),
	.w3(32'h39949f3f),
	.w4(32'h3982b4d8),
	.w5(32'h38df9282),
	.w6(32'h39a94c14),
	.w7(32'h398d796a),
	.w8(32'h38b96963),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94486d4),
	.w1(32'hb9d421e1),
	.w2(32'h3b083422),
	.w3(32'h39ae57b8),
	.w4(32'h3a80d673),
	.w5(32'h3b254ce5),
	.w6(32'hb9daf4c8),
	.w7(32'h39bf0820),
	.w8(32'h3b07686d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c605e),
	.w1(32'h3ac926de),
	.w2(32'h3b848648),
	.w3(32'h3b33fb33),
	.w4(32'h3a538acb),
	.w5(32'h3b57fc53),
	.w6(32'h388d3cac),
	.w7(32'h398240e6),
	.w8(32'h3b44fd59),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b98ea),
	.w1(32'h3996fa26),
	.w2(32'h3aaecfc5),
	.w3(32'h3b3b9ea9),
	.w4(32'h3ab87b86),
	.w5(32'h3ab6df96),
	.w6(32'h3b3a2290),
	.w7(32'h3aad9bd9),
	.w8(32'h3ac8f17f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca1507),
	.w1(32'hbb25a429),
	.w2(32'hba31d123),
	.w3(32'h397c08f3),
	.w4(32'hbaf498f7),
	.w5(32'h38c802ad),
	.w6(32'h39e0d7f3),
	.w7(32'hbada8513),
	.w8(32'hb84c6c76),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa889b0),
	.w1(32'hb93329e3),
	.w2(32'h3ae5f16d),
	.w3(32'h3a107b8c),
	.w4(32'hba95e56e),
	.w5(32'h3aa58a12),
	.w6(32'h39edf3ab),
	.w7(32'hbad02e7c),
	.w8(32'h3a0996e8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb357b),
	.w1(32'hb7a89fa7),
	.w2(32'hb78c2eb2),
	.w3(32'hb90d238f),
	.w4(32'hb7845b39),
	.w5(32'hb702fd9c),
	.w6(32'hb7b33c73),
	.w7(32'hb73ffccb),
	.w8(32'hb823c8d5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81689ce),
	.w1(32'hb7e5b0ef),
	.w2(32'hb736a3ab),
	.w3(32'hb80d78bb),
	.w4(32'h3779ebdd),
	.w5(32'h37b26888),
	.w6(32'hb805ed6f),
	.w7(32'hb6643259),
	.w8(32'hb781b5b6),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10bc98),
	.w1(32'hb93bead3),
	.w2(32'hb924cbd3),
	.w3(32'hb7d31e37),
	.w4(32'h398f904b),
	.w5(32'h39398f57),
	.w6(32'h380d6771),
	.w7(32'h398ff1c1),
	.w8(32'hb8c779d6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e90f7d),
	.w1(32'h37f69551),
	.w2(32'hb843d416),
	.w3(32'hb90ac596),
	.w4(32'h37efe465),
	.w5(32'hb8743f1a),
	.w6(32'hb5c12926),
	.w7(32'h360346e9),
	.w8(32'hb78edcc6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e107f),
	.w1(32'h38d4ef84),
	.w2(32'h39e47e36),
	.w3(32'hb8f0ab39),
	.w4(32'h39970df9),
	.w5(32'h39e2ed65),
	.w6(32'hb8693b58),
	.w7(32'h399ce5d9),
	.w8(32'h39a8efeb),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e9de),
	.w1(32'h39303946),
	.w2(32'h3ac7cbf7),
	.w3(32'hb8fadfbb),
	.w4(32'hba6aa9b8),
	.w5(32'h3a444b05),
	.w6(32'hba92fbc5),
	.w7(32'hba93514b),
	.w8(32'h3a28a80e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3dbada),
	.w1(32'h3842c0ae),
	.w2(32'h3a9690c0),
	.w3(32'h3a3027d6),
	.w4(32'hb984ea32),
	.w5(32'h3a8519be),
	.w6(32'hb98302dd),
	.w7(32'hba3e4365),
	.w8(32'h3a22d313),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901a37e),
	.w1(32'hb8e66a5e),
	.w2(32'h36ae3285),
	.w3(32'hb901ade1),
	.w4(32'hb77f85cb),
	.w5(32'h38b7f0aa),
	.w6(32'hb895c0f8),
	.w7(32'hb7950517),
	.w8(32'hb87fe116),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a097a6c),
	.w1(32'h389107f3),
	.w2(32'h3b267ce8),
	.w3(32'h3b0abba8),
	.w4(32'h3a2d4a04),
	.w5(32'h3b19ce3e),
	.w6(32'h3ae6dfe0),
	.w7(32'h3a1e9b8c),
	.w8(32'h3b37c40e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c8ab3),
	.w1(32'h3a159244),
	.w2(32'h3a5a6629),
	.w3(32'h3a4d4762),
	.w4(32'h39f6e8ca),
	.w5(32'h3a158f49),
	.w6(32'h39d9c2d4),
	.w7(32'h39fec6cf),
	.w8(32'h3a1f7be5),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ed6a3),
	.w1(32'h38a445f3),
	.w2(32'hb795f984),
	.w3(32'h384d61ee),
	.w4(32'h38f8ecf5),
	.w5(32'h37959e1d),
	.w6(32'h3909663f),
	.w7(32'h38875cc9),
	.w8(32'h36dda3f4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984e568),
	.w1(32'h394cad47),
	.w2(32'h3a4d6dbc),
	.w3(32'h3a133487),
	.w4(32'h39e47208),
	.w5(32'h3a20748c),
	.w6(32'h39cf4943),
	.w7(32'h39a424e4),
	.w8(32'h3a11402d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8008180),
	.w1(32'hb81d6673),
	.w2(32'hb8562948),
	.w3(32'hb7b58fcd),
	.w4(32'hb7bf86d5),
	.w5(32'hb82956f1),
	.w6(32'hb78c24e1),
	.w7(32'hb66fe206),
	.w8(32'hb858cab1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70fdcc3),
	.w1(32'h383d02e4),
	.w2(32'h3882d9d5),
	.w3(32'hb87258a9),
	.w4(32'hb793f1dd),
	.w5(32'h35eee788),
	.w6(32'hb6237cdc),
	.w7(32'hb78b4a12),
	.w8(32'h378ff496),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7633db5),
	.w1(32'h35d50ba7),
	.w2(32'hb80461e7),
	.w3(32'hb79a346a),
	.w4(32'h3742cc98),
	.w5(32'hb7747421),
	.w6(32'h3642bcb4),
	.w7(32'hb707dd18),
	.w8(32'hb719b4aa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c6c66f),
	.w1(32'hb68bde6f),
	.w2(32'hb7efcebd),
	.w3(32'hb78905b3),
	.w4(32'h35e5f14f),
	.w5(32'hb7b4ddbf),
	.w6(32'hb6caea05),
	.w7(32'h367d7946),
	.w8(32'hb7219e62),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba203433),
	.w1(32'hba8159c5),
	.w2(32'hb995194e),
	.w3(32'hb9220240),
	.w4(32'hba4d4925),
	.w5(32'h388d1393),
	.w6(32'h38000d9d),
	.w7(32'hba5024b1),
	.w8(32'h37ce3b80),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f495),
	.w1(32'h3b06b9ec),
	.w2(32'h3b610dbd),
	.w3(32'h3a0e2fb9),
	.w4(32'hb8998ab7),
	.w5(32'h3aa0ba5d),
	.w6(32'h39ea968b),
	.w7(32'h38747c31),
	.w8(32'h3ac01986),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb82f3),
	.w1(32'h3906864c),
	.w2(32'h3aa5447e),
	.w3(32'hb979bbfc),
	.w4(32'hba25af76),
	.w5(32'h39d543ae),
	.w6(32'hba320eaa),
	.w7(32'hba4a727c),
	.w8(32'h39d482cb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a946bcb),
	.w1(32'h3b0385f4),
	.w2(32'h3b4dc0cd),
	.w3(32'h3adb3990),
	.w4(32'h3aadca65),
	.w5(32'h3b0c5a54),
	.w6(32'h3a94d041),
	.w7(32'h3ab61634),
	.w8(32'h3ae70dc3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77d53c6),
	.w1(32'hb7e92cc8),
	.w2(32'hb7a52caf),
	.w3(32'hb63a6672),
	.w4(32'hb7e0e47a),
	.w5(32'hb7e5b7d6),
	.w6(32'h386908de),
	.w7(32'hb66f2c15),
	.w8(32'h380b8586),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f75137),
	.w1(32'h3939a899),
	.w2(32'h379b363f),
	.w3(32'h38cd3259),
	.w4(32'h3929a166),
	.w5(32'hb7a96114),
	.w6(32'h38c27456),
	.w7(32'h38ff4f61),
	.w8(32'h386ffb5c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77746ca),
	.w1(32'hb6a808b3),
	.w2(32'hb81aa4f5),
	.w3(32'h32b90c05),
	.w4(32'h3757f35b),
	.w5(32'hb7d2c637),
	.w6(32'hb5094224),
	.w7(32'hb74c183e),
	.w8(32'hb7812281),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8018364),
	.w1(32'hb71a4eae),
	.w2(32'hb8664f80),
	.w3(32'hb7c98c16),
	.w4(32'h36cb0ce3),
	.w5(32'hb811ade5),
	.w6(32'hb778dc27),
	.w7(32'hb773379c),
	.w8(32'hb788f251),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a6d9),
	.w1(32'h3a7adb67),
	.w2(32'h3ab9d816),
	.w3(32'h399c7a47),
	.w4(32'hb96b43b0),
	.w5(32'h39d5a86c),
	.w6(32'h390156d5),
	.w7(32'hb99b1e66),
	.w8(32'h3a73e9ee),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fdf504),
	.w1(32'h35b2504d),
	.w2(32'h374e9bf6),
	.w3(32'hb6ce9320),
	.w4(32'h366ad2a3),
	.w5(32'h37eddba6),
	.w6(32'hb6d0bae0),
	.w7(32'h37e77fe3),
	.w8(32'hb85e0d6c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea5220),
	.w1(32'hba6beeec),
	.w2(32'h39aefa21),
	.w3(32'hb9fcb2e6),
	.w4(32'hba32d33f),
	.w5(32'h395189fd),
	.w6(32'hb98a6928),
	.w7(32'hba43843d),
	.w8(32'h3985468a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd191d),
	.w1(32'h38cf9203),
	.w2(32'h398bf4e8),
	.w3(32'h3965410c),
	.w4(32'hb8de5efa),
	.w5(32'h371fd9a0),
	.w6(32'h39db61fa),
	.w7(32'hb8464991),
	.w8(32'h37c0c9a7),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb740b352),
	.w1(32'h34155b48),
	.w2(32'hb7f9b12d),
	.w3(32'h36aa600d),
	.w4(32'h379585c0),
	.w5(32'hb78289c0),
	.w6(32'h37669e70),
	.w7(32'hb707c9d6),
	.w8(32'hb4054182),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392573c5),
	.w1(32'hb8079232),
	.w2(32'h397eed9a),
	.w3(32'h39a348d1),
	.w4(32'h3838b5c1),
	.w5(32'h39bd022f),
	.w6(32'hb8e87fa7),
	.w7(32'h39351dbe),
	.w8(32'h3a17aa6b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38af242a),
	.w1(32'h38d3c290),
	.w2(32'h33461bd4),
	.w3(32'h38818e6d),
	.w4(32'h3897733f),
	.w5(32'hb7891a1e),
	.w6(32'h38d5aa84),
	.w7(32'h38f73a0e),
	.w8(32'h38ce93d1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21b8c),
	.w1(32'h3b1e2e89),
	.w2(32'h3b3c33e6),
	.w3(32'h3a6088b5),
	.w4(32'h39fb79ac),
	.w5(32'h3a0e82da),
	.w6(32'h3abab049),
	.w7(32'h3a062552),
	.w8(32'h3998208f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f2dc13),
	.w1(32'h396e5ed3),
	.w2(32'h393db461),
	.w3(32'hb7a47f18),
	.w4(32'h38f326a6),
	.w5(32'hb84f279e),
	.w6(32'h38a4d0c1),
	.w7(32'hb8201b21),
	.w8(32'h378e30e0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39973a3c),
	.w1(32'hbb0b51b9),
	.w2(32'hbb10f5f2),
	.w3(32'hba5a527f),
	.w4(32'hbb37025b),
	.w5(32'hbb0d50c9),
	.w6(32'h3ab5cd5b),
	.w7(32'hbaa2de6b),
	.w8(32'hba1ea747),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule