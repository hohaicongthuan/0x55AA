module layer_10_featuremap_5(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8ae84),
	.w1(32'hbc47c65f),
	.w2(32'hba7fedb6),
	.w3(32'h3b0da8d0),
	.w4(32'h3bdb4bdf),
	.w5(32'hb9afea56),
	.w6(32'h3ba1506c),
	.w7(32'h3c34e3c2),
	.w8(32'hbaca0044),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd709b1),
	.w1(32'h3c9158fa),
	.w2(32'hba02ebcb),
	.w3(32'h3b52ef1b),
	.w4(32'h3c86b09c),
	.w5(32'hbb49e303),
	.w6(32'hba8ea52a),
	.w7(32'hb8c425a8),
	.w8(32'hbab7e28e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7315da),
	.w1(32'hbb0b1a89),
	.w2(32'h3b98fc66),
	.w3(32'h3bf4dc52),
	.w4(32'hbb152b7a),
	.w5(32'h3b4f179c),
	.w6(32'hbb8a6296),
	.w7(32'hbbfc81b4),
	.w8(32'hbb1de816),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45a353),
	.w1(32'hbadfb047),
	.w2(32'h3b523ba3),
	.w3(32'h3a270b07),
	.w4(32'hba9bfc01),
	.w5(32'h3a8d2268),
	.w6(32'h3bb4cd23),
	.w7(32'h3b234b6d),
	.w8(32'hbb65543f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e5ad),
	.w1(32'h3bb35e79),
	.w2(32'hbc3c8e80),
	.w3(32'h3ba84a5a),
	.w4(32'h3b2f11db),
	.w5(32'hbc1f2b2b),
	.w6(32'hbb878f3e),
	.w7(32'hbb5f9df0),
	.w8(32'hbc488008),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd54b9e),
	.w1(32'hbb713b2a),
	.w2(32'h392de0e7),
	.w3(32'hbb6afe76),
	.w4(32'hbb9658b6),
	.w5(32'hba89b4d8),
	.w6(32'hbc573384),
	.w7(32'hbc433017),
	.w8(32'hbadeebb1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b05ce),
	.w1(32'h3964b69a),
	.w2(32'hbc07da4d),
	.w3(32'hba135b7d),
	.w4(32'hba120cda),
	.w5(32'hbbb8279a),
	.w6(32'h39ad9d85),
	.w7(32'h38bfe8b0),
	.w8(32'hb9a64900),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf714),
	.w1(32'h3bcba5c0),
	.w2(32'hbbc740a6),
	.w3(32'h3a8b03cc),
	.w4(32'h3c0b1e64),
	.w5(32'hbbba0180),
	.w6(32'hbafafd6c),
	.w7(32'hbb17cfd2),
	.w8(32'hbb94855f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34335c),
	.w1(32'h3b5ff190),
	.w2(32'h3c36d724),
	.w3(32'hbc024e66),
	.w4(32'hb949a9b9),
	.w5(32'h3c860be7),
	.w6(32'hbb94103b),
	.w7(32'hbaed8cb1),
	.w8(32'h3c882934),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0ab6a),
	.w1(32'hbca9eb62),
	.w2(32'h3969a9bf),
	.w3(32'hbb033096),
	.w4(32'hbc8ac15b),
	.w5(32'h3bbd5d7e),
	.w6(32'h3c4074b2),
	.w7(32'h3aa4995c),
	.w8(32'h3bd50b4c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb269cb1),
	.w1(32'hbc0f2e9a),
	.w2(32'h3a1cc027),
	.w3(32'h3af03252),
	.w4(32'hbc0fa57e),
	.w5(32'hbb1709a0),
	.w6(32'h3bb9a76c),
	.w7(32'hb8d991c9),
	.w8(32'hbb97d9ab),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab73a73),
	.w1(32'hbc0aed43),
	.w2(32'hbbdd0ec7),
	.w3(32'hb8f943b2),
	.w4(32'h3bae03bf),
	.w5(32'hbc36eb98),
	.w6(32'h3bff1517),
	.w7(32'h3aa9fc9f),
	.w8(32'hbc1b4951),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee54e6),
	.w1(32'h3b0e44d3),
	.w2(32'hbb254e6b),
	.w3(32'hbc580a6b),
	.w4(32'h391a6d7d),
	.w5(32'hba93db06),
	.w6(32'hbc46dd21),
	.w7(32'hbb0f03ec),
	.w8(32'hbb4b3706),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1407d5),
	.w1(32'h3b32ad02),
	.w2(32'hbbef3338),
	.w3(32'hbabc2595),
	.w4(32'h3afae4d7),
	.w5(32'hbbb7bab4),
	.w6(32'hbbafcbb4),
	.w7(32'h3a8f6a89),
	.w8(32'hb983013f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390496c9),
	.w1(32'hb9f54855),
	.w2(32'hba9cce0c),
	.w3(32'hbbce763d),
	.w4(32'hbc04d874),
	.w5(32'h3a9bf680),
	.w6(32'hbb804de9),
	.w7(32'hbbac6f66),
	.w8(32'hbbb64a42),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96c526),
	.w1(32'hbb160f3d),
	.w2(32'h38bc8c61),
	.w3(32'h3b641463),
	.w4(32'h3bbad809),
	.w5(32'h3b78c2a1),
	.w6(32'hbaa18907),
	.w7(32'h3bc0870a),
	.w8(32'h3bab36f4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9498363),
	.w1(32'hbb8f6004),
	.w2(32'hba2799c5),
	.w3(32'h3ae845a4),
	.w4(32'hbb872851),
	.w5(32'hbb2f8519),
	.w6(32'h3b94f078),
	.w7(32'h3abb330e),
	.w8(32'hbb19a3d6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf41bf4),
	.w1(32'hbb7d85b3),
	.w2(32'hbc05c995),
	.w3(32'hbb97ac36),
	.w4(32'hbb115d5b),
	.w5(32'hbbc184c1),
	.w6(32'h3b94263f),
	.w7(32'h3b03ace8),
	.w8(32'hbba812a0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315295),
	.w1(32'hbaf21502),
	.w2(32'hbb29d6ce),
	.w3(32'hbb9da00a),
	.w4(32'h38cb93b7),
	.w5(32'h3b16d7e8),
	.w6(32'hbb36c596),
	.w7(32'h3a400ccd),
	.w8(32'hba00592e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0dbe5),
	.w1(32'hbc381177),
	.w2(32'hb91a5944),
	.w3(32'hba1eeb41),
	.w4(32'hbc256743),
	.w5(32'hbb9b9070),
	.w6(32'hb96c829c),
	.w7(32'hbb0f7167),
	.w8(32'hbb7f9ec7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9208d7),
	.w1(32'h3bff2013),
	.w2(32'h3915e6c5),
	.w3(32'h3b50ab02),
	.w4(32'h3c05c25d),
	.w5(32'h3b835476),
	.w6(32'hbbb61a79),
	.w7(32'hbad5ff9a),
	.w8(32'hbb12bbef),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca959),
	.w1(32'hba95f0fc),
	.w2(32'h3a514982),
	.w3(32'hbb814877),
	.w4(32'hbb9e8883),
	.w5(32'hbb0386c5),
	.w6(32'hb91b48c6),
	.w7(32'h3b32214c),
	.w8(32'h3b6d4ca1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b78fb),
	.w1(32'h3b20ef26),
	.w2(32'hbc73f6ad),
	.w3(32'hbbc90b15),
	.w4(32'h3b9d8cb7),
	.w5(32'hbc960d26),
	.w6(32'hba946cc8),
	.w7(32'h3c27b988),
	.w8(32'hbc1434f8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcaeff),
	.w1(32'h3bc03b0c),
	.w2(32'h3ba7ec70),
	.w3(32'hbbd74ffe),
	.w4(32'h3b840463),
	.w5(32'h3b934fbc),
	.w6(32'hbb9cf036),
	.w7(32'h3b86c8a6),
	.w8(32'h39e6fb98),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bce63),
	.w1(32'h3bf57174),
	.w2(32'h3abf2197),
	.w3(32'hba7988ba),
	.w4(32'h3bb7fa44),
	.w5(32'h3b9c5437),
	.w6(32'hbb56ecfb),
	.w7(32'h3a7c4456),
	.w8(32'h3c167734),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badf3c0),
	.w1(32'h3bdbcbb7),
	.w2(32'h3bc6e03f),
	.w3(32'hb9c820e7),
	.w4(32'h3be3d546),
	.w5(32'h3b5136a9),
	.w6(32'h3aa95b44),
	.w7(32'h3bbbc431),
	.w8(32'h3c07330b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545b1e),
	.w1(32'hba5c2836),
	.w2(32'hbb92872c),
	.w3(32'h3bc003ec),
	.w4(32'hbafe632a),
	.w5(32'hbab9d283),
	.w6(32'h3b34bf9a),
	.w7(32'hbb3cef32),
	.w8(32'hbb25de36),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31996a),
	.w1(32'h37400244),
	.w2(32'h3cac0ce1),
	.w3(32'h3ad6bb5b),
	.w4(32'h3b408ae4),
	.w5(32'h3c9d4d7b),
	.w6(32'hba9181d5),
	.w7(32'hb93e98fa),
	.w8(32'h3c6530e3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2fc03),
	.w1(32'h3bfe7b14),
	.w2(32'hbaa6af13),
	.w3(32'h3c81b6c2),
	.w4(32'h3aa048a1),
	.w5(32'hbbba2dd3),
	.w6(32'h3bf6e136),
	.w7(32'hbbef3d61),
	.w8(32'h3afe895b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf53cc8),
	.w1(32'hba3a34d1),
	.w2(32'hbc114ef1),
	.w3(32'hbc1e017f),
	.w4(32'h3a52c092),
	.w5(32'h3c64ec99),
	.w6(32'hbc01a37d),
	.w7(32'hbb226f21),
	.w8(32'h3b4c7bdb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09767c),
	.w1(32'h3b06492e),
	.w2(32'h3aab1080),
	.w3(32'h3d370a6e),
	.w4(32'h3d105882),
	.w5(32'h3bb6a8f6),
	.w6(32'h3cfd203e),
	.w7(32'h3cbc79f6),
	.w8(32'h3bdb36e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bb3b5),
	.w1(32'h3be7f078),
	.w2(32'h3acbbcac),
	.w3(32'h3badd05f),
	.w4(32'h3b7c0d24),
	.w5(32'h3c0ee1a0),
	.w6(32'h3c1cb7c7),
	.w7(32'h3c1db418),
	.w8(32'h3c5e7aa6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf39c2),
	.w1(32'h393a4946),
	.w2(32'hbd18cede),
	.w3(32'h3c0839d5),
	.w4(32'h3bbc556d),
	.w5(32'hbc9b291e),
	.w6(32'h3c96b820),
	.w7(32'h3c37b33f),
	.w8(32'hbceb6122),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb49bc6),
	.w1(32'hbcf399d3),
	.w2(32'hbbaef755),
	.w3(32'h3b81493f),
	.w4(32'hbbe15f00),
	.w5(32'hbb4b50be),
	.w6(32'hbc0d7564),
	.w7(32'hbc9abc0a),
	.w8(32'hbb434796),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30fb25),
	.w1(32'hbc4f751f),
	.w2(32'h3a6fb5b4),
	.w3(32'hbbf89704),
	.w4(32'hbba68204),
	.w5(32'hbc84906e),
	.w6(32'hba8138e5),
	.w7(32'hbbb1a063),
	.w8(32'hbc1b67ec),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ead7b),
	.w1(32'hbc27d4b4),
	.w2(32'h3843d6fe),
	.w3(32'hbd2176b3),
	.w4(32'hbd077c4e),
	.w5(32'h3aac74a1),
	.w6(32'hbce114ae),
	.w7(32'hbcb2e42c),
	.w8(32'h3bc85bc8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a45bb),
	.w1(32'hbbad74ce),
	.w2(32'hbcbc24c2),
	.w3(32'hbc30fd21),
	.w4(32'hbc12f0c7),
	.w5(32'hbc978c2a),
	.w6(32'hbbb12227),
	.w7(32'hba9497d7),
	.w8(32'hbce3dac5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a88d5),
	.w1(32'hbc81c066),
	.w2(32'h3c1f7d2a),
	.w3(32'hbc3b7b6b),
	.w4(32'hbc51815b),
	.w5(32'h3b80ad39),
	.w6(32'hbce89c34),
	.w7(32'hbcdfaca0),
	.w8(32'hba4b54cc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fc166),
	.w1(32'h3c2c768d),
	.w2(32'h3c4684ee),
	.w3(32'h3a79bb53),
	.w4(32'h3bdd0dd3),
	.w5(32'h3b98ac3d),
	.w6(32'hbb7f291a),
	.w7(32'h3a5613d7),
	.w8(32'h3bbfacad),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f53b),
	.w1(32'h3be12634),
	.w2(32'h39804a0c),
	.w3(32'h3b20f753),
	.w4(32'hbb62522e),
	.w5(32'h3b0e2d68),
	.w6(32'hb999b5a7),
	.w7(32'hbb635b86),
	.w8(32'h3b07c4e7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1417d0),
	.w1(32'h3abd9c14),
	.w2(32'hbbb72a32),
	.w3(32'h3ab17549),
	.w4(32'h3bc6b7ff),
	.w5(32'hbbc2ea00),
	.w6(32'h3ba2a395),
	.w7(32'h3bbf7a10),
	.w8(32'hba3de0c9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c5daf),
	.w1(32'hbbbdf2d0),
	.w2(32'h3aa39356),
	.w3(32'hba772bf6),
	.w4(32'hbb8ee151),
	.w5(32'h3adb651e),
	.w6(32'h3a205267),
	.w7(32'h3a193f3c),
	.w8(32'h3b613e35),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba715b1),
	.w1(32'h3bf2f7b5),
	.w2(32'h3c3a65fa),
	.w3(32'h3bb940f2),
	.w4(32'h3ab5d3f6),
	.w5(32'hbc72c9f0),
	.w6(32'h3b42a502),
	.w7(32'h3b6cfa31),
	.w8(32'hbb33d5ad),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d587c),
	.w1(32'hbb8b5718),
	.w2(32'hbb3eff71),
	.w3(32'hbd452358),
	.w4(32'hbd1523db),
	.w5(32'hbb5e903d),
	.w6(32'hbcf7adc3),
	.w7(32'hbc9666b4),
	.w8(32'hbb9d4f60),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb066592),
	.w1(32'h3aa13262),
	.w2(32'hba5767c8),
	.w3(32'h3b5f01b6),
	.w4(32'h3bbf4f9a),
	.w5(32'h3ab2d48b),
	.w6(32'hbb632a9b),
	.w7(32'h3b077be5),
	.w8(32'h3a3a3a77),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407e28),
	.w1(32'h3b76764e),
	.w2(32'h3bbe1c53),
	.w3(32'hbbc6498a),
	.w4(32'hbbbd4025),
	.w5(32'h3baa3f96),
	.w6(32'hbbaf54ac),
	.w7(32'hbbb02c22),
	.w8(32'h3bd33757),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10309d),
	.w1(32'h3b980f29),
	.w2(32'h3985b6d9),
	.w3(32'h3c5cb1f0),
	.w4(32'h3c196ec1),
	.w5(32'h3a29cbc9),
	.w6(32'h3bc0ed37),
	.w7(32'h3c0ae526),
	.w8(32'hbb28c093),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5776fa),
	.w1(32'hbc82e204),
	.w2(32'hbc5c3212),
	.w3(32'hbbb220e0),
	.w4(32'hbc1719d7),
	.w5(32'hbd2cef3f),
	.w6(32'h3be51460),
	.w7(32'h39ab5613),
	.w8(32'hbcd9241d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01b55a),
	.w1(32'hbcc5392f),
	.w2(32'h3c046268),
	.w3(32'hbd9b5175),
	.w4(32'hbd81b07b),
	.w5(32'h3bda0c12),
	.w6(32'hbd7f6caa),
	.w7(32'hbd51b357),
	.w8(32'h3b97a4a6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a7475),
	.w1(32'h3b8cf8e5),
	.w2(32'hbb70012b),
	.w3(32'h3be07376),
	.w4(32'h3c1fcb38),
	.w5(32'hbbcdacb6),
	.w6(32'h3bc53c0f),
	.w7(32'h3c014318),
	.w8(32'hbb2f451d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93bc8c),
	.w1(32'hba6e8f72),
	.w2(32'h3a8f87b0),
	.w3(32'hbbf053c5),
	.w4(32'hb89e7d7c),
	.w5(32'h3ac32080),
	.w6(32'h3b36c3ce),
	.w7(32'h393d77dc),
	.w8(32'h3b4aac62),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be7937),
	.w1(32'h3b00b182),
	.w2(32'hbab60f81),
	.w3(32'h3c23abc8),
	.w4(32'h3b90e38f),
	.w5(32'hbb10ab89),
	.w6(32'h3b9c442f),
	.w7(32'h3906aad0),
	.w8(32'h3b1d59ce),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51f914),
	.w1(32'h388c9e45),
	.w2(32'hbb70d50f),
	.w3(32'hba5a3131),
	.w4(32'hbbc4dca0),
	.w5(32'h3add479e),
	.w6(32'h3b89ffd2),
	.w7(32'hbb394e8f),
	.w8(32'h3a654495),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20624f),
	.w1(32'hbc0a950f),
	.w2(32'h3a5fb029),
	.w3(32'h3b1020fe),
	.w4(32'h3966f503),
	.w5(32'h3a54b3e1),
	.w6(32'h3b801d5c),
	.w7(32'h3b8ac9d9),
	.w8(32'hbab976ff),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60645c),
	.w1(32'h3bf4ebfb),
	.w2(32'hbc4395f3),
	.w3(32'h3bf0cafd),
	.w4(32'h3c64e697),
	.w5(32'hbc413d14),
	.w6(32'h3b4f5cc1),
	.w7(32'h3b8ce8f0),
	.w8(32'hbc058ca3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c61cd),
	.w1(32'hbbb88136),
	.w2(32'h3acb4556),
	.w3(32'hbc16cf2a),
	.w4(32'hbc220bdd),
	.w5(32'h3b8a6119),
	.w6(32'hbc0dae72),
	.w7(32'hbaef966f),
	.w8(32'h3c16561a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baafaf8),
	.w1(32'h3b84715b),
	.w2(32'h3cbf2cbf),
	.w3(32'h3bc5d1d4),
	.w4(32'hba832e64),
	.w5(32'h3c8ffb58),
	.w6(32'h3c1897bd),
	.w7(32'h3be9bf6b),
	.w8(32'h3c6dc8fa),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab1105),
	.w1(32'h3c572581),
	.w2(32'h3b47c86a),
	.w3(32'h3c8055ee),
	.w4(32'h3b4522fe),
	.w5(32'h3b606968),
	.w6(32'h3c25b8da),
	.w7(32'h3a8f6344),
	.w8(32'h3b7714f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b925996),
	.w1(32'h3bb6c93c),
	.w2(32'h3c264875),
	.w3(32'h3bb0428d),
	.w4(32'h3be1ede0),
	.w5(32'h3bdc4715),
	.w6(32'h3b71aa7d),
	.w7(32'h3ba81df4),
	.w8(32'h3b020d04),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a42b7),
	.w1(32'h3c3e5146),
	.w2(32'h3c16530b),
	.w3(32'h3c678721),
	.w4(32'h3c1d89db),
	.w5(32'h3b2fc4e8),
	.w6(32'h3b166dac),
	.w7(32'h3a850108),
	.w8(32'h3ab5bcb1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189951),
	.w1(32'h3bc5c7f3),
	.w2(32'hbb37004c),
	.w3(32'hba9d704a),
	.w4(32'h3b4516dd),
	.w5(32'hbb6b4940),
	.w6(32'h3b1983c2),
	.w7(32'h3b1b5093),
	.w8(32'hbb4bc2d2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b665c42),
	.w1(32'h3c070f7d),
	.w2(32'hbb893117),
	.w3(32'h3b13569b),
	.w4(32'h3c0817b8),
	.w5(32'h3ab0ce98),
	.w6(32'h3b535230),
	.w7(32'h39884fe8),
	.w8(32'hbb476b41),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b5cf),
	.w1(32'h3a3a1773),
	.w2(32'h3a488689),
	.w3(32'h3a432896),
	.w4(32'hba7e2abf),
	.w5(32'hbc2ae7ac),
	.w6(32'hb9ca4d80),
	.w7(32'hbb36a107),
	.w8(32'hb8f6a731),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b4630),
	.w1(32'h3ab8802b),
	.w2(32'hbad11412),
	.w3(32'hbc28c7dc),
	.w4(32'hbc198cdc),
	.w5(32'hb9558e05),
	.w6(32'h3b0daf85),
	.w7(32'h3b7a56ab),
	.w8(32'h3b605208),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f8c05),
	.w1(32'h3a7779d7),
	.w2(32'h3bba87dc),
	.w3(32'hbbb489ca),
	.w4(32'hbb81296d),
	.w5(32'h3c18fe70),
	.w6(32'h3a8b3a90),
	.w7(32'hbaf2d6b6),
	.w8(32'h3c3cf025),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4703cd),
	.w1(32'hbb79897e),
	.w2(32'hbbbaf108),
	.w3(32'h3b8197d6),
	.w4(32'hbb487171),
	.w5(32'hbc11cacd),
	.w6(32'h3bef9099),
	.w7(32'hb9fd0dc7),
	.w8(32'hbbe74aaf),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e7d0),
	.w1(32'hbc085290),
	.w2(32'hba2adc46),
	.w3(32'hbc2d2ae7),
	.w4(32'hbc371c90),
	.w5(32'hb8f3f584),
	.w6(32'hbc04c0a5),
	.w7(32'hbbb1babf),
	.w8(32'h3b9aa1ae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9939380),
	.w1(32'h3b1a8efb),
	.w2(32'h3ad76eb3),
	.w3(32'h3b0ac28b),
	.w4(32'h3b943e75),
	.w5(32'h3bcecfab),
	.w6(32'h3b8e17e7),
	.w7(32'h3bef985a),
	.w8(32'h3bf722b4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92d334),
	.w1(32'hb995f249),
	.w2(32'hbaf7b007),
	.w3(32'h37bd948a),
	.w4(32'h3b967fdb),
	.w5(32'hba1c045e),
	.w6(32'h3b1aaa51),
	.w7(32'h3bac276c),
	.w8(32'h3b0bc63f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219b18),
	.w1(32'h3c41e93c),
	.w2(32'h3c8c6abc),
	.w3(32'hbb52813e),
	.w4(32'h3c243dfd),
	.w5(32'h3c08403b),
	.w6(32'hbb72f0ee),
	.w7(32'h3c26fb14),
	.w8(32'h3c31d5d3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78a292),
	.w1(32'h3c5864ed),
	.w2(32'hbaf872df),
	.w3(32'h3c68bc0e),
	.w4(32'h3c39f960),
	.w5(32'h3aec3177),
	.w6(32'h3c7abd29),
	.w7(32'h3c4f3145),
	.w8(32'h3ad8138f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed4f1f),
	.w1(32'h3b9148aa),
	.w2(32'h3afd0274),
	.w3(32'h3c0e9aa4),
	.w4(32'h3b881417),
	.w5(32'h3b20e9a4),
	.w6(32'h3bb38dad),
	.w7(32'h3b25c553),
	.w8(32'hba033e9b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6bcc1),
	.w1(32'h3a52dbf0),
	.w2(32'hba34fef8),
	.w3(32'h3a4e8937),
	.w4(32'h3ba73bf7),
	.w5(32'h3a4eaf3d),
	.w6(32'hbb0f8a23),
	.w7(32'h3b2c64a5),
	.w8(32'hbacaae67),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8faa95),
	.w1(32'hbb305a0c),
	.w2(32'hbacbe1b8),
	.w3(32'hbbb67093),
	.w4(32'hbc03e658),
	.w5(32'hbc8e4968),
	.w6(32'hbc03d1be),
	.w7(32'hbba34827),
	.w8(32'hbc2a1100),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69b6af),
	.w1(32'hbc5c57fa),
	.w2(32'h3bf0a530),
	.w3(32'hbd181192),
	.w4(32'hbd0e138e),
	.w5(32'h3c1bb572),
	.w6(32'hbce4cf84),
	.w7(32'hbcd00457),
	.w8(32'h3c3c3984),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be26d),
	.w1(32'h3a55f048),
	.w2(32'hb9e85d29),
	.w3(32'h3c2a17ef),
	.w4(32'h3b938a4a),
	.w5(32'hbc0b4335),
	.w6(32'h3c742196),
	.w7(32'h3c2b965e),
	.w8(32'hbacf9c67),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b729),
	.w1(32'hbb6a890d),
	.w2(32'hbc426742),
	.w3(32'hbb980cdc),
	.w4(32'hbbbbfd02),
	.w5(32'hbb74d9cb),
	.w6(32'h3bb782d3),
	.w7(32'h3bdb058e),
	.w8(32'hbb87ed36),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c917ca),
	.w1(32'hbb3f3cbb),
	.w2(32'h3c260e11),
	.w3(32'hbab1e919),
	.w4(32'h3b749fa1),
	.w5(32'h3c24f5ce),
	.w6(32'hbb41b688),
	.w7(32'h3b30d79b),
	.w8(32'h3bf2f640),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b4be),
	.w1(32'h3b15ae82),
	.w2(32'hbbd579b9),
	.w3(32'h3c75843a),
	.w4(32'h3bfdad12),
	.w5(32'hb97098ed),
	.w6(32'h3bfaaf51),
	.w7(32'h3c0986b9),
	.w8(32'hbb9b5c37),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbe50),
	.w1(32'hbbba1aa7),
	.w2(32'hbb2887b4),
	.w3(32'h3882811a),
	.w4(32'h3b265648),
	.w5(32'hbb1231c1),
	.w6(32'hbb83b58b),
	.w7(32'hbb13e359),
	.w8(32'h3996823c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b4d68),
	.w1(32'hb9ff774b),
	.w2(32'hbcbdd9fc),
	.w3(32'h3b56cdea),
	.w4(32'h3b95702c),
	.w5(32'hbbf5a36f),
	.w6(32'h3b27193e),
	.w7(32'h3b751b0c),
	.w8(32'hbc3c7ac2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3afaf0),
	.w1(32'hbca470dd),
	.w2(32'hbc07f56f),
	.w3(32'h3c737a8c),
	.w4(32'h3afbff79),
	.w5(32'hbc4d239c),
	.w6(32'h3bf9d278),
	.w7(32'hba884213),
	.w8(32'hbc357d73),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58798d),
	.w1(32'hbb4fb7f7),
	.w2(32'h3b924cda),
	.w3(32'hbc322ea2),
	.w4(32'hbb54a719),
	.w5(32'h3ac70659),
	.w6(32'hbc49154f),
	.w7(32'hbaea4be0),
	.w8(32'hbac6dcec),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea274f),
	.w1(32'h3c345598),
	.w2(32'hbabda8fc),
	.w3(32'h3be4186a),
	.w4(32'h3c4ca533),
	.w5(32'h3b0477dd),
	.w6(32'h3af87288),
	.w7(32'h3c0cd60b),
	.w8(32'hba572a22),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb3458),
	.w1(32'hbb5f722b),
	.w2(32'hbb2d2dfd),
	.w3(32'h3b908fda),
	.w4(32'h3b243547),
	.w5(32'hb9818dd4),
	.w6(32'h3a919761),
	.w7(32'hbaf560fd),
	.w8(32'hbaf6cc84),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099896),
	.w1(32'h3902ac3e),
	.w2(32'h3b5175c6),
	.w3(32'h3b52752b),
	.w4(32'hbb67cb30),
	.w5(32'h3baeb215),
	.w6(32'h39a04d00),
	.w7(32'hbb885e3f),
	.w8(32'h3bb008f5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9d8d),
	.w1(32'hbacd28a7),
	.w2(32'h3ac5e271),
	.w3(32'h3b051e8a),
	.w4(32'hbb6d05cb),
	.w5(32'h38372a27),
	.w6(32'h3a3fed17),
	.w7(32'hbb00d5f0),
	.w8(32'hba85e5c1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42c659),
	.w1(32'h3af1ddb7),
	.w2(32'h39aebac9),
	.w3(32'hbb1cdacb),
	.w4(32'h3a381a7c),
	.w5(32'h3b31d1bf),
	.w6(32'hbae39d78),
	.w7(32'hba2cafaf),
	.w8(32'hbadda5f8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefbe5),
	.w1(32'h3ab5e3c2),
	.w2(32'h3be3aabe),
	.w3(32'hba95a345),
	.w4(32'h3b5ada2e),
	.w5(32'h3a1eed96),
	.w6(32'h3b1f82e3),
	.w7(32'h3a78b485),
	.w8(32'h3b720cf1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53725e),
	.w1(32'hb9ae94a0),
	.w2(32'hbb1ce955),
	.w3(32'hbb8ffb56),
	.w4(32'hba6e55d2),
	.w5(32'hbb21769e),
	.w6(32'hbb167576),
	.w7(32'hbb046c9c),
	.w8(32'h3c0b56e0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff1eb1),
	.w1(32'hbb566148),
	.w2(32'h3c579a67),
	.w3(32'hbc03847e),
	.w4(32'hbc223403),
	.w5(32'h3b135d0f),
	.w6(32'h3b5856d4),
	.w7(32'h3b64bd4a),
	.w8(32'h3b7cc202),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e860),
	.w1(32'h3bef226b),
	.w2(32'hbb7cb89c),
	.w3(32'hbc749cd0),
	.w4(32'hbc2a2339),
	.w5(32'hbbc22331),
	.w6(32'hbc05f36b),
	.w7(32'hbbe1add7),
	.w8(32'hbaaea64f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00bbd),
	.w1(32'h3b944149),
	.w2(32'h39091aa8),
	.w3(32'hbbe1f971),
	.w4(32'h3b06506b),
	.w5(32'hbb8e64f2),
	.w6(32'hbbc2057f),
	.w7(32'h3b2ab7f7),
	.w8(32'hbb14b475),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44e63),
	.w1(32'h38370fab),
	.w2(32'h3b85faa8),
	.w3(32'hbc008c0a),
	.w4(32'hbb6f6989),
	.w5(32'h3b05ce37),
	.w6(32'hbb3f0191),
	.w7(32'h3a9ac6af),
	.w8(32'h3ba0b499),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c275b),
	.w1(32'h3bb0a481),
	.w2(32'hbc018c52),
	.w3(32'hbaa7e2e4),
	.w4(32'h3a4c0b9c),
	.w5(32'hbc25a557),
	.w6(32'h3b22e185),
	.w7(32'h3aea7cfb),
	.w8(32'hbb82f31a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc625bba),
	.w1(32'hbbda200b),
	.w2(32'h3c7ceae9),
	.w3(32'hbc45d243),
	.w4(32'hbc133aba),
	.w5(32'h3c926b89),
	.w6(32'hbc7fc66d),
	.w7(32'hbba77483),
	.w8(32'h3c684cf9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85eb57),
	.w1(32'h3c0e3bdb),
	.w2(32'hbc117a14),
	.w3(32'h3c97d3f1),
	.w4(32'h3c5bddc9),
	.w5(32'h3968faa5),
	.w6(32'h3c2dcf7d),
	.w7(32'h3c3bca86),
	.w8(32'hbb4721a3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2ee8f),
	.w1(32'hbbde8c91),
	.w2(32'h395c1c6f),
	.w3(32'hbb380a51),
	.w4(32'hbbac03b1),
	.w5(32'h3c3f7108),
	.w6(32'hbbbc739d),
	.w7(32'hba105dff),
	.w8(32'h3c120cc5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99f426),
	.w1(32'h3be3d03b),
	.w2(32'hbbe53fc8),
	.w3(32'h3c44d5ce),
	.w4(32'h3c387e16),
	.w5(32'hbc7b3821),
	.w6(32'h3c8acb3d),
	.w7(32'h3c6b0dbe),
	.w8(32'hbc850009),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0965c5),
	.w1(32'h3997e061),
	.w2(32'hbbe0da6e),
	.w3(32'hbc731a4c),
	.w4(32'hbb22f90b),
	.w5(32'h3b4fc464),
	.w6(32'hbc511758),
	.w7(32'h3a39ec1f),
	.w8(32'hbba0852b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81c907),
	.w1(32'h3bfcb6da),
	.w2(32'hba01085a),
	.w3(32'h3c005df9),
	.w4(32'h3bcba99b),
	.w5(32'h39930056),
	.w6(32'h39e712a0),
	.w7(32'h3b2b8166),
	.w8(32'h3b58e07d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2ece9),
	.w1(32'hbb09f6a6),
	.w2(32'h3c27aa38),
	.w3(32'h37f34b9d),
	.w4(32'hbba8f0b6),
	.w5(32'h3c04faeb),
	.w6(32'hba4304ba),
	.w7(32'h3b284ba1),
	.w8(32'h3b9d2c5c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c208),
	.w1(32'hbb9af2c9),
	.w2(32'hbb9f4944),
	.w3(32'hba9b5c89),
	.w4(32'hbb506edd),
	.w5(32'hbaca53f1),
	.w6(32'hbafe3ebc),
	.w7(32'h3a738431),
	.w8(32'hba49e277),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b45d),
	.w1(32'hbb0413da),
	.w2(32'h3b517f45),
	.w3(32'h3b7c9fa6),
	.w4(32'h3b05c118),
	.w5(32'h3c25f876),
	.w6(32'h3b76925f),
	.w7(32'h3927fc23),
	.w8(32'h3bac380b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c248ea6),
	.w1(32'h3c081cea),
	.w2(32'hbb6ffa23),
	.w3(32'h3bd86a3b),
	.w4(32'h3be42701),
	.w5(32'hbb315947),
	.w6(32'h3c2ef854),
	.w7(32'h3c421866),
	.w8(32'hba4d1738),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f101a),
	.w1(32'h3a526493),
	.w2(32'h3c34ea9b),
	.w3(32'h3bc4d9b8),
	.w4(32'h3b801a3c),
	.w5(32'h3c7807f5),
	.w6(32'h3bba1f63),
	.w7(32'h3acb99bb),
	.w8(32'h3c83900e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0549da),
	.w1(32'h3b2eed3e),
	.w2(32'h3b4aeeaf),
	.w3(32'h3c4cd0ab),
	.w4(32'h3b389c8b),
	.w5(32'h3a2d2857),
	.w6(32'h3c61fadc),
	.w7(32'h3b6ae4a6),
	.w8(32'h3a65bc3f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0c607),
	.w1(32'h3b275d75),
	.w2(32'h3b5fe02a),
	.w3(32'h3bf00b27),
	.w4(32'h3be87ef8),
	.w5(32'h3bf88753),
	.w6(32'h3b56cf67),
	.w7(32'h3a8afd88),
	.w8(32'h3b4bd884),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b494cde),
	.w1(32'hbaaef0f7),
	.w2(32'h3b00bafa),
	.w3(32'h3b9217d6),
	.w4(32'h3a3e3746),
	.w5(32'h3bae525b),
	.w6(32'h3b988517),
	.w7(32'h3b6b4015),
	.w8(32'h3a21ca09),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96bcf7),
	.w1(32'h3bdb30b4),
	.w2(32'h3b6304f6),
	.w3(32'h3b88094b),
	.w4(32'h3b66de84),
	.w5(32'hbb004e86),
	.w6(32'h3bda013b),
	.w7(32'h3be248b9),
	.w8(32'h3b271889),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cb278),
	.w1(32'hbae19d5d),
	.w2(32'h3a1df396),
	.w3(32'hba308011),
	.w4(32'hbb5ff4a1),
	.w5(32'h3aae89ff),
	.w6(32'hbae8543f),
	.w7(32'hba9e320c),
	.w8(32'h3b1f75f1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9659),
	.w1(32'hbb2e5b32),
	.w2(32'hbae22d1f),
	.w3(32'hbafcee60),
	.w4(32'hb94535bb),
	.w5(32'h3b0806ce),
	.w6(32'h3ba48b95),
	.w7(32'h3b287d33),
	.w8(32'h3aa69ff9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b7f8),
	.w1(32'hbbc716a2),
	.w2(32'h3bbe3f3a),
	.w3(32'hbc260623),
	.w4(32'h3a757892),
	.w5(32'h3c0f458a),
	.w6(32'hbb427a33),
	.w7(32'h3c578bbd),
	.w8(32'h3c5ef941),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917f5f),
	.w1(32'h3bf89fac),
	.w2(32'hbc3739bb),
	.w3(32'h3c46e9b4),
	.w4(32'h3b94048b),
	.w5(32'hbbf06c01),
	.w6(32'h3c50b36d),
	.w7(32'h3c31bfce),
	.w8(32'hbaa010e9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb957671),
	.w1(32'hba2164c7),
	.w2(32'h3c08bf3f),
	.w3(32'hbaadec68),
	.w4(32'h3b87d0df),
	.w5(32'h3b5853b0),
	.w6(32'h3a147fe7),
	.w7(32'h3c05d5ef),
	.w8(32'hbba78bd0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b8a04),
	.w1(32'h3c19f996),
	.w2(32'hb9e0f341),
	.w3(32'h3b8ae5b6),
	.w4(32'h3ba7fa4a),
	.w5(32'h3c269257),
	.w6(32'hbbdec87b),
	.w7(32'hbbc953f2),
	.w8(32'h3c60315d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843168),
	.w1(32'hba8fe8b3),
	.w2(32'h3c0af398),
	.w3(32'h3c0c5d28),
	.w4(32'h3c122d98),
	.w5(32'hb99a383b),
	.w6(32'h3c7d16d7),
	.w7(32'h3c16092b),
	.w8(32'hbb069f59),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40ddf8),
	.w1(32'h3c1701e1),
	.w2(32'h3be9a5d2),
	.w3(32'h3b5d1d08),
	.w4(32'h3a68ac30),
	.w5(32'h3bb48422),
	.w6(32'hbb000d0f),
	.w7(32'hbb4fda53),
	.w8(32'h3b96787c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9922b),
	.w1(32'h3b3a6d4a),
	.w2(32'hbac6f3fb),
	.w3(32'h3ba22784),
	.w4(32'h3bff9ee6),
	.w5(32'h3a69d6ad),
	.w6(32'h3c3f2452),
	.w7(32'h3bcc6c81),
	.w8(32'hb8b795ad),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3273),
	.w1(32'hbaad2183),
	.w2(32'h3b914dcb),
	.w3(32'h3ba9525d),
	.w4(32'h393e125e),
	.w5(32'h3bfb8250),
	.w6(32'h39a74492),
	.w7(32'h3bd58f9f),
	.w8(32'h3c0ec2ab),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80194d),
	.w1(32'h3aac6fda),
	.w2(32'hbc4296b3),
	.w3(32'h3b1a76be),
	.w4(32'h3b378c30),
	.w5(32'hbc337b3f),
	.w6(32'h3b51f79b),
	.w7(32'h3b87dfc7),
	.w8(32'hbc31440a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a7518),
	.w1(32'hbc1ec123),
	.w2(32'h3c03b59a),
	.w3(32'hbc09c9bb),
	.w4(32'hbbe2c9cb),
	.w5(32'h3cb11d12),
	.w6(32'hbbc34066),
	.w7(32'hbb542668),
	.w8(32'h3c9a6615),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb44400),
	.w1(32'h3cba9c24),
	.w2(32'h3ba67b4e),
	.w3(32'h3d276547),
	.w4(32'h3d1cc186),
	.w5(32'h3b99e4fb),
	.w6(32'h3d0bccb2),
	.w7(32'h3d0295cc),
	.w8(32'h3c178cbe),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7c70b),
	.w1(32'h3c054d67),
	.w2(32'h3c445c3a),
	.w3(32'h3b8abdca),
	.w4(32'h3b7a9729),
	.w5(32'h3c1ff3cd),
	.w6(32'h3b768b8c),
	.w7(32'h3bda3d2b),
	.w8(32'h3bad08ad),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00381c),
	.w1(32'h3a08f88e),
	.w2(32'h3c70e4de),
	.w3(32'h3bba3346),
	.w4(32'hbb7d1916),
	.w5(32'h3c51ae69),
	.w6(32'hbb1790d2),
	.w7(32'hbc2105e1),
	.w8(32'h3bf629d5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27f6c4),
	.w1(32'h3c420b7d),
	.w2(32'hbb8c9ac1),
	.w3(32'h3c3d4227),
	.w4(32'h3c80ceea),
	.w5(32'hbbb62947),
	.w6(32'h3c2b7a1d),
	.w7(32'h3c5f5d9f),
	.w8(32'hbbca98bf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1fbd),
	.w1(32'hbab02d18),
	.w2(32'hbb9ba8ce),
	.w3(32'h3b63ba91),
	.w4(32'h3b8fe5ee),
	.w5(32'hbb40827c),
	.w6(32'hbb38d132),
	.w7(32'h3b70f414),
	.w8(32'hbb067375),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99e8a9),
	.w1(32'hbbedf3a7),
	.w2(32'hbbcf455e),
	.w3(32'h3b3f95d5),
	.w4(32'hbb167f75),
	.w5(32'hbb245bce),
	.w6(32'h3b4a0e9b),
	.w7(32'hb9882e96),
	.w8(32'hbb878ab6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945117),
	.w1(32'hbbadfcf1),
	.w2(32'h3b7caa81),
	.w3(32'hbadfb9ee),
	.w4(32'hbbc19835),
	.w5(32'h3b1a3e06),
	.w6(32'hbc06177a),
	.w7(32'hbc1db848),
	.w8(32'h3af17b3d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3e129),
	.w1(32'h3b8305ac),
	.w2(32'hba837427),
	.w3(32'hba91546c),
	.w4(32'h3adadccf),
	.w5(32'hba8313c8),
	.w6(32'h3b699be7),
	.w7(32'h391b8733),
	.w8(32'hbbd9857f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfd472),
	.w1(32'hbaaa8091),
	.w2(32'hb9aaf47d),
	.w3(32'hbc2cc862),
	.w4(32'hbc33e9c3),
	.w5(32'hbb49e2f8),
	.w6(32'hbc24aa8d),
	.w7(32'hbba25ea1),
	.w8(32'h3b5ccf83),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00bd7f),
	.w1(32'hbab5786a),
	.w2(32'h3bfec269),
	.w3(32'h3b969160),
	.w4(32'hbad49981),
	.w5(32'h3c16032d),
	.w6(32'h3afc5d8a),
	.w7(32'h3aaeabc8),
	.w8(32'h3b039ccc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a8fee),
	.w1(32'h3bd9e151),
	.w2(32'hbae49f6c),
	.w3(32'h3c1d925b),
	.w4(32'h3bcde423),
	.w5(32'hbae8c915),
	.w6(32'h3b941b85),
	.w7(32'h3b20b00c),
	.w8(32'hbc02192f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98dfcb),
	.w1(32'hbb924b40),
	.w2(32'h3c4abcd0),
	.w3(32'hbc586292),
	.w4(32'hbbf253b5),
	.w5(32'hbb1c7f5b),
	.w6(32'hbc43e86b),
	.w7(32'hbc2caa35),
	.w8(32'h3b800516),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9077e),
	.w1(32'hbbbd72c2),
	.w2(32'h3a2528fc),
	.w3(32'hbce5f65a),
	.w4(32'hbcce082b),
	.w5(32'hbb04de90),
	.w6(32'hbc2dcb45),
	.w7(32'hbc0515eb),
	.w8(32'h39d18a0c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becf29e),
	.w1(32'h3be69f6d),
	.w2(32'h3c2bbb23),
	.w3(32'h3c314fd2),
	.w4(32'h3bc794d8),
	.w5(32'h3c4a4d31),
	.w6(32'hba8b28fb),
	.w7(32'hbb086959),
	.w8(32'h3c73a7e9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec7cda),
	.w1(32'h389faf2d),
	.w2(32'h3bd6528c),
	.w3(32'h3c2861c1),
	.w4(32'h3b334941),
	.w5(32'h3c139aef),
	.w6(32'h3bcf1e4b),
	.w7(32'h3b4095c4),
	.w8(32'h3bb6239c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7918),
	.w1(32'h3b2b27b1),
	.w2(32'h3bb6995c),
	.w3(32'h3b1f271c),
	.w4(32'h3b58990c),
	.w5(32'h3cbf161d),
	.w6(32'h3c242ee0),
	.w7(32'h3bf28ac6),
	.w8(32'h3c994eb8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3db18),
	.w1(32'h3cb16a65),
	.w2(32'hba8b0738),
	.w3(32'h3d4a2ffe),
	.w4(32'h3d2cd12d),
	.w5(32'hba8001c8),
	.w6(32'h3d1f211c),
	.w7(32'h3d08f53a),
	.w8(32'h3b3a4cb9),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fbde7),
	.w1(32'h3a0bc9a4),
	.w2(32'hbb81e74f),
	.w3(32'hbad29ee5),
	.w4(32'h3b2cbcf6),
	.w5(32'hbc0d4384),
	.w6(32'hb9d68a94),
	.w7(32'hba86268d),
	.w8(32'hbbeb28dc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf63eee),
	.w1(32'hbbc008dd),
	.w2(32'hbc71ef25),
	.w3(32'hbc7c3907),
	.w4(32'hbc55d4d4),
	.w5(32'hbc45a729),
	.w6(32'hbc5d4b23),
	.w7(32'hbc42bbaa),
	.w8(32'hbc43ef63),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc887dc8),
	.w1(32'hbb15946c),
	.w2(32'h3b1b1320),
	.w3(32'hbca0b4c3),
	.w4(32'hbc15c2d8),
	.w5(32'h3b4b2a1c),
	.w6(32'hbc550d36),
	.w7(32'hbbb247cd),
	.w8(32'hbc13edbc),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aaa9c),
	.w1(32'hbb9e0875),
	.w2(32'hb9a7ab00),
	.w3(32'hbaead103),
	.w4(32'hbaf0364f),
	.w5(32'hbbc83191),
	.w6(32'hbba6b3dd),
	.w7(32'hbc01d6e0),
	.w8(32'hbbfee3be),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6e4e2),
	.w1(32'h3b0d8e0c),
	.w2(32'h3bc20367),
	.w3(32'hbb455af5),
	.w4(32'hbb29e542),
	.w5(32'h3c89feff),
	.w6(32'hbbd90d64),
	.w7(32'hbb326610),
	.w8(32'h3c4caddf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c812fb2),
	.w1(32'h3c507b20),
	.w2(32'h3c01a6db),
	.w3(32'h3d083a2c),
	.w4(32'h3cdefebd),
	.w5(32'h3b334d07),
	.w6(32'h3cd8d557),
	.w7(32'h3caec5fa),
	.w8(32'hba7bb994),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88fdce),
	.w1(32'h3b54ad0d),
	.w2(32'hbc0b6886),
	.w3(32'hba1bcabe),
	.w4(32'hba2703a9),
	.w5(32'hbc10116a),
	.w6(32'hbc0427fb),
	.w7(32'hbc2344d6),
	.w8(32'hbc0e5ef1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d7750),
	.w1(32'hbbb25654),
	.w2(32'hbbc4196a),
	.w3(32'hbc4997fe),
	.w4(32'hbc17c24f),
	.w5(32'hbb7e9e66),
	.w6(32'hbc3df715),
	.w7(32'hbb5ef055),
	.w8(32'hbacabd4b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b9e6f),
	.w1(32'h3910745a),
	.w2(32'h3bc34ca9),
	.w3(32'hba953e07),
	.w4(32'hbb853f91),
	.w5(32'h3b84187a),
	.w6(32'hbb11b04c),
	.w7(32'hb718291f),
	.w8(32'h3b3a4089),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b658dc7),
	.w1(32'h3aed7fef),
	.w2(32'hbb9c813e),
	.w3(32'h3b88e497),
	.w4(32'h3b18324e),
	.w5(32'h3933c7ba),
	.w6(32'h3b069aba),
	.w7(32'hba944ae7),
	.w8(32'hbbbf3a5f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1d781),
	.w1(32'hbbedd46a),
	.w2(32'hba3503e3),
	.w3(32'hbb84758c),
	.w4(32'hbb9f692b),
	.w5(32'h3a4e9e25),
	.w6(32'hbbc2dabd),
	.w7(32'hbb8c24e7),
	.w8(32'hba8aa886),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42f838),
	.w1(32'h39d51485),
	.w2(32'hbc8bd6c5),
	.w3(32'hba9d7424),
	.w4(32'h3ae81a17),
	.w5(32'hbb914424),
	.w6(32'hb8e3cb46),
	.w7(32'hbb1226da),
	.w8(32'hbc27688d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31c114),
	.w1(32'hbc5b9f8b),
	.w2(32'hbbed0b95),
	.w3(32'h3bddf109),
	.w4(32'h3ad41adb),
	.w5(32'hbc35d4fd),
	.w6(32'h3b97de0a),
	.w7(32'h3b4747cc),
	.w8(32'hbbc0bfd9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67bc10),
	.w1(32'hbad54751),
	.w2(32'h3ba3e875),
	.w3(32'hbc621661),
	.w4(32'hbc3bb12a),
	.w5(32'h3bcaad7f),
	.w6(32'hbc6f2670),
	.w7(32'hbb9f6a7f),
	.w8(32'h3bbea42f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c302968),
	.w1(32'h3c434398),
	.w2(32'hbba6a5a1),
	.w3(32'h3bf97dd1),
	.w4(32'h3c2ffdc6),
	.w5(32'hbb331771),
	.w6(32'hbafa503c),
	.w7(32'h3b4eb935),
	.w8(32'hbb0df7cc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c726f),
	.w1(32'hbbc8bbeb),
	.w2(32'h3883e205),
	.w3(32'h3a8aeff4),
	.w4(32'h39ff597f),
	.w5(32'h3a1c533f),
	.w6(32'h3950c0f6),
	.w7(32'hbaca7cfc),
	.w8(32'h3a4616dc),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe6333),
	.w1(32'h3ab17739),
	.w2(32'h39a49f3b),
	.w3(32'hba8ce7e5),
	.w4(32'h3accb3ad),
	.w5(32'h39f9e624),
	.w6(32'h3a8e431c),
	.w7(32'h3aea2bb8),
	.w8(32'h39cdcb0a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf834e2),
	.w1(32'h3ae3af89),
	.w2(32'h3b22cb12),
	.w3(32'h3b9aeedb),
	.w4(32'h3c1b6e4a),
	.w5(32'h3c491d43),
	.w6(32'hbbfaf015),
	.w7(32'hba24be56),
	.w8(32'h3b6dda59),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55286),
	.w1(32'h3c819f85),
	.w2(32'hbaa8d29b),
	.w3(32'hbced6b42),
	.w4(32'hbc0065a5),
	.w5(32'hb949567b),
	.w6(32'h3ba02c20),
	.w7(32'h3b9c3fab),
	.w8(32'h3bad3347),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c6407),
	.w1(32'hbb741669),
	.w2(32'hb9b01e6a),
	.w3(32'hbb0b3077),
	.w4(32'hbb926478),
	.w5(32'hba7a19ee),
	.w6(32'h3b76b49e),
	.w7(32'hba460b59),
	.w8(32'hbc006a6a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d8c9f),
	.w1(32'hbb4b1e15),
	.w2(32'hbc00ed2d),
	.w3(32'h3c025426),
	.w4(32'hbc8b3f1f),
	.w5(32'hb9f5e251),
	.w6(32'h3c822613),
	.w7(32'h3a953c30),
	.w8(32'h3b6c87cf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91bf7a),
	.w1(32'hbba0308c),
	.w2(32'h3b454cde),
	.w3(32'hbc8f3667),
	.w4(32'hbc9869b4),
	.w5(32'h3aa1a892),
	.w6(32'h3c42d711),
	.w7(32'hbb7125a6),
	.w8(32'h3b3f6af6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad14708),
	.w1(32'hb94653bc),
	.w2(32'hba96a918),
	.w3(32'h39f5be26),
	.w4(32'hbb1cddc5),
	.w5(32'h3be9b600),
	.w6(32'h3b1db6dc),
	.w7(32'hbae244c2),
	.w8(32'h3b22b5bd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fa007),
	.w1(32'h3cd30b58),
	.w2(32'hb9c3aae6),
	.w3(32'hbc2441e1),
	.w4(32'h3cca90a0),
	.w5(32'hbb8ac923),
	.w6(32'hbca73f8a),
	.w7(32'hbbd6e5dc),
	.w8(32'hbb58a045),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb731f35),
	.w1(32'hbb51fdf8),
	.w2(32'hbc448335),
	.w3(32'hbb6b1225),
	.w4(32'hbb0f01d1),
	.w5(32'h3d0c2392),
	.w6(32'hbb18e75b),
	.w7(32'hba06d3a7),
	.w8(32'h3c872bcb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1cbfc4),
	.w1(32'h3be44e83),
	.w2(32'h3c1388c2),
	.w3(32'h3c1c6d3a),
	.w4(32'hbc3e6a7a),
	.w5(32'h3b1e5392),
	.w6(32'h3caf1f13),
	.w7(32'hbbd9492d),
	.w8(32'h3a975e15),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b389c98),
	.w1(32'h3952ca01),
	.w2(32'hbb367226),
	.w3(32'hbb250918),
	.w4(32'hbbb54f95),
	.w5(32'hbb7c96e6),
	.w6(32'hbb65264d),
	.w7(32'hbbb1fc13),
	.w8(32'hbbc829ca),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b989d),
	.w1(32'hbbf17226),
	.w2(32'hbc19e956),
	.w3(32'hb83f719a),
	.w4(32'h3c94db34),
	.w5(32'hbc452afb),
	.w6(32'hbb146bdb),
	.w7(32'h3a0dc7e6),
	.w8(32'hbbaa4332),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d608b),
	.w1(32'h3c8fe048),
	.w2(32'h3ac41f2e),
	.w3(32'hbc834b45),
	.w4(32'h3c109cdc),
	.w5(32'hbb195656),
	.w6(32'hbcc925fe),
	.w7(32'h3a12db57),
	.w8(32'hbb58ece6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9d22),
	.w1(32'hba3b6b4f),
	.w2(32'hbb18c895),
	.w3(32'hbc2f6690),
	.w4(32'hbb2b33d3),
	.w5(32'hbc6140a2),
	.w6(32'hbc2ae411),
	.w7(32'hbbcd1a1f),
	.w8(32'h3b281a8b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9bd54),
	.w1(32'hba54c098),
	.w2(32'hbb10068e),
	.w3(32'hbba7253a),
	.w4(32'h3bd42985),
	.w5(32'h3c5b7711),
	.w6(32'h3be2fa79),
	.w7(32'h3c4d2bfd),
	.w8(32'h3b980a52),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6944d8),
	.w1(32'hbbd50237),
	.w2(32'h3b1aaff4),
	.w3(32'hbc5680a2),
	.w4(32'hbc5ec739),
	.w5(32'h3b1cdcee),
	.w6(32'hbbd1235c),
	.w7(32'hbc1dc15c),
	.w8(32'hb9d5809a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98efe9),
	.w1(32'h3b6a3d49),
	.w2(32'h3b9247ee),
	.w3(32'h3b284904),
	.w4(32'h3b92c008),
	.w5(32'hbcff57cc),
	.w6(32'hbab40ca1),
	.w7(32'h3b1877f8),
	.w8(32'hbb8a6e9c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a9f16),
	.w1(32'h3ca48514),
	.w2(32'h3bbd9355),
	.w3(32'hbc730432),
	.w4(32'h3cbbda61),
	.w5(32'hbceedf44),
	.w6(32'hbd1305f7),
	.w7(32'hbb69e9b2),
	.w8(32'hbcd21a8b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d011325),
	.w1(32'h3cb445b8),
	.w2(32'h3b6b2b98),
	.w3(32'h3ac93b10),
	.w4(32'h3d04fc56),
	.w5(32'h3b11f03d),
	.w6(32'hbcac735b),
	.w7(32'h3c637a2f),
	.w8(32'h3b35deae),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed16f9),
	.w1(32'hbc0f911e),
	.w2(32'h3a3599fd),
	.w3(32'hbc6b7125),
	.w4(32'hbc496b7a),
	.w5(32'hbaae6b4e),
	.w6(32'h3bf9ebc2),
	.w7(32'hbc1400a4),
	.w8(32'hbbb618b1),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37ca70),
	.w1(32'hbbf53c47),
	.w2(32'h38e08706),
	.w3(32'hbb7c0802),
	.w4(32'hbc471558),
	.w5(32'h3aa3e5d3),
	.w6(32'h3c4933d9),
	.w7(32'hbb879c4a),
	.w8(32'hbb13f6b0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6b278),
	.w1(32'hbb25c097),
	.w2(32'h3b96e632),
	.w3(32'hba88298f),
	.w4(32'h3b608e82),
	.w5(32'hba856f49),
	.w6(32'hbb4a4f52),
	.w7(32'h3b5a7398),
	.w8(32'hbc4fc61e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc072a),
	.w1(32'hbbb7c067),
	.w2(32'hbc5653c0),
	.w3(32'h3ca83d49),
	.w4(32'hbc0325b7),
	.w5(32'hbc9a120d),
	.w6(32'hbbaa1e20),
	.w7(32'hbc1d4e97),
	.w8(32'h3b8c1e46),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2be728),
	.w1(32'h3c85552f),
	.w2(32'hbb5ad1e7),
	.w3(32'hbc94222d),
	.w4(32'h3cb817df),
	.w5(32'hbbcf70e1),
	.w6(32'hbd0c37c2),
	.w7(32'hbb9f3247),
	.w8(32'hbc48c8f0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c671a3b),
	.w1(32'h3b6c158d),
	.w2(32'hbc6200ec),
	.w3(32'h3c48b032),
	.w4(32'h3c871ae8),
	.w5(32'hbd09a756),
	.w6(32'hbc3e06ed),
	.w7(32'h3b978d6f),
	.w8(32'hbc531332),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81384d),
	.w1(32'h3c47ea09),
	.w2(32'h3bbaeede),
	.w3(32'hbcab7fe8),
	.w4(32'h3cc3c14e),
	.w5(32'hbaa3fc73),
	.w6(32'hbd219fa3),
	.w7(32'hbb3db9d7),
	.w8(32'hbbc61ae4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9259f),
	.w1(32'hbb17a147),
	.w2(32'h3bc0ebc1),
	.w3(32'h3bca58c1),
	.w4(32'hba4043e0),
	.w5(32'h3c5355e7),
	.w6(32'h3ba7b487),
	.w7(32'h3baecf27),
	.w8(32'h3b084ccc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4bdf62),
	.w1(32'h3b8b39a9),
	.w2(32'hba8249e0),
	.w3(32'h3a8f4a35),
	.w4(32'h3c2a4dcc),
	.w5(32'h3c2f024f),
	.w6(32'h3bd0d346),
	.w7(32'hbb0bafcf),
	.w8(32'h3c2a2581),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc812c14),
	.w1(32'hba254f47),
	.w2(32'h3b5b8f82),
	.w3(32'h3c2db9cd),
	.w4(32'hbc17cf22),
	.w5(32'hbc1f128a),
	.w6(32'h3d2a4ef2),
	.w7(32'h3c66eaad),
	.w8(32'hbb906b5a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bf670),
	.w1(32'h3bd0a630),
	.w2(32'hbb18df58),
	.w3(32'hbc89ae03),
	.w4(32'h3c413748),
	.w5(32'hbb828f00),
	.w6(32'hbc15829b),
	.w7(32'hbbf410a5),
	.w8(32'hbbc54be6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd27b56),
	.w1(32'hbc0a1115),
	.w2(32'hb9de0f96),
	.w3(32'h39d45f6b),
	.w4(32'hbb132759),
	.w5(32'hbb462e78),
	.w6(32'h3b2bf9fe),
	.w7(32'h3bd7d76c),
	.w8(32'h3b9645b7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd52c56),
	.w1(32'h398df229),
	.w2(32'h3b33ac1c),
	.w3(32'hbc146988),
	.w4(32'hbb8d7987),
	.w5(32'hbb52a14f),
	.w6(32'h356f2e10),
	.w7(32'h3b2053bc),
	.w8(32'hbbd8fd55),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c51d),
	.w1(32'hbb72f210),
	.w2(32'hb9e12197),
	.w3(32'hbba0606b),
	.w4(32'hbc314bfb),
	.w5(32'hbb2b85e5),
	.w6(32'h3bbc49d9),
	.w7(32'hbb57f288),
	.w8(32'h3bc3ecd0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace10b),
	.w1(32'h3bb554c1),
	.w2(32'h3bc7ed60),
	.w3(32'h3b95cc54),
	.w4(32'h3b97b935),
	.w5(32'h3bca8325),
	.w6(32'hbb9d4822),
	.w7(32'h3b506c26),
	.w8(32'h3b099249),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4290c9),
	.w1(32'h3b7a8859),
	.w2(32'hb9dc08f6),
	.w3(32'hbbdc9ef3),
	.w4(32'hbbcf3dc6),
	.w5(32'h3c14b1be),
	.w6(32'hbb9d86bd),
	.w7(32'hbb7b490e),
	.w8(32'h3aace1b9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1564a),
	.w1(32'hbb8e4543),
	.w2(32'h38d271d5),
	.w3(32'hbb91d1c2),
	.w4(32'h3a6870ef),
	.w5(32'hbae488f2),
	.w6(32'hba056537),
	.w7(32'h3bb3aada),
	.w8(32'hbb80bd5c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0899bf),
	.w1(32'hbae61d02),
	.w2(32'h3b88089c),
	.w3(32'hbb9f7fc8),
	.w4(32'hbb53b4ad),
	.w5(32'h3c0801f4),
	.w6(32'hb9b3e365),
	.w7(32'h3ba10595),
	.w8(32'hbbf430f7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f718),
	.w1(32'hbc39e549),
	.w2(32'hbbc07d32),
	.w3(32'h3c7bd15c),
	.w4(32'hbc25211e),
	.w5(32'hbc31930f),
	.w6(32'h3ce36308),
	.w7(32'h3c68bf99),
	.w8(32'hbbc6f23e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeca524),
	.w1(32'hbb04fdde),
	.w2(32'hbb031fdf),
	.w3(32'hbbc8ba46),
	.w4(32'hbb02b6f9),
	.w5(32'hba1982d2),
	.w6(32'hbb934c80),
	.w7(32'hba1ee57b),
	.w8(32'h3b827c6c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83dc5),
	.w1(32'h3b95846b),
	.w2(32'hbc44452a),
	.w3(32'h3a992b62),
	.w4(32'h3bbc5ddd),
	.w5(32'hbc516954),
	.w6(32'h3b6dcbce),
	.w7(32'h3bec8d19),
	.w8(32'h3c77d484),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808199),
	.w1(32'h3c18f905),
	.w2(32'hba3e3a20),
	.w3(32'hbcb4cbdd),
	.w4(32'h3afb0a2e),
	.w5(32'hbc52679d),
	.w6(32'hbc3669ae),
	.w7(32'hbbeeb87a),
	.w8(32'hbc5cfe96),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11d638),
	.w1(32'h3c232d04),
	.w2(32'hbaf39676),
	.w3(32'hba54d984),
	.w4(32'h3c84f23b),
	.w5(32'hbb19e646),
	.w6(32'hbccbbffd),
	.w7(32'hbb1d1b1f),
	.w8(32'hb9b755af),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc569),
	.w1(32'hbb8eee20),
	.w2(32'hbc7721b2),
	.w3(32'hbbc63df6),
	.w4(32'hbba29c40),
	.w5(32'hbb08a5b1),
	.w6(32'hb93b936e),
	.w7(32'hb9331d30),
	.w8(32'h3c2df704),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70aba5),
	.w1(32'h3bcccab4),
	.w2(32'h3b8114d1),
	.w3(32'hbbd8635d),
	.w4(32'h3c0d0f3b),
	.w5(32'hba44d662),
	.w6(32'hbacf34e5),
	.w7(32'hbac955af),
	.w8(32'h3c3e464e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be769ae),
	.w1(32'hb8e62291),
	.w2(32'h3a8a5c56),
	.w3(32'hb97470a5),
	.w4(32'h3b8a5c1b),
	.w5(32'hbac3c168),
	.w6(32'hbb2d3e62),
	.w7(32'hbb550a84),
	.w8(32'h3c2f3e7c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc395bdd),
	.w1(32'hbaaa3b34),
	.w2(32'hba1172b7),
	.w3(32'hbc4a7c2e),
	.w4(32'hbc36a897),
	.w5(32'hbbf14a27),
	.w6(32'h3cbacc62),
	.w7(32'h3b583714),
	.w8(32'hbd2865ae),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33fff5),
	.w1(32'hbc728a6b),
	.w2(32'h3ab02eff),
	.w3(32'h3d02500f),
	.w4(32'h3c8447ad),
	.w5(32'hbb244f55),
	.w6(32'hbce32e99),
	.w7(32'h3b610b14),
	.w8(32'hbb22103b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16d1bd),
	.w1(32'hbb59544f),
	.w2(32'hbb75af67),
	.w3(32'hbbe4d398),
	.w4(32'hbba6e235),
	.w5(32'hbbcf863f),
	.w6(32'hbbc3454d),
	.w7(32'hb8828e98),
	.w8(32'hbb9a5ee9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83107ff),
	.w1(32'hb9ef17a6),
	.w2(32'h3c3d6800),
	.w3(32'hbb1a6617),
	.w4(32'hba90c078),
	.w5(32'hbbb9e89a),
	.w6(32'hbbb531cb),
	.w7(32'hbb4a67d4),
	.w8(32'hbcf8c26f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c511e32),
	.w1(32'h3ba260c2),
	.w2(32'h3b412df7),
	.w3(32'h3cc2a9a8),
	.w4(32'h3cea6f3b),
	.w5(32'hbb8d153d),
	.w6(32'hbc55cb85),
	.w7(32'h3c9bb984),
	.w8(32'hbce4d686),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2415e),
	.w1(32'hbc1cf33a),
	.w2(32'hbb100db1),
	.w3(32'h3cc82b04),
	.w4(32'h3c8ccfbf),
	.w5(32'hbb706f60),
	.w6(32'hbc16faf9),
	.w7(32'h3c745b94),
	.w8(32'h3a88a29c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a9ac1),
	.w1(32'h3ba4e074),
	.w2(32'h3b49044c),
	.w3(32'hbc3ab9e3),
	.w4(32'hbb567280),
	.w5(32'h3b8b3fc5),
	.w6(32'h3b1218ef),
	.w7(32'h3ab73387),
	.w8(32'h3bac33d6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d857d0),
	.w1(32'h3b007fec),
	.w2(32'hbc232faf),
	.w3(32'hbaf29077),
	.w4(32'h3a8a2f2a),
	.w5(32'hbbbf6e93),
	.w6(32'h3aaec8fa),
	.w7(32'h3b23241d),
	.w8(32'h3b83ec1d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20d2ed),
	.w1(32'h39a1b8c4),
	.w2(32'hbbc84bfb),
	.w3(32'hbbd70507),
	.w4(32'hbab42f75),
	.w5(32'hbbe65c32),
	.w6(32'h3aba6d73),
	.w7(32'hbaf0f85b),
	.w8(32'h3b36c2f1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd645b2),
	.w1(32'hbbc10a3f),
	.w2(32'h3c6076b3),
	.w3(32'hbc0d0b76),
	.w4(32'hbbf17857),
	.w5(32'h3c941a36),
	.w6(32'hbb0e7bc2),
	.w7(32'hbb72fbd7),
	.w8(32'h3bb6a27e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a4c12),
	.w1(32'h3ba40ad5),
	.w2(32'hbab7b570),
	.w3(32'hbb0e372a),
	.w4(32'hbcaa90a0),
	.w5(32'h399a3501),
	.w6(32'h3c720c6c),
	.w7(32'hbc959242),
	.w8(32'hbab9b516),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc134e2a),
	.w1(32'hbc636018),
	.w2(32'hbb36c25d),
	.w3(32'h3b3bb9dc),
	.w4(32'hbc992ed1),
	.w5(32'h3bdf6f4d),
	.w6(32'h3bbc6397),
	.w7(32'hbbaaa016),
	.w8(32'hbb92d26d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb33d57),
	.w1(32'hbb7fddda),
	.w2(32'hbc087e61),
	.w3(32'hbc0e6861),
	.w4(32'hbc090ec6),
	.w5(32'hbc3f8b47),
	.w6(32'h3bea49dd),
	.w7(32'h3b9b7f43),
	.w8(32'h38f83484),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf18bc),
	.w1(32'h3b99666c),
	.w2(32'hbb95850d),
	.w3(32'hbc122b41),
	.w4(32'h3b9250c3),
	.w5(32'hbb7674c6),
	.w6(32'hbbedc8e9),
	.w7(32'hbbfffc3b),
	.w8(32'hbb865223),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9523c31),
	.w1(32'hbb2ff4c9),
	.w2(32'hbbeca59d),
	.w3(32'hbb3bd529),
	.w4(32'h3a9c664c),
	.w5(32'hbae7ec60),
	.w6(32'hba7ba5d5),
	.w7(32'h3a5fb946),
	.w8(32'hba960aef),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e7bd1),
	.w1(32'h3a21ba2e),
	.w2(32'hbbc5f6ee),
	.w3(32'hbadbcb2f),
	.w4(32'h3bae69b9),
	.w5(32'hbc9c7190),
	.w6(32'h3a94e236),
	.w7(32'h3b8ee9f2),
	.w8(32'hbc7ff777),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c213df6),
	.w1(32'h3c64b643),
	.w2(32'hbbc04b6d),
	.w3(32'hbbb47dbc),
	.w4(32'h3ce94ad0),
	.w5(32'h3a357151),
	.w6(32'hbd28e5d2),
	.w7(32'hbbdf2ecc),
	.w8(32'h3c2d6182),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc365ea8),
	.w1(32'hbc0220e5),
	.w2(32'h3b61dad9),
	.w3(32'hbacdbba5),
	.w4(32'h3b368ae7),
	.w5(32'hbc2d3488),
	.w6(32'h3c95b798),
	.w7(32'h3cc726c3),
	.w8(32'h3a3db041),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb593ec4),
	.w1(32'hbb9cf15f),
	.w2(32'hbaf3050f),
	.w3(32'hbc126edb),
	.w4(32'hbbc52e7a),
	.w5(32'hbb90eea8),
	.w6(32'hbc1f445e),
	.w7(32'hbb85cdb6),
	.w8(32'h3aecf157),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafa6b9),
	.w1(32'hbc505ea2),
	.w2(32'hbadfc5ce),
	.w3(32'hbb892e75),
	.w4(32'hbb242344),
	.w5(32'hbb9ac082),
	.w6(32'hbb55e5e4),
	.w7(32'hbaefc4a1),
	.w8(32'hbbc17981),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8c9ba),
	.w1(32'h3b309241),
	.w2(32'h3a2587da),
	.w3(32'hbbb6317f),
	.w4(32'hbb1e8a44),
	.w5(32'h3aa8dc51),
	.w6(32'hbb9218d4),
	.w7(32'h391db94f),
	.w8(32'hb9a80175),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf4d66),
	.w1(32'h3bd522a2),
	.w2(32'hbb19bcbf),
	.w3(32'hbaa142c7),
	.w4(32'h3bc2729b),
	.w5(32'hbc66d715),
	.w6(32'hbb1d7c37),
	.w7(32'h3b4611dc),
	.w8(32'hbc80d6ec),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd680c2),
	.w1(32'h3c0d28f0),
	.w2(32'h3c952bad),
	.w3(32'hbb5a643e),
	.w4(32'h3cb56663),
	.w5(32'hbc91cee1),
	.w6(32'hbce54619),
	.w7(32'hba5f1ad9),
	.w8(32'hbca8ceda),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6e329),
	.w1(32'hbc88c5b8),
	.w2(32'hbb06a1c8),
	.w3(32'h3cf87e72),
	.w4(32'h3caab338),
	.w5(32'h3b10b387),
	.w6(32'hbb76fd3a),
	.w7(32'h3c24491d),
	.w8(32'hbb957adb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565d52),
	.w1(32'h3bef6984),
	.w2(32'h3c4b37d0),
	.w3(32'h3b502bd4),
	.w4(32'hbbde014e),
	.w5(32'h3c3ee91c),
	.w6(32'h3ab39e98),
	.w7(32'hbbe55fc9),
	.w8(32'hbc049174),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b9b0bf),
	.w1(32'h3c157b6f),
	.w2(32'h3bc9f4c5),
	.w3(32'hbb08d8ec),
	.w4(32'hba0749e5),
	.w5(32'hbbb0047b),
	.w6(32'hbbd80fbf),
	.w7(32'hbb823e74),
	.w8(32'hbcb01e5b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dbd67),
	.w1(32'hbb78c0dd),
	.w2(32'h3b8b8f08),
	.w3(32'h3cb279bf),
	.w4(32'h3c2f5b6c),
	.w5(32'hbb20dc5f),
	.w6(32'hbafa4a2b),
	.w7(32'h3c130dfb),
	.w8(32'h3b457f8a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6640e5),
	.w1(32'hbb889529),
	.w2(32'h3b45cb09),
	.w3(32'hbb515cbd),
	.w4(32'h3af36022),
	.w5(32'h3ba7ecd7),
	.w6(32'hbbec282a),
	.w7(32'hbbc506e7),
	.w8(32'h3c0a840c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fefd3),
	.w1(32'hbccac175),
	.w2(32'h3c3b6c41),
	.w3(32'h3c6959f7),
	.w4(32'hbce10b5d),
	.w5(32'h38335669),
	.w6(32'h3cbf14fd),
	.w7(32'h3c3eb0d3),
	.w8(32'h3b89bf0d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc644c79),
	.w1(32'hbcda9283),
	.w2(32'hba884539),
	.w3(32'h3c95c3b5),
	.w4(32'hbc943eb5),
	.w5(32'hbb5a7c68),
	.w6(32'h3d12e9e6),
	.w7(32'h3c51b182),
	.w8(32'h3a9fba03),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa468dc),
	.w1(32'hbc0ff42b),
	.w2(32'hbc1e2957),
	.w3(32'h3b12a9df),
	.w4(32'hbb288932),
	.w5(32'hbaafbc1e),
	.w6(32'h3bfa311f),
	.w7(32'h3c80135c),
	.w8(32'h3b8a3061),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23cd4e),
	.w1(32'hbbcfd666),
	.w2(32'hbba04906),
	.w3(32'h3a44222b),
	.w4(32'hbb7bd346),
	.w5(32'hbc24a45a),
	.w6(32'h3c2086b7),
	.w7(32'h3be0cf63),
	.w8(32'h3c1d2c6a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9401a4),
	.w1(32'h3c35a146),
	.w2(32'hbb87a709),
	.w3(32'hbcac0eb4),
	.w4(32'h3b914cc1),
	.w5(32'h3a8dc701),
	.w6(32'hbc7bf4ee),
	.w7(32'hbb9e20bc),
	.w8(32'hbaba115e),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b7f7),
	.w1(32'hbaadced1),
	.w2(32'hbb8f722c),
	.w3(32'h3addd5b9),
	.w4(32'h3b28b0f6),
	.w5(32'hba869c04),
	.w6(32'hba38b168),
	.w7(32'hbb0ea372),
	.w8(32'h3be51ece),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba95952),
	.w1(32'hbabfbc94),
	.w2(32'h39382fe2),
	.w3(32'h396bdca8),
	.w4(32'h3b4f7911),
	.w5(32'hbba13144),
	.w6(32'hba3de0c4),
	.w7(32'h39f91564),
	.w8(32'h3bd01709),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf813a5),
	.w1(32'h39844dc1),
	.w2(32'hbc1416a1),
	.w3(32'hbc12c559),
	.w4(32'hbadcb2d7),
	.w5(32'h3bec1568),
	.w6(32'hbb139140),
	.w7(32'hbc1d38c6),
	.w8(32'h3bf1c56e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8c74),
	.w1(32'hbbb06908),
	.w2(32'h3bf44939),
	.w3(32'hbc2d7e56),
	.w4(32'h3be1f796),
	.w5(32'h3c231aa6),
	.w6(32'h3b8e25fe),
	.w7(32'h3c1b7602),
	.w8(32'h3b7ee101),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06cc25),
	.w1(32'hbc6f1e98),
	.w2(32'h3bb3e28e),
	.w3(32'h3c8b487a),
	.w4(32'hbc60d991),
	.w5(32'hbade490d),
	.w6(32'h3c9a70a9),
	.w7(32'h3c0afed0),
	.w8(32'hbb507ed3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3609c),
	.w1(32'h3b107905),
	.w2(32'hbc19a76c),
	.w3(32'hbbfdd8e2),
	.w4(32'h3a9f84e5),
	.w5(32'hbc01f0ed),
	.w6(32'hbc200c9b),
	.w7(32'hbaa0f703),
	.w8(32'h3c29a0ab),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06dad2),
	.w1(32'h3c6270ab),
	.w2(32'h3b1e1c7c),
	.w3(32'hbb9fe977),
	.w4(32'h3c16d935),
	.w5(32'h3c4adb30),
	.w6(32'hbc15447c),
	.w7(32'hbb071f5e),
	.w8(32'h3c7ef015),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf498c7),
	.w1(32'h3c7266b4),
	.w2(32'hb991d667),
	.w3(32'hbc8d57a3),
	.w4(32'h3c1e829f),
	.w5(32'h3bdd415a),
	.w6(32'hbc073db6),
	.w7(32'hbc57ebed),
	.w8(32'h3c2e70c7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c9a8),
	.w1(32'hbb2f83ff),
	.w2(32'hbbcff78e),
	.w3(32'hbc017cc5),
	.w4(32'hbc524912),
	.w5(32'h3b90e49e),
	.w6(32'h3c404997),
	.w7(32'hbc1815b8),
	.w8(32'hbc219628),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bc6b0),
	.w1(32'hbc195e62),
	.w2(32'hbb694961),
	.w3(32'h3c246a22),
	.w4(32'hb984c2d5),
	.w5(32'hbbd28727),
	.w6(32'h3b72e2a7),
	.w7(32'h3c1ac90d),
	.w8(32'hbbedddd3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e864c),
	.w1(32'hba2d942b),
	.w2(32'h3bacb4b4),
	.w3(32'hbbbe1a50),
	.w4(32'hbb3cc0ff),
	.w5(32'hbb8a4c2b),
	.w6(32'hbbca7194),
	.w7(32'hbaec02d8),
	.w8(32'hba87bc8c),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9219d16),
	.w1(32'h3a9b3f35),
	.w2(32'h3a725049),
	.w3(32'hba5131c0),
	.w4(32'h3ac5d1db),
	.w5(32'hbaf14339),
	.w6(32'h3b6d5339),
	.w7(32'h3b871146),
	.w8(32'h3b1168b3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869335b),
	.w1(32'hbb26be07),
	.w2(32'h3c0b2c39),
	.w3(32'hbb4d0054),
	.w4(32'hbbf89749),
	.w5(32'hbbb526df),
	.w6(32'h3bf9509f),
	.w7(32'h3b988c89),
	.w8(32'hbca1999b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b567a5e),
	.w1(32'hbc482ef3),
	.w2(32'h3bf3e361),
	.w3(32'h3c9b90c2),
	.w4(32'hbbcc80c7),
	.w5(32'h3c7eac14),
	.w6(32'h3c34b5da),
	.w7(32'h3c2bb578),
	.w8(32'h3c4dd580),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ee6da),
	.w1(32'hbcabcd31),
	.w2(32'h3b86fad2),
	.w3(32'h3c6d5fa8),
	.w4(32'hbd0c6bfb),
	.w5(32'h3b0333bb),
	.w6(32'h3ce9482b),
	.w7(32'h3b852484),
	.w8(32'h3a06a855),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192727),
	.w1(32'hbb0deda5),
	.w2(32'hbb713aaa),
	.w3(32'hbb136cdd),
	.w4(32'hbb746d5b),
	.w5(32'hbb818c6f),
	.w6(32'hbb56fce8),
	.w7(32'hbbd01c3b),
	.w8(32'h396f8b00),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba665e9),
	.w1(32'hbb8d67d3),
	.w2(32'hbb0147df),
	.w3(32'hbb5e5845),
	.w4(32'h39a2aff8),
	.w5(32'hbb3d8197),
	.w6(32'hbaa3a274),
	.w7(32'h3ae5e8af),
	.w8(32'h3adff07b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad25aa5),
	.w1(32'h3a022e58),
	.w2(32'hbb31ae72),
	.w3(32'hba7be426),
	.w4(32'hbaa17bab),
	.w5(32'h3c927d39),
	.w6(32'h3a1c8e5a),
	.w7(32'h3a1607f5),
	.w8(32'h3c36afee),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee309f),
	.w1(32'hbc1c1ef6),
	.w2(32'hbb0ae043),
	.w3(32'hbb9834f3),
	.w4(32'hbbe6d57d),
	.w5(32'h3ad69e71),
	.w6(32'h3c0e88a5),
	.w7(32'hbc10c961),
	.w8(32'h3bb7529e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3940fb3f),
	.w1(32'hbbe06f2d),
	.w2(32'h3b13fd6d),
	.w3(32'h3b4a073d),
	.w4(32'hbb730221),
	.w5(32'hbc42fb95),
	.w6(32'h3b4f4d89),
	.w7(32'h3aa9c6aa),
	.w8(32'hba82ae1d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6d2ca),
	.w1(32'h3c00367a),
	.w2(32'hbc0c08ca),
	.w3(32'hbc4cf608),
	.w4(32'h3c294a3d),
	.w5(32'hbc8a13bb),
	.w6(32'hbcbd0205),
	.w7(32'hbbbe65de),
	.w8(32'h3cb1678f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0d057),
	.w1(32'h3c8baeb2),
	.w2(32'hbbe8842f),
	.w3(32'hbcf1f9ec),
	.w4(32'h3ab3f91e),
	.w5(32'hbc01d1da),
	.w6(32'hbc1110ff),
	.w7(32'hbc95094f),
	.w8(32'h3c8334ab),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1691b),
	.w1(32'h3c1772b3),
	.w2(32'hbc1302ee),
	.w3(32'hbcd8fcdc),
	.w4(32'hbc05dfc6),
	.w5(32'hbc528d0f),
	.w6(32'hba5b730c),
	.w7(32'hbc06826c),
	.w8(32'h3b574bc2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule