module layer_10_featuremap_447(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2835fb),
	.w1(32'h3a8d6ba9),
	.w2(32'h3b58120c),
	.w3(32'hbbb4a775),
	.w4(32'hbb87c970),
	.w5(32'hbb68f2d2),
	.w6(32'hbbad5d3f),
	.w7(32'hbbc1d299),
	.w8(32'hbba8e9ba),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ead64),
	.w1(32'hba99e926),
	.w2(32'h3a24438b),
	.w3(32'hba44a7d5),
	.w4(32'hba751f48),
	.w5(32'hbbe88068),
	.w6(32'hbb645ceb),
	.w7(32'h3a4fdf40),
	.w8(32'hbc170393),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0def32),
	.w1(32'h3b2fc4ee),
	.w2(32'hbb9bd099),
	.w3(32'hbb1e9024),
	.w4(32'hbbb7c7ec),
	.w5(32'hbbb447bd),
	.w6(32'hbbb380be),
	.w7(32'hbb1bb4dc),
	.w8(32'hbbde39a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3a0d),
	.w1(32'h3b2c5683),
	.w2(32'h3b262a1a),
	.w3(32'hbc814943),
	.w4(32'h3bb1069c),
	.w5(32'hbc13ef31),
	.w6(32'hbc655e87),
	.w7(32'h3b4eff69),
	.w8(32'h3bc59213),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeda188),
	.w1(32'hbb9e57da),
	.w2(32'hbb041986),
	.w3(32'h3b0a31b6),
	.w4(32'hbb34ec5d),
	.w5(32'hbb67601b),
	.w6(32'h3a9f632a),
	.w7(32'hba08d79d),
	.w8(32'h3b5d7508),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a645a9a),
	.w1(32'hba8ed829),
	.w2(32'hbadc3fbb),
	.w3(32'hba49def2),
	.w4(32'h3ace343f),
	.w5(32'h3c261365),
	.w6(32'h3ab6b5e3),
	.w7(32'h3a51227c),
	.w8(32'h3bf3cf2d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d7da),
	.w1(32'hba7bd3b6),
	.w2(32'hbba9a757),
	.w3(32'h3ba9b1b6),
	.w4(32'hbb5909c7),
	.w5(32'h3c6b96a8),
	.w6(32'h3bc510e4),
	.w7(32'hbad50d80),
	.w8(32'hbb9389cc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6a32a),
	.w1(32'h3be1bd74),
	.w2(32'h3c0b7c0a),
	.w3(32'hbc2d712d),
	.w4(32'h3be5a860),
	.w5(32'h3cba8f83),
	.w6(32'hbc2d1394),
	.w7(32'h3bd0b5df),
	.w8(32'h3b91d514),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54c009),
	.w1(32'hbbfedbca),
	.w2(32'hbbefa7cf),
	.w3(32'h3b414ebb),
	.w4(32'hbbaf8b55),
	.w5(32'hbbe75d5f),
	.w6(32'h3b1ae782),
	.w7(32'h3b0d825d),
	.w8(32'hbaa6d67e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0c44f),
	.w1(32'h3b293a54),
	.w2(32'h3ad28429),
	.w3(32'hbbdf88d4),
	.w4(32'h3b117ace),
	.w5(32'hbc21d46d),
	.w6(32'hbc1b3087),
	.w7(32'h3aba6d35),
	.w8(32'h3bfb0f64),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76c6ef),
	.w1(32'hbb04a108),
	.w2(32'hbb80a6c3),
	.w3(32'hbacdb751),
	.w4(32'h3b5415c0),
	.w5(32'hbae96a38),
	.w6(32'hba88123a),
	.w7(32'h3b258d82),
	.w8(32'h3bb49ce6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a14d2),
	.w1(32'hbb200e41),
	.w2(32'h3aa5f959),
	.w3(32'hb9f9884d),
	.w4(32'hbc0df4e0),
	.w5(32'h3b4d5017),
	.w6(32'hbb60963c),
	.w7(32'hbc13816b),
	.w8(32'hbc2f3c15),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b600234),
	.w1(32'hbbb7a311),
	.w2(32'hbbee458a),
	.w3(32'hbb3195dd),
	.w4(32'hbb94556f),
	.w5(32'hbc8933f2),
	.w6(32'hbc2510f6),
	.w7(32'hbb6726ff),
	.w8(32'hbc64a219),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc33ea2),
	.w1(32'hbb540813),
	.w2(32'h3af2cf4b),
	.w3(32'hbadec914),
	.w4(32'hbbf50c96),
	.w5(32'hbc0e5457),
	.w6(32'hbb5ded93),
	.w7(32'hbb420cd7),
	.w8(32'hbbfc1b30),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba359338),
	.w1(32'h39fdadb1),
	.w2(32'hbab4cb83),
	.w3(32'h3a99e13f),
	.w4(32'h3bb14336),
	.w5(32'hbb087c77),
	.w6(32'hbb0f97b7),
	.w7(32'hbbcf0be0),
	.w8(32'h3b388e55),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a679b),
	.w1(32'h3b544e59),
	.w2(32'hbba1e48e),
	.w3(32'h3aa53f04),
	.w4(32'h3b7fa143),
	.w5(32'h3be1fb6c),
	.w6(32'h390081b4),
	.w7(32'hbb45d751),
	.w8(32'h3a2dd751),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a49db),
	.w1(32'hba07a323),
	.w2(32'hbb14c85f),
	.w3(32'hbb2e545e),
	.w4(32'h3b3cf49c),
	.w5(32'h3bc9176e),
	.w6(32'hbb5da667),
	.w7(32'hbbd0b020),
	.w8(32'hbad3bf76),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb803a1b),
	.w1(32'h3bf2e16e),
	.w2(32'h3ba9c540),
	.w3(32'hbb28fe85),
	.w4(32'hbbc8d49d),
	.w5(32'h3a2f98d1),
	.w6(32'hbb9b69bb),
	.w7(32'hbc2f0c66),
	.w8(32'hbbb3212a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40845e),
	.w1(32'hba35caaa),
	.w2(32'h3ad8ed2c),
	.w3(32'hbaa015ac),
	.w4(32'hbbb61d17),
	.w5(32'h3bb91f06),
	.w6(32'hbbb801fa),
	.w7(32'hbbefd553),
	.w8(32'hb99a8bb6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fe593),
	.w1(32'hbb1be547),
	.w2(32'hbb90efdc),
	.w3(32'hbbaacc62),
	.w4(32'hbaa5bb58),
	.w5(32'hbc48af16),
	.w6(32'hbc1397f5),
	.w7(32'h3b4b9533),
	.w8(32'hbc0f73f2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c29d1),
	.w1(32'h3b57f3d0),
	.w2(32'h3b5bec83),
	.w3(32'hbafc40da),
	.w4(32'h3b15374e),
	.w5(32'h3bca5b55),
	.w6(32'hbc11bd54),
	.w7(32'h3c3f7911),
	.w8(32'h3b7928eb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba713cb1),
	.w1(32'h3afa1ba2),
	.w2(32'hba9879b8),
	.w3(32'h3a4da80a),
	.w4(32'h3a12c927),
	.w5(32'h3c018cba),
	.w6(32'h3c326b1d),
	.w7(32'h3af39826),
	.w8(32'h3bd8e8b2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0aef1e),
	.w1(32'h3b6509e6),
	.w2(32'hbb004c5c),
	.w3(32'hbbca4bb5),
	.w4(32'hb99bd085),
	.w5(32'hbc264965),
	.w6(32'h3b1cfe6b),
	.w7(32'hbb9b2fcd),
	.w8(32'h3af9c546),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b251e05),
	.w1(32'h3b879bf5),
	.w2(32'h3c16044c),
	.w3(32'h3c22b94d),
	.w4(32'h3b9b870a),
	.w5(32'h3baf76b3),
	.w6(32'hb98294c1),
	.w7(32'hba91beba),
	.w8(32'h3b97afb4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e062),
	.w1(32'h3b9285b0),
	.w2(32'h3bcadc0d),
	.w3(32'h3b7dd0b8),
	.w4(32'hbbb0a732),
	.w5(32'h3841187c),
	.w6(32'h3b906e2f),
	.w7(32'h3aec099f),
	.w8(32'h3ba53d23),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9993b6),
	.w1(32'h3acda81b),
	.w2(32'h3a83e76b),
	.w3(32'hbbc25d65),
	.w4(32'h3c061529),
	.w5(32'hbba82d50),
	.w6(32'hbb306c55),
	.w7(32'h3c59ab2c),
	.w8(32'h3c4238d0),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c237711),
	.w1(32'h3a719b32),
	.w2(32'hbb0e9e9b),
	.w3(32'h3c8bf543),
	.w4(32'h39dc071b),
	.w5(32'h3bc0839c),
	.w6(32'h3c5a31b8),
	.w7(32'h3aba2f63),
	.w8(32'hbb83a279),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0354ef),
	.w1(32'hb9fdced4),
	.w2(32'hbac22a82),
	.w3(32'h39ae3581),
	.w4(32'h3b15a773),
	.w5(32'hbc11a05a),
	.w6(32'hbb620c1b),
	.w7(32'hbb240262),
	.w8(32'hbbb79490),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8046a1),
	.w1(32'h3b17d16d),
	.w2(32'hbba96bf9),
	.w3(32'hbae9608c),
	.w4(32'hbc0c7ec7),
	.w5(32'hbc46d58e),
	.w6(32'hbb788044),
	.w7(32'hbc5b200d),
	.w8(32'hbc429536),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c63b6),
	.w1(32'h3b4c301b),
	.w2(32'h382a72a7),
	.w3(32'hbc02a106),
	.w4(32'h3740da17),
	.w5(32'hbb6c8b49),
	.w6(32'hbb18500d),
	.w7(32'h3b74b0ee),
	.w8(32'h3b5d3c34),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85188f),
	.w1(32'hbb8b03c2),
	.w2(32'hbc1780fe),
	.w3(32'hbb8c721e),
	.w4(32'hb7b62d49),
	.w5(32'h3aca89bf),
	.w6(32'h3b9e0909),
	.w7(32'hbbb604a1),
	.w8(32'hbb2adf49),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64edc),
	.w1(32'h3baaf13d),
	.w2(32'hbb7f3bc9),
	.w3(32'hbbca21fb),
	.w4(32'h3a94e40e),
	.w5(32'hbb26e01a),
	.w6(32'hbb9c8bf4),
	.w7(32'hba76ac3a),
	.w8(32'h3af420d1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bec9),
	.w1(32'h3a24ffd2),
	.w2(32'hbb21da2c),
	.w3(32'hb630c28a),
	.w4(32'hbb0db793),
	.w5(32'h3b18b204),
	.w6(32'h3b44d94f),
	.w7(32'hb79a7f95),
	.w8(32'h3b7b86cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd233c9),
	.w1(32'hbb898cdd),
	.w2(32'hbb340a70),
	.w3(32'hbbf31087),
	.w4(32'h3b0dd4b9),
	.w5(32'h3bdb2758),
	.w6(32'hbb8d66f7),
	.w7(32'hbb12b9ea),
	.w8(32'hbb58e638),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30c882),
	.w1(32'hbb6ab89f),
	.w2(32'h3ae509fd),
	.w3(32'hbaad11b5),
	.w4(32'h399afea6),
	.w5(32'h3938ed5a),
	.w6(32'hbb3e3659),
	.w7(32'h3b588f25),
	.w8(32'h3a01023d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d0b92),
	.w1(32'hbb038e33),
	.w2(32'hba844565),
	.w3(32'hbb39c059),
	.w4(32'hbb749f22),
	.w5(32'h3abd0931),
	.w6(32'hbaaf13a1),
	.w7(32'hbbf76916),
	.w8(32'h3b1cf3a4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc6e5d),
	.w1(32'h3b21fcb3),
	.w2(32'hba87e165),
	.w3(32'h3ba232cf),
	.w4(32'h3a246e3d),
	.w5(32'hbbcc1bf8),
	.w6(32'h3af5f383),
	.w7(32'h3bc3139d),
	.w8(32'h3bc785d7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66773b),
	.w1(32'hbc0c0abf),
	.w2(32'hbbc8835f),
	.w3(32'h3a295170),
	.w4(32'hba7d8c75),
	.w5(32'h3a355978),
	.w6(32'hbb46dda5),
	.w7(32'hbb3b0306),
	.w8(32'h3a1f7d21),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb386c69),
	.w1(32'hbb90f75d),
	.w2(32'hb9dc355b),
	.w3(32'h3a6dbcd7),
	.w4(32'hbbca96f7),
	.w5(32'hbbae02ed),
	.w6(32'h3b69ea1a),
	.w7(32'hbbb29013),
	.w8(32'hbc01ba69),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb824),
	.w1(32'h3bce1261),
	.w2(32'h3b47d5ed),
	.w3(32'h3a3a65a8),
	.w4(32'h3b3ceace),
	.w5(32'hbb8e02da),
	.w6(32'hbb8081b0),
	.w7(32'h3b942862),
	.w8(32'h3bcf4e32),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb408378),
	.w1(32'hbb9737c4),
	.w2(32'h3c02a3e2),
	.w3(32'h3bae68dd),
	.w4(32'h3bae7f95),
	.w5(32'hbc26b4c8),
	.w6(32'h3c04b722),
	.w7(32'hba4e01da),
	.w8(32'hbc1eb02f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5474),
	.w1(32'hbb598496),
	.w2(32'hbc06e329),
	.w3(32'hbb95e7a5),
	.w4(32'hbb544637),
	.w5(32'hbb1060e8),
	.w6(32'hb95f1fc1),
	.w7(32'hbb1081d0),
	.w8(32'h3bc34d4c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b9d21),
	.w1(32'h38c6135e),
	.w2(32'h3b43d141),
	.w3(32'hbba14d7b),
	.w4(32'hbb3fa7ba),
	.w5(32'hbbe9affd),
	.w6(32'hbb3b513a),
	.w7(32'hbb2aec5d),
	.w8(32'hbbab1707),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a25dc),
	.w1(32'h3b741991),
	.w2(32'h3be7698b),
	.w3(32'h3b2b59e8),
	.w4(32'h3bfea764),
	.w5(32'h3af3b27d),
	.w6(32'hba6028ae),
	.w7(32'h3b7221ce),
	.w8(32'h3aa8e9ed),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91f7c1d),
	.w1(32'h3a2b4fa3),
	.w2(32'hbaf49cb3),
	.w3(32'h394849ca),
	.w4(32'hbb122519),
	.w5(32'hba4cff29),
	.w6(32'h39445e3d),
	.w7(32'hba883e13),
	.w8(32'h3b877ec8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963519d),
	.w1(32'hb8acf872),
	.w2(32'hbbc63b5f),
	.w3(32'h3b50f82a),
	.w4(32'h3b44723e),
	.w5(32'h3b1646ce),
	.w6(32'h3bb6bc0b),
	.w7(32'hbb45369d),
	.w8(32'hbac3c07b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab1e4a),
	.w1(32'hbc0a8b2e),
	.w2(32'hbb8ff43b),
	.w3(32'h3b3b212d),
	.w4(32'h3b01804d),
	.w5(32'hbbcb231e),
	.w6(32'hbbcb1198),
	.w7(32'hba16675e),
	.w8(32'hbc03a5a5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd810af),
	.w1(32'hbacbe43a),
	.w2(32'hbb00d8a9),
	.w3(32'hb827357e),
	.w4(32'h3b502ff2),
	.w5(32'hbb0e184f),
	.w6(32'hbb1b7e47),
	.w7(32'hb9a3b206),
	.w8(32'hbb3b9440),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6a6ca),
	.w1(32'hbbbd5f5e),
	.w2(32'hbbcdc903),
	.w3(32'h3b7217d8),
	.w4(32'hba962f50),
	.w5(32'h3ba1427e),
	.w6(32'h3b22ede2),
	.w7(32'h3afb6f49),
	.w8(32'h3a804ce3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d8286),
	.w1(32'h3b7dbbda),
	.w2(32'hb9e5d2ec),
	.w3(32'hbb104999),
	.w4(32'hbac1863a),
	.w5(32'h3bd23e60),
	.w6(32'h3a035fb8),
	.w7(32'hbb7ef5de),
	.w8(32'h3c11b321),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98121bc),
	.w1(32'hbb47b776),
	.w2(32'h3b41615f),
	.w3(32'h3a90fd38),
	.w4(32'hbb7c388e),
	.w5(32'hba1fc39c),
	.w6(32'h3be434bb),
	.w7(32'hbbaad377),
	.w8(32'hbc3a4c20),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c228e),
	.w1(32'h3b7f82db),
	.w2(32'hba5c2941),
	.w3(32'h3a1a622e),
	.w4(32'h3ab889e4),
	.w5(32'h3bdba78f),
	.w6(32'hbb9830c1),
	.w7(32'h3bf35ca8),
	.w8(32'h3c1bf687),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2fe6d),
	.w1(32'hbbe55184),
	.w2(32'h3a8fb588),
	.w3(32'hba408bc4),
	.w4(32'hbb96fa23),
	.w5(32'h3c78f17e),
	.w6(32'hbafa107a),
	.w7(32'h3a12db0d),
	.w8(32'h3bbb31e3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b20c),
	.w1(32'h3bfbb594),
	.w2(32'h3c735e3c),
	.w3(32'h3b55e0df),
	.w4(32'h3b00f683),
	.w5(32'h3ca2a8dd),
	.w6(32'h39cacfe6),
	.w7(32'hb84344be),
	.w8(32'hbb3d0007),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c8343),
	.w1(32'h3b874503),
	.w2(32'hbbf7d34c),
	.w3(32'h3b9b5ec2),
	.w4(32'h3b479d50),
	.w5(32'hbae8594d),
	.w6(32'h3b84aaba),
	.w7(32'h3b24f14f),
	.w8(32'hba612551),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad3bf5),
	.w1(32'hbbbc9458),
	.w2(32'hba885671),
	.w3(32'hbba4c092),
	.w4(32'hbbbce2b9),
	.w5(32'hbbd9dd61),
	.w6(32'hbb0c0138),
	.w7(32'hbb20fddf),
	.w8(32'hbbed33c6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb726faf),
	.w1(32'h39a3c2c0),
	.w2(32'h3bcdc0ae),
	.w3(32'hbbe082fa),
	.w4(32'hbbcefb37),
	.w5(32'hbab94d84),
	.w6(32'hbbfec740),
	.w7(32'hbab271aa),
	.w8(32'hbae35324),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223597),
	.w1(32'h3af6e74a),
	.w2(32'hbbcdc5cc),
	.w3(32'hbb1b1ac6),
	.w4(32'h3b07dbea),
	.w5(32'hbc243c22),
	.w6(32'h3b2fdc63),
	.w7(32'h3b07c492),
	.w8(32'h3bd71172),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed2ecb),
	.w1(32'h3bbb9a87),
	.w2(32'h3bbe1cd8),
	.w3(32'h379fdad0),
	.w4(32'h3c39c04e),
	.w5(32'h3ba562a6),
	.w6(32'h3af66973),
	.w7(32'h3ba1df7f),
	.w8(32'h3be4602d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3170a1),
	.w1(32'hba87e577),
	.w2(32'h3b1ed756),
	.w3(32'hbba9f6e2),
	.w4(32'h3b527ce7),
	.w5(32'h3c532e89),
	.w6(32'hbb255cb2),
	.w7(32'h3c75001a),
	.w8(32'h3b9c0102),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7e1e),
	.w1(32'h3b219437),
	.w2(32'h3b62487e),
	.w3(32'h3bacfeb4),
	.w4(32'h3bb1e489),
	.w5(32'h3b1e6bf7),
	.w6(32'h3a70e02a),
	.w7(32'h3758d6e5),
	.w8(32'hbb137c1e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3caf5),
	.w1(32'h3ad34b35),
	.w2(32'h3a6a4beb),
	.w3(32'hbb15895c),
	.w4(32'h3af1a891),
	.w5(32'hbbfac3c3),
	.w6(32'hba7ecf55),
	.w7(32'hbb0b1593),
	.w8(32'hbbe6f661),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6edf21),
	.w1(32'h3bf0dded),
	.w2(32'h3a83952e),
	.w3(32'h3b2d09c1),
	.w4(32'h3a36ec0e),
	.w5(32'hbc2677eb),
	.w6(32'hbba2810e),
	.w7(32'hb97395fd),
	.w8(32'hbbc7c6db),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15278e),
	.w1(32'h3ace5f90),
	.w2(32'h3baefca4),
	.w3(32'hbc80f4fa),
	.w4(32'hbbadf990),
	.w5(32'h3b9210f3),
	.w6(32'hbc8aaead),
	.w7(32'hbbc1c772),
	.w8(32'hbbb5a55f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d325b),
	.w1(32'hba9e235d),
	.w2(32'hb9d6bc9a),
	.w3(32'h3b68049c),
	.w4(32'hbb8572ee),
	.w5(32'hbabd43ee),
	.w6(32'hbb6d7437),
	.w7(32'hbbab57dd),
	.w8(32'hba800db4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5425c),
	.w1(32'hbb04b4b6),
	.w2(32'h3ac159ea),
	.w3(32'hbb63b238),
	.w4(32'hbb2ebcd6),
	.w5(32'h3bb44ff3),
	.w6(32'hbb57b140),
	.w7(32'h3b58df10),
	.w8(32'h3b7d8b21),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15efc6),
	.w1(32'h3c104c75),
	.w2(32'h3b3cd78b),
	.w3(32'h3aafd059),
	.w4(32'hbb1a0ca1),
	.w5(32'hbae718f8),
	.w6(32'hbb8f341e),
	.w7(32'hbb0bd378),
	.w8(32'hbbb3c044),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67e7dc),
	.w1(32'h3bdb38ba),
	.w2(32'h3af47a31),
	.w3(32'hbba6cc00),
	.w4(32'h3bbec3d3),
	.w5(32'h3c0a23d9),
	.w6(32'hbb7286f7),
	.w7(32'h3b1ab950),
	.w8(32'hb9f50878),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f8e1c),
	.w1(32'hbb1f75cc),
	.w2(32'hbaff57e0),
	.w3(32'h3b1014ec),
	.w4(32'hb9a8fafd),
	.w5(32'hbb5af4fa),
	.w6(32'hbbbad146),
	.w7(32'hbaa130e1),
	.w8(32'hbc1275ed),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a51ef),
	.w1(32'h3b1df933),
	.w2(32'h3bad417c),
	.w3(32'hba256bea),
	.w4(32'hbbaec808),
	.w5(32'hbbf62f48),
	.w6(32'hbb5f939e),
	.w7(32'hbb83545b),
	.w8(32'hbc34c4a6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6814000),
	.w1(32'h3c05c26b),
	.w2(32'h3b8c5958),
	.w3(32'h3ba6bb56),
	.w4(32'h3c863bcc),
	.w5(32'h3c54a097),
	.w6(32'h3b19c357),
	.w7(32'h3c14b387),
	.w8(32'h38b509db),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d2e4a),
	.w1(32'hb9aab903),
	.w2(32'h3b26df96),
	.w3(32'h3c20f7d2),
	.w4(32'hbbde712c),
	.w5(32'h3c4280f7),
	.w6(32'h3b0e1e99),
	.w7(32'h3b35c196),
	.w8(32'h3bf0958e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53b31c),
	.w1(32'hbbe64c8e),
	.w2(32'hbb69d7d1),
	.w3(32'h3acf95e9),
	.w4(32'hbbcb6d7b),
	.w5(32'hbb35b99f),
	.w6(32'h3c9dc1e7),
	.w7(32'h3af956ed),
	.w8(32'h3a7807c7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c220e50),
	.w1(32'hbb1b2494),
	.w2(32'hbaac2daa),
	.w3(32'hbba23f97),
	.w4(32'hba9ad0f2),
	.w5(32'hbc151aae),
	.w6(32'hbb8e6afd),
	.w7(32'hbbca04e5),
	.w8(32'h3b22707a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7bfa8),
	.w1(32'h3b514b4c),
	.w2(32'hbbe500d0),
	.w3(32'hbb2ac624),
	.w4(32'hbc9b8ada),
	.w5(32'hbc935a54),
	.w6(32'hbb7d3580),
	.w7(32'hbba9211c),
	.w8(32'h3b1ec51c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8e906),
	.w1(32'hbba4d457),
	.w2(32'h3bdf07cc),
	.w3(32'hbc139ef6),
	.w4(32'hbc158918),
	.w5(32'hbc642477),
	.w6(32'hb8249a53),
	.w7(32'hbb83cc15),
	.w8(32'h39e605fa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221657),
	.w1(32'h3bc57a4b),
	.w2(32'h3af5ec0c),
	.w3(32'hbbfbfed3),
	.w4(32'h3ba57c9a),
	.w5(32'hbae7807e),
	.w6(32'hbc06dd05),
	.w7(32'hbba66674),
	.w8(32'h3ad81755),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bf66d),
	.w1(32'hbcc41414),
	.w2(32'hbc807436),
	.w3(32'h3a89a20c),
	.w4(32'hbd04a5bc),
	.w5(32'hbd1c4592),
	.w6(32'h3b549810),
	.w7(32'hbce75d9a),
	.w8(32'hbc14a91d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87ab10),
	.w1(32'hbb59205e),
	.w2(32'h3b067cf4),
	.w3(32'hbc206166),
	.w4(32'hbba09676),
	.w5(32'hbc7c9003),
	.w6(32'hbcd6b77f),
	.w7(32'h3b60ffd4),
	.w8(32'hbab470ff),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff3a82),
	.w1(32'h3b87cc7f),
	.w2(32'hbb912a3d),
	.w3(32'hbc22ae7b),
	.w4(32'hbac0e8e2),
	.w5(32'h3baf448c),
	.w6(32'hbc55a3e1),
	.w7(32'hbade02ce),
	.w8(32'h3b0b09cf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84120f2),
	.w1(32'h3c29d2e1),
	.w2(32'h3c9f2110),
	.w3(32'hbaae624b),
	.w4(32'h3c251f16),
	.w5(32'h3c01049f),
	.w6(32'h391844ae),
	.w7(32'h36ed0004),
	.w8(32'h3ba55b57),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c968e),
	.w1(32'hbbb14cc8),
	.w2(32'h3b7148b7),
	.w3(32'h3c4015f4),
	.w4(32'hbaadf34f),
	.w5(32'h3b5b84b4),
	.w6(32'h3bc01622),
	.w7(32'hbb72b6be),
	.w8(32'h3ad90968),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f3dc),
	.w1(32'hbc1d0176),
	.w2(32'hbb20ab02),
	.w3(32'h3b6d9f62),
	.w4(32'h3afdfd32),
	.w5(32'h3ccd7ca5),
	.w6(32'hbbae65cd),
	.w7(32'hbaba74bc),
	.w8(32'hbb98fdca),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b5db9),
	.w1(32'h3a998291),
	.w2(32'hbb60e653),
	.w3(32'h3aa45c9b),
	.w4(32'hbb030b08),
	.w5(32'h3c107815),
	.w6(32'hbc4d5cfb),
	.w7(32'h3b7a4486),
	.w8(32'h3b97cf0f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b370371),
	.w1(32'hbc14eadb),
	.w2(32'hbbdda353),
	.w3(32'h3b02dfae),
	.w4(32'hbbb26778),
	.w5(32'hba0e3267),
	.w6(32'hbab3144e),
	.w7(32'h3b08cc5e),
	.w8(32'h3b6bda6d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3fb08),
	.w1(32'h3bbcfa52),
	.w2(32'h3b3db07d),
	.w3(32'hbc185301),
	.w4(32'h3b835074),
	.w5(32'h3c2e7a08),
	.w6(32'hbad9e7ea),
	.w7(32'hbb297c4e),
	.w8(32'hbb139ea7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9ca8),
	.w1(32'h3bb85a5c),
	.w2(32'h3bf017d0),
	.w3(32'hbc2bddb3),
	.w4(32'h3c8596ff),
	.w5(32'h3c140944),
	.w6(32'hbb4d3cea),
	.w7(32'h3bafe574),
	.w8(32'h3c4142f7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7960),
	.w1(32'h3b641214),
	.w2(32'hbbc5640d),
	.w3(32'h3c937ae9),
	.w4(32'h3c58f2af),
	.w5(32'hbb425181),
	.w6(32'h3c1eb231),
	.w7(32'h3b050505),
	.w8(32'h3a15642e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46e38e),
	.w1(32'hb935960e),
	.w2(32'hbbb09ea5),
	.w3(32'h3bdbbdc0),
	.w4(32'hbacc2932),
	.w5(32'h3c3c3782),
	.w6(32'hbb3c9baf),
	.w7(32'h3c04e064),
	.w8(32'h3bb15ccb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa0e45),
	.w1(32'hbc67c82c),
	.w2(32'hbc523404),
	.w3(32'h3c0501a4),
	.w4(32'h3b04e773),
	.w5(32'hbae52752),
	.w6(32'hbab9a9ee),
	.w7(32'h3ac7ce1e),
	.w8(32'hbb873817),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f8e74),
	.w1(32'hbb78efab),
	.w2(32'hbb1ccfba),
	.w3(32'hb8bc3e92),
	.w4(32'h3a9938bc),
	.w5(32'h3b8f0533),
	.w6(32'hbba3cf8a),
	.w7(32'hbac5e32d),
	.w8(32'hbaa8a6cf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cd15e),
	.w1(32'h3b3d4273),
	.w2(32'h38193959),
	.w3(32'h3b04c41c),
	.w4(32'h3c2082d7),
	.w5(32'hbb2c0737),
	.w6(32'h3a93a533),
	.w7(32'hbb0ffd90),
	.w8(32'hbbd2cdd3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0403c8),
	.w1(32'hbb000598),
	.w2(32'h3ad7476d),
	.w3(32'h3aa74d29),
	.w4(32'h3b1246f0),
	.w5(32'h3cb2c293),
	.w6(32'hba800f05),
	.w7(32'hbb68faaa),
	.w8(32'h3c1aaf5a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc8f31),
	.w1(32'h3a828eda),
	.w2(32'h3bf672a6),
	.w3(32'hbbb70759),
	.w4(32'h3c31e604),
	.w5(32'h3c682545),
	.w6(32'hbc2eb44b),
	.w7(32'h3ba60081),
	.w8(32'h3c03021a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac285ae),
	.w1(32'h3a5a5b42),
	.w2(32'hbb954013),
	.w3(32'h3bf4ffe9),
	.w4(32'hbab9047d),
	.w5(32'h3c26b918),
	.w6(32'h3aed3b4a),
	.w7(32'h3bb7fa99),
	.w8(32'hbb21c956),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e94f4),
	.w1(32'hbcaf1249),
	.w2(32'hbc964e40),
	.w3(32'h3c05d92d),
	.w4(32'hbc7889e9),
	.w5(32'hbc7be6cd),
	.w6(32'h3c68c8b5),
	.w7(32'hbcc2d345),
	.w8(32'hbc25e212),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e228),
	.w1(32'h3ab8d2d6),
	.w2(32'h3bbccd27),
	.w3(32'hbc1aa535),
	.w4(32'h3c40fe2b),
	.w5(32'hb866efd4),
	.w6(32'hbbb8d3c3),
	.w7(32'hbb354f6c),
	.w8(32'hbb004802),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c558ec3),
	.w1(32'hba62c5a1),
	.w2(32'hbc164153),
	.w3(32'h3bcb49b9),
	.w4(32'h3b45a388),
	.w5(32'hbbad037b),
	.w6(32'h3babd82c),
	.w7(32'hb812fff4),
	.w8(32'hbb4e8bc1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c921),
	.w1(32'hbbf3f06f),
	.w2(32'hbc4f84c3),
	.w3(32'hbb272990),
	.w4(32'hbb369f07),
	.w5(32'hbbb05d8e),
	.w6(32'hbb4014c3),
	.w7(32'hbb23dc23),
	.w8(32'hbc14fdef),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e7a1d),
	.w1(32'h3b0bf8e1),
	.w2(32'hba8d48ca),
	.w3(32'hbbf4c744),
	.w4(32'hbbc0cb3d),
	.w5(32'hbca6e849),
	.w6(32'hbbd697c0),
	.w7(32'h3b533a55),
	.w8(32'h3b43f0b1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcba056),
	.w1(32'h3b9df730),
	.w2(32'h3acbdf11),
	.w3(32'hbbed147e),
	.w4(32'h3c66d75c),
	.w5(32'h3cc020b1),
	.w6(32'hbba34c37),
	.w7(32'h3c0904af),
	.w8(32'h3bc85a9b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12f92c),
	.w1(32'hbbcc3dcd),
	.w2(32'h3bb81b2d),
	.w3(32'h3c8273b3),
	.w4(32'hbc2ef339),
	.w5(32'hbc2b8a9b),
	.w6(32'h3aa4bb18),
	.w7(32'hbb22fa7e),
	.w8(32'h3bbe9ae3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b474230),
	.w1(32'hbbb68692),
	.w2(32'hbc295903),
	.w3(32'hbba100a4),
	.w4(32'h3c6a4fac),
	.w5(32'h3afd08f2),
	.w6(32'hbbb80bec),
	.w7(32'hbbd809cd),
	.w8(32'h3a3eb63c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc19b17),
	.w1(32'hbc479308),
	.w2(32'hbbcf9d55),
	.w3(32'h3b94dc84),
	.w4(32'hbc06ce29),
	.w5(32'hbc38046f),
	.w6(32'hbc0c44ec),
	.w7(32'hb89a8c6d),
	.w8(32'h3b146067),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12dd3),
	.w1(32'hbc03b1f5),
	.w2(32'hbb7c29f3),
	.w3(32'hbc7ce0b6),
	.w4(32'hbc1e63a2),
	.w5(32'h3d16ef95),
	.w6(32'hbc12ef48),
	.w7(32'hbc2c3fb6),
	.w8(32'hbc2e6a00),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a555d),
	.w1(32'h3b119366),
	.w2(32'hb9e893e8),
	.w3(32'hbbd13e2e),
	.w4(32'hbb223301),
	.w5(32'h3c30a7ff),
	.w6(32'hbbe7115a),
	.w7(32'h3ac9837c),
	.w8(32'h3a18cedf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba585a2f),
	.w1(32'hbb38d2ec),
	.w2(32'h3b42f85b),
	.w3(32'hb9d01bdb),
	.w4(32'hba3c7015),
	.w5(32'hbc39942c),
	.w6(32'h3a37d37e),
	.w7(32'hbb57ef1f),
	.w8(32'hbc6a134b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc28c8c),
	.w1(32'hbb8b3394),
	.w2(32'hbb9c82e1),
	.w3(32'hbbac5834),
	.w4(32'hba14363a),
	.w5(32'hbb3eeb65),
	.w6(32'hbc5215b4),
	.w7(32'h3a028842),
	.w8(32'hbb8cb1cf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb84ae),
	.w1(32'h3b4c453b),
	.w2(32'hbaaff5e1),
	.w3(32'hb99c2df6),
	.w4(32'hb985e2d4),
	.w5(32'h3d198c9c),
	.w6(32'h3c11758c),
	.w7(32'hbbcbf3ee),
	.w8(32'hbc3c2726),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c7925),
	.w1(32'hbc4a4497),
	.w2(32'hbc5514ad),
	.w3(32'hba9e9e34),
	.w4(32'hbcbab659),
	.w5(32'h3d0bbcc3),
	.w6(32'hb99422c7),
	.w7(32'hbc7099d8),
	.w8(32'hbc3b8845),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a6883),
	.w1(32'h3be324fa),
	.w2(32'h3c2ff8b6),
	.w3(32'hbc9a1073),
	.w4(32'h3af317dc),
	.w5(32'h3b79618d),
	.w6(32'hbc47da40),
	.w7(32'h3ab2e0c1),
	.w8(32'h3b302519),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c81b6),
	.w1(32'hbb3451af),
	.w2(32'h3b4f97bd),
	.w3(32'hb8addfc3),
	.w4(32'h3b37c3dd),
	.w5(32'h3b1c61f7),
	.w6(32'h3b5a960f),
	.w7(32'h3b99ce34),
	.w8(32'hba1b8743),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b5a46),
	.w1(32'h3c177883),
	.w2(32'hbb9e7123),
	.w3(32'hbaf29bd3),
	.w4(32'h3b9fa0c0),
	.w5(32'hbc81e328),
	.w6(32'hb9da89fb),
	.w7(32'h3b4ea734),
	.w8(32'h3ce13f40),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd236d),
	.w1(32'hbc263692),
	.w2(32'hbc05dbb8),
	.w3(32'h3a81b488),
	.w4(32'h3b3b147a),
	.w5(32'h3ca288a0),
	.w6(32'h3ca59253),
	.w7(32'h3b50152c),
	.w8(32'h3c1497f0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7565),
	.w1(32'hbb1de159),
	.w2(32'hbb844270),
	.w3(32'hbb22bfb9),
	.w4(32'hbad88128),
	.w5(32'h3c164728),
	.w6(32'hbc47dfe5),
	.w7(32'h3b9351b1),
	.w8(32'h3c096f42),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f577e),
	.w1(32'h3aebe7cb),
	.w2(32'h39c2985e),
	.w3(32'h3c52883b),
	.w4(32'h3bf190ed),
	.w5(32'h3b4e8d25),
	.w6(32'h3a87bd06),
	.w7(32'h3c06f4d3),
	.w8(32'h3bd0666a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08efa4),
	.w1(32'hbb81885d),
	.w2(32'hbbf79acc),
	.w3(32'hb8b01ae5),
	.w4(32'hbb6c6839),
	.w5(32'h3c2aa697),
	.w6(32'hbb4d3e8f),
	.w7(32'h3b3b7386),
	.w8(32'h3bf4447b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5547),
	.w1(32'hba1b9c08),
	.w2(32'h3c4c2588),
	.w3(32'hbc7f39d6),
	.w4(32'h39bf793b),
	.w5(32'h3c14747c),
	.w6(32'hbb6e7045),
	.w7(32'h3c46d300),
	.w8(32'h3b923b0c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21a1ec),
	.w1(32'hbca4c74a),
	.w2(32'hbcda143f),
	.w3(32'hba0040c5),
	.w4(32'hbca82122),
	.w5(32'hbc8d662f),
	.w6(32'hbbacaa8d),
	.w7(32'hbcf3442e),
	.w8(32'hbcb8ed95),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce5348f),
	.w1(32'hbb828f1e),
	.w2(32'hbc0b64ab),
	.w3(32'hbc9c3382),
	.w4(32'hbc33fd3b),
	.w5(32'hbc449b02),
	.w6(32'hbcca238f),
	.w7(32'hbc34c500),
	.w8(32'hbb81eace),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba11c32),
	.w1(32'hbb12012a),
	.w2(32'hbaf601cf),
	.w3(32'h3ba1e7b7),
	.w4(32'hba8ddb3b),
	.w5(32'h3b10b8cc),
	.w6(32'h3b119764),
	.w7(32'hbc267708),
	.w8(32'hb9596ca2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bafb9),
	.w1(32'hbb00de31),
	.w2(32'hbbaa019e),
	.w3(32'hbba8bcf2),
	.w4(32'hbb055c58),
	.w5(32'hbbce001a),
	.w6(32'hbc16970f),
	.w7(32'hbb23d9a5),
	.w8(32'hbc1bfce9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed5827),
	.w1(32'h3ba773f9),
	.w2(32'hbba9ee7f),
	.w3(32'hbbcb0de1),
	.w4(32'h3c6fa733),
	.w5(32'h3bc546be),
	.w6(32'hbaa8d3d6),
	.w7(32'h3bf291ce),
	.w8(32'h3c4379ef),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf14bcd),
	.w1(32'h3b794f90),
	.w2(32'h3c45386a),
	.w3(32'h3c766322),
	.w4(32'hbaca591d),
	.w5(32'h3c3c5683),
	.w6(32'h3b812b15),
	.w7(32'hbc0078a1),
	.w8(32'h3c178645),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6ac5),
	.w1(32'h3bcbe606),
	.w2(32'h3c11797d),
	.w3(32'h3c3831f2),
	.w4(32'hbaf1bed0),
	.w5(32'h3bffc454),
	.w6(32'h3c4bd6fc),
	.w7(32'h3c7df414),
	.w8(32'h3c829558),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39861b53),
	.w1(32'hbbfc404a),
	.w2(32'hbc925c26),
	.w3(32'hbc2cbbe3),
	.w4(32'hbc4a307e),
	.w5(32'h3b8eccfb),
	.w6(32'h3c2d4528),
	.w7(32'hbb8b5553),
	.w8(32'h3c0a4060),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e988e),
	.w1(32'hbb0500fe),
	.w2(32'hbb452f86),
	.w3(32'hbccf7176),
	.w4(32'hbab15ed8),
	.w5(32'hbbcbbd17),
	.w6(32'hbbddc2e9),
	.w7(32'hbc3e394f),
	.w8(32'hbc1ead84),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908759),
	.w1(32'h3c36fb56),
	.w2(32'h3b9e8b33),
	.w3(32'hbbddb06c),
	.w4(32'hbaa27c60),
	.w5(32'h3bf7e845),
	.w6(32'hbc6bc00e),
	.w7(32'hbbe8874c),
	.w8(32'h3b8d8f7e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd82e60),
	.w1(32'h3b889ae7),
	.w2(32'h3addaca6),
	.w3(32'h3c13713d),
	.w4(32'h3b7cf632),
	.w5(32'h3c2b2ec2),
	.w6(32'h3b07e5b3),
	.w7(32'h3b28d0fc),
	.w8(32'h3b484b2f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af162e3),
	.w1(32'hbb9332fc),
	.w2(32'hbc69a825),
	.w3(32'h3ba20e07),
	.w4(32'hbaae3753),
	.w5(32'h3bc0d1ef),
	.w6(32'h3b102500),
	.w7(32'h3ad7ce55),
	.w8(32'h3c2bb651),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6dfaa),
	.w1(32'hbb838b91),
	.w2(32'hbb5e3e2f),
	.w3(32'h39dc711b),
	.w4(32'hbab22e43),
	.w5(32'h3cd6102a),
	.w6(32'h3baaecc1),
	.w7(32'hbc2e8a14),
	.w8(32'hb9ff6f4a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318ad7),
	.w1(32'h3c27197b),
	.w2(32'h3ca83cda),
	.w3(32'h3bc6d86a),
	.w4(32'h3aae29cd),
	.w5(32'hbb74c846),
	.w6(32'hbc3d3864),
	.w7(32'h3bc75679),
	.w8(32'h3c46dcfc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a292f),
	.w1(32'h3aa8a7a0),
	.w2(32'h3c06df6e),
	.w3(32'hbba138a7),
	.w4(32'hbba24760),
	.w5(32'hbb9f195f),
	.w6(32'h3c36cd17),
	.w7(32'hba79e19f),
	.w8(32'hbc153571),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b501272),
	.w1(32'hbb4df96c),
	.w2(32'hbbebcb62),
	.w3(32'h3aed2e8e),
	.w4(32'hbb74d47f),
	.w5(32'hbb3e7ff2),
	.w6(32'h3b12b547),
	.w7(32'h3ac15a1f),
	.w8(32'h3c36e04e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d101),
	.w1(32'h3bdbed1b),
	.w2(32'h3c4e0349),
	.w3(32'hbb2c3762),
	.w4(32'h3ad1c497),
	.w5(32'hbc8ee217),
	.w6(32'hbb629d35),
	.w7(32'hbc05ab94),
	.w8(32'h3bc99309),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c5aa),
	.w1(32'h3a827d28),
	.w2(32'h3af95173),
	.w3(32'h3b96d2ad),
	.w4(32'h3bd8239a),
	.w5(32'hbc2c64d0),
	.w6(32'hbac11ebf),
	.w7(32'hba97b17a),
	.w8(32'h3b283ff8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870703),
	.w1(32'hbb2a8c78),
	.w2(32'hbb83df28),
	.w3(32'hbbc90bbd),
	.w4(32'hbc23dfb2),
	.w5(32'hbc8ade03),
	.w6(32'hbc1d0ff7),
	.w7(32'hbc1ab317),
	.w8(32'hbc779548),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ab57),
	.w1(32'h3b195eed),
	.w2(32'h3a3328cf),
	.w3(32'hbbe9b929),
	.w4(32'hbc1ea099),
	.w5(32'hb91f7da6),
	.w6(32'h3ba730be),
	.w7(32'hbb7ba749),
	.w8(32'hbc0d8b4d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6abf),
	.w1(32'hbae839b3),
	.w2(32'hbb34d335),
	.w3(32'hbbea5393),
	.w4(32'hbbeb4bd6),
	.w5(32'h3bb0e8ae),
	.w6(32'h3a1aa277),
	.w7(32'hbc1e2983),
	.w8(32'hbc980d21),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992d69),
	.w1(32'hbb676f6e),
	.w2(32'h3a5e2cb5),
	.w3(32'hbbc42888),
	.w4(32'hba704731),
	.w5(32'h3bef237d),
	.w6(32'hbb553ca8),
	.w7(32'h3ae5ea23),
	.w8(32'h3bc76156),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d5044),
	.w1(32'hbbe93388),
	.w2(32'hbc86fd89),
	.w3(32'h38df4987),
	.w4(32'hbbe7c367),
	.w5(32'hbb461399),
	.w6(32'hba24d8c5),
	.w7(32'hbc819c73),
	.w8(32'hbacda740),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062146),
	.w1(32'hbc30cdd6),
	.w2(32'hbc35a4cb),
	.w3(32'h3ae18857),
	.w4(32'hbb01b34b),
	.w5(32'h3cefdeca),
	.w6(32'hbc248479),
	.w7(32'hbc662c9c),
	.w8(32'hbbf9bde7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec34a3),
	.w1(32'h3a62af8e),
	.w2(32'h3c02954a),
	.w3(32'hbb61238d),
	.w4(32'hba93d251),
	.w5(32'h3b901d8e),
	.w6(32'hbbc7a044),
	.w7(32'h3bcc298b),
	.w8(32'h3acd018d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f4418),
	.w1(32'hbbc8a7f9),
	.w2(32'h3bd7e39f),
	.w3(32'hbbb17cb4),
	.w4(32'hbac5db4d),
	.w5(32'h3b0e5601),
	.w6(32'hbadf2840),
	.w7(32'hbac777ff),
	.w8(32'h3bd3714a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba666582),
	.w1(32'hbc3eff47),
	.w2(32'hbbe2c50d),
	.w3(32'h3bddbd19),
	.w4(32'hbc0ba660),
	.w5(32'hbc6861ec),
	.w6(32'h3b6a8ca0),
	.w7(32'h3ba95532),
	.w8(32'hba8fa967),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3967a873),
	.w1(32'hbb482e6e),
	.w2(32'hbb67eaf1),
	.w3(32'hbc5a6183),
	.w4(32'h3b737eff),
	.w5(32'h3bff273c),
	.w6(32'hbbef27f7),
	.w7(32'hbb99f740),
	.w8(32'hbb9a4242),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2465d4),
	.w1(32'hbac4cb59),
	.w2(32'h393de262),
	.w3(32'hbaab9dbe),
	.w4(32'hba417591),
	.w5(32'h3bc3d887),
	.w6(32'hbbb82a4d),
	.w7(32'h3b452c5b),
	.w8(32'h3bd47619),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f3aa6),
	.w1(32'hbc477829),
	.w2(32'hbb4a0f2b),
	.w3(32'h3b69bb11),
	.w4(32'hbba86fe0),
	.w5(32'hbbf51ad3),
	.w6(32'h3b36dd43),
	.w7(32'h3bc1f1ba),
	.w8(32'h3ae2cd0d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c198d64),
	.w1(32'h3ba94ab4),
	.w2(32'h3b87a9b5),
	.w3(32'hbbed1597),
	.w4(32'h3c0a0584),
	.w5(32'h3c012f1a),
	.w6(32'hbb8a12c3),
	.w7(32'h3b6e73a6),
	.w8(32'h3bbadd36),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d55ce),
	.w1(32'hbacfa0f3),
	.w2(32'hbbb2cf3a),
	.w3(32'h3a80b442),
	.w4(32'h3bb5b6db),
	.w5(32'h3ba312f0),
	.w6(32'h394893ad),
	.w7(32'h3b070523),
	.w8(32'h3c032c37),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5c54b),
	.w1(32'h3bc5c54e),
	.w2(32'h3a2ab49d),
	.w3(32'h3a92c98e),
	.w4(32'hbc12fab9),
	.w5(32'hbc9f2fe9),
	.w6(32'h3a357cfc),
	.w7(32'hbb2f9b57),
	.w8(32'h3ba9fb74),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bca48),
	.w1(32'h3bfd8f90),
	.w2(32'h3b894dc3),
	.w3(32'hbac0a4af),
	.w4(32'h39cacb70),
	.w5(32'hbb05c90e),
	.w6(32'hbac18729),
	.w7(32'hbbb5eb18),
	.w8(32'h3aec8518),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a1a4),
	.w1(32'hbb4697a8),
	.w2(32'h3c00a571),
	.w3(32'h3a6f3221),
	.w4(32'h3b4dc7c2),
	.w5(32'h3bd5eab2),
	.w6(32'hba07267c),
	.w7(32'hb9ea5dda),
	.w8(32'h3bc70837),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba73f7f),
	.w1(32'h3bb2f8b4),
	.w2(32'h3c1a1f7d),
	.w3(32'h3b589d80),
	.w4(32'h3bb1a8be),
	.w5(32'hbc23f64b),
	.w6(32'h3b3ba3c1),
	.w7(32'h3b3acd2d),
	.w8(32'hbb3f3dfb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbbf06),
	.w1(32'hbc198241),
	.w2(32'h3be587aa),
	.w3(32'h3b847e37),
	.w4(32'h3b13b2a1),
	.w5(32'h3b0cc867),
	.w6(32'hba94b931),
	.w7(32'h3a2e507a),
	.w8(32'h3bcd6b93),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc65722),
	.w1(32'hbb8a8802),
	.w2(32'hbbb7c51a),
	.w3(32'hba576731),
	.w4(32'hbb869b61),
	.w5(32'hbb0e636f),
	.w6(32'h3c14fbe0),
	.w7(32'hbb505121),
	.w8(32'h3ac0df1d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f22b4),
	.w1(32'hbbcff8c6),
	.w2(32'hbc3b2c97),
	.w3(32'h3b1e4212),
	.w4(32'hbc0c63e2),
	.w5(32'hbc47fac9),
	.w6(32'hbb60c624),
	.w7(32'hbc0c5d1c),
	.w8(32'hb97e8d63),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb99179),
	.w1(32'hbc31a2c3),
	.w2(32'hbbb64535),
	.w3(32'h3bad6fed),
	.w4(32'hbb803bf3),
	.w5(32'hbbdefdbb),
	.w6(32'h3a53005c),
	.w7(32'h3a294c44),
	.w8(32'hbb941f16),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39eaab),
	.w1(32'h3abb4dc8),
	.w2(32'h3a001e8b),
	.w3(32'hbbca899f),
	.w4(32'h3a72f2be),
	.w5(32'h3b9f74c9),
	.w6(32'hbc61d169),
	.w7(32'hbc0efea9),
	.w8(32'hbaa5a1e0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d83817),
	.w1(32'hbc16b9bb),
	.w2(32'hbb9dc8b2),
	.w3(32'hbb3c1a44),
	.w4(32'hbc478389),
	.w5(32'hbc3b1774),
	.w6(32'h3b87d4f3),
	.w7(32'hbbf2c5fa),
	.w8(32'hbc093c16),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839e2c),
	.w1(32'hbb0b707c),
	.w2(32'h3b8f4fde),
	.w3(32'hbb8f79bd),
	.w4(32'h3c2192d7),
	.w5(32'h3bd008b8),
	.w6(32'hbc43e98a),
	.w7(32'h3b569911),
	.w8(32'h3c22d19c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49d29e),
	.w1(32'hbb22fd6e),
	.w2(32'hbb63aef1),
	.w3(32'h3c594bc7),
	.w4(32'h3a7be29e),
	.w5(32'hbbcf16a0),
	.w6(32'h3a463638),
	.w7(32'h3bbecabc),
	.w8(32'h3cedd393),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39586b6d),
	.w1(32'h3a7b21c5),
	.w2(32'h3c06e0aa),
	.w3(32'h3b913aeb),
	.w4(32'h3b11a2ca),
	.w5(32'h3c2e5e98),
	.w6(32'h3b8ee8e2),
	.w7(32'hb9b388ec),
	.w8(32'h3b33503f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78cf1),
	.w1(32'h3b4a1024),
	.w2(32'h3c1bb1ab),
	.w3(32'h3b2ee6e9),
	.w4(32'h3a4a7fdc),
	.w5(32'h3b9c8a5e),
	.w6(32'hbacabed8),
	.w7(32'h3c5c800f),
	.w8(32'h3bca0814),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b247700),
	.w1(32'h3ba10b45),
	.w2(32'hba4b8e71),
	.w3(32'h39a677e5),
	.w4(32'h3c3a6af4),
	.w5(32'h3a67dd5a),
	.w6(32'h3b2a39a4),
	.w7(32'h3b8abca4),
	.w8(32'hbaa52e52),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2255ab),
	.w1(32'hba7d1ddd),
	.w2(32'h3b924901),
	.w3(32'hbbcf99b8),
	.w4(32'hbb1ee9fd),
	.w5(32'hbc8afd7d),
	.w6(32'hbaaca85c),
	.w7(32'hbb99289b),
	.w8(32'hbc6ad455),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d1c93),
	.w1(32'hbb8d2f26),
	.w2(32'hbc1ffc80),
	.w3(32'hbb3c5628),
	.w4(32'hbc3d4e88),
	.w5(32'hbac318d2),
	.w6(32'hbc97de7c),
	.w7(32'hbc9f490d),
	.w8(32'hbc65ff4a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4f3c),
	.w1(32'h3c43c400),
	.w2(32'h3c883230),
	.w3(32'hb9d9a329),
	.w4(32'h3c03fcef),
	.w5(32'hbb06bb14),
	.w6(32'h3bb7087e),
	.w7(32'h3bef6771),
	.w8(32'hb9cae4a5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baffad1),
	.w1(32'hbb084bcc),
	.w2(32'hbb87e236),
	.w3(32'h3b95cbc8),
	.w4(32'hbbd48af8),
	.w5(32'h3c02a0f2),
	.w6(32'hbb1ff48c),
	.w7(32'hbc705064),
	.w8(32'h3c26a994),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33962b),
	.w1(32'hbbf8eb55),
	.w2(32'hba52bcd2),
	.w3(32'hbc26b211),
	.w4(32'h3a9415fe),
	.w5(32'hbb7ce1d3),
	.w6(32'hbc1e6b52),
	.w7(32'h3b3c0d70),
	.w8(32'hbc1fa4f9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc9555),
	.w1(32'hbbacea3c),
	.w2(32'hbc4bb0d7),
	.w3(32'hbb444a6a),
	.w4(32'hbc1058ed),
	.w5(32'hbc2f59f8),
	.w6(32'hbbb274c4),
	.w7(32'h3b2425ea),
	.w8(32'h3c10f675),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc537579),
	.w1(32'h3bec8566),
	.w2(32'h3c0ccc6e),
	.w3(32'hbbbd968d),
	.w4(32'h3b488ef2),
	.w5(32'hbb1cdccb),
	.w6(32'hba16c7c7),
	.w7(32'hbaaab4ed),
	.w8(32'h3c0f3fed),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fe502),
	.w1(32'h3b50e9ae),
	.w2(32'hb8469266),
	.w3(32'hbb5d074c),
	.w4(32'h3c309646),
	.w5(32'h3c2bdd9c),
	.w6(32'h3ba1cb9b),
	.w7(32'h3ba46b3c),
	.w8(32'h3c208358),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13ebcb),
	.w1(32'hbb20c419),
	.w2(32'h3aeec887),
	.w3(32'h3c3b81b3),
	.w4(32'h3bb2723a),
	.w5(32'hbc19ec87),
	.w6(32'h3b9c1b33),
	.w7(32'hbafb7e65),
	.w8(32'hbb6d0d63),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dbc3b),
	.w1(32'h3a294234),
	.w2(32'hbb5162ee),
	.w3(32'h3a8d332a),
	.w4(32'hbbb8418d),
	.w5(32'h3ccff50d),
	.w6(32'h3bf50b43),
	.w7(32'hbbe95463),
	.w8(32'hbc1ae8e4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc066afd),
	.w1(32'h3bcfc35b),
	.w2(32'h3addb1db),
	.w3(32'hbb374d36),
	.w4(32'h38806ba7),
	.w5(32'hbb6c2932),
	.w6(32'hbc202d47),
	.w7(32'hbb14e4b9),
	.w8(32'hbb36dea4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc0248),
	.w1(32'h3b4f2523),
	.w2(32'h3c034db4),
	.w3(32'hba108ac6),
	.w4(32'hbb219ce2),
	.w5(32'h3bbb414d),
	.w6(32'h39d4f863),
	.w7(32'hbb6fb529),
	.w8(32'h3bb9b8bb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3896),
	.w1(32'h3bc4f1e7),
	.w2(32'h3bd92ae0),
	.w3(32'hba40dbe8),
	.w4(32'hbbc34c0d),
	.w5(32'hbb1fac42),
	.w6(32'h3bf4a436),
	.w7(32'h3b979095),
	.w8(32'h3c218fd5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91f91d),
	.w1(32'h3affb8a9),
	.w2(32'h396e198b),
	.w3(32'hbb1d4d06),
	.w4(32'h3b602dc3),
	.w5(32'h3a8ea137),
	.w6(32'hbbe122ef),
	.w7(32'hbb3761de),
	.w8(32'h3b50451e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29382e),
	.w1(32'h39c867f1),
	.w2(32'h3a626b53),
	.w3(32'hbb067e8c),
	.w4(32'hbb0232f5),
	.w5(32'h3a2e634a),
	.w6(32'hbb9205a5),
	.w7(32'hbb88257f),
	.w8(32'hbba1b6bf),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf37e),
	.w1(32'h3bea61b2),
	.w2(32'hbbcaa9a6),
	.w3(32'hbb4d6320),
	.w4(32'hbc1a2b1c),
	.w5(32'hbc8fff2c),
	.w6(32'h3b08839d),
	.w7(32'hbc0aed1b),
	.w8(32'h388d08a4),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf15a83),
	.w1(32'h3b07af36),
	.w2(32'hbab8eacb),
	.w3(32'h3ab141fc),
	.w4(32'h39b37735),
	.w5(32'hbcac1a43),
	.w6(32'hbc23a98c),
	.w7(32'h3c2c6674),
	.w8(32'h3bd9cd0e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c258837),
	.w1(32'h3a853bf4),
	.w2(32'h3ba93210),
	.w3(32'h3b174ba1),
	.w4(32'hbc193a1f),
	.w5(32'hbc57e50d),
	.w6(32'hbaf959fe),
	.w7(32'hbc648e4a),
	.w8(32'hbc7cc4bc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab61097),
	.w1(32'h3a9bf224),
	.w2(32'hbb5394c6),
	.w3(32'h3b40a8e2),
	.w4(32'hbb541f70),
	.w5(32'hbbdc3a42),
	.w6(32'hbb28af97),
	.w7(32'h3bcf43d1),
	.w8(32'h3baebbd3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeac683),
	.w1(32'h3aa571fd),
	.w2(32'h3b8e4aeb),
	.w3(32'h3bbc1232),
	.w4(32'h3a035bd1),
	.w5(32'hbb537fc0),
	.w6(32'h3b253c3f),
	.w7(32'hbaf92ebf),
	.w8(32'h3b1b15d7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa70a93),
	.w1(32'hbbcd7214),
	.w2(32'hbb846d3d),
	.w3(32'hb9f59818),
	.w4(32'hb9946527),
	.w5(32'hbbfe4507),
	.w6(32'h39a5a8eb),
	.w7(32'h3b618d80),
	.w8(32'hbbb4af3b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9706b0),
	.w1(32'h3c3dcecd),
	.w2(32'hbbc317a6),
	.w3(32'hb9ae984f),
	.w4(32'h3aaad4c6),
	.w5(32'hbb75503e),
	.w6(32'hbb9a2017),
	.w7(32'h3a89ad9e),
	.w8(32'h3b8da060),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebddde),
	.w1(32'hb8a33164),
	.w2(32'h3c4071a4),
	.w3(32'h3ad79500),
	.w4(32'h3aa2c80b),
	.w5(32'h3aef09c0),
	.w6(32'h3b2278fe),
	.w7(32'h3b8aebed),
	.w8(32'hbc379f45),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeafb6),
	.w1(32'h3a9000a6),
	.w2(32'h3b08050b),
	.w3(32'h3996bad3),
	.w4(32'hb97b4815),
	.w5(32'h3ba0e9b3),
	.w6(32'h3bcd8ed5),
	.w7(32'hbb8659d1),
	.w8(32'hbc1f64d6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb417),
	.w1(32'hbb35fea0),
	.w2(32'hbbbad1c3),
	.w3(32'hb9fd2d4d),
	.w4(32'hb91682df),
	.w5(32'h3c12b88a),
	.w6(32'h3bdd291a),
	.w7(32'hba5f82b7),
	.w8(32'h3ad1a967),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66bf30),
	.w1(32'h3bd0ef73),
	.w2(32'h3afedf09),
	.w3(32'h39601ad0),
	.w4(32'hbb3d37e8),
	.w5(32'hbc24833a),
	.w6(32'h3c1957c2),
	.w7(32'h38b7add4),
	.w8(32'h3b1b8b4c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3185c0),
	.w1(32'h3b016674),
	.w2(32'hbac42303),
	.w3(32'hbbd4df61),
	.w4(32'h3a2048c1),
	.w5(32'h3c08382d),
	.w6(32'hbb510216),
	.w7(32'h3a9295be),
	.w8(32'h3c002a48),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75f896),
	.w1(32'h3bd60c3d),
	.w2(32'h3c45542e),
	.w3(32'hba392503),
	.w4(32'hbad38d1e),
	.w5(32'hbb822d81),
	.w6(32'h3b20ff5f),
	.w7(32'hbb239135),
	.w8(32'hbbd96086),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bcf90),
	.w1(32'hbbc04d93),
	.w2(32'hbbeedef2),
	.w3(32'hbb2fa56e),
	.w4(32'hbbdb7ab9),
	.w5(32'hbc6395f7),
	.w6(32'hbbbce700),
	.w7(32'hbcab1b82),
	.w8(32'hbc468a7e),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409dbd),
	.w1(32'hbbccc496),
	.w2(32'hbc07b5c4),
	.w3(32'hbb954b5b),
	.w4(32'h3c83c4a9),
	.w5(32'h3c94f1ed),
	.w6(32'h3b98da2f),
	.w7(32'h3c7617c0),
	.w8(32'h3bea3fa6),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd91c7b),
	.w1(32'h3b24ea35),
	.w2(32'hbc1a79c9),
	.w3(32'hbb1eab43),
	.w4(32'h3c43a8e6),
	.w5(32'h3bd31920),
	.w6(32'h3bb0d572),
	.w7(32'h3c1342de),
	.w8(32'h3a4c12c0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba84df7),
	.w1(32'h3a6755d8),
	.w2(32'hbab38a13),
	.w3(32'h3b54af21),
	.w4(32'h3ac5f047),
	.w5(32'h3b01aa67),
	.w6(32'h3bb4c29f),
	.w7(32'h3b6ce05b),
	.w8(32'h3b5e12e8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ae6c9),
	.w1(32'h39a11b7e),
	.w2(32'hbbd5141d),
	.w3(32'h3ba2623d),
	.w4(32'h3b1712cb),
	.w5(32'hbc23a274),
	.w6(32'h3ab5637e),
	.w7(32'h3a4aacf5),
	.w8(32'hbc1a364d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf11f43),
	.w1(32'h3b93ce21),
	.w2(32'h3b7dcb10),
	.w3(32'h3c1a8b91),
	.w4(32'h3bbba94c),
	.w5(32'h3ac9383b),
	.w6(32'h3c406b4b),
	.w7(32'hbbf7a5b2),
	.w8(32'hbc9206a2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038aa5),
	.w1(32'hb99e173d),
	.w2(32'h3c932558),
	.w3(32'hbc5567dc),
	.w4(32'h3bf8ce67),
	.w5(32'h3cc5741c),
	.w6(32'hbbf8d6be),
	.w7(32'h3ba438b8),
	.w8(32'hbb237663),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b3a95),
	.w1(32'hbac9caa8),
	.w2(32'h3a8cf5ac),
	.w3(32'hbbced181),
	.w4(32'hba1f57b8),
	.w5(32'h39cbce06),
	.w6(32'h3c40d100),
	.w7(32'hbb650a14),
	.w8(32'hbb573fc5),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be25c11),
	.w1(32'hbc594689),
	.w2(32'hbc1d8889),
	.w3(32'h3beac4fe),
	.w4(32'hbc3af097),
	.w5(32'h3c2b87f3),
	.w6(32'hbb7634f8),
	.w7(32'hbbc5da16),
	.w8(32'h3ce63853),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1b39),
	.w1(32'h3b1cedc5),
	.w2(32'h3b9f4de1),
	.w3(32'h3cda6eb3),
	.w4(32'h3b9d1753),
	.w5(32'h3c06ca15),
	.w6(32'hbad65220),
	.w7(32'h3c4f4641),
	.w8(32'h3b971d60),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf8891),
	.w1(32'hbb22d8c3),
	.w2(32'hbbc6b2dd),
	.w3(32'h3a889dee),
	.w4(32'hbc20b605),
	.w5(32'hbcd64d49),
	.w6(32'hbb4e253b),
	.w7(32'hbc0b92dd),
	.w8(32'hbba05441),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50e0f),
	.w1(32'h3b6a0cd7),
	.w2(32'hbadf3ea8),
	.w3(32'hbb8c7588),
	.w4(32'h3ac34f85),
	.w5(32'hbbe8fda2),
	.w6(32'hbc7ed689),
	.w7(32'h3a806d57),
	.w8(32'hbab64cc5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b208f0b),
	.w1(32'h3b10c7a3),
	.w2(32'hbc5172b6),
	.w3(32'h3b930375),
	.w4(32'h3c37b34a),
	.w5(32'h3b45865e),
	.w6(32'hba8deac7),
	.w7(32'hbb88fcbe),
	.w8(32'h3c17a282),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45fa95),
	.w1(32'h3b741336),
	.w2(32'h3b82564a),
	.w3(32'hbc679d9b),
	.w4(32'h3b491fe0),
	.w5(32'h3bebbf74),
	.w6(32'hbb8dffd6),
	.w7(32'h3b3cb617),
	.w8(32'hbb30ad95),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb425cc1),
	.w1(32'hbb089298),
	.w2(32'hbbfc0121),
	.w3(32'hbbca7437),
	.w4(32'h3b9b2a03),
	.w5(32'hbc2093fa),
	.w6(32'hbbbf3572),
	.w7(32'h3b326ef6),
	.w8(32'hbbb7597d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fa94e),
	.w1(32'h3b2e2542),
	.w2(32'h3af72293),
	.w3(32'hbb83fdd0),
	.w4(32'h3bef5e30),
	.w5(32'h3c79a1fd),
	.w6(32'hbbf5983b),
	.w7(32'h3c08bcb3),
	.w8(32'h3babb3f6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42d758),
	.w1(32'hbc041bc1),
	.w2(32'h3b1c2710),
	.w3(32'h3ae81e10),
	.w4(32'hbc938892),
	.w5(32'h3b37d55a),
	.w6(32'h3c224e9d),
	.w7(32'hbc2393ca),
	.w8(32'h3b26c4d7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce1e02),
	.w1(32'h3bb82b18),
	.w2(32'h3ca09100),
	.w3(32'h3c5e687a),
	.w4(32'h3c46b636),
	.w5(32'h3c584e40),
	.w6(32'h3bc52082),
	.w7(32'hbb932094),
	.w8(32'hbcd12a21),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dbefd),
	.w1(32'h3c213759),
	.w2(32'hbb4cf334),
	.w3(32'hbce4417a),
	.w4(32'hba3c1fe8),
	.w5(32'hbc05c752),
	.w6(32'hbc1cdd8a),
	.w7(32'hbb3cc540),
	.w8(32'h3c0f3aae),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca34e5),
	.w1(32'hbc1adc27),
	.w2(32'h3c8d028c),
	.w3(32'hb9cb9ffa),
	.w4(32'hbb7341e1),
	.w5(32'h3d06f23b),
	.w6(32'h3bd0f20f),
	.w7(32'h3c04408c),
	.w8(32'h3c3f80b7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2700d),
	.w1(32'h3b6df214),
	.w2(32'h3a3628ff),
	.w3(32'h3ca46bd5),
	.w4(32'hbbbe6445),
	.w5(32'h39c5bd3a),
	.w6(32'h3b5c66f2),
	.w7(32'h3b409c09),
	.w8(32'h3ba7fe3b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998a1a),
	.w1(32'hbc0a3f7b),
	.w2(32'hbb5209fa),
	.w3(32'h3ad54434),
	.w4(32'hbbabca84),
	.w5(32'hba99e48d),
	.w6(32'hbc11d74a),
	.w7(32'hbc17f028),
	.w8(32'h3a1a4903),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39803e),
	.w1(32'hbbb04877),
	.w2(32'hbc6c937a),
	.w3(32'hbbd122b0),
	.w4(32'hbc2cb3eb),
	.w5(32'hbc3c9c22),
	.w6(32'hbc606b14),
	.w7(32'hbc5a5e0f),
	.w8(32'h3b0b2707),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcedd0d),
	.w1(32'h3af0de85),
	.w2(32'hbb8ac208),
	.w3(32'hbbab5e29),
	.w4(32'hbbba1d60),
	.w5(32'hbb9c4f22),
	.w6(32'hbbdea386),
	.w7(32'hbc0c2838),
	.w8(32'hbc0d000d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9590d7),
	.w1(32'hbc0e9a0b),
	.w2(32'hbc69c16e),
	.w3(32'hbc054575),
	.w4(32'hbb0dfba9),
	.w5(32'hbc830c2c),
	.w6(32'hbc1414d5),
	.w7(32'hbb9aaf48),
	.w8(32'hbc1ff3ad),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85225b),
	.w1(32'hbbb0dbd3),
	.w2(32'hbacced46),
	.w3(32'hbc7fdc6f),
	.w4(32'hba52041a),
	.w5(32'hbc946730),
	.w6(32'hbc8d2dc1),
	.w7(32'hbb9ef16c),
	.w8(32'hbc503d46),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a861a6a),
	.w1(32'h3adf0510),
	.w2(32'h3ac3ccc8),
	.w3(32'h3a6d9b3b),
	.w4(32'h3a512397),
	.w5(32'hbae86301),
	.w6(32'hbb4588ce),
	.w7(32'hbb9cb623),
	.w8(32'h3b7de628),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed943e),
	.w1(32'hbc297f49),
	.w2(32'h3c54650d),
	.w3(32'h3be6b37a),
	.w4(32'hbbfb2691),
	.w5(32'h3c8b1886),
	.w6(32'hbc0bc3db),
	.w7(32'hbc67d530),
	.w8(32'hbc27883f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab5a36),
	.w1(32'hba626849),
	.w2(32'hbcc292a8),
	.w3(32'h3b81f212),
	.w4(32'h3c141dc1),
	.w5(32'h3b34a9ef),
	.w6(32'h3bf92c4e),
	.w7(32'hba4b79ca),
	.w8(32'h3c668120),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1cd50),
	.w1(32'h3aa9addf),
	.w2(32'h3b85324c),
	.w3(32'hbb871d2d),
	.w4(32'hbc08d2b5),
	.w5(32'hbc4a4edc),
	.w6(32'hbc605a9c),
	.w7(32'hba3478b3),
	.w8(32'h3b01d619),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db83a),
	.w1(32'hbc11ffee),
	.w2(32'h3a7730fa),
	.w3(32'hbb3af267),
	.w4(32'hbbfc24b4),
	.w5(32'h3c8aa798),
	.w6(32'hbaa29fc3),
	.w7(32'hbab09984),
	.w8(32'hba8a12fd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4da484),
	.w1(32'h3c7bbafd),
	.w2(32'hba81ec8d),
	.w3(32'h3bf0ba39),
	.w4(32'hbb8376c1),
	.w5(32'hbb15ced6),
	.w6(32'hbcceab1e),
	.w7(32'hbb20745d),
	.w8(32'h3cce7731),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376746),
	.w1(32'h388ec8cf),
	.w2(32'h39c32860),
	.w3(32'h3d1164d5),
	.w4(32'h3be001ea),
	.w5(32'hbbadbff0),
	.w6(32'h3bf13971),
	.w7(32'h385d7963),
	.w8(32'hbaeb5476),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fdace),
	.w1(32'h3a673183),
	.w2(32'hbb23a8e4),
	.w3(32'hbbdc35d6),
	.w4(32'hbbc753da),
	.w5(32'hbcacd0ca),
	.w6(32'hbbcfa234),
	.w7(32'h3c0b9ab8),
	.w8(32'h3bb0b705),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e2445),
	.w1(32'hbacf2b45),
	.w2(32'h3ad617ca),
	.w3(32'h3bfd274d),
	.w4(32'hbaad59cb),
	.w5(32'hbbe5be6d),
	.w6(32'hbb80f987),
	.w7(32'h3bb8edd5),
	.w8(32'h3bb7c0b2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcaf65),
	.w1(32'h3be1d671),
	.w2(32'hbb3bf1d4),
	.w3(32'h3ac4e458),
	.w4(32'h3c23bea8),
	.w5(32'h3c4f5565),
	.w6(32'h3a23c7ed),
	.w7(32'h3c2c984c),
	.w8(32'h3d1b252f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d625d),
	.w1(32'hbb80f6fd),
	.w2(32'h3a857d86),
	.w3(32'h3c529bdc),
	.w4(32'hbb5e1819),
	.w5(32'h3c49a388),
	.w6(32'hbbda0482),
	.w7(32'hbae4af73),
	.w8(32'hbc6398e2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d6b20),
	.w1(32'hb9467371),
	.w2(32'h3c837232),
	.w3(32'h3c842530),
	.w4(32'h3bd3a6e7),
	.w5(32'hbbcc7e0c),
	.w6(32'hbc4d7626),
	.w7(32'hbaeec34b),
	.w8(32'hbce5ab88),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ede8ba),
	.w1(32'hbbd25e07),
	.w2(32'h3bc1037b),
	.w3(32'hbc43d2ef),
	.w4(32'hbcd4f6f4),
	.w5(32'h3ca0deba),
	.w6(32'h3bb5ec4d),
	.w7(32'hb9c1e904),
	.w8(32'hbbfc649c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb309fb),
	.w1(32'hbc1bac5b),
	.w2(32'h3ba049d5),
	.w3(32'h3cd80617),
	.w4(32'hbb5eb18c),
	.w5(32'h3b9d75c9),
	.w6(32'hbbbf710f),
	.w7(32'hbbd163cc),
	.w8(32'hbcae17d1),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af6d2),
	.w1(32'hbc7a119a),
	.w2(32'hbbe880da),
	.w3(32'hbbf3e4cc),
	.w4(32'hbc6246c3),
	.w5(32'h3aa92d52),
	.w6(32'hbb8fd29e),
	.w7(32'h3bc5cf08),
	.w8(32'h3c87b54f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2def42),
	.w1(32'h3c935634),
	.w2(32'hbb846aff),
	.w3(32'h3c96f354),
	.w4(32'h3ce31228),
	.w5(32'hbc685372),
	.w6(32'h3c2ccb67),
	.w7(32'h3c45678d),
	.w8(32'hbc47d935),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabcd67),
	.w1(32'hbb9a907a),
	.w2(32'h3978e9d6),
	.w3(32'hbd3240a8),
	.w4(32'hba7873e8),
	.w5(32'hbbc65751),
	.w6(32'hbcb485f0),
	.w7(32'hbc2cdb80),
	.w8(32'hbbb89f9a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a457),
	.w1(32'hbbeb00b7),
	.w2(32'h3b4b204e),
	.w3(32'hbac66160),
	.w4(32'hbc4ad381),
	.w5(32'hbb89ba78),
	.w6(32'h3a190917),
	.w7(32'h3b7af35a),
	.w8(32'hbbe08d29),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3228),
	.w1(32'h3c43604c),
	.w2(32'h3b46040f),
	.w3(32'h3b0b51e8),
	.w4(32'h3c483c9d),
	.w5(32'h3cc78f73),
	.w6(32'h3c4df15a),
	.w7(32'h3b376dce),
	.w8(32'h3baf6766),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e4f76),
	.w1(32'h3c2171eb),
	.w2(32'hbb97effb),
	.w3(32'h3b63dc76),
	.w4(32'hbc3f2f08),
	.w5(32'hbca007e6),
	.w6(32'h3a721209),
	.w7(32'hbbe9658b),
	.w8(32'hbc11c221),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bfce5),
	.w1(32'h3a0991ad),
	.w2(32'h3a9ff167),
	.w3(32'hbba31e53),
	.w4(32'hbbf9459a),
	.w5(32'hbc1c4365),
	.w6(32'hbc05676c),
	.w7(32'h3bcf9e11),
	.w8(32'hb9882e11),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7c289),
	.w1(32'hbc172384),
	.w2(32'hbc2072e3),
	.w3(32'h3c8b27a6),
	.w4(32'hbc26eb11),
	.w5(32'hbc49a9c7),
	.w6(32'h3be1d18a),
	.w7(32'hbac059c3),
	.w8(32'h3b78aee9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace18df),
	.w1(32'hbbce0d38),
	.w2(32'hbc296998),
	.w3(32'h3c30febd),
	.w4(32'hbb22f838),
	.w5(32'hbcc296e1),
	.w6(32'hb9b87c0a),
	.w7(32'hbad7d9b2),
	.w8(32'hbbb083e2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33fc8d),
	.w1(32'h3c43964f),
	.w2(32'hbb3de5f2),
	.w3(32'h3c2d6034),
	.w4(32'h3c820789),
	.w5(32'hbc113193),
	.w6(32'hbc8619cd),
	.w7(32'h3c6cb6e3),
	.w8(32'h3bda9343),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb471cd),
	.w1(32'hbb98c5a7),
	.w2(32'h3c084897),
	.w3(32'hbc48819d),
	.w4(32'hbafd7378),
	.w5(32'h3cb668f5),
	.w6(32'hbb04af8f),
	.w7(32'h365971d8),
	.w8(32'h3bd0d655),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862187),
	.w1(32'h3c430423),
	.w2(32'h3b8047b7),
	.w3(32'h3bc70d4f),
	.w4(32'h3b4978bf),
	.w5(32'hbc6ada94),
	.w6(32'h3a9b0faa),
	.w7(32'h3c64f809),
	.w8(32'h3a156b81),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd60d62),
	.w1(32'h3ba58798),
	.w2(32'hbb3b378d),
	.w3(32'h3b99b95b),
	.w4(32'hb909dd4b),
	.w5(32'hbb0fe333),
	.w6(32'h3aa91800),
	.w7(32'hbba37308),
	.w8(32'hb9d82cea),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be6a8),
	.w1(32'hbbea0b2b),
	.w2(32'hbbc01ec6),
	.w3(32'hbbec10e2),
	.w4(32'h39974a26),
	.w5(32'h3bfcfc42),
	.w6(32'hbc78f622),
	.w7(32'hbc643084),
	.w8(32'h3be0d892),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805cc8),
	.w1(32'h3bcbb713),
	.w2(32'hb9739ca5),
	.w3(32'h3b5d773c),
	.w4(32'h3d16d093),
	.w5(32'hbb8d3d6f),
	.w6(32'hbc553fde),
	.w7(32'h3b845163),
	.w8(32'hbb3a578c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb39460),
	.w1(32'h3b9c90a1),
	.w2(32'h3adaaf11),
	.w3(32'hbcdde387),
	.w4(32'h3b3df70e),
	.w5(32'h3c07c5c8),
	.w6(32'hbc2117ca),
	.w7(32'hbb5f991c),
	.w8(32'hbb806e4f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01794),
	.w1(32'hbb0eee9a),
	.w2(32'h3c378d32),
	.w3(32'hbc271c46),
	.w4(32'h3b929ff6),
	.w5(32'hbad95dd4),
	.w6(32'hbc0ef3f4),
	.w7(32'h3b03c7e6),
	.w8(32'hbbeb7bff),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb63ebf),
	.w1(32'hbba166fa),
	.w2(32'hbc4f0d3e),
	.w3(32'hbb23f8cd),
	.w4(32'hbbe99c1a),
	.w5(32'hbc87d4c6),
	.w6(32'h3bcc2545),
	.w7(32'hbc8efda6),
	.w8(32'hbc9c4e19),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64ca64),
	.w1(32'hbc80ca78),
	.w2(32'h3bd0fdc9),
	.w3(32'hbc86703c),
	.w4(32'hbd12804b),
	.w5(32'h3c736a40),
	.w6(32'hbc729db1),
	.w7(32'hbca7b2f0),
	.w8(32'h3b9dace5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85f788),
	.w1(32'h3b67e774),
	.w2(32'h3c822887),
	.w3(32'h3d127e0d),
	.w4(32'hbbb6b0e6),
	.w5(32'h3b2819c6),
	.w6(32'h3c7d23e2),
	.w7(32'hbbf93867),
	.w8(32'hbcccf0cd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ee292),
	.w1(32'h3c4239b9),
	.w2(32'h3b9c71fc),
	.w3(32'hbb79c1b1),
	.w4(32'h3b08faa0),
	.w5(32'h3b28818a),
	.w6(32'h3a0d96ba),
	.w7(32'h3b0d5780),
	.w8(32'hbbe9eb50),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b2713),
	.w1(32'hba3c9212),
	.w2(32'hbafa1274),
	.w3(32'hbbdd1cb1),
	.w4(32'hbaaf5ffe),
	.w5(32'hbc786e84),
	.w6(32'hbc625b61),
	.w7(32'hbb0dc4ca),
	.w8(32'hbb00d944),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35f146),
	.w1(32'h3c416c2e),
	.w2(32'h3b75268c),
	.w3(32'hbc1c0134),
	.w4(32'h3bb15c4a),
	.w5(32'hbc0081fe),
	.w6(32'hbc6aafe2),
	.w7(32'h39a817b8),
	.w8(32'hbba8afc7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule