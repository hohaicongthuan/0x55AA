module layer_10_featuremap_222(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc371cb1),
	.w1(32'hb962b001),
	.w2(32'hbc19edc4),
	.w3(32'h3b5ff060),
	.w4(32'h3b0cf09b),
	.w5(32'hbd36c774),
	.w6(32'h3c3c9f23),
	.w7(32'hbb691140),
	.w8(32'hbbbe132c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc8312),
	.w1(32'hbaaed38d),
	.w2(32'h3984c60a),
	.w3(32'h3a9261a2),
	.w4(32'hbc3eaab4),
	.w5(32'hbc81132e),
	.w6(32'hbb1ec7f2),
	.w7(32'hb91443a8),
	.w8(32'hbb3e5c2c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc429713),
	.w1(32'hbc6ee9b4),
	.w2(32'hbbc3e0ac),
	.w3(32'hb821c012),
	.w4(32'hbc0da228),
	.w5(32'h3c0f97c9),
	.w6(32'hbc2bb9cc),
	.w7(32'h3b279f5e),
	.w8(32'h3c0f452b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d436b),
	.w1(32'hbbbacfbd),
	.w2(32'hbbb3a2fa),
	.w3(32'hbbe52b15),
	.w4(32'hbbab2053),
	.w5(32'hbb7bf003),
	.w6(32'h3bf78c27),
	.w7(32'hbc749a22),
	.w8(32'h3983c193),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e5c59),
	.w1(32'h3c57bb13),
	.w2(32'h37e1668d),
	.w3(32'h3baaa916),
	.w4(32'hbc05a4c2),
	.w5(32'hbabf63f9),
	.w6(32'hbbc3759f),
	.w7(32'hbbf2cf3c),
	.w8(32'hbb5c4172),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc55a),
	.w1(32'h3ab31c1a),
	.w2(32'hbb62a89b),
	.w3(32'hbc058519),
	.w4(32'h3b91a1cc),
	.w5(32'hbd3c7235),
	.w6(32'hbc91a263),
	.w7(32'h3c069012),
	.w8(32'hbc0beed0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ef719),
	.w1(32'hbcf19d03),
	.w2(32'hbcbd2438),
	.w3(32'h3c42aebf),
	.w4(32'hbc941ba4),
	.w5(32'hbb12ab96),
	.w6(32'hbc18782a),
	.w7(32'hbaaa163b),
	.w8(32'hbd05135e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdabf538),
	.w1(32'h38ec4b54),
	.w2(32'h3c09cdb5),
	.w3(32'hbd16f4c1),
	.w4(32'hbccaa211),
	.w5(32'h3cbe5913),
	.w6(32'hbcedb70a),
	.w7(32'h3bd905a5),
	.w8(32'h3b8ad00f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d09bd),
	.w1(32'h3bd93899),
	.w2(32'hbbdf9e26),
	.w3(32'h3a36f49e),
	.w4(32'hbb678b4a),
	.w5(32'h3c2543bf),
	.w6(32'h3bfe8a4c),
	.w7(32'hbb854b7c),
	.w8(32'hb84a76b5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ca097),
	.w1(32'hbc3056d1),
	.w2(32'hbb9fca1b),
	.w3(32'h3b8a25ce),
	.w4(32'h3b7575f6),
	.w5(32'h3c9fe6b6),
	.w6(32'hbb47b0eb),
	.w7(32'h3c2f0e45),
	.w8(32'h3d0db025),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95471e),
	.w1(32'h3c498b2a),
	.w2(32'h3a318549),
	.w3(32'h3c2919ff),
	.w4(32'hbbba2579),
	.w5(32'hbbf1c2fb),
	.w6(32'h398a7bb8),
	.w7(32'h3bdc6696),
	.w8(32'h3c714e41),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc963c13),
	.w1(32'hbd0d495d),
	.w2(32'hbc415628),
	.w3(32'h3c530c98),
	.w4(32'hbb623f2a),
	.w5(32'hbbbdb3ef),
	.w6(32'hbb9a6043),
	.w7(32'hbb7bafed),
	.w8(32'hbcce5f54),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71209),
	.w1(32'hbc4fdab0),
	.w2(32'h3baee141),
	.w3(32'h39b8f786),
	.w4(32'h3bae9263),
	.w5(32'h3ce6a8bb),
	.w6(32'hbce50c3e),
	.w7(32'h3b15151b),
	.w8(32'h3bdfbe1c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a238144),
	.w1(32'hbc43b77b),
	.w2(32'hbcad55a0),
	.w3(32'h3aba9ffe),
	.w4(32'h3bc6c684),
	.w5(32'h3c25042f),
	.w6(32'hbb877d74),
	.w7(32'hbc245833),
	.w8(32'h3c73508a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad61c5),
	.w1(32'h3bace9ef),
	.w2(32'hbb3baaf0),
	.w3(32'hbc1478fa),
	.w4(32'hbc51376e),
	.w5(32'hbb322077),
	.w6(32'h3d8e3c34),
	.w7(32'h3c0ae050),
	.w8(32'h3ba71a86),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0f689),
	.w1(32'hbbc37783),
	.w2(32'h3c8a92c6),
	.w3(32'hbcbad774),
	.w4(32'h3c91292f),
	.w5(32'h3cfc8393),
	.w6(32'h3c0996ef),
	.w7(32'h3b38b917),
	.w8(32'h3cfe3811),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb983677),
	.w1(32'h39f6b845),
	.w2(32'hbc6843c5),
	.w3(32'hbb749d97),
	.w4(32'h38fcd652),
	.w5(32'h3bc3bdd1),
	.w6(32'hbbbbdacd),
	.w7(32'hba0134e7),
	.w8(32'hbb47b877),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14cb18),
	.w1(32'hbb58c63a),
	.w2(32'h3c08bf62),
	.w3(32'h3bc2332d),
	.w4(32'h3c247507),
	.w5(32'h3d2e5c22),
	.w6(32'hbc8e4dfc),
	.w7(32'h3c803209),
	.w8(32'h3b1983c2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eac23),
	.w1(32'h3b4b429c),
	.w2(32'h3c4d37c8),
	.w3(32'hbc2754f2),
	.w4(32'h3c0e378a),
	.w5(32'h3c8459fb),
	.w6(32'hbb20d59a),
	.w7(32'h3c74b779),
	.w8(32'hbc0bfbac),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ea6d2),
	.w1(32'h3b5f9590),
	.w2(32'hbbfc9a6f),
	.w3(32'h3c36c3e6),
	.w4(32'h3b43a370),
	.w5(32'h3ad7c302),
	.w6(32'h3c98be33),
	.w7(32'h3b90e4f2),
	.w8(32'hbc0208c4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c734f54),
	.w1(32'hbbc9318f),
	.w2(32'hbb0fa5e1),
	.w3(32'hb9976ffa),
	.w4(32'hba62d147),
	.w5(32'h3cd444c5),
	.w6(32'hbb624254),
	.w7(32'hbbdeeee3),
	.w8(32'hbbd1de6b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0299c2),
	.w1(32'h3b33c47b),
	.w2(32'h3b7091b3),
	.w3(32'hb9d5a82f),
	.w4(32'hbb2faa11),
	.w5(32'hbbffdff3),
	.w6(32'hb9d999b1),
	.w7(32'h3aedcaa5),
	.w8(32'hbbda56e1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd39292d),
	.w1(32'hbd1a314c),
	.w2(32'h3caa3bba),
	.w3(32'hbc45fd34),
	.w4(32'h3ca7b596),
	.w5(32'h3c851bc4),
	.w6(32'hbc975c86),
	.w7(32'h3bcbac6e),
	.w8(32'h3c7fa600),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98600c),
	.w1(32'h375fda7c),
	.w2(32'hbb8d92f4),
	.w3(32'h3bd33b0f),
	.w4(32'hbb9c03d2),
	.w5(32'hbb954835),
	.w6(32'h3b7ff6ac),
	.w7(32'h3ba33b62),
	.w8(32'h3b37040b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6e45aa),
	.w1(32'h3cf97c59),
	.w2(32'h3c423b7c),
	.w3(32'hbba5cdab),
	.w4(32'hbb6d85c5),
	.w5(32'hbcb26a15),
	.w6(32'h3cd2889b),
	.w7(32'h3c88f46a),
	.w8(32'h3bc70a84),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060711),
	.w1(32'h3bff02f5),
	.w2(32'h3bf0d657),
	.w3(32'hbbdad352),
	.w4(32'h3cd51292),
	.w5(32'hbc4320ff),
	.w6(32'hbbd50c7d),
	.w7(32'hb98590c0),
	.w8(32'hbbbfd288),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b2201),
	.w1(32'hbafbea4b),
	.w2(32'hbc6f5d17),
	.w3(32'hbbdc4f9c),
	.w4(32'h39bd425c),
	.w5(32'h3af032c9),
	.w6(32'hbc13a68e),
	.w7(32'hbb254c53),
	.w8(32'h3bda433b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6040f5),
	.w1(32'hbd1116ba),
	.w2(32'hbcc59002),
	.w3(32'h3d523278),
	.w4(32'hbcc7de5a),
	.w5(32'h3c0100ba),
	.w6(32'h3db1e364),
	.w7(32'hbbe25645),
	.w8(32'h3d378950),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36bc18),
	.w1(32'h3ba28afe),
	.w2(32'h3c80c9bd),
	.w3(32'hba0cd810),
	.w4(32'hbbc749ab),
	.w5(32'hbbf0a5d2),
	.w6(32'hb9a2fdbb),
	.w7(32'h3b5cddbc),
	.w8(32'h3b943157),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd09600),
	.w1(32'h3ce6307e),
	.w2(32'h3c516f8c),
	.w3(32'h3d917dca),
	.w4(32'hbc510088),
	.w5(32'hbd1fe6a5),
	.w6(32'h3db500e6),
	.w7(32'h3b47a181),
	.w8(32'h3b7d5fe3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea4b45),
	.w1(32'h3c2909da),
	.w2(32'h3bfd8770),
	.w3(32'hbb365225),
	.w4(32'h3b9fc064),
	.w5(32'h3c2346d4),
	.w6(32'h3c1fa650),
	.w7(32'hba401bb9),
	.w8(32'hbb92cb82),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb664599),
	.w1(32'h3b93f548),
	.w2(32'h3c2365ea),
	.w3(32'hbc375114),
	.w4(32'h3c496b81),
	.w5(32'h3c2252a0),
	.w6(32'hbc58d3b1),
	.w7(32'h3bf11c7b),
	.w8(32'h3b8fd29f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55de4),
	.w1(32'h3bb4e4b5),
	.w2(32'h3bbe43e4),
	.w3(32'h3bf083bd),
	.w4(32'h3becceef),
	.w5(32'h3c312f4b),
	.w6(32'hbc2be612),
	.w7(32'hbc2f35f5),
	.w8(32'h3b3d8106),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7a963),
	.w1(32'hbb3bb21b),
	.w2(32'h3bc95e73),
	.w3(32'h3b3dd337),
	.w4(32'hbb70444a),
	.w5(32'hbbf3e1b5),
	.w6(32'h3bbbe6e1),
	.w7(32'h3ba8e983),
	.w8(32'h3b4de4d4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeb36f),
	.w1(32'hbc5e4e33),
	.w2(32'h3caec9af),
	.w3(32'hba1f3943),
	.w4(32'h3b934055),
	.w5(32'h3b9216de),
	.w6(32'hbc0f56d5),
	.w7(32'h3a381087),
	.w8(32'h3bd5da84),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a12cc),
	.w1(32'hbc45150a),
	.w2(32'hba915c65),
	.w3(32'h3c520d15),
	.w4(32'hbc8e7e0c),
	.w5(32'hbb0d6af6),
	.w6(32'h3a9fa186),
	.w7(32'h3cdd59e7),
	.w8(32'hba8d7fb9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7e392b),
	.w1(32'hbcf8d175),
	.w2(32'hbd1d29cf),
	.w3(32'h3b76d405),
	.w4(32'h3c2310de),
	.w5(32'hbd041f0c),
	.w6(32'hbc184bca),
	.w7(32'hbccef1c8),
	.w8(32'hbd174da0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc6caa2),
	.w1(32'h3c733aab),
	.w2(32'h3be6b95f),
	.w3(32'h3cc62d92),
	.w4(32'hbce72cc7),
	.w5(32'hbd3e8b80),
	.w6(32'h3d88561f),
	.w7(32'h3c273a59),
	.w8(32'hbc7178d6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd335cc),
	.w1(32'hbbb0ac5c),
	.w2(32'hbc8ff297),
	.w3(32'h3ca6925b),
	.w4(32'hbd55c0aa),
	.w5(32'hbd6f8be3),
	.w6(32'h3dde2527),
	.w7(32'hbb8552f9),
	.w8(32'hbc319b36),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c512cd1),
	.w1(32'h3c99499c),
	.w2(32'h3b671f7e),
	.w3(32'h3a504166),
	.w4(32'hbb438842),
	.w5(32'h3b3b7852),
	.w6(32'h3c95df6d),
	.w7(32'hbb52890c),
	.w8(32'hbb31c603),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86118d6),
	.w1(32'hbcf1a22e),
	.w2(32'h3cb3b4b8),
	.w3(32'hbb5ed9fc),
	.w4(32'h3d4c5954),
	.w5(32'h3b3a0f16),
	.w6(32'hb9a056c7),
	.w7(32'h39e1c89c),
	.w8(32'h3bc8520d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00d96f),
	.w1(32'hbb7add4b),
	.w2(32'hbbf03477),
	.w3(32'hbc107008),
	.w4(32'hba213353),
	.w5(32'hbb9ff57a),
	.w6(32'hbc271a3a),
	.w7(32'h3baa0565),
	.w8(32'hbc4f3ec8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7dd3),
	.w1(32'h39b74ff6),
	.w2(32'h3b2ba751),
	.w3(32'hba02e32f),
	.w4(32'h3c46ba10),
	.w5(32'h3c61ed73),
	.w6(32'h3c0c03ab),
	.w7(32'h3c8b5618),
	.w8(32'h3c2537db),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeef8ec),
	.w1(32'hbc4d226f),
	.w2(32'hbc1c05d4),
	.w3(32'h3abf18b5),
	.w4(32'h3ce4a2e5),
	.w5(32'h3d15273e),
	.w6(32'hbc178ea4),
	.w7(32'h3bcb67bb),
	.w8(32'h3cc9dd6c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9281c5),
	.w1(32'h3c5fa5ff),
	.w2(32'h3c19c417),
	.w3(32'h3bcb8856),
	.w4(32'hbbaeea79),
	.w5(32'hbb6fe043),
	.w6(32'h3cde2bef),
	.w7(32'h3cacba9c),
	.w8(32'h3bd6711d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c04ed),
	.w1(32'h3c278e02),
	.w2(32'h3c4dd840),
	.w3(32'h3b841b10),
	.w4(32'h3bc557cc),
	.w5(32'hbc2e94e5),
	.w6(32'h3b98301f),
	.w7(32'h3bcdec2a),
	.w8(32'h3be69fe1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a7f0),
	.w1(32'h3bbe7e79),
	.w2(32'h3bc06e30),
	.w3(32'h3c2b371f),
	.w4(32'h3c4790dd),
	.w5(32'h3c56c0f7),
	.w6(32'h3c8b60aa),
	.w7(32'h3c327e7e),
	.w8(32'h3c6bfc2a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd183256),
	.w1(32'hbcc3eacb),
	.w2(32'h3b892d73),
	.w3(32'h3c9fc813),
	.w4(32'h3ccc725c),
	.w5(32'h3d0441f0),
	.w6(32'hbb3bbc97),
	.w7(32'hbb2b7380),
	.w8(32'h3bf52bf1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fd8f9),
	.w1(32'h3cc63c45),
	.w2(32'hbb834940),
	.w3(32'hbb933726),
	.w4(32'hbc841447),
	.w5(32'h3c6f6868),
	.w6(32'h3bd3e6aa),
	.w7(32'h3b05367d),
	.w8(32'h3c609dfb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b4d81),
	.w1(32'hbbadee61),
	.w2(32'hbc0d4817),
	.w3(32'h3b432ee2),
	.w4(32'h3c4036bc),
	.w5(32'hbb85cf80),
	.w6(32'hb9d85b08),
	.w7(32'hba6aae6d),
	.w8(32'h3a7fe7b1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9441ea6),
	.w1(32'h3c0997cb),
	.w2(32'h3a25a049),
	.w3(32'h39525482),
	.w4(32'h3b52cc54),
	.w5(32'hb9c092bd),
	.w6(32'hb939655e),
	.w7(32'h3c4658cd),
	.w8(32'hbb0176b7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48cb11),
	.w1(32'h3aec429f),
	.w2(32'h3c767df3),
	.w3(32'h3c042263),
	.w4(32'hba7e2e95),
	.w5(32'hbbfa55cc),
	.w6(32'h3be7e49b),
	.w7(32'hbba3fa35),
	.w8(32'h3bde5786),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc13a56),
	.w1(32'h3ba4a76a),
	.w2(32'h3c9eca34),
	.w3(32'hbc65be92),
	.w4(32'h3c09c68c),
	.w5(32'h3bf3f77d),
	.w6(32'h3bcee052),
	.w7(32'hb9756a13),
	.w8(32'h3c92876c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01e5de),
	.w1(32'hbb7c51c1),
	.w2(32'h39caf3ca),
	.w3(32'h3bdb7b63),
	.w4(32'h3d06cc27),
	.w5(32'h3cefd9b8),
	.w6(32'hbb4ed9ea),
	.w7(32'hb91a6d1c),
	.w8(32'hbafe5d04),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b897a76),
	.w1(32'h3c072bbc),
	.w2(32'h3b1168db),
	.w3(32'hbbf6e460),
	.w4(32'hbb604ae4),
	.w5(32'h3c6d560f),
	.w6(32'h3be2919c),
	.w7(32'h3b0ad244),
	.w8(32'hbb463c81),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecfb2b),
	.w1(32'hbaf22fd3),
	.w2(32'h39b59b3f),
	.w3(32'h3be2214e),
	.w4(32'hbbd53c7a),
	.w5(32'h3c17c2cb),
	.w6(32'h3a45b815),
	.w7(32'h3bad07a4),
	.w8(32'h3ba075e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5ee11),
	.w1(32'h3b7ec608),
	.w2(32'hba3bc02b),
	.w3(32'h3bcdbfdb),
	.w4(32'hba5baf05),
	.w5(32'hbc0f9375),
	.w6(32'hbbf1198a),
	.w7(32'h3c73ace4),
	.w8(32'h3b019e5a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3ebad),
	.w1(32'h3c760c4c),
	.w2(32'h3bc2e90d),
	.w3(32'hbb9c2b23),
	.w4(32'h3aa01721),
	.w5(32'hbb846fa3),
	.w6(32'h3b44e9a8),
	.w7(32'h3bc20cd7),
	.w8(32'hbb542af2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f676a),
	.w1(32'hbbfc438a),
	.w2(32'h3b82193a),
	.w3(32'h3bb5b1ca),
	.w4(32'hbb7b4321),
	.w5(32'h3b56abe4),
	.w6(32'h3c1465d2),
	.w7(32'h3b128458),
	.w8(32'hbc21242e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cb918),
	.w1(32'hbc2e1629),
	.w2(32'h3bb0d402),
	.w3(32'h3bd61d1a),
	.w4(32'h3b2ca062),
	.w5(32'h3c8936dd),
	.w6(32'h3be2c16b),
	.w7(32'hbc2717cc),
	.w8(32'hbb998d5f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b15b9),
	.w1(32'hbb8b81a2),
	.w2(32'h3c6955c3),
	.w3(32'hbb84d445),
	.w4(32'h3c785fd5),
	.w5(32'h3bb80e7d),
	.w6(32'hbc7196ac),
	.w7(32'h3be53a2f),
	.w8(32'h3bd05cfb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52569c),
	.w1(32'hbca06c16),
	.w2(32'h3c0560fc),
	.w3(32'h3c203dc3),
	.w4(32'hbc370ad9),
	.w5(32'h3d0f6bc3),
	.w6(32'h3bdc5894),
	.w7(32'h3c5b91c7),
	.w8(32'h3c5e2731),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fb51c),
	.w1(32'hbac6bbae),
	.w2(32'h3aae4d1d),
	.w3(32'hbb9fead4),
	.w4(32'h3b10d3ce),
	.w5(32'hbbf09438),
	.w6(32'h3b8a1bcc),
	.w7(32'h3af5a227),
	.w8(32'h3ac3b20c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9796fd),
	.w1(32'hb9bce9a4),
	.w2(32'h39b0dc81),
	.w3(32'h3aa4f32a),
	.w4(32'h3bc416de),
	.w5(32'h3a6d197c),
	.w6(32'hbbfaab0a),
	.w7(32'hbbcbc7ce),
	.w8(32'h3d0f8b09),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff60cc),
	.w1(32'h3aa0f8a1),
	.w2(32'h3a4e2ba1),
	.w3(32'h3a3e8c69),
	.w4(32'h3b154df1),
	.w5(32'hbbe67636),
	.w6(32'h3a254c25),
	.w7(32'hba123f9c),
	.w8(32'hb8ff2aea),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9890),
	.w1(32'hbb62c44d),
	.w2(32'h3b6210d8),
	.w3(32'h3c297a44),
	.w4(32'h3bc4e893),
	.w5(32'hbab47f21),
	.w6(32'hbb8adadb),
	.w7(32'hbba8b677),
	.w8(32'hbc0bed85),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd590ed7),
	.w1(32'hbd019748),
	.w2(32'hbbb4523f),
	.w3(32'hbaa36bdf),
	.w4(32'h3d6c9e04),
	.w5(32'h3dcf0f35),
	.w6(32'h3c0955f0),
	.w7(32'h3c92dfff),
	.w8(32'h3d97eae5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fccb9),
	.w1(32'h3d0584b5),
	.w2(32'h3d7f51d2),
	.w3(32'hbc8d6aa4),
	.w4(32'h3b77a901),
	.w5(32'h3abca81d),
	.w6(32'hbcb60682),
	.w7(32'h3ccab2c0),
	.w8(32'h3cb28fbd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6dba),
	.w1(32'h3ba3e8c7),
	.w2(32'h3cd2c288),
	.w3(32'h3ae09835),
	.w4(32'h3cb5d76a),
	.w5(32'h3c976cb3),
	.w6(32'hbab3f030),
	.w7(32'h3ceb1b91),
	.w8(32'h3c2ab44f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dbccce5),
	.w1(32'h3d2f6952),
	.w2(32'h3c9dcba3),
	.w3(32'h3cee0fcb),
	.w4(32'hbc862335),
	.w5(32'hbcc0fbaf),
	.w6(32'h3d2c636d),
	.w7(32'h3bd5fed3),
	.w8(32'h3a843064),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0054d),
	.w1(32'hbbb112ad),
	.w2(32'h3c84315b),
	.w3(32'h3ac4f521),
	.w4(32'hb9c80ac5),
	.w5(32'h3c0d7716),
	.w6(32'hb93e1a5d),
	.w7(32'hbc0558a0),
	.w8(32'hbb97c1b8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa65c26),
	.w1(32'h3b8fbd39),
	.w2(32'hbc5087aa),
	.w3(32'h38273690),
	.w4(32'hbc452d9f),
	.w5(32'hb919b2e7),
	.w6(32'hbba7b769),
	.w7(32'hbba931ab),
	.w8(32'hbc415154),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1249bd),
	.w1(32'h3ba62abc),
	.w2(32'h39caecef),
	.w3(32'h3a99c3f5),
	.w4(32'h3b9d514b),
	.w5(32'h3c58a516),
	.w6(32'hbaafffe9),
	.w7(32'h3c2bf9a2),
	.w8(32'h3b9f75c1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc551047),
	.w1(32'hba368617),
	.w2(32'h3bda361c),
	.w3(32'h3ad1336f),
	.w4(32'h3ca20d09),
	.w5(32'h3c1e0ce9),
	.w6(32'hbb8ae3a4),
	.w7(32'h3c7a36c8),
	.w8(32'h3b175d16),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba997522),
	.w1(32'h3bb6b0ce),
	.w2(32'hba5c8451),
	.w3(32'hbbf73726),
	.w4(32'h3c8e61d3),
	.w5(32'h3b13c707),
	.w6(32'h3baf1131),
	.w7(32'h3c0c61f5),
	.w8(32'h3c1affdb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ca932),
	.w1(32'hbbff859f),
	.w2(32'hbc792dd3),
	.w3(32'h3ab731f2),
	.w4(32'h3a3499c5),
	.w5(32'h3c958973),
	.w6(32'hba9613a9),
	.w7(32'hbbffa29b),
	.w8(32'h3b9ea352),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdafdc8),
	.w1(32'hbcdcadd4),
	.w2(32'h3c2c79aa),
	.w3(32'h3a2e8cf8),
	.w4(32'h3b215f25),
	.w5(32'h3cd91c1c),
	.w6(32'hbbab71b0),
	.w7(32'h3b069228),
	.w8(32'h3c064708),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca66459),
	.w1(32'h3c1f0ac8),
	.w2(32'h3bad213b),
	.w3(32'hbbad9f3e),
	.w4(32'hba59bb7d),
	.w5(32'hbb82c60f),
	.w6(32'h3cc72a31),
	.w7(32'hbafbd8e5),
	.w8(32'h3b81c7a9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900a29),
	.w1(32'h3bac5767),
	.w2(32'h3be2e0ee),
	.w3(32'hbb77f765),
	.w4(32'h3c04bd9e),
	.w5(32'h3ca45a2f),
	.w6(32'hbb5e6b6c),
	.w7(32'h3b2510a0),
	.w8(32'h3c6916dc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e4d5a),
	.w1(32'hbb9067fa),
	.w2(32'hbcac5242),
	.w3(32'h3c3f3568),
	.w4(32'h3c4229c2),
	.w5(32'h3cd78cbc),
	.w6(32'h3c31d065),
	.w7(32'h3bd02f8c),
	.w8(32'h3c4fa00b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fc923),
	.w1(32'h3c156674),
	.w2(32'hba9033ca),
	.w3(32'h3b88a45c),
	.w4(32'h3b399eb9),
	.w5(32'h3c0e65b0),
	.w6(32'h3cb644f3),
	.w7(32'h39b36a4b),
	.w8(32'h3be3ca61),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af37de5),
	.w1(32'hbb3b7399),
	.w2(32'h3bae02b2),
	.w3(32'hbb499ccc),
	.w4(32'h3b47f38e),
	.w5(32'h3b916afe),
	.w6(32'hbbd0bbd8),
	.w7(32'h3c036a69),
	.w8(32'hbc0f2746),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ee9fa),
	.w1(32'hbc85910e),
	.w2(32'h3c382fbc),
	.w3(32'h3bca6cd7),
	.w4(32'h3c8ca632),
	.w5(32'h3ba2438c),
	.w6(32'h3b58f194),
	.w7(32'h3a9f23ce),
	.w8(32'h3c2efb4b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83bba1),
	.w1(32'hbb692576),
	.w2(32'h3c0bd0bd),
	.w3(32'h3bdb8083),
	.w4(32'h3ba1485a),
	.w5(32'hba1850fd),
	.w6(32'hbac7a604),
	.w7(32'hbc7c0489),
	.w8(32'hbc57b429),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb811eba),
	.w1(32'hbcba93e6),
	.w2(32'h3bc8a642),
	.w3(32'h3b57abd4),
	.w4(32'hbab3426d),
	.w5(32'hbc0ae6dc),
	.w6(32'hbbb6412a),
	.w7(32'hbca1c049),
	.w8(32'hbcce99f0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84882f),
	.w1(32'hbca4e0bb),
	.w2(32'hbd35aa63),
	.w3(32'h3c46b643),
	.w4(32'hbc5ddb53),
	.w5(32'hbbbb0633),
	.w6(32'h3ba4b33f),
	.w7(32'hbc2a8b1f),
	.w8(32'hbb97f1c5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aa4fc),
	.w1(32'h3ba944a4),
	.w2(32'hbb8a3088),
	.w3(32'h3c1d9eee),
	.w4(32'hbcec3060),
	.w5(32'hbcab38a0),
	.w6(32'hbc055a67),
	.w7(32'h3c243e21),
	.w8(32'h3bb195d8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43f5c9),
	.w1(32'h3cb1ff66),
	.w2(32'hbc39dfe0),
	.w3(32'hbb8871dd),
	.w4(32'hbbd919c7),
	.w5(32'h3a88aeb4),
	.w6(32'h3c805850),
	.w7(32'h3ba215e4),
	.w8(32'hbc9cc435),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca714b0),
	.w1(32'h3d50175c),
	.w2(32'h3c7a2071),
	.w3(32'hbc057055),
	.w4(32'h3b3f7c27),
	.w5(32'hbb0fbe8a),
	.w6(32'hbc241d95),
	.w7(32'h3c8d2714),
	.w8(32'h3b1aade4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de8f7),
	.w1(32'hbbda5ef9),
	.w2(32'h3c0d03c3),
	.w3(32'h3c5559b2),
	.w4(32'h3b9a5724),
	.w5(32'h3cf37c27),
	.w6(32'hbc360a9c),
	.w7(32'hbc8e5ec0),
	.w8(32'hbb5b76b0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e3adf),
	.w1(32'hbb71ec06),
	.w2(32'hbd071ba8),
	.w3(32'h3d0117ee),
	.w4(32'hbd1bda99),
	.w5(32'hbd03e99e),
	.w6(32'h3d3e3efb),
	.w7(32'h3c7bb23f),
	.w8(32'hbca796cf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8448f1),
	.w1(32'hbd68e13c),
	.w2(32'hbb80b251),
	.w3(32'h3d580694),
	.w4(32'h3be3500c),
	.w5(32'h3d27943d),
	.w6(32'hbd00104f),
	.w7(32'h3cd1644f),
	.w8(32'hbc9a73c4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac15452),
	.w1(32'hbc0ec9c2),
	.w2(32'h3c884c9f),
	.w3(32'hbb02789c),
	.w4(32'h3c1636e7),
	.w5(32'hbcd15903),
	.w6(32'h3bd09308),
	.w7(32'hbc319324),
	.w8(32'hbd3a0d20),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc741436),
	.w1(32'hb99e6908),
	.w2(32'h3c6141bb),
	.w3(32'hbc98063b),
	.w4(32'h3d6d6991),
	.w5(32'h3dfae022),
	.w6(32'hbc0d8f1b),
	.w7(32'h3bb0d59c),
	.w8(32'h3d23cbc5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300eea),
	.w1(32'hbb9b9ddf),
	.w2(32'h3b488cee),
	.w3(32'h3beeee34),
	.w4(32'h3b7c3fe2),
	.w5(32'h3c4a6ce5),
	.w6(32'h3ca86179),
	.w7(32'h3bc4409d),
	.w8(32'h3cd853c6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ae2c7),
	.w1(32'h3bb2a068),
	.w2(32'hbb48644d),
	.w3(32'hbaa92d40),
	.w4(32'h3ce5e687),
	.w5(32'hbd090530),
	.w6(32'h3dad4313),
	.w7(32'h3bf16e0f),
	.w8(32'hbbbb666f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26eea1),
	.w1(32'hbbb15263),
	.w2(32'h3b8eb515),
	.w3(32'h3a3482f5),
	.w4(32'hbc1724e0),
	.w5(32'h3c8c6d27),
	.w6(32'h3c8b4776),
	.w7(32'h3b2b40a8),
	.w8(32'hb8a2ab4a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68ffed),
	.w1(32'hbc65f67f),
	.w2(32'h3c2800c9),
	.w3(32'h3a3e7da1),
	.w4(32'hbb451b60),
	.w5(32'h3cdd2230),
	.w6(32'hbc121923),
	.w7(32'hbb28d006),
	.w8(32'h3cb102b2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd125d47),
	.w1(32'hbd0460dc),
	.w2(32'hbce2b4f4),
	.w3(32'h3b3b32c4),
	.w4(32'h3cd17c44),
	.w5(32'h3d5860fd),
	.w6(32'h3b3890d8),
	.w7(32'hb9c10518),
	.w8(32'h3c8c2b4f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd6803),
	.w1(32'hbd8bc729),
	.w2(32'hbd32bd2e),
	.w3(32'hbd1da53c),
	.w4(32'h3be78987),
	.w5(32'hbba2c8e0),
	.w6(32'hbd293e5f),
	.w7(32'h3b162c5a),
	.w8(32'h3a3c3d9c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3dce21),
	.w1(32'h3be60bf9),
	.w2(32'hbb90d862),
	.w3(32'hbc0f294e),
	.w4(32'hbd3c6d20),
	.w5(32'hbd50922c),
	.w6(32'h3d359926),
	.w7(32'hbb2b7b77),
	.w8(32'hbc5fe721),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbfdbaa),
	.w1(32'h3cde09e9),
	.w2(32'h3b662a5f),
	.w3(32'h3bda2628),
	.w4(32'hbc13ee99),
	.w5(32'hbc1c47f5),
	.w6(32'h3c6b93eb),
	.w7(32'h3bd31746),
	.w8(32'h3c0db2d8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7a466),
	.w1(32'hbd475c31),
	.w2(32'hbcceca61),
	.w3(32'h3cb2c51d),
	.w4(32'h3d2467f1),
	.w5(32'h3b9256b4),
	.w6(32'h3b79c1b4),
	.w7(32'hbb610b4d),
	.w8(32'h3caa0ad0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b22e9),
	.w1(32'h3b6539bc),
	.w2(32'hbc5b0c5f),
	.w3(32'h3b1d388d),
	.w4(32'h3b14ab66),
	.w5(32'hbbb316c0),
	.w6(32'hbc33cf61),
	.w7(32'h3b06bbee),
	.w8(32'h3b00dc95),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20651d),
	.w1(32'hbc7d70c6),
	.w2(32'hbd162f44),
	.w3(32'hbd1a87dc),
	.w4(32'hbcab7f4e),
	.w5(32'h3c666d74),
	.w6(32'hbd1b7be0),
	.w7(32'h3b9c6026),
	.w8(32'hbcb2f712),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a3cf2),
	.w1(32'h3acbf652),
	.w2(32'hbd052e57),
	.w3(32'h3c3dd70a),
	.w4(32'h3cad5831),
	.w5(32'hbcd0da6d),
	.w6(32'hbc8e8907),
	.w7(32'hbcea3790),
	.w8(32'hbcdd7077),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e319c),
	.w1(32'hbbf5c65f),
	.w2(32'hbc07947b),
	.w3(32'hbbf72086),
	.w4(32'hb7cc0a84),
	.w5(32'h3bf234ff),
	.w6(32'h3c189811),
	.w7(32'hbc9f073f),
	.w8(32'h39f0cad1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d798),
	.w1(32'h3d019f1a),
	.w2(32'h3b8d52ef),
	.w3(32'hbc9af3a9),
	.w4(32'hbb902472),
	.w5(32'hbc15e688),
	.w6(32'h3cad98d1),
	.w7(32'h3b9a4f65),
	.w8(32'h3a29052e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f7c03),
	.w1(32'hbcb181d0),
	.w2(32'hbc6ff0e0),
	.w3(32'h3cc0f606),
	.w4(32'hbc1d63f6),
	.w5(32'h3b26ec1c),
	.w6(32'h3c27367f),
	.w7(32'hbc0187db),
	.w8(32'hbc6404c7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c865a78),
	.w1(32'h3c77ff26),
	.w2(32'hbc1c3645),
	.w3(32'h3bd85ce9),
	.w4(32'hbc0868dc),
	.w5(32'hbc2ead44),
	.w6(32'h3cb59952),
	.w7(32'h3c47fcb5),
	.w8(32'h3ab345a0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d46166e),
	.w1(32'h3ccd3639),
	.w2(32'hbd488e07),
	.w3(32'h3c75707d),
	.w4(32'hbcae8e7b),
	.w5(32'hbdea1803),
	.w6(32'h3d1c524f),
	.w7(32'hb8a0bbe8),
	.w8(32'h3b2a1a9a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2bd83),
	.w1(32'hbc2f1f74),
	.w2(32'hbc4fef67),
	.w3(32'h3c9d8bdb),
	.w4(32'h3bc2ef1d),
	.w5(32'h39006b66),
	.w6(32'h3bcfef46),
	.w7(32'h3c8812b7),
	.w8(32'hbcc6b47f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b4e3c),
	.w1(32'h3d13fd2a),
	.w2(32'h3d508ef9),
	.w3(32'hbb3ac14e),
	.w4(32'h3c8c7f89),
	.w5(32'h3cc549fd),
	.w6(32'hbc4d4b56),
	.w7(32'hbb21b563),
	.w8(32'h3c794543),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93307f),
	.w1(32'hbcccef80),
	.w2(32'hbc94d599),
	.w3(32'hbc0f3551),
	.w4(32'h3d7c34ea),
	.w5(32'h3d2524ce),
	.w6(32'h3c4cf007),
	.w7(32'h3bbc398b),
	.w8(32'h3d174276),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c082edf),
	.w1(32'h3c6f557e),
	.w2(32'hbc08506f),
	.w3(32'h3abea4ba),
	.w4(32'h3cb45d2d),
	.w5(32'hb9ff132c),
	.w6(32'hbb8f9eac),
	.w7(32'h3c64e918),
	.w8(32'hbc536cbe),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befdad3),
	.w1(32'hbc81598d),
	.w2(32'h385448d6),
	.w3(32'h3cb94282),
	.w4(32'h3b6dca59),
	.w5(32'h3c4573e6),
	.w6(32'h3ccff8a7),
	.w7(32'hbc32489b),
	.w8(32'h3cc6250e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3552ed),
	.w1(32'h3a00c8cf),
	.w2(32'h3a9875a7),
	.w3(32'hbc83ae16),
	.w4(32'hbc08807f),
	.w5(32'hba1abede),
	.w6(32'h3c881bf5),
	.w7(32'hbb4f3412),
	.w8(32'hbc10cd3d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979a5a1),
	.w1(32'h396a7aef),
	.w2(32'h3c03300a),
	.w3(32'hbc12fd9f),
	.w4(32'h3c0e24d7),
	.w5(32'h3d02c799),
	.w6(32'hbc52cdf4),
	.w7(32'h3b44719c),
	.w8(32'h3aeae81c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf856b4),
	.w1(32'h3b25f23c),
	.w2(32'hbae82f4c),
	.w3(32'hbaaf134d),
	.w4(32'hbb5bf5fe),
	.w5(32'h3b707ce6),
	.w6(32'hbc0cfe36),
	.w7(32'h3baa1af1),
	.w8(32'hbca24962),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0331a),
	.w1(32'h3bdd9c26),
	.w2(32'h3cd8551e),
	.w3(32'h3ccd6611),
	.w4(32'hbc0ff226),
	.w5(32'h3ac33feb),
	.w6(32'h3beebcc7),
	.w7(32'h3c402cab),
	.w8(32'hbc84c436),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e842),
	.w1(32'h3a46f942),
	.w2(32'hbb53f7d2),
	.w3(32'hbc3b3054),
	.w4(32'h3c55c9dc),
	.w5(32'h3d7f893e),
	.w6(32'h3c1e9052),
	.w7(32'hbb9f6b9f),
	.w8(32'hbc20e478),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc848b5e),
	.w1(32'hbd00763e),
	.w2(32'hbc953935),
	.w3(32'h3bcebef0),
	.w4(32'hbad11d1f),
	.w5(32'h3c8d5803),
	.w6(32'hbc4731f0),
	.w7(32'hbb5f6f37),
	.w8(32'h3b562bcc),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d430072),
	.w1(32'h3c5bec8a),
	.w2(32'h3c879800),
	.w3(32'hbb2eacc9),
	.w4(32'hbc78130b),
	.w5(32'hbceaef42),
	.w6(32'h3d345075),
	.w7(32'h3c6f3415),
	.w8(32'hb9a10084),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8384d),
	.w1(32'h3b99dcd9),
	.w2(32'h3bc16935),
	.w3(32'hb7522630),
	.w4(32'hbc11c398),
	.w5(32'hbc680a33),
	.w6(32'hb8b0ffac),
	.w7(32'h3c1b1931),
	.w8(32'h3c0be96c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca90fb6),
	.w1(32'hba1c7ca5),
	.w2(32'hbb09e7f6),
	.w3(32'h3b045b17),
	.w4(32'hbb8ce21b),
	.w5(32'hbb327e22),
	.w6(32'h3a6340d0),
	.w7(32'h3b279603),
	.w8(32'hbc852f06),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78302a),
	.w1(32'h360a1119),
	.w2(32'hbcf41ef1),
	.w3(32'h3cae73bf),
	.w4(32'h3b89e166),
	.w5(32'hbc95fe02),
	.w6(32'h3ab146a8),
	.w7(32'h3af16e5d),
	.w8(32'hbb9a3d03),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0bf0c),
	.w1(32'hbc1b5122),
	.w2(32'hbbbef9c0),
	.w3(32'h3ba1a107),
	.w4(32'hbcfb2d18),
	.w5(32'hbb3bd35d),
	.w6(32'hba18db85),
	.w7(32'hbc999930),
	.w8(32'hbae25045),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c990eb5),
	.w1(32'hbc16c94b),
	.w2(32'h3c7013a6),
	.w3(32'h3cd5aaf0),
	.w4(32'hbb58dd1b),
	.w5(32'h3cb74c83),
	.w6(32'hbc906da1),
	.w7(32'h3c8045a7),
	.w8(32'h3c97f4bd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc980931),
	.w1(32'hbc821ebc),
	.w2(32'h3c310e7c),
	.w3(32'hba9a8873),
	.w4(32'h3bec6eae),
	.w5(32'h3c7bfff5),
	.w6(32'hbc830402),
	.w7(32'hbcb855fd),
	.w8(32'h3c178fc2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b911b29),
	.w1(32'hbae56c1f),
	.w2(32'hba79ca81),
	.w3(32'h3b81031c),
	.w4(32'hbaaa70d7),
	.w5(32'h3a525293),
	.w6(32'h3a4535d6),
	.w7(32'hbc2d5008),
	.w8(32'hbae17b05),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f272a),
	.w1(32'h3b4cb409),
	.w2(32'h3c5efd7e),
	.w3(32'hb9b3dbeb),
	.w4(32'h3c3c285a),
	.w5(32'h3baa8875),
	.w6(32'hb8911dfb),
	.w7(32'h3c15ac21),
	.w8(32'hbb1b7065),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac92ed),
	.w1(32'h3961d367),
	.w2(32'hbb419896),
	.w3(32'h3c2d4d46),
	.w4(32'hbafe4a16),
	.w5(32'h3cc42266),
	.w6(32'h3c854221),
	.w7(32'h39374880),
	.w8(32'hbbc92d5a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad094e),
	.w1(32'h3bacf283),
	.w2(32'hb899bd87),
	.w3(32'h3be85386),
	.w4(32'hbc3fe5a5),
	.w5(32'h3c27361e),
	.w6(32'h3c8f0944),
	.w7(32'h3b76fead),
	.w8(32'hbc332272),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcc38b),
	.w1(32'h3c8c07c8),
	.w2(32'h3bc40924),
	.w3(32'hbb04c6f1),
	.w4(32'h3cf9f434),
	.w5(32'h3c1ea4dc),
	.w6(32'h3c1cf65a),
	.w7(32'h3917815e),
	.w8(32'h3d3fd2bf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ee447),
	.w1(32'hbd1565f3),
	.w2(32'hbbaac232),
	.w3(32'hbbf8ca7e),
	.w4(32'h3b856b97),
	.w5(32'h3ccda78a),
	.w6(32'hbc3548aa),
	.w7(32'h3cb14f4c),
	.w8(32'h3c184edf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc52d9b),
	.w1(32'h3c295e60),
	.w2(32'h3b9f4fbf),
	.w3(32'hbc72af44),
	.w4(32'hbc175851),
	.w5(32'hbc7650e8),
	.w6(32'h3c306921),
	.w7(32'h3b602f85),
	.w8(32'h3bbcdfa6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29f4b8),
	.w1(32'hbc844e6c),
	.w2(32'h3c5b79fe),
	.w3(32'hba9f89a5),
	.w4(32'h3c58eadd),
	.w5(32'h3cc6fac6),
	.w6(32'hbb03eb14),
	.w7(32'h3ca4da38),
	.w8(32'h3c72dbfc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6b688),
	.w1(32'hbc8e3e97),
	.w2(32'hbbc23023),
	.w3(32'h3cd9e1ad),
	.w4(32'h3d0f3286),
	.w5(32'h3cfb4a0f),
	.w6(32'h3afa05c4),
	.w7(32'hbbfdb165),
	.w8(32'h3ca05106),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d27598d),
	.w1(32'h3c7d7e21),
	.w2(32'h3c8c2c2c),
	.w3(32'hbc9ce097),
	.w4(32'h3cee8faa),
	.w5(32'h3ba8ed71),
	.w6(32'hbc9ff5d0),
	.w7(32'hbb0cf7ef),
	.w8(32'h3c31df68),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc015fa4),
	.w1(32'h3cbd8868),
	.w2(32'hbc8f9005),
	.w3(32'hbc2b7ec8),
	.w4(32'h3c4894ad),
	.w5(32'h3cd3fa52),
	.w6(32'hbc37bab1),
	.w7(32'h3c50b5c1),
	.w8(32'h3bc9a0c6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c0123),
	.w1(32'hbc66589c),
	.w2(32'h3b4e3fb6),
	.w3(32'h39a83eab),
	.w4(32'hbb1a50a6),
	.w5(32'h3a6ac790),
	.w6(32'h3c287bda),
	.w7(32'hbb697f85),
	.w8(32'h3aaabe8e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3df80e91),
	.w1(32'h3c7a1e54),
	.w2(32'h3d18db4e),
	.w3(32'h3d4af30a),
	.w4(32'hbd260f39),
	.w5(32'hbc36a066),
	.w6(32'h3da7b0a0),
	.w7(32'hbbbe53db),
	.w8(32'hbbf7d1ac),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1728f),
	.w1(32'h3c03c30a),
	.w2(32'h3c9518df),
	.w3(32'h3c988150),
	.w4(32'h3b1e3d51),
	.w5(32'h3b7e5ade),
	.w6(32'h3c1b031b),
	.w7(32'h3cf324e0),
	.w8(32'h3c1d269e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe238b0),
	.w1(32'h3a9c183d),
	.w2(32'h3c89edc6),
	.w3(32'h39cc9125),
	.w4(32'hbc119132),
	.w5(32'hbbf9e005),
	.w6(32'hba8b2a58),
	.w7(32'h3bf3423f),
	.w8(32'hba9efbb9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f2e1),
	.w1(32'hbb5ca751),
	.w2(32'hbc43d3b6),
	.w3(32'hbc03dae4),
	.w4(32'hbb847081),
	.w5(32'h3a54e74c),
	.w6(32'h3b2d0ed5),
	.w7(32'h3c3ff5cb),
	.w8(32'h3b2578d6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83845f),
	.w1(32'hbc11e0e5),
	.w2(32'hbbec0592),
	.w3(32'h3bcf565d),
	.w4(32'h3bd58707),
	.w5(32'h3a80caa5),
	.w6(32'hbc04bc3d),
	.w7(32'h3b8c7d86),
	.w8(32'hb919953e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd2cc),
	.w1(32'h3c987d66),
	.w2(32'h3c361d9a),
	.w3(32'h3c1a4f63),
	.w4(32'h3b66441f),
	.w5(32'hbc0a08b0),
	.w6(32'h3bf927a6),
	.w7(32'hbb723e79),
	.w8(32'hbc246c62),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18698a),
	.w1(32'h3c388a2c),
	.w2(32'h3bc93197),
	.w3(32'hba4027ef),
	.w4(32'hbb4a2200),
	.w5(32'h3afc09d5),
	.w6(32'h3c3918fc),
	.w7(32'hbb1a030c),
	.w8(32'h3bb9164b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54f0d2),
	.w1(32'h394d5e86),
	.w2(32'hba31418c),
	.w3(32'hbb56a5ea),
	.w4(32'hbbb12261),
	.w5(32'h3ce26baa),
	.w6(32'h3abebfe4),
	.w7(32'h3bdf330e),
	.w8(32'h3b1212f3),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfc168),
	.w1(32'hbc2c5756),
	.w2(32'h3b5192c4),
	.w3(32'hbc0fc8a0),
	.w4(32'h3bfb5ae2),
	.w5(32'h3c95abd2),
	.w6(32'hbb1d0e9e),
	.w7(32'h3cc1b0b3),
	.w8(32'h3b32ee6b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2901d7),
	.w1(32'h3bbabf54),
	.w2(32'h3b93e344),
	.w3(32'hbb0442f7),
	.w4(32'hbb81165f),
	.w5(32'h3b29700e),
	.w6(32'h3a36ac65),
	.w7(32'h3b84c67d),
	.w8(32'hbb4f267a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd84709),
	.w1(32'hbcd27290),
	.w2(32'h39e53bf9),
	.w3(32'h3b86c354),
	.w4(32'h3b87b496),
	.w5(32'h3d0e534d),
	.w6(32'hbb18cdf1),
	.w7(32'h3c350585),
	.w8(32'h3bf4840e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9d4443),
	.w1(32'h3cad4c64),
	.w2(32'hb9de8aeb),
	.w3(32'h3d86ce26),
	.w4(32'h3c0a2d48),
	.w5(32'hbc6e06c5),
	.w6(32'h3dbac61e),
	.w7(32'h3b928e95),
	.w8(32'h3c1f3d78),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0ce57),
	.w1(32'h3b11ba4f),
	.w2(32'hbaede8e8),
	.w3(32'h39b83410),
	.w4(32'hbb52c5f5),
	.w5(32'hbaddf518),
	.w6(32'h3b28ca66),
	.w7(32'h3ab74c73),
	.w8(32'hb8947812),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa392e0),
	.w1(32'h3bfdb5ee),
	.w2(32'h3bc42de5),
	.w3(32'hbc6d3dfb),
	.w4(32'h3b6e154d),
	.w5(32'h3c0c8790),
	.w6(32'hbc3023b5),
	.w7(32'h39d70605),
	.w8(32'h3ad045eb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc60a97),
	.w1(32'h3ca871f2),
	.w2(32'h3c20f504),
	.w3(32'h3c2ffb58),
	.w4(32'hbc38a1dc),
	.w5(32'h3b058089),
	.w6(32'h3c7497b0),
	.w7(32'h3bd96fde),
	.w8(32'hbbe99551),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2990),
	.w1(32'h3bbc32e2),
	.w2(32'hbc5bcbae),
	.w3(32'h3b1d1f01),
	.w4(32'hbb74ec97),
	.w5(32'h3b28d4e7),
	.w6(32'h3c669783),
	.w7(32'h38d4e1ce),
	.w8(32'h3c589b45),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb6b8f),
	.w1(32'h3bc0c6de),
	.w2(32'h3ba9e27c),
	.w3(32'h3b7178bf),
	.w4(32'hbbce6151),
	.w5(32'h3a43a082),
	.w6(32'h3c41d377),
	.w7(32'h3c2d7ec2),
	.w8(32'hbc239a61),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0907c1),
	.w1(32'hbbbc70e4),
	.w2(32'hbb3fd0bb),
	.w3(32'hbba0ac09),
	.w4(32'h3b625773),
	.w5(32'h3c81e41e),
	.w6(32'hbbcddfef),
	.w7(32'h399b039b),
	.w8(32'h3c10f7b2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e27e98),
	.w1(32'h3b3771d4),
	.w2(32'hb9555d08),
	.w3(32'hbbaa31ee),
	.w4(32'hbc8b593e),
	.w5(32'h3acb17bc),
	.w6(32'hbb1d5e3d),
	.w7(32'hbb652549),
	.w8(32'hbc1de4d8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7fa51),
	.w1(32'hbcc7318c),
	.w2(32'hbc2ac503),
	.w3(32'h3c9d815b),
	.w4(32'h3c8af4f8),
	.w5(32'h3cdf7062),
	.w6(32'hba5f4261),
	.w7(32'hb850f911),
	.w8(32'h3be0cbf4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58167f),
	.w1(32'h3c221bf2),
	.w2(32'hbc4db7f4),
	.w3(32'h3c3191c8),
	.w4(32'hbbe424f6),
	.w5(32'hbb8fe203),
	.w6(32'hba1a253b),
	.w7(32'hbb446d63),
	.w8(32'h3a09a9be),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5eb0a),
	.w1(32'h3ca04448),
	.w2(32'h3beab7ad),
	.w3(32'h3c641517),
	.w4(32'hbb5d21b6),
	.w5(32'h3a63b8e2),
	.w6(32'h3c8572b9),
	.w7(32'h3c88805e),
	.w8(32'hbc71d338),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b692e58),
	.w1(32'hb91757b2),
	.w2(32'h3aef1f7e),
	.w3(32'hbbf451af),
	.w4(32'hbb2c68f8),
	.w5(32'hb9a335ef),
	.w6(32'hbbe702cc),
	.w7(32'h3b703aa7),
	.w8(32'h3be49003),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf63fe5),
	.w1(32'h3c60944f),
	.w2(32'h3b4c038a),
	.w3(32'h3bd9d2f5),
	.w4(32'hbb94afdc),
	.w5(32'hbb7232c1),
	.w6(32'hbb0ff557),
	.w7(32'hbab88293),
	.w8(32'h3b55d23b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026f24),
	.w1(32'hb98bc14e),
	.w2(32'hbbe68bc7),
	.w3(32'hbb06a3ac),
	.w4(32'hbb27c861),
	.w5(32'hbab2b736),
	.w6(32'h3b599e23),
	.w7(32'h3b3605b4),
	.w8(32'h3bd66d07),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35e5d7),
	.w1(32'h3c0b44e6),
	.w2(32'hbc71561d),
	.w3(32'h3c827063),
	.w4(32'h3bc88ff3),
	.w5(32'hba25f3c6),
	.w6(32'hbbdff8fa),
	.w7(32'hbc6fe299),
	.w8(32'h3bab4d2c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f9982),
	.w1(32'hbbf982aa),
	.w2(32'hbc75051a),
	.w3(32'hbb6df900),
	.w4(32'hbb8fa601),
	.w5(32'hbc03150f),
	.w6(32'h3ba04224),
	.w7(32'h3b4ba6c6),
	.w8(32'hbc68dcc7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3ff89),
	.w1(32'hbb1d2ab0),
	.w2(32'h3bbe1265),
	.w3(32'h3c63a446),
	.w4(32'hbbc49796),
	.w5(32'h3c266982),
	.w6(32'h3c9dd542),
	.w7(32'hb90c1098),
	.w8(32'h3b03af62),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532801),
	.w1(32'hbbe009c1),
	.w2(32'hbbecdfe1),
	.w3(32'hbae48fb8),
	.w4(32'hbae38b73),
	.w5(32'hbc451b65),
	.w6(32'hbbfdf4cb),
	.w7(32'hbc388dcd),
	.w8(32'h3c1a76e9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d766155),
	.w1(32'h3c14c493),
	.w2(32'h3bb00f55),
	.w3(32'h3bba59ac),
	.w4(32'hbadcc74e),
	.w5(32'hbbf0ec06),
	.w6(32'h3cb9da08),
	.w7(32'h3c3b0d57),
	.w8(32'hbd264055),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c878d83),
	.w1(32'hbc273ead),
	.w2(32'h3c9c2e2d),
	.w3(32'h3c8cd9a4),
	.w4(32'h3c8f7471),
	.w5(32'h3bfaaf4d),
	.w6(32'h3c9e169a),
	.w7(32'hb9f09559),
	.w8(32'h3c3aa11b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9564ab),
	.w1(32'hbc779239),
	.w2(32'h3b4638ed),
	.w3(32'hbbc86a2c),
	.w4(32'h3c65f6fd),
	.w5(32'h3c6e1ed1),
	.w6(32'h3a6bcd01),
	.w7(32'h3b0abcc0),
	.w8(32'h3cc23257),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e4a3f),
	.w1(32'hbbca4767),
	.w2(32'hbbcfa538),
	.w3(32'hbc0d7243),
	.w4(32'h3c143d13),
	.w5(32'h3c5fefd7),
	.w6(32'h3be9eb4b),
	.w7(32'h3b6313a0),
	.w8(32'h3c856dcd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc176916),
	.w1(32'hbc5205a1),
	.w2(32'h3c6d9a7b),
	.w3(32'hbc7b5c01),
	.w4(32'h3c8c2058),
	.w5(32'h3bbb12b5),
	.w6(32'hbbfcd57e),
	.w7(32'h3b3e4400),
	.w8(32'h3c15f335),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d71604),
	.w1(32'h3b0e505c),
	.w2(32'hbbc04571),
	.w3(32'hbbfa2990),
	.w4(32'hbab7d08c),
	.w5(32'hbba4dcbd),
	.w6(32'hbb93f9e9),
	.w7(32'hbbf293af),
	.w8(32'h3b35924b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c943659),
	.w1(32'hbb59ff8a),
	.w2(32'h3b18817e),
	.w3(32'h3be8ffdc),
	.w4(32'h3ba7874b),
	.w5(32'h3cc31e6c),
	.w6(32'h3c30fd01),
	.w7(32'h3b873ca9),
	.w8(32'h3c2b22a4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914c234),
	.w1(32'hba160ec2),
	.w2(32'hbb691505),
	.w3(32'h3aa62bfb),
	.w4(32'h3d3ae994),
	.w5(32'hbb2c7fac),
	.w6(32'hbb84644b),
	.w7(32'hbb32db4a),
	.w8(32'hbbec710b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf79902),
	.w1(32'hbb18da17),
	.w2(32'hbbfb4354),
	.w3(32'hb75f1c58),
	.w4(32'h3abf1b51),
	.w5(32'hba4ddf81),
	.w6(32'h3c30257e),
	.w7(32'hbbc4d231),
	.w8(32'h3c09c638),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90ded3),
	.w1(32'h3c055d68),
	.w2(32'hbbfb7849),
	.w3(32'hbc255ece),
	.w4(32'hbbc0a465),
	.w5(32'hbc0cc755),
	.w6(32'hba92d45b),
	.w7(32'hbb5c3889),
	.w8(32'h3c7892da),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29d529),
	.w1(32'hbbb205bd),
	.w2(32'h3bb2c30b),
	.w3(32'hbc17425e),
	.w4(32'h3c1acb96),
	.w5(32'h3ca5c4d5),
	.w6(32'h3b135258),
	.w7(32'h3b4e6150),
	.w8(32'h3cf9db98),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f014),
	.w1(32'h3bcfe66a),
	.w2(32'hbb8d653c),
	.w3(32'hbc235b4b),
	.w4(32'hbd01977b),
	.w5(32'hbb6700da),
	.w6(32'h3a250db9),
	.w7(32'hbb6a5fcd),
	.w8(32'hbabb4cd4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c6e18),
	.w1(32'hbbdfe346),
	.w2(32'hbbecd71d),
	.w3(32'hb9f87448),
	.w4(32'hbb4c5d2b),
	.w5(32'hbb6d8cab),
	.w6(32'hb73c1cc9),
	.w7(32'hbc03d5e6),
	.w8(32'h3c2e360a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a6d98),
	.w1(32'h3c739e3d),
	.w2(32'hbca7daed),
	.w3(32'h3c0f5de7),
	.w4(32'hbad3ea47),
	.w5(32'hbb51f4c7),
	.w6(32'h3bd439ea),
	.w7(32'hbbadba15),
	.w8(32'h3c9606b8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0923a),
	.w1(32'h3b477f6b),
	.w2(32'hbc73cc7c),
	.w3(32'h3ca8dbc2),
	.w4(32'h3d0cd828),
	.w5(32'hbb2b1c12),
	.w6(32'hbc4d9ad3),
	.w7(32'h3c62c66b),
	.w8(32'h3c3e5c23),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff3d99),
	.w1(32'hbca6775b),
	.w2(32'hbca6731c),
	.w3(32'h3ac80169),
	.w4(32'hbc6a33f9),
	.w5(32'hbbcca215),
	.w6(32'hbc127366),
	.w7(32'hbc5a5486),
	.w8(32'hbced2288),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf35cf2),
	.w1(32'hbbd354f6),
	.w2(32'h3b0f21e1),
	.w3(32'h3a44e1f6),
	.w4(32'h3b82832f),
	.w5(32'h3bc3bce3),
	.w6(32'hb9e1e20a),
	.w7(32'hbd22ca80),
	.w8(32'hbb9d289a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd14d96),
	.w1(32'hbc475098),
	.w2(32'h3c4be1ac),
	.w3(32'hbbc76c2d),
	.w4(32'h3c33238b),
	.w5(32'h3d0a477c),
	.w6(32'hbcda409a),
	.w7(32'h3b12a10e),
	.w8(32'h3b2a7f6d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc86cf2),
	.w1(32'hbc868e26),
	.w2(32'hbc0e1dec),
	.w3(32'h3d016618),
	.w4(32'h3cf9abdc),
	.w5(32'h3cad7dfd),
	.w6(32'h3d6a2797),
	.w7(32'h3cbde3b3),
	.w8(32'h3d168e95),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc0441),
	.w1(32'hbc1fdca8),
	.w2(32'hbc63b681),
	.w3(32'h3b8414fd),
	.w4(32'hbc7ee430),
	.w5(32'h3b8346b2),
	.w6(32'hbbbb62a5),
	.w7(32'hbc3a8c32),
	.w8(32'hbc32bc91),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac609b8),
	.w1(32'hbb0faced),
	.w2(32'h3a8d2643),
	.w3(32'h3c8b6ce8),
	.w4(32'h3beb83c0),
	.w5(32'hbab055c5),
	.w6(32'hbad9c493),
	.w7(32'h3c4a417e),
	.w8(32'h3bd4babe),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33c05a),
	.w1(32'hbbe2665b),
	.w2(32'h3a40fa23),
	.w3(32'hbb5b3f8d),
	.w4(32'hbb78e101),
	.w5(32'h3a6a9ff6),
	.w6(32'hbbf25f28),
	.w7(32'h3bd7c7af),
	.w8(32'h3d0b7eb3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f055e),
	.w1(32'hb9dafdd9),
	.w2(32'hbb680fd9),
	.w3(32'hbb9419f8),
	.w4(32'hbb3e7e17),
	.w5(32'hbbe66564),
	.w6(32'h37a2b90b),
	.w7(32'hbb2b3bc8),
	.w8(32'hb8e63135),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060508),
	.w1(32'hbd6e8124),
	.w2(32'hbccc2014),
	.w3(32'h3b86b930),
	.w4(32'hbca720ff),
	.w5(32'hba8eb164),
	.w6(32'hbbb1f186),
	.w7(32'h3c66344c),
	.w8(32'hbb81374c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade7bb7),
	.w1(32'hba063f85),
	.w2(32'h3c121ede),
	.w3(32'h3abc3e07),
	.w4(32'h3ad009e3),
	.w5(32'hbb32919a),
	.w6(32'hbc53bb87),
	.w7(32'hbb383682),
	.w8(32'h3a7bec5e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8d84c),
	.w1(32'h3be26a14),
	.w2(32'h3b0b1c77),
	.w3(32'h3c979d67),
	.w4(32'hbc0bd5e0),
	.w5(32'hbb7c2153),
	.w6(32'h3cc259e2),
	.w7(32'h3cdae46b),
	.w8(32'h3bb28da2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2f417),
	.w1(32'h3bcea82f),
	.w2(32'hbac933be),
	.w3(32'h3ba9715d),
	.w4(32'h3b0ffa6c),
	.w5(32'h3ae7f323),
	.w6(32'hbb47d897),
	.w7(32'h3bca0b59),
	.w8(32'hbc1a2f47),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bc6aa),
	.w1(32'hbc98897f),
	.w2(32'h3bbf3f5b),
	.w3(32'h3b963464),
	.w4(32'h3bc19673),
	.w5(32'h3cdeb01b),
	.w6(32'hbbd15f06),
	.w7(32'hbbeb801d),
	.w8(32'hbba2d263),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf750d),
	.w1(32'hbc261f2a),
	.w2(32'hbcb03bd4),
	.w3(32'hbb3714b5),
	.w4(32'hbbfa061a),
	.w5(32'hbbbb462d),
	.w6(32'hb8cc1906),
	.w7(32'h3c00714f),
	.w8(32'hbc8f0bd3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819802),
	.w1(32'hba2fb88f),
	.w2(32'hbc0f2aa9),
	.w3(32'h3a1c0b29),
	.w4(32'hbc297227),
	.w5(32'h3b860919),
	.w6(32'hba3fc5ef),
	.w7(32'hba81d3a6),
	.w8(32'hbae0a11c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b0bf4),
	.w1(32'hbc735d86),
	.w2(32'h3bfd9fa3),
	.w3(32'hbca70552),
	.w4(32'h3c48ead5),
	.w5(32'h3c93997f),
	.w6(32'h3b6c9642),
	.w7(32'h3cb00315),
	.w8(32'h3c32ee82),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada067a),
	.w1(32'hbbdff84b),
	.w2(32'h3b3834d9),
	.w3(32'h3bcc9520),
	.w4(32'hbc1074c5),
	.w5(32'h3a914f64),
	.w6(32'h398edb18),
	.w7(32'h3cf4d654),
	.w8(32'hbb50df50),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21407b),
	.w1(32'hbc83c6c4),
	.w2(32'hbbf46dfe),
	.w3(32'hbc2d53c4),
	.w4(32'h3c164d9e),
	.w5(32'h3b9b5f95),
	.w6(32'hbb22e8e1),
	.w7(32'h3a0b9c7b),
	.w8(32'hbc2c410e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a491f),
	.w1(32'h3bcf248f),
	.w2(32'h3af511b5),
	.w3(32'h3c5631b8),
	.w4(32'h3b5284ae),
	.w5(32'hbc3bc571),
	.w6(32'h3c44e61a),
	.w7(32'hbb062468),
	.w8(32'h3b635a98),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc3966),
	.w1(32'h3ce05581),
	.w2(32'h3c56ab63),
	.w3(32'hbba22c9c),
	.w4(32'h3b93d923),
	.w5(32'hbb92c74b),
	.w6(32'h3b3f0ac7),
	.w7(32'h3bc9d998),
	.w8(32'h3d48ca62),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f868),
	.w1(32'h3c2b6e40),
	.w2(32'hb980bc8d),
	.w3(32'hb9a90241),
	.w4(32'hbd8a5da7),
	.w5(32'h3bbe81b5),
	.w6(32'h3a4bc603),
	.w7(32'hbc296ca7),
	.w8(32'h3b7f2ba3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d18e228),
	.w1(32'h3c7cb056),
	.w2(32'hb9f8f506),
	.w3(32'h3be14248),
	.w4(32'h3af535fd),
	.w5(32'h3b99b237),
	.w6(32'h3d0283a2),
	.w7(32'h3c7dca9f),
	.w8(32'h3b0150aa),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba339300),
	.w1(32'h3a1496c7),
	.w2(32'hbaf8bda2),
	.w3(32'h3c0e1874),
	.w4(32'hb94694cb),
	.w5(32'h3d093060),
	.w6(32'hbc62e7ff),
	.w7(32'hbd2910c6),
	.w8(32'h3bfa93eb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a942921),
	.w1(32'h3c82735e),
	.w2(32'h3bd67f7f),
	.w3(32'h3c2f8ef3),
	.w4(32'h3b8cd329),
	.w5(32'hbcbb56d3),
	.w6(32'h3b668c09),
	.w7(32'h3b1c8542),
	.w8(32'hbbb73146),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc034580),
	.w1(32'h3c95029e),
	.w2(32'hbb323971),
	.w3(32'hbbb07a45),
	.w4(32'hbb7ccbab),
	.w5(32'hbc0db150),
	.w6(32'h3be145de),
	.w7(32'h3b9f6d31),
	.w8(32'hbc116199),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2afb95),
	.w1(32'h3a0565e6),
	.w2(32'h39c4d5e2),
	.w3(32'h3b325160),
	.w4(32'hbb1c87f8),
	.w5(32'hbad6f0ef),
	.w6(32'hbb8f2643),
	.w7(32'h3b0adc48),
	.w8(32'hbb679b1c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccc1e9d),
	.w1(32'h3c64883a),
	.w2(32'h3c8ddc88),
	.w3(32'h3c866364),
	.w4(32'hbb5054aa),
	.w5(32'h3b19d5bf),
	.w6(32'hbbd495e6),
	.w7(32'h3c8251e9),
	.w8(32'h3c9e1903),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92d0a),
	.w1(32'hbb1dcded),
	.w2(32'h3cef5081),
	.w3(32'h3b05a7dd),
	.w4(32'hba9b73a8),
	.w5(32'h3d2ec13e),
	.w6(32'hbcb3fb10),
	.w7(32'h3c30339c),
	.w8(32'h3c025469),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83cf9b),
	.w1(32'h3cc6a3c0),
	.w2(32'h3cf5eb64),
	.w3(32'h3c4b8291),
	.w4(32'h3b6a7a97),
	.w5(32'hbc09f6f5),
	.w6(32'h3c04c765),
	.w7(32'hbb03255b),
	.w8(32'h3c81be5c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc994f4),
	.w1(32'hbca0ff7b),
	.w2(32'hbcafb762),
	.w3(32'h3affb0ad),
	.w4(32'h3ca72eb2),
	.w5(32'h3cbebe68),
	.w6(32'h3c7cfe41),
	.w7(32'h3c035a3f),
	.w8(32'h3c19de4b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2195fb),
	.w1(32'hbb4e6f83),
	.w2(32'hbc25a836),
	.w3(32'hbc52aab2),
	.w4(32'h3bf3aab3),
	.w5(32'hbc17caeb),
	.w6(32'hbb6fcbda),
	.w7(32'h3ae2e61b),
	.w8(32'h3a6b31df),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e03b3),
	.w1(32'hbc55ca30),
	.w2(32'h3c35fe70),
	.w3(32'h3c68e817),
	.w4(32'h3b263c40),
	.w5(32'h3c56b442),
	.w6(32'hbc22720e),
	.w7(32'h3bae666d),
	.w8(32'h3be44442),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e5e0),
	.w1(32'hbcb68cc3),
	.w2(32'h3c37e1d7),
	.w3(32'h3c2299e5),
	.w4(32'hbb9d4c17),
	.w5(32'hbcea5c5d),
	.w6(32'hbcde6675),
	.w7(32'hbc607441),
	.w8(32'hbcb71b87),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1bfb0c),
	.w1(32'hbcaf7983),
	.w2(32'h3bcea85b),
	.w3(32'h3b1f4cd6),
	.w4(32'hbb69d9fc),
	.w5(32'h3cd75e4e),
	.w6(32'hbca70900),
	.w7(32'hbb674b16),
	.w8(32'h3a93429c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc954a31),
	.w1(32'hbcf4132a),
	.w2(32'hbc5532ae),
	.w3(32'h3c9a3f16),
	.w4(32'h3b8b890a),
	.w5(32'h3c576d21),
	.w6(32'hbca1b8d8),
	.w7(32'h3c41e72f),
	.w8(32'hbb34f54b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d39ee51),
	.w1(32'h3c977045),
	.w2(32'h3bde35c2),
	.w3(32'h3cd32721),
	.w4(32'hbc22277e),
	.w5(32'hbca8e25a),
	.w6(32'h3cafe1bb),
	.w7(32'h3ab2b399),
	.w8(32'hba9b67ab),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0ea086),
	.w1(32'h3c518c2c),
	.w2(32'hbc55dcc5),
	.w3(32'h3a4ff042),
	.w4(32'hbbc2aff0),
	.w5(32'hbc8dad67),
	.w6(32'h3cdbdb12),
	.w7(32'h3bb9ebb6),
	.w8(32'hbbc8ddc0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc62d0d),
	.w1(32'hbb9b1d5a),
	.w2(32'h3bb0c7bb),
	.w3(32'h3c11cd65),
	.w4(32'hbbbfe8f4),
	.w5(32'h3c88f1f1),
	.w6(32'h3bcf859a),
	.w7(32'h3bdb3855),
	.w8(32'h3bb8e23c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1367),
	.w1(32'hba57e81c),
	.w2(32'h3b76612a),
	.w3(32'hba66043d),
	.w4(32'h3c487f5b),
	.w5(32'hb982c83e),
	.w6(32'h3bd68474),
	.w7(32'h3c3ccd3a),
	.w8(32'h3b7d472e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7534d9),
	.w1(32'h3b61f74e),
	.w2(32'h3b7dccbe),
	.w3(32'h3c010ab0),
	.w4(32'h3cbf0943),
	.w5(32'hbc205ee6),
	.w6(32'hba42378d),
	.w7(32'h3c4cb268),
	.w8(32'hbc2155a8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a472),
	.w1(32'h3b9785ce),
	.w2(32'hbc0167a2),
	.w3(32'h3d09274f),
	.w4(32'h3b4069a7),
	.w5(32'h3ae94d89),
	.w6(32'hbac479da),
	.w7(32'hbb3b31d1),
	.w8(32'hbac99142),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51ec5e),
	.w1(32'hbc2c53ea),
	.w2(32'hbcaf93a4),
	.w3(32'hbc6e6008),
	.w4(32'hbbadb51a),
	.w5(32'hbbf48dc2),
	.w6(32'h3abae27b),
	.w7(32'hbbd56309),
	.w8(32'h3c31b3f6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6715a0),
	.w1(32'hbba4d08c),
	.w2(32'h3cb73df6),
	.w3(32'h3b1fb27f),
	.w4(32'h3be9c709),
	.w5(32'hbc0c3b96),
	.w6(32'hbc86c9a7),
	.w7(32'h3b21124c),
	.w8(32'h3c4df371),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43626),
	.w1(32'h3c3a9a55),
	.w2(32'h3b543493),
	.w3(32'hbbb01f34),
	.w4(32'h3af51a22),
	.w5(32'hbbad73f5),
	.w6(32'h3b987b75),
	.w7(32'hbd734f29),
	.w8(32'hbc103d4e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a712c),
	.w1(32'hbb41a66c),
	.w2(32'h3ac461f6),
	.w3(32'h3b90d3f9),
	.w4(32'h3a393513),
	.w5(32'h3af2f947),
	.w6(32'h3c3fe987),
	.w7(32'hbb3772f8),
	.w8(32'hb8143bd4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6196d0),
	.w1(32'hbd1b9952),
	.w2(32'hbcdaef89),
	.w3(32'h3bc7b791),
	.w4(32'h3a108c3c),
	.w5(32'h3c897ef6),
	.w6(32'hbd43d6dc),
	.w7(32'hba1336ee),
	.w8(32'hbbeb04b9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f2e92),
	.w1(32'hbc0297da),
	.w2(32'hbc1b1550),
	.w3(32'h3bb5a71e),
	.w4(32'hbbae1aa0),
	.w5(32'h3c2d5cf4),
	.w6(32'hbc2bb135),
	.w7(32'hbb8316df),
	.w8(32'h3b796d0b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a2b8),
	.w1(32'h39874523),
	.w2(32'hbb200c12),
	.w3(32'h3ba533ab),
	.w4(32'hbb4604bc),
	.w5(32'h3b9a573c),
	.w6(32'h3a7a59f2),
	.w7(32'hba0ccfa9),
	.w8(32'hbc2f6ea0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38d716),
	.w1(32'hbcb31841),
	.w2(32'hbc259c15),
	.w3(32'hbaf8e287),
	.w4(32'h3b8b9cdf),
	.w5(32'h3c6711dc),
	.w6(32'hbbcf0987),
	.w7(32'hbc054d0f),
	.w8(32'h3a90fa0f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc670aef),
	.w1(32'h3c616145),
	.w2(32'hba3face4),
	.w3(32'hbbabd2cb),
	.w4(32'h3c580f41),
	.w5(32'hbc4a5d37),
	.w6(32'h3b5fa2ef),
	.w7(32'h3a888acb),
	.w8(32'hbb6df622),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f2682),
	.w1(32'h3b094b5c),
	.w2(32'hbb546fbe),
	.w3(32'h3b65d0e7),
	.w4(32'h3c1568bf),
	.w5(32'hbc160719),
	.w6(32'h3ba56173),
	.w7(32'hbb0bcbf9),
	.w8(32'h3c20b897),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed8366),
	.w1(32'h3a04b5b1),
	.w2(32'h3b0b3239),
	.w3(32'hbb9c622a),
	.w4(32'h3b021b94),
	.w5(32'hbc36afa9),
	.w6(32'h38ab9af1),
	.w7(32'h3c2ec6a6),
	.w8(32'hb8b5f045),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4650f0),
	.w1(32'hbbb1b303),
	.w2(32'hbbf05808),
	.w3(32'hbc11a493),
	.w4(32'hbb9a6ce2),
	.w5(32'h3a20de64),
	.w6(32'h3bf7f9c1),
	.w7(32'h3b4b7821),
	.w8(32'h3aa8d06b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c534890),
	.w1(32'hbbb6bb59),
	.w2(32'hbab21990),
	.w3(32'h3b34ee0c),
	.w4(32'hbbf56c8b),
	.w5(32'hbc185e1f),
	.w6(32'h3c0b770a),
	.w7(32'h3c2c0f26),
	.w8(32'hba88a11f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c631b82),
	.w1(32'hbc53a7cc),
	.w2(32'hbb8c5d06),
	.w3(32'h3ad1c99e),
	.w4(32'h3cf19e86),
	.w5(32'h3d444459),
	.w6(32'h3c80dc9f),
	.w7(32'h3ba97eea),
	.w8(32'h3ca500a0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc990aaf),
	.w1(32'h3a37c63d),
	.w2(32'hbc5b91be),
	.w3(32'hbb0f25d9),
	.w4(32'hbb030028),
	.w5(32'h3c95022f),
	.w6(32'hbb87698f),
	.w7(32'h3d008e3b),
	.w8(32'hbbb1b7a3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd57ee94),
	.w1(32'hbce24d7b),
	.w2(32'hbc16d552),
	.w3(32'h3a690126),
	.w4(32'h3cb39da9),
	.w5(32'h3ccb9b3b),
	.w6(32'hbc0faf12),
	.w7(32'hbca95348),
	.w8(32'h3cc3952c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd2320),
	.w1(32'h39e3a9e6),
	.w2(32'hbc11d489),
	.w3(32'hbb8f08d4),
	.w4(32'h395e4613),
	.w5(32'h3b2004eb),
	.w6(32'h3b0aaaa6),
	.w7(32'h38fe70ff),
	.w8(32'h3a520ea9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872e9a),
	.w1(32'hbba58560),
	.w2(32'h3bc63ae0),
	.w3(32'hbb68186a),
	.w4(32'h3c84d5eb),
	.w5(32'h39cfe323),
	.w6(32'h3ae0d8a5),
	.w7(32'h3b9522ce),
	.w8(32'h3bba5e6d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c76251),
	.w1(32'hbc82ae7c),
	.w2(32'hb938dc29),
	.w3(32'hbc04cb3b),
	.w4(32'hbaa68ffc),
	.w5(32'hbb1f8aa5),
	.w6(32'hbb58f3fd),
	.w7(32'hbc541a19),
	.w8(32'hbcbc71a6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e87d9),
	.w1(32'h378ca0bd),
	.w2(32'h3c015128),
	.w3(32'h3c37194b),
	.w4(32'hba3b6f81),
	.w5(32'hbc026b54),
	.w6(32'hbb83823e),
	.w7(32'hbbd94d72),
	.w8(32'h3c05a7e7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4818d4),
	.w1(32'hbc0c31e1),
	.w2(32'h3bd659f2),
	.w3(32'h3a2a6e62),
	.w4(32'h3ca57211),
	.w5(32'h3d128334),
	.w6(32'h3bbaf22d),
	.w7(32'hbc687105),
	.w8(32'h3c9bead5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc781737),
	.w1(32'h3bc556ad),
	.w2(32'hbb8400af),
	.w3(32'hbb45a929),
	.w4(32'hbbba0535),
	.w5(32'h3b4e1359),
	.w6(32'hbbf34ca0),
	.w7(32'hbc134ceb),
	.w8(32'hbb02ae9b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99476b),
	.w1(32'hba7d3fec),
	.w2(32'hba8e85f0),
	.w3(32'hbb246164),
	.w4(32'hbb8e6e4d),
	.w5(32'hbc221854),
	.w6(32'hbc93f578),
	.w7(32'h3c371e46),
	.w8(32'h3b90e079),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e1f83),
	.w1(32'hbb18d7e6),
	.w2(32'h3b013f7e),
	.w3(32'hbc301598),
	.w4(32'h3b59d119),
	.w5(32'hb816f4c0),
	.w6(32'h3b48fe44),
	.w7(32'h3c133625),
	.w8(32'h3ba93c73),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b455),
	.w1(32'hbc72322b),
	.w2(32'h3baa589b),
	.w3(32'hba4babd5),
	.w4(32'hbbaf180f),
	.w5(32'h3b2e4679),
	.w6(32'hbd695211),
	.w7(32'hbc8481e3),
	.w8(32'h3b911e19),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20e68d),
	.w1(32'h39e1e3e0),
	.w2(32'hba755049),
	.w3(32'hba3e2786),
	.w4(32'hbb3100ba),
	.w5(32'h3bd42502),
	.w6(32'hbbdcc25e),
	.w7(32'hbac9585c),
	.w8(32'h3abb26e9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f65c9),
	.w1(32'h3bb82740),
	.w2(32'hba60468a),
	.w3(32'hbb9f8cfb),
	.w4(32'hbcbd8b83),
	.w5(32'hbb42aeed),
	.w6(32'h3afb11b9),
	.w7(32'hb99ba958),
	.w8(32'hbc1a8189),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc681a7c),
	.w1(32'hbc925910),
	.w2(32'hbb7de327),
	.w3(32'hbb6c9475),
	.w4(32'h3d0736cb),
	.w5(32'h3d681b4e),
	.w6(32'h3caa687e),
	.w7(32'h3b7feabd),
	.w8(32'h3d30b43e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61e963),
	.w1(32'hba2c89b2),
	.w2(32'hbb45e39b),
	.w3(32'hb9e1706e),
	.w4(32'hbbfd98e7),
	.w5(32'hbb9565d7),
	.w6(32'hbb745b8b),
	.w7(32'hbb0c492a),
	.w8(32'hbbc08bf3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b647f),
	.w1(32'h3d1b8dea),
	.w2(32'h3cae69a9),
	.w3(32'hbb194515),
	.w4(32'h3a247223),
	.w5(32'hbc0116f4),
	.w6(32'hbc761ba3),
	.w7(32'h3ccb18f1),
	.w8(32'hbbd53cc9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule