module layer_10_featuremap_243(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3d3a9),
	.w1(32'h3a40ac05),
	.w2(32'h3b880656),
	.w3(32'h3ace8e49),
	.w4(32'h3b823791),
	.w5(32'hbb3a7677),
	.w6(32'hbac1d237),
	.w7(32'h3b5cedbe),
	.w8(32'hbbbebb63),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e846),
	.w1(32'hbb55000c),
	.w2(32'hbb5dc7ac),
	.w3(32'hbaf601f9),
	.w4(32'hbb9b86a0),
	.w5(32'h394b8de7),
	.w6(32'hbad0567e),
	.w7(32'hbb5362d6),
	.w8(32'h3aaec089),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b3b11),
	.w1(32'h3ba8dba4),
	.w2(32'h3bbd9521),
	.w3(32'h3ad69f17),
	.w4(32'h3ab8c3da),
	.w5(32'h3ab71164),
	.w6(32'h3ba91300),
	.w7(32'h3b9c7ec7),
	.w8(32'h3b0e5990),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a451),
	.w1(32'h39d27eb6),
	.w2(32'h3a9c584a),
	.w3(32'hb9f47a14),
	.w4(32'h38d579a3),
	.w5(32'h3b9a9c24),
	.w6(32'hba218827),
	.w7(32'h39f061c6),
	.w8(32'hbb9501fa),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398108d5),
	.w1(32'hbb519d02),
	.w2(32'hbb5500f7),
	.w3(32'h3ab1d781),
	.w4(32'h398c1c74),
	.w5(32'h3ba64616),
	.w6(32'hbc18e84b),
	.w7(32'hbbc482f6),
	.w8(32'h3b772579),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18c3e8),
	.w1(32'h3b40b7ff),
	.w2(32'h3ad4477d),
	.w3(32'h3bb12379),
	.w4(32'h3b8ed686),
	.w5(32'h3b4c6de8),
	.w6(32'h3b34d8d7),
	.w7(32'h3b1c6e13),
	.w8(32'h3b170d25),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b049218),
	.w1(32'h3904b175),
	.w2(32'hba9e0904),
	.w3(32'h3b03db9d),
	.w4(32'h3a30c729),
	.w5(32'h3aa6d7e8),
	.w6(32'h3bd280bf),
	.w7(32'h3b21ea9c),
	.w8(32'hba5ee590),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec0aec),
	.w1(32'h3b0956f7),
	.w2(32'h3bc2ffaa),
	.w3(32'h3bcd3aaf),
	.w4(32'h3b0f00f9),
	.w5(32'h3baa1b9e),
	.w6(32'h3c1e0f82),
	.w7(32'h3c108768),
	.w8(32'h3b919d0a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2645ab),
	.w1(32'hb8511689),
	.w2(32'h3abf6bc8),
	.w3(32'h39aa7e15),
	.w4(32'h3b3bfa4f),
	.w5(32'h3b058467),
	.w6(32'h3a3bd585),
	.w7(32'h3b2d2518),
	.w8(32'h3abd45a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae92c97),
	.w1(32'hbbc6d4ad),
	.w2(32'hbc00a53c),
	.w3(32'h3b0d1ea0),
	.w4(32'hbbb703e3),
	.w5(32'hbba06e7c),
	.w6(32'h3b43da7c),
	.w7(32'hbad1836a),
	.w8(32'h3a6e8c5f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e4704),
	.w1(32'h3a88d8f1),
	.w2(32'h3ac74fde),
	.w3(32'h3b205593),
	.w4(32'h3b4d42ee),
	.w5(32'hbb730439),
	.w6(32'h3a0f76e5),
	.w7(32'h3b037016),
	.w8(32'hbac284d2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290f15),
	.w1(32'hba1b5051),
	.w2(32'hbae78b53),
	.w3(32'h3a1a6023),
	.w4(32'hbbbcb3b3),
	.w5(32'hbc448831),
	.w6(32'h3c034f72),
	.w7(32'hba7a134a),
	.w8(32'hbc352400),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30acad),
	.w1(32'hbc85944a),
	.w2(32'hbc465dcb),
	.w3(32'hbbafb341),
	.w4(32'hbc2757bf),
	.w5(32'hbbf32ed0),
	.w6(32'hbbfee75b),
	.w7(32'hbc09c7fb),
	.w8(32'hbae62a80),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b504727),
	.w1(32'hbb0e6003),
	.w2(32'hbb44c553),
	.w3(32'hbaa43948),
	.w4(32'hbb5b3a87),
	.w5(32'hbb3d8a50),
	.w6(32'h3aa6aaf5),
	.w7(32'hbbae57cd),
	.w8(32'hbb8787b6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d7c8a),
	.w1(32'hbbff07ce),
	.w2(32'hbbc19cba),
	.w3(32'hbb86d58e),
	.w4(32'hbbba5a2c),
	.w5(32'hbba44d28),
	.w6(32'hbb95b76a),
	.w7(32'hbba9f420),
	.w8(32'hbb1b9723),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a288c),
	.w1(32'hbc6125c5),
	.w2(32'hbc38ec20),
	.w3(32'hbbb9e2b0),
	.w4(32'hbc21c421),
	.w5(32'hbaeb1a6a),
	.w6(32'hbb6c1b79),
	.w7(32'hbbf0bbdd),
	.w8(32'hbb139b2c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33272b),
	.w1(32'hba60ba15),
	.w2(32'hbad6f2ea),
	.w3(32'h3ac23b54),
	.w4(32'h3b0513a2),
	.w5(32'hbb18bccc),
	.w6(32'hba526cac),
	.w7(32'hb886fd8a),
	.w8(32'hbb147506),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30561),
	.w1(32'h3a2273f0),
	.w2(32'h3b341adc),
	.w3(32'h3bb28056),
	.w4(32'h3b040c70),
	.w5(32'h3b15350e),
	.w6(32'h3c43322f),
	.w7(32'h3bea989a),
	.w8(32'h3c09bb97),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c85864),
	.w1(32'hbb71a8e9),
	.w2(32'hbb1582e7),
	.w3(32'hb9da12b0),
	.w4(32'hbb35c8aa),
	.w5(32'hbb542a5e),
	.w6(32'h3b6d0d88),
	.w7(32'h3b0e26d1),
	.w8(32'hbb2a7d26),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e917),
	.w1(32'hbb1c1ebe),
	.w2(32'h3ab11f23),
	.w3(32'h3956c617),
	.w4(32'h39a9e737),
	.w5(32'hbb32bd10),
	.w6(32'h3a204c49),
	.w7(32'h3995c1fa),
	.w8(32'hbb293c85),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09222),
	.w1(32'hbbbc6937),
	.w2(32'hbbb9e6ea),
	.w3(32'hbb9da630),
	.w4(32'hbbadcc5c),
	.w5(32'h3bc5f1a9),
	.w6(32'hbba43e65),
	.w7(32'hbb6e16a3),
	.w8(32'h3bc20537),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f6c15),
	.w1(32'h3c0180f2),
	.w2(32'h3bc91895),
	.w3(32'h3bbe9a10),
	.w4(32'h3bcb5a07),
	.w5(32'h3a83b5c7),
	.w6(32'h3b687d70),
	.w7(32'h3b835a08),
	.w8(32'h3aeec3d0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f74c),
	.w1(32'h3c0c6704),
	.w2(32'h39c3a922),
	.w3(32'h3c50918e),
	.w4(32'h3c2ec37d),
	.w5(32'h3bec819a),
	.w6(32'h3cd54753),
	.w7(32'h3ca74051),
	.w8(32'h3c901d13),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb5d5c),
	.w1(32'hbc306ca1),
	.w2(32'hbc76272e),
	.w3(32'hbb8b984a),
	.w4(32'hbc19f623),
	.w5(32'hbc3aef02),
	.w6(32'h39672a29),
	.w7(32'hbc1110a5),
	.w8(32'hbbd43669),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610128),
	.w1(32'hba001983),
	.w2(32'hbb00541a),
	.w3(32'hb9afe34d),
	.w4(32'hbbe74999),
	.w5(32'hba78cdf7),
	.w6(32'hbb9bf6c2),
	.w7(32'hbbb10fef),
	.w8(32'hbb345e0b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa2180),
	.w1(32'hba914b16),
	.w2(32'hbb21c0ae),
	.w3(32'h390a53e3),
	.w4(32'hbad7e19e),
	.w5(32'hbb7ce71e),
	.w6(32'hba556ed4),
	.w7(32'hbb152f10),
	.w8(32'hbb0884db),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad72fa8),
	.w1(32'hbaa99825),
	.w2(32'hbba89cfd),
	.w3(32'hbb109c33),
	.w4(32'hbb8f3e96),
	.w5(32'h3b96407c),
	.w6(32'h3a956096),
	.w7(32'hbb837b25),
	.w8(32'h3b28f104),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45e220),
	.w1(32'h3b926f4b),
	.w2(32'h3bc45198),
	.w3(32'hb8c399eb),
	.w4(32'h3b3aed78),
	.w5(32'h3c002fe4),
	.w6(32'hbc267cce),
	.w7(32'hbb1bae05),
	.w8(32'h3c21c700),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44a1a6),
	.w1(32'h3bf3e4fd),
	.w2(32'h3a36fb1b),
	.w3(32'h3b9a630a),
	.w4(32'h3b977ee9),
	.w5(32'h3b76fe6c),
	.w6(32'h3bdf0851),
	.w7(32'h3b8cc15c),
	.w8(32'h3b88b35d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca839),
	.w1(32'hbb381eb2),
	.w2(32'hbaa3c649),
	.w3(32'h3a2e3ebe),
	.w4(32'hbb28250e),
	.w5(32'h3b1f935d),
	.w6(32'hbb8cb30d),
	.w7(32'hbbab1dd0),
	.w8(32'h3a4dbb21),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e82f1),
	.w1(32'hba8e7191),
	.w2(32'hbb4fa3fd),
	.w3(32'h39ed8035),
	.w4(32'hba202e1a),
	.w5(32'h3a908fa4),
	.w6(32'hbab82a65),
	.w7(32'hbb1ab4b3),
	.w8(32'h3b9639ee),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6738ff),
	.w1(32'h3bc5fb86),
	.w2(32'h3b4fa83a),
	.w3(32'h3ad7d4e9),
	.w4(32'hbac46ef1),
	.w5(32'hbb3c4c35),
	.w6(32'h3b0fd00a),
	.w7(32'h39bf2263),
	.w8(32'hbb1520b1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba99b02),
	.w1(32'hbb40804d),
	.w2(32'hbba70244),
	.w3(32'hbaf42153),
	.w4(32'hbb69bf1b),
	.w5(32'hbb8f4c43),
	.w6(32'hba987e4c),
	.w7(32'hbb16eb75),
	.w8(32'hbae58ff4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63865a),
	.w1(32'hbbd84e77),
	.w2(32'hbbfe7f05),
	.w3(32'hbba5e1a3),
	.w4(32'hbbd81e8c),
	.w5(32'h39bd5162),
	.w6(32'hbbb66428),
	.w7(32'hbc07ab39),
	.w8(32'h3ab98c94),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafd4bd),
	.w1(32'h3a4023a3),
	.w2(32'hba22ccec),
	.w3(32'h3a6de181),
	.w4(32'h39963be4),
	.w5(32'hbbb21c6d),
	.w6(32'hb8b4b720),
	.w7(32'h39664cc7),
	.w8(32'hbb8ed202),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9110d69),
	.w1(32'h3b2d2f3f),
	.w2(32'h3abde4ea),
	.w3(32'hbb172b1c),
	.w4(32'h3a61c2fd),
	.w5(32'hb9b8a16d),
	.w6(32'h3bb3e322),
	.w7(32'h3bb6b527),
	.w8(32'h3a64247f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3623f),
	.w1(32'h3bfce8e6),
	.w2(32'hbb772500),
	.w3(32'hbae7b6df),
	.w4(32'h3bea21d2),
	.w5(32'hbbad1d3d),
	.w6(32'h3b9e4d87),
	.w7(32'h3c7de3e9),
	.w8(32'hbb27a0d7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acafff1),
	.w1(32'h3a29124e),
	.w2(32'h3a5b376e),
	.w3(32'h3a8ff982),
	.w4(32'h3b0707da),
	.w5(32'hbb277d1c),
	.w6(32'h3b42f873),
	.w7(32'h3bd25676),
	.w8(32'h3b3f9053),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574336),
	.w1(32'hbaa37406),
	.w2(32'h3a83f784),
	.w3(32'hbafd7769),
	.w4(32'h378c6de8),
	.w5(32'h3c07b1f6),
	.w6(32'hbb604c7c),
	.w7(32'hbb9e8bae),
	.w8(32'h3bbcd4e7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69426),
	.w1(32'h3bb8e332),
	.w2(32'h3bcc3b5c),
	.w3(32'h3ba89273),
	.w4(32'h3bc764bb),
	.w5(32'h3b0cb23a),
	.w6(32'h3b957d72),
	.w7(32'h3be38f00),
	.w8(32'h3b86d324),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b578d5e),
	.w1(32'hba119283),
	.w2(32'hbb155d41),
	.w3(32'hbb3252cf),
	.w4(32'hbb90e79b),
	.w5(32'h3b87d61d),
	.w6(32'hba836f1f),
	.w7(32'hbb2be2a2),
	.w8(32'h3b2ee06b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8855d8),
	.w1(32'h39ed9720),
	.w2(32'hbb3470d0),
	.w3(32'h3b037e1e),
	.w4(32'hba18c360),
	.w5(32'hbbe93c5b),
	.w6(32'h397595a2),
	.w7(32'hbaa87e41),
	.w8(32'hbb9145a8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2c4a6),
	.w1(32'hbb7692a7),
	.w2(32'hb84b518b),
	.w3(32'hbbea249f),
	.w4(32'hbb9afb47),
	.w5(32'hba8a8d4c),
	.w6(32'hbb8b1444),
	.w7(32'hbb09afa7),
	.w8(32'hbb34e60f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef7cec),
	.w1(32'hbc62660a),
	.w2(32'hbc49fab1),
	.w3(32'hbac36f8b),
	.w4(32'hbc415562),
	.w5(32'h3be8db5f),
	.w6(32'h3b9a5abf),
	.w7(32'hbbcbda51),
	.w8(32'h3c18ad46),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab9c65),
	.w1(32'hbae084a8),
	.w2(32'hbaef8e23),
	.w3(32'h3ab7c904),
	.w4(32'hbb0be41b),
	.w5(32'hbaa24658),
	.w6(32'hbac9445a),
	.w7(32'hba8a8902),
	.w8(32'hbb313777),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00af03),
	.w1(32'hbbe6e37f),
	.w2(32'hbc1c3efa),
	.w3(32'h3b3e3692),
	.w4(32'hbb918002),
	.w5(32'hbb55efb0),
	.w6(32'hbad423de),
	.w7(32'hbba55629),
	.w8(32'hba6862f9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c2d14),
	.w1(32'hbbe43d9c),
	.w2(32'hbc209570),
	.w3(32'hba7bd0cf),
	.w4(32'hbbfc2d44),
	.w5(32'h3b36d894),
	.w6(32'hbb47eb15),
	.w7(32'hbbeb2f78),
	.w8(32'h3b858a1e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63707f),
	.w1(32'h3c6a5ffd),
	.w2(32'h3c1ed012),
	.w3(32'h3ca29f79),
	.w4(32'h3c92f0ff),
	.w5(32'hbbe599fc),
	.w6(32'h3cea20f8),
	.w7(32'h3cabb304),
	.w8(32'hbb06f95b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc55d49),
	.w1(32'hbb8c300c),
	.w2(32'hbb016a21),
	.w3(32'hbb8890f2),
	.w4(32'hbaa86aba),
	.w5(32'h3bda4f2a),
	.w6(32'hbba3bafb),
	.w7(32'hbb2b6152),
	.w8(32'h3b9ba072),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fd63),
	.w1(32'h3b82ae0a),
	.w2(32'h3b137875),
	.w3(32'h3b9a77b8),
	.w4(32'h3b379189),
	.w5(32'h39e43405),
	.w6(32'h3b50de38),
	.w7(32'h3ae91fec),
	.w8(32'hbb4da8f1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe705),
	.w1(32'h3b60118b),
	.w2(32'h3b062b7d),
	.w3(32'h3b4609de),
	.w4(32'h3b9f9dda),
	.w5(32'hbb3b0b34),
	.w6(32'h3a9c0533),
	.w7(32'h3b03ac91),
	.w8(32'hbb1c0a0b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fd0f7),
	.w1(32'hbbf631c4),
	.w2(32'hbba91372),
	.w3(32'hbb6f566d),
	.w4(32'hbbe9b0e2),
	.w5(32'h3bad1ef4),
	.w6(32'hbae6bfb1),
	.w7(32'hbba8aa5d),
	.w8(32'h3c1b3293),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79fab),
	.w1(32'h39d8ef56),
	.w2(32'hbb00b288),
	.w3(32'h3b52e7ff),
	.w4(32'h3a3dcac9),
	.w5(32'h3b446ea5),
	.w6(32'h3baea723),
	.w7(32'h3ae2d0c4),
	.w8(32'h3b3e8302),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab88e15),
	.w1(32'hbb594e30),
	.w2(32'hbacce4ea),
	.w3(32'h3bf05257),
	.w4(32'hbb883df0),
	.w5(32'hbb4943d3),
	.w6(32'h3c975ede),
	.w7(32'h3b8779aa),
	.w8(32'hba7aab3a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc014c31),
	.w1(32'hbb78c33a),
	.w2(32'h39bc4dbf),
	.w3(32'h397238f3),
	.w4(32'hbadba943),
	.w5(32'h3b97cbcd),
	.w6(32'hba13ef6a),
	.w7(32'h3921405d),
	.w8(32'h3ba72d22),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dd1bf),
	.w1(32'h39821fad),
	.w2(32'h38a53b12),
	.w3(32'h3a837a3a),
	.w4(32'h3ae2f592),
	.w5(32'hb92fbc27),
	.w6(32'hbb7594aa),
	.w7(32'hba9861b0),
	.w8(32'h3978f1c2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2afa21),
	.w1(32'hb9114262),
	.w2(32'hbad73c88),
	.w3(32'hbb6258eb),
	.w4(32'hbabfe53b),
	.w5(32'h3b9c88a6),
	.w6(32'hbb8f6388),
	.w7(32'hbb19ccaa),
	.w8(32'h3b84559a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e8d9b),
	.w1(32'h3b333474),
	.w2(32'h3b7462c8),
	.w3(32'h3b1f7c4f),
	.w4(32'h3bacdb07),
	.w5(32'h3bda68a2),
	.w6(32'h3b913bc2),
	.w7(32'h3b87fa89),
	.w8(32'h3ba61d54),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea6d69),
	.w1(32'h3bb9dcfc),
	.w2(32'h3b6a69b5),
	.w3(32'h3b9f8077),
	.w4(32'h3b9d67f7),
	.w5(32'h39908ed6),
	.w6(32'h3b8bcf50),
	.w7(32'h3b828f2b),
	.w8(32'hbb3921c3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2028),
	.w1(32'h3a6035e5),
	.w2(32'h3bbac0a7),
	.w3(32'h3ab960bc),
	.w4(32'h3b97efa9),
	.w5(32'hba6ede3f),
	.w6(32'hbbc5b918),
	.w7(32'h3b1e6376),
	.w8(32'hb9e09ae9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ec516),
	.w1(32'hbaa3a991),
	.w2(32'hbb494987),
	.w3(32'hbab08cae),
	.w4(32'hb949737a),
	.w5(32'h3a0e4c2f),
	.w6(32'h3b0dee0c),
	.w7(32'hbb33ee49),
	.w8(32'hbb3704d8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5e682),
	.w1(32'hbb910c16),
	.w2(32'hbaeb9936),
	.w3(32'h3a2e3acb),
	.w4(32'hbab37b04),
	.w5(32'h3b8dabc5),
	.w6(32'hbb9ec7e3),
	.w7(32'hbb38c932),
	.w8(32'h39b17030),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd533cf),
	.w1(32'hbba11299),
	.w2(32'hbbc2b5a3),
	.w3(32'hb94fe01b),
	.w4(32'hba155e55),
	.w5(32'h3b0b41d2),
	.w6(32'hbb76c6f4),
	.w7(32'hbb91d087),
	.w8(32'h3b1cb35b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b426ce9),
	.w1(32'hba708305),
	.w2(32'hbac7aedd),
	.w3(32'hbab891e3),
	.w4(32'hba36fb50),
	.w5(32'hb8d2b428),
	.w6(32'hbb077402),
	.w7(32'hbacb44ff),
	.w8(32'hba062d50),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ee047),
	.w1(32'hba801ba0),
	.w2(32'hbaacc9f9),
	.w3(32'hba0c2dc9),
	.w4(32'hba162e5b),
	.w5(32'hba20131b),
	.w6(32'h3a0bb8c5),
	.w7(32'hbb03133a),
	.w8(32'hbb0fc903),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012ced),
	.w1(32'hbbac63a7),
	.w2(32'hbb7d1a0d),
	.w3(32'h3af43b62),
	.w4(32'hbb4ec630),
	.w5(32'h3bcd5505),
	.w6(32'hbae9da43),
	.w7(32'hbb0a651f),
	.w8(32'h3b4fb7c2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36779),
	.w1(32'h3932c892),
	.w2(32'h3b067a8b),
	.w3(32'h3bd12f63),
	.w4(32'hbafbc250),
	.w5(32'hbb2a9c82),
	.w6(32'h3b93f2e2),
	.w7(32'h3a2ea02c),
	.w8(32'hbb95366a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab0742),
	.w1(32'hbc1c387e),
	.w2(32'hbc24c340),
	.w3(32'h3b6fbebd),
	.w4(32'hbbc380f3),
	.w5(32'hbb976165),
	.w6(32'h3bcc34fa),
	.w7(32'hbadf0305),
	.w8(32'hb9d16aa1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900006d),
	.w1(32'h3a41fbdb),
	.w2(32'hba813ae5),
	.w3(32'h3bcf4dad),
	.w4(32'h3b09f05b),
	.w5(32'h3bd621e0),
	.w6(32'h3c446fbc),
	.w7(32'h3bc8a8e5),
	.w8(32'h3bc94e6b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e49a5),
	.w1(32'hbc38045b),
	.w2(32'hbc197ff4),
	.w3(32'hba3ce75a),
	.w4(32'hbc5a70e2),
	.w5(32'hbc52177e),
	.w6(32'hb9eeeb0d),
	.w7(32'hbc1e3d81),
	.w8(32'hbbcf53f7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ef156),
	.w1(32'hbaae44c6),
	.w2(32'hba1fe154),
	.w3(32'hbb715f9d),
	.w4(32'hbb370266),
	.w5(32'h3a518782),
	.w6(32'hbace5c6e),
	.w7(32'hba1c9f17),
	.w8(32'hba42700e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa43d9),
	.w1(32'h3a20cf92),
	.w2(32'hba7449db),
	.w3(32'hb8ccda2e),
	.w4(32'hba80c061),
	.w5(32'hbb46807a),
	.w6(32'h3b491997),
	.w7(32'h39ca3d76),
	.w8(32'hbb643589),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b39a2),
	.w1(32'hb7f8d138),
	.w2(32'hba9c9b43),
	.w3(32'hbb5db0a0),
	.w4(32'hb9317757),
	.w5(32'hbb704b93),
	.w6(32'hbacce561),
	.w7(32'h3ade07a2),
	.w8(32'hbb6b44f3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc48ab0),
	.w1(32'hbbd49e16),
	.w2(32'hbbcd4f0e),
	.w3(32'hbb786f11),
	.w4(32'hbb75c3dd),
	.w5(32'h3b686623),
	.w6(32'hbb093f1a),
	.w7(32'hbb74e787),
	.w8(32'h3b83e2cc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affe826),
	.w1(32'h3a44b641),
	.w2(32'h3a95bb03),
	.w3(32'h3bae4f07),
	.w4(32'h3b0cd4ec),
	.w5(32'hbc382c34),
	.w6(32'h3b11fdf3),
	.w7(32'h3a9ee9e8),
	.w8(32'hbc28dcf5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfd054),
	.w1(32'hbbac8fd0),
	.w2(32'hbb09b511),
	.w3(32'hbb883c9b),
	.w4(32'hbac6e73d),
	.w5(32'h3b5b9f82),
	.w6(32'h39bb82b6),
	.w7(32'h3af2d980),
	.w8(32'h3b9be769),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c076036),
	.w1(32'h3ad8f25d),
	.w2(32'h3a9b9bd1),
	.w3(32'h3b9d6168),
	.w4(32'h3bbb75da),
	.w5(32'h3b05522d),
	.w6(32'h3c7cce8f),
	.w7(32'h3c32ac3a),
	.w8(32'h3b6df365),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7fb1b),
	.w1(32'hbc1ea7c1),
	.w2(32'hbc323a8e),
	.w3(32'hbba805d4),
	.w4(32'hbc21a1bc),
	.w5(32'hbc23efd2),
	.w6(32'hbc103bf0),
	.w7(32'hbc373e4b),
	.w8(32'hbc142c77),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b6a7),
	.w1(32'hbbefc2f7),
	.w2(32'hbb2baad6),
	.w3(32'hbb2fb874),
	.w4(32'hbb5939b6),
	.w5(32'h3b07b21f),
	.w6(32'hbb2908aa),
	.w7(32'hb9a69c79),
	.w8(32'h3a8ec694),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b253dc4),
	.w1(32'h3ad61a61),
	.w2(32'hb9992282),
	.w3(32'h3ba151b5),
	.w4(32'h3b93e5e2),
	.w5(32'hbbf779c7),
	.w6(32'h3b1da043),
	.w7(32'h3a6e00e1),
	.w8(32'hbc0bc204),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba631cc),
	.w1(32'hbb9b3b25),
	.w2(32'hbb15cea9),
	.w3(32'hbba9de8f),
	.w4(32'hbbd4aa7d),
	.w5(32'hbbc9e29a),
	.w6(32'hbbb42160),
	.w7(32'hbb3bdf9a),
	.w8(32'hbbe8bfbb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfc98),
	.w1(32'hbb40c52e),
	.w2(32'hbad7c3f4),
	.w3(32'hbaffbaba),
	.w4(32'hbaf8b74f),
	.w5(32'hb8440534),
	.w6(32'h3a780903),
	.w7(32'h39b4071c),
	.w8(32'h3ae424ae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77da9f),
	.w1(32'hb97f3f8b),
	.w2(32'hba3301e1),
	.w3(32'hbb80734c),
	.w4(32'hbb99fa50),
	.w5(32'h3b9ea1b9),
	.w6(32'hb99cf66c),
	.w7(32'hb77643d9),
	.w8(32'h3be0f1f5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1b193),
	.w1(32'hb98131f7),
	.w2(32'hbb5f4780),
	.w3(32'h3ae90ee4),
	.w4(32'hba983a88),
	.w5(32'hbb11563d),
	.w6(32'h3afe3b80),
	.w7(32'hbb73e6ca),
	.w8(32'hbab4a713),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f3709),
	.w1(32'hbb27af37),
	.w2(32'hba80b650),
	.w3(32'hbb301ea5),
	.w4(32'hbb7d28f5),
	.w5(32'h3ab41d7d),
	.w6(32'hba419e8b),
	.w7(32'h39bab43b),
	.w8(32'hba92945c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb253453),
	.w1(32'hb8be8b6d),
	.w2(32'hbae0661b),
	.w3(32'h3b073c17),
	.w4(32'hbb12f405),
	.w5(32'h39da2b6a),
	.w6(32'hbb3d99a4),
	.w7(32'hbb64e112),
	.w8(32'hbad7912f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc73033),
	.w1(32'hbc084671),
	.w2(32'hbc13b181),
	.w3(32'hbb7c6ce5),
	.w4(32'hbbd7f5e6),
	.w5(32'hbb1bbb2b),
	.w6(32'hba4e898f),
	.w7(32'hbbb09f22),
	.w8(32'hbb9ced7f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58588f),
	.w1(32'hbaa46f6a),
	.w2(32'hba6a20d1),
	.w3(32'h3a36e451),
	.w4(32'h38eece32),
	.w5(32'h3ad7f793),
	.w6(32'hbab37636),
	.w7(32'hba8e5c86),
	.w8(32'hb9d9561f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5b1de),
	.w1(32'hbb5be4ad),
	.w2(32'hbb64c116),
	.w3(32'h3ba8e8b0),
	.w4(32'h3b28d6f3),
	.w5(32'h3bbae43e),
	.w6(32'h3b8cbba6),
	.w7(32'h3b057f46),
	.w8(32'h3c067721),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6676c4),
	.w1(32'h3c439f37),
	.w2(32'h3c701228),
	.w3(32'h3c8e8716),
	.w4(32'h3c951f77),
	.w5(32'h3b9a801f),
	.w6(32'h3cbcd836),
	.w7(32'h3cbf3b34),
	.w8(32'h3be3bfe1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a0de6),
	.w1(32'h3afe4d21),
	.w2(32'h3a1a8e18),
	.w3(32'hbb6cdfbc),
	.w4(32'h3a95a717),
	.w5(32'h3b2c3885),
	.w6(32'h3b489c2d),
	.w7(32'hbafbc961),
	.w8(32'h3acee86f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ace2e),
	.w1(32'h3b9c2099),
	.w2(32'hbbde4c17),
	.w3(32'h3c0d4c32),
	.w4(32'hbae69881),
	.w5(32'hbb42c464),
	.w6(32'h3c89a90f),
	.w7(32'hb9f105d1),
	.w8(32'h3a832113),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7b488),
	.w1(32'hbb1fa5cf),
	.w2(32'hbb84b69e),
	.w3(32'hbb40d4dc),
	.w4(32'hbb5e8beb),
	.w5(32'hbb05265f),
	.w6(32'hbb8d6ff9),
	.w7(32'hbb80adf8),
	.w8(32'h39c8229a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6b4be),
	.w1(32'hbc1b0806),
	.w2(32'hbb9dc019),
	.w3(32'hba439c4f),
	.w4(32'hbb5353ec),
	.w5(32'hbb61b552),
	.w6(32'h3be04b08),
	.w7(32'h3b3ee176),
	.w8(32'hbaf03f9b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29215f),
	.w1(32'hbb3a8006),
	.w2(32'hbb10c5f9),
	.w3(32'hbb0733b8),
	.w4(32'hbb79e7af),
	.w5(32'hb9bcd7d3),
	.w6(32'h3ae781aa),
	.w7(32'hbab53526),
	.w8(32'h3b1ca064),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd728),
	.w1(32'hbb31ee10),
	.w2(32'hba34606d),
	.w3(32'hbb8b2f08),
	.w4(32'hbc0a7c01),
	.w5(32'hbba3a3df),
	.w6(32'hb93ad147),
	.w7(32'hbb584d17),
	.w8(32'hbb481211),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeec51),
	.w1(32'h37eb19b6),
	.w2(32'h3b88bad9),
	.w3(32'hbb5b0e26),
	.w4(32'h3b18d6b3),
	.w5(32'h3bdac352),
	.w6(32'hbb6bc367),
	.w7(32'h3b63a134),
	.w8(32'h3b9a1c04),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd077),
	.w1(32'hbb670cd9),
	.w2(32'hbaa3d461),
	.w3(32'h3b90e0a4),
	.w4(32'h3b745e57),
	.w5(32'hbbaa7395),
	.w6(32'h3be9e6a3),
	.w7(32'h3c04cde8),
	.w8(32'h3a524f70),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2ebe0),
	.w1(32'h3b12d78a),
	.w2(32'hbb356803),
	.w3(32'hb983fca5),
	.w4(32'h3987b15b),
	.w5(32'hbb8a8ab1),
	.w6(32'h3c1860c3),
	.w7(32'h3b58e951),
	.w8(32'hbbdc7660),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c578d),
	.w1(32'h3b59459e),
	.w2(32'h37991f01),
	.w3(32'h3baa3a46),
	.w4(32'h3c00518c),
	.w5(32'hbb70b862),
	.w6(32'h3c8a0dcf),
	.w7(32'h3c806c5e),
	.w8(32'h3b638488),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ec83f),
	.w1(32'hbc42df37),
	.w2(32'hbb9c5d8e),
	.w3(32'hbc50163b),
	.w4(32'hbbac0df7),
	.w5(32'h3bdad089),
	.w6(32'hbb860549),
	.w7(32'hbb610954),
	.w8(32'h3b6d95a2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb800b8c8),
	.w1(32'hbb75411a),
	.w2(32'hbba9e78f),
	.w3(32'h3bd2b85a),
	.w4(32'hbb4b02d0),
	.w5(32'hbb52737c),
	.w6(32'hbad67ca5),
	.w7(32'hbc128510),
	.w8(32'hbae3299f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaceae75),
	.w1(32'h3ab253b9),
	.w2(32'hb9c152e5),
	.w3(32'hbac5409b),
	.w4(32'h3aad33b6),
	.w5(32'hbc0bc9a8),
	.w6(32'h3c149016),
	.w7(32'h3be82c6a),
	.w8(32'hbb1ef3d5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b0952),
	.w1(32'hba955e59),
	.w2(32'h3ab036af),
	.w3(32'hbb812ed8),
	.w4(32'h3ad4fad3),
	.w5(32'h3c03bcf3),
	.w6(32'hbb32a864),
	.w7(32'hbac0bae3),
	.w8(32'hbad0b8ff),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5bef),
	.w1(32'h3bdb9905),
	.w2(32'h3bd61aeb),
	.w3(32'h3be0bc8f),
	.w4(32'h3c31c6ec),
	.w5(32'h3b3747a6),
	.w6(32'h3c6489bf),
	.w7(32'h3c917397),
	.w8(32'h3bf681d5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38baa2ba),
	.w1(32'hba066ef8),
	.w2(32'hbb5a848c),
	.w3(32'hbb973a3f),
	.w4(32'hbb8d9951),
	.w5(32'hbab9ce3a),
	.w6(32'hbaf46527),
	.w7(32'hbb66bca1),
	.w8(32'hbbd3cb23),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f2dc8),
	.w1(32'hbabc5b50),
	.w2(32'hbb5a5775),
	.w3(32'hbba58ab4),
	.w4(32'hbac856e6),
	.w5(32'h3b710188),
	.w6(32'hbb4df62e),
	.w7(32'h3ac4c73c),
	.w8(32'h3a271086),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae061c6),
	.w1(32'h3b2ab701),
	.w2(32'h3aa4be8c),
	.w3(32'h3b831658),
	.w4(32'hbb900eb9),
	.w5(32'hb89377e5),
	.w6(32'h3c3b1b62),
	.w7(32'h3af434bc),
	.w8(32'h3a04a673),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987f09),
	.w1(32'h3aaed8d2),
	.w2(32'h3913a62d),
	.w3(32'h3b3f02bc),
	.w4(32'h3b3ee94a),
	.w5(32'h3b00c990),
	.w6(32'h3bb5a27e),
	.w7(32'h3b96ede8),
	.w8(32'h3bbc96dd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf95533),
	.w1(32'h3bca9590),
	.w2(32'h3b3da6ed),
	.w3(32'h3c41a2b8),
	.w4(32'h3b3f780d),
	.w5(32'hbc2d0013),
	.w6(32'h3c0ab727),
	.w7(32'h3b8ce2ad),
	.w8(32'hbc7243b7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37ebea),
	.w1(32'hbc8061ab),
	.w2(32'hbc101258),
	.w3(32'hbc5880d2),
	.w4(32'hbc5413c5),
	.w5(32'h3bc283df),
	.w6(32'hbc9ad64c),
	.w7(32'hbc418ca6),
	.w8(32'h3b41e010),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25d133),
	.w1(32'hbbd295f2),
	.w2(32'hb9480776),
	.w3(32'hbb48163a),
	.w4(32'hbb93eb9b),
	.w5(32'hbb8d215f),
	.w6(32'hbb86912d),
	.w7(32'hba808182),
	.w8(32'hbb91b329),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4d411),
	.w1(32'h3addb172),
	.w2(32'hbb83b0af),
	.w3(32'h3ab9ba34),
	.w4(32'h3a11d497),
	.w5(32'hbb5d162d),
	.w6(32'h3aa2893d),
	.w7(32'h3bafd532),
	.w8(32'h3a1f2de6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1a57e),
	.w1(32'h3acf6dd5),
	.w2(32'h3b6e0f39),
	.w3(32'h392ba964),
	.w4(32'hba190de6),
	.w5(32'h3aa9a548),
	.w6(32'h3b8231ef),
	.w7(32'h3ab29849),
	.w8(32'h3ab15b3f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b57f4),
	.w1(32'hb9074740),
	.w2(32'h3a00efde),
	.w3(32'h3b4c7c51),
	.w4(32'h3aa86c36),
	.w5(32'h3b353442),
	.w6(32'h3babe7cd),
	.w7(32'h3b63609f),
	.w8(32'hba101c99),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb914c14),
	.w1(32'hbaa833e6),
	.w2(32'h3a9e6882),
	.w3(32'hb89b7360),
	.w4(32'hbb9a2498),
	.w5(32'h39e4e7ff),
	.w6(32'hbb708ee4),
	.w7(32'hbba4df84),
	.w8(32'h3b0a046f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad77fbc),
	.w1(32'hbab02dfc),
	.w2(32'hba9ed59c),
	.w3(32'h39a677de),
	.w4(32'hba36ea5f),
	.w5(32'hba536366),
	.w6(32'hb9e31e48),
	.w7(32'hbaaab2a0),
	.w8(32'hbb4eb159),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5bcc),
	.w1(32'hbb36561a),
	.w2(32'hbb0d45fa),
	.w3(32'hbb621818),
	.w4(32'h3aabb59b),
	.w5(32'hbc0cebf7),
	.w6(32'h3aaaeaa3),
	.w7(32'hba7c56c5),
	.w8(32'hbb8dc2e4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb04b6),
	.w1(32'h3a9c304e),
	.w2(32'hbb219a17),
	.w3(32'hbaa00f8f),
	.w4(32'hbafb19cd),
	.w5(32'h3ae6e955),
	.w6(32'h3b1ff2a3),
	.w7(32'h38ca3245),
	.w8(32'h3b4365b4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53f6b2),
	.w1(32'h3a4c7adf),
	.w2(32'h3b202949),
	.w3(32'h3a9b7f0d),
	.w4(32'h3b5d45ae),
	.w5(32'h3a8c19c5),
	.w6(32'h3b4bb351),
	.w7(32'h3bbac85f),
	.w8(32'h3a13605c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb130312),
	.w1(32'hbb2943b1),
	.w2(32'h3b023bde),
	.w3(32'hbb5404f1),
	.w4(32'hbb525225),
	.w5(32'hbaab1ad0),
	.w6(32'hbb1bd94c),
	.w7(32'hbaa25cec),
	.w8(32'h3a60e06a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c3f62),
	.w1(32'hbc00c4c1),
	.w2(32'hba8fb81b),
	.w3(32'hbaf8ea7b),
	.w4(32'hbb526dff),
	.w5(32'hbb89a689),
	.w6(32'hbba1d490),
	.w7(32'hba9d69c3),
	.w8(32'h3bcf6121),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa81157),
	.w1(32'hbaca70f4),
	.w2(32'hbb7f73bf),
	.w3(32'h3b107797),
	.w4(32'h3bb86a17),
	.w5(32'hbbb51cf0),
	.w6(32'hba78268a),
	.w7(32'hbbae9602),
	.w8(32'hbc334f2f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd22d54),
	.w1(32'hbc0e242d),
	.w2(32'hbc008b17),
	.w3(32'hbbf56296),
	.w4(32'hbc363c13),
	.w5(32'hbbec22c2),
	.w6(32'hbc716bfc),
	.w7(32'hbc2d1bb9),
	.w8(32'h3b0cf8ab),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b0be),
	.w1(32'h399e371f),
	.w2(32'hbb69f24f),
	.w3(32'h3a44e372),
	.w4(32'h3af4a2b2),
	.w5(32'h3613ad5d),
	.w6(32'h3b6a92aa),
	.w7(32'h3b322dbc),
	.w8(32'hbb8af8b4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb356295),
	.w1(32'hbb91ff3f),
	.w2(32'hbaeef8f7),
	.w3(32'hbb02d1d5),
	.w4(32'hbaa2ccf4),
	.w5(32'h3af8b774),
	.w6(32'hbb993dee),
	.w7(32'hbb12f7cd),
	.w8(32'h3bb24618),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b6001),
	.w1(32'h3b6e1a7c),
	.w2(32'h3b979007),
	.w3(32'h3b5015e9),
	.w4(32'h3add5370),
	.w5(32'hbb9719b0),
	.w6(32'h3bf0829c),
	.w7(32'h3bde16a9),
	.w8(32'hbb40a9f9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a217ce5),
	.w1(32'hb960a058),
	.w2(32'hbb721861),
	.w3(32'h3b8cf757),
	.w4(32'h3a00d533),
	.w5(32'hbb342643),
	.w6(32'h3c2585a4),
	.w7(32'h3b5d3b71),
	.w8(32'h3c354384),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd34da4),
	.w1(32'h3c07ff50),
	.w2(32'h3b910d57),
	.w3(32'h3bebaad2),
	.w4(32'h3ab770d1),
	.w5(32'hbc175db0),
	.w6(32'h3c6db326),
	.w7(32'h3c89f2d1),
	.w8(32'hbab4f7ff),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a872b),
	.w1(32'hba0f7c13),
	.w2(32'hbb268a74),
	.w3(32'h3957f299),
	.w4(32'h3aa0d796),
	.w5(32'h393bca36),
	.w6(32'h3b8c7dd9),
	.w7(32'h3b393abf),
	.w8(32'h3ab60562),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3031c9),
	.w1(32'h3a739b07),
	.w2(32'hbb000153),
	.w3(32'h3b493162),
	.w4(32'hb9fd724d),
	.w5(32'hb9fd1985),
	.w6(32'h3bcd6a85),
	.w7(32'h3ab85a2a),
	.w8(32'hbac4f153),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb0c98),
	.w1(32'hbb8bc16e),
	.w2(32'h3941bd37),
	.w3(32'hbb24ff06),
	.w4(32'hb9f5b56e),
	.w5(32'h367f6ee2),
	.w6(32'hbb6c2fb0),
	.w7(32'h39f60f25),
	.w8(32'hbbd6390e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09d379),
	.w1(32'h3b374dc0),
	.w2(32'h3bab717b),
	.w3(32'h3bad03df),
	.w4(32'h3b92ae71),
	.w5(32'h3b965517),
	.w6(32'hbbc4b298),
	.w7(32'hba6b3c50),
	.w8(32'h3bf22209),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803030),
	.w1(32'h39b7edd3),
	.w2(32'h3b8ef9c8),
	.w3(32'h3a80f542),
	.w4(32'h3a6faa5d),
	.w5(32'h3b73f61e),
	.w6(32'h3b48df32),
	.w7(32'h3b99e9eb),
	.w8(32'h3bb7b44f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea474e),
	.w1(32'h3b18928f),
	.w2(32'h3be26642),
	.w3(32'h3c1e5623),
	.w4(32'h3bb55a67),
	.w5(32'h3bac9792),
	.w6(32'h3c849c86),
	.w7(32'h3c8540a0),
	.w8(32'h3c7727c3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b9bfb),
	.w1(32'h3c02ea8a),
	.w2(32'h3ab35c05),
	.w3(32'h3c0b756b),
	.w4(32'h3c045fe5),
	.w5(32'hbb44a9a9),
	.w6(32'h3c6da097),
	.w7(32'h3c51ac1d),
	.w8(32'hba4c30d6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2832b7),
	.w1(32'hba2a6edd),
	.w2(32'hbb72b5fe),
	.w3(32'h3a82b333),
	.w4(32'hbb4063fd),
	.w5(32'h3b6b0a92),
	.w6(32'h3ba6270f),
	.w7(32'h3b491114),
	.w8(32'h3c1602f9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3a8d8),
	.w1(32'h3b4576a0),
	.w2(32'h3bb17b25),
	.w3(32'h3bc7134e),
	.w4(32'h3be5398c),
	.w5(32'h3b59b0c0),
	.w6(32'h3c5e06d5),
	.w7(32'h3c4d0ddc),
	.w8(32'h3c079c8b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b89b7),
	.w1(32'hbbb36d69),
	.w2(32'h3b281117),
	.w3(32'hbb281616),
	.w4(32'h39cf4814),
	.w5(32'hbb1f143d),
	.w6(32'h3a950554),
	.w7(32'h3bd3c32e),
	.w8(32'hbae1169a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc04ee),
	.w1(32'hbb61fe81),
	.w2(32'hbb1ffd8e),
	.w3(32'hbafff1e7),
	.w4(32'hbb488772),
	.w5(32'hbb72407d),
	.w6(32'h3b6a81e9),
	.w7(32'hbb228d84),
	.w8(32'hbb569069),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7aec6),
	.w1(32'hbac5981d),
	.w2(32'hbb941db1),
	.w3(32'hbb997eb4),
	.w4(32'hbaaf88e8),
	.w5(32'h3ab0a2e2),
	.w6(32'hbbaac7a1),
	.w7(32'hbbbfb3a9),
	.w8(32'h3a95d549),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b6309),
	.w1(32'hb5a946e8),
	.w2(32'hbb7056fb),
	.w3(32'h3ae2f16b),
	.w4(32'hbb63a608),
	.w5(32'hbc24cc0c),
	.w6(32'hbba879e1),
	.w7(32'hbb1d11a1),
	.w8(32'hbc1b7be5),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08e21),
	.w1(32'hbc142097),
	.w2(32'hbb2c6e55),
	.w3(32'hbc35d192),
	.w4(32'hbbd08290),
	.w5(32'h3b6c330f),
	.w6(32'hbc78b5d0),
	.w7(32'hbbc45dc4),
	.w8(32'h3b9cecbb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e83aa),
	.w1(32'h3aa96ab6),
	.w2(32'h3b9fb4b5),
	.w3(32'hbb149b33),
	.w4(32'h3b45b512),
	.w5(32'h3ab41247),
	.w6(32'hbc1e210b),
	.w7(32'h3af20588),
	.w8(32'hbaf54ddd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad9a1e),
	.w1(32'h3c12f128),
	.w2(32'h3b9e5ba9),
	.w3(32'h3b17b4cc),
	.w4(32'hbb8cf7f4),
	.w5(32'hba56d5c5),
	.w6(32'h3c318bbd),
	.w7(32'h3b1fc365),
	.w8(32'hb882de77),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b303d),
	.w1(32'h3aeaef49),
	.w2(32'hbb1c89a3),
	.w3(32'hba1878bb),
	.w4(32'hbb7d7945),
	.w5(32'hbb910b24),
	.w6(32'h3b33604b),
	.w7(32'hbacacc76),
	.w8(32'hbbae76d9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee5e80),
	.w1(32'hbb87d218),
	.w2(32'hbae7d40f),
	.w3(32'hbbba125a),
	.w4(32'hbbc29438),
	.w5(32'hbbc3bf4c),
	.w6(32'hbb77f941),
	.w7(32'hbba1ffcf),
	.w8(32'hbbb81bb7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc34a0f),
	.w1(32'hbb8b57ce),
	.w2(32'hbbe2b95e),
	.w3(32'h3aef95e7),
	.w4(32'hbbd33c6b),
	.w5(32'hbbc11d25),
	.w6(32'h3b5072e1),
	.w7(32'hbb0f7809),
	.w8(32'hbb81b882),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238e93),
	.w1(32'hbb3b8a73),
	.w2(32'hba822091),
	.w3(32'hbb252701),
	.w4(32'hb79ce41c),
	.w5(32'hbad9ea7f),
	.w6(32'hbc3fa5a8),
	.w7(32'hbb922bd5),
	.w8(32'hbb0de4a2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06db3c),
	.w1(32'hbb9b1c93),
	.w2(32'hbbd30bf4),
	.w3(32'hb9926d5e),
	.w4(32'hbbf70296),
	.w5(32'hbb51df92),
	.w6(32'h3b2822f8),
	.w7(32'hbb417f41),
	.w8(32'hbb6f6fb9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6fee9),
	.w1(32'hb908543b),
	.w2(32'hb92b98f5),
	.w3(32'h3b77af3c),
	.w4(32'hbb817e46),
	.w5(32'h3b03a9ff),
	.w6(32'h3b45c29d),
	.w7(32'h3996191f),
	.w8(32'h3beb022c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0ff46),
	.w1(32'hb926636b),
	.w2(32'h39955a62),
	.w3(32'hbb83a044),
	.w4(32'h3b8a2c90),
	.w5(32'hba2c87bf),
	.w6(32'h3b1b286f),
	.w7(32'h3c232344),
	.w8(32'hbbe4355a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ffcdc),
	.w1(32'hbb600634),
	.w2(32'h3a5923c3),
	.w3(32'hbafe63e3),
	.w4(32'hbb4dcedf),
	.w5(32'h3bce4b29),
	.w6(32'hbbd73f69),
	.w7(32'hbc053861),
	.w8(32'hba86f7f5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08ef8b),
	.w1(32'hbb8d59e9),
	.w2(32'h3af4df70),
	.w3(32'hbc0218f6),
	.w4(32'hbbe61add),
	.w5(32'h39dec8da),
	.w6(32'hbc254d91),
	.w7(32'hbb808c34),
	.w8(32'h38d4d6c9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84efeb),
	.w1(32'hbb1efce9),
	.w2(32'h3b6089ff),
	.w3(32'hbaaf0962),
	.w4(32'h3b78c16b),
	.w5(32'h3b833699),
	.w6(32'hbb32c5e8),
	.w7(32'h3b8a84b6),
	.w8(32'h3ba9b6e5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92fa9e),
	.w1(32'h3b42406c),
	.w2(32'hbb4c37f6),
	.w3(32'h38f32047),
	.w4(32'hbbb6f831),
	.w5(32'hbb4a8df6),
	.w6(32'hbb259135),
	.w7(32'hbba98d2b),
	.w8(32'hbb6a3516),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f676),
	.w1(32'h3a301145),
	.w2(32'h3a5965e2),
	.w3(32'hbb441f2a),
	.w4(32'hbbb92c5b),
	.w5(32'h3a096349),
	.w6(32'hbb119533),
	.w7(32'hbb600746),
	.w8(32'hb78782f6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27e716),
	.w1(32'h3903a7c0),
	.w2(32'h3b992bb2),
	.w3(32'h3a9f6f8d),
	.w4(32'hb91d2be0),
	.w5(32'hb9d7e830),
	.w6(32'hbb68e050),
	.w7(32'h382d562a),
	.w8(32'h3bbaa04d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a833723),
	.w1(32'hbba38b89),
	.w2(32'hba1121ef),
	.w3(32'h3c307f12),
	.w4(32'h3c4a6a68),
	.w5(32'hbb337c64),
	.w6(32'h3b40219a),
	.w7(32'hb9a3544d),
	.w8(32'hbb488408),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af27f42),
	.w1(32'hbb8749f9),
	.w2(32'hbb50c9f0),
	.w3(32'hbbaa3f5b),
	.w4(32'hbbfb9a56),
	.w5(32'h3ac6c8e4),
	.w6(32'hbbc4ec35),
	.w7(32'hbc030d25),
	.w8(32'hbb6cd30b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb881c85),
	.w1(32'h3a7cd93f),
	.w2(32'hbad28046),
	.w3(32'h3a64bb6b),
	.w4(32'hbb47ff8e),
	.w5(32'hba9549e4),
	.w6(32'h3b78e4d6),
	.w7(32'h3b06927e),
	.w8(32'h3a066860),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96acd67),
	.w1(32'h3bb81bbe),
	.w2(32'h3b0e1a79),
	.w3(32'hb96decd4),
	.w4(32'hba932c24),
	.w5(32'h3a16d376),
	.w6(32'h3b124354),
	.w7(32'h393c6b7b),
	.w8(32'hbb5f5b20),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99446dd),
	.w1(32'h3abe16fc),
	.w2(32'h3a99abe8),
	.w3(32'hbb45f129),
	.w4(32'hbbf2e161),
	.w5(32'h3b0d725b),
	.w6(32'hbb21195b),
	.w7(32'hbb805690),
	.w8(32'h3b6b1a0c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a3ad1),
	.w1(32'h3b6977eb),
	.w2(32'h3b6a9435),
	.w3(32'hb954167d),
	.w4(32'hbb74d249),
	.w5(32'h39f43e3a),
	.w6(32'h3b22310e),
	.w7(32'h3ae75317),
	.w8(32'hbbeb6341),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19afbe),
	.w1(32'h3aa03564),
	.w2(32'hba852c0f),
	.w3(32'h3b513973),
	.w4(32'hba62e706),
	.w5(32'hbae78948),
	.w6(32'h3b87cebd),
	.w7(32'hbb068fb1),
	.w8(32'h3b2531ed),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac54b5c),
	.w1(32'hbc01b6cf),
	.w2(32'h3a8e7556),
	.w3(32'hbbdab3ae),
	.w4(32'h3b3b9b26),
	.w5(32'hbb01fadb),
	.w6(32'hbc2ea226),
	.w7(32'h3a94fcfc),
	.w8(32'hbb390d1b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e907bc),
	.w1(32'hb9c79b46),
	.w2(32'hbb997fba),
	.w3(32'h3b7e411a),
	.w4(32'h39c7dbfb),
	.w5(32'hbb8450dd),
	.w6(32'h3a910bc7),
	.w7(32'h3b520148),
	.w8(32'hbb5d9e60),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf88fdd),
	.w1(32'hbb8d1326),
	.w2(32'hbb67d06c),
	.w3(32'hbb67b619),
	.w4(32'hbbb45483),
	.w5(32'hbb02d1f4),
	.w6(32'h39ba2aca),
	.w7(32'h3a2d7ce3),
	.w8(32'hba435afe),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96db4d0),
	.w1(32'h39a94e33),
	.w2(32'hbad683fa),
	.w3(32'h3bbd62e2),
	.w4(32'hbb96d448),
	.w5(32'h3b797423),
	.w6(32'h3c5ab977),
	.w7(32'h3ad4baaa),
	.w8(32'h3c058d93),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad89f8),
	.w1(32'h3b90ed6f),
	.w2(32'h3b968b57),
	.w3(32'h3a88a69a),
	.w4(32'h3aeb040a),
	.w5(32'h3abe7850),
	.w6(32'h3bb83bc6),
	.w7(32'h3b944362),
	.w8(32'h3bda27c9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e724b),
	.w1(32'hbc0ab792),
	.w2(32'hbbd1c2dc),
	.w3(32'h3ab854bf),
	.w4(32'h3b70da88),
	.w5(32'h3a8aca9d),
	.w6(32'h3b1e9189),
	.w7(32'h3b2e0acb),
	.w8(32'h3bf32394),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a9c1b),
	.w1(32'h3b6cc7a1),
	.w2(32'h3a81fc93),
	.w3(32'h3aa3dc4d),
	.w4(32'h3b0664ac),
	.w5(32'hbb937535),
	.w6(32'h3b85ac83),
	.w7(32'h3b4e736d),
	.w8(32'hbb8bde1f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1c5e),
	.w1(32'hbc0da7d2),
	.w2(32'hbbd4977b),
	.w3(32'hbbae250e),
	.w4(32'hbc19d911),
	.w5(32'hbb5abde2),
	.w6(32'hbafe4c4d),
	.w7(32'hbbcee73a),
	.w8(32'hbb13ba8f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3fe3),
	.w1(32'hbb69a802),
	.w2(32'h39b3ba41),
	.w3(32'h3b921213),
	.w4(32'hbbacf031),
	.w5(32'hbba41701),
	.w6(32'h3c5a313e),
	.w7(32'h3b70d214),
	.w8(32'hbb09db4f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb497d26),
	.w1(32'hbbd59f28),
	.w2(32'hbb59c942),
	.w3(32'hbb815e17),
	.w4(32'hbb829012),
	.w5(32'hbb257b61),
	.w6(32'h3ade1c82),
	.w7(32'h39f2d0da),
	.w8(32'hbb4cdc52),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090ee2),
	.w1(32'h399cc322),
	.w2(32'hb9b68a3f),
	.w3(32'h39b0f8ac),
	.w4(32'hba838ec9),
	.w5(32'hbab0b80f),
	.w6(32'hbb0d78de),
	.w7(32'h3a188fc2),
	.w8(32'h3bddf277),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebe413),
	.w1(32'hbba949b8),
	.w2(32'hbbe2892d),
	.w3(32'hbae3ab1b),
	.w4(32'hbbc8a2d2),
	.w5(32'hbbe29839),
	.w6(32'h3a65a91d),
	.w7(32'hbbbc5ce3),
	.w8(32'hbc047d3a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc34e),
	.w1(32'hbb726290),
	.w2(32'hbb0577cf),
	.w3(32'hbba2ada9),
	.w4(32'hbb18cb42),
	.w5(32'h3ba6b732),
	.w6(32'hbc1f9ccd),
	.w7(32'hbb5b2dfb),
	.w8(32'h3af39dc6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d712a),
	.w1(32'h3b4f079e),
	.w2(32'h3987f638),
	.w3(32'h3b9e08a4),
	.w4(32'hbb24e84c),
	.w5(32'hbb62c778),
	.w6(32'h3b4938b9),
	.w7(32'hbb610d60),
	.w8(32'hbb1a20cc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a463),
	.w1(32'hbabcf565),
	.w2(32'hbb077782),
	.w3(32'hbb46ca6e),
	.w4(32'hba924468),
	.w5(32'h3b9f58a5),
	.w6(32'hbac0d59c),
	.w7(32'hba677f4e),
	.w8(32'h3b9820b4),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa28ec5),
	.w1(32'hbc1bafa3),
	.w2(32'hbaf66738),
	.w3(32'hbb7f7c94),
	.w4(32'hbbdd8c8e),
	.w5(32'hbac146f6),
	.w6(32'hba8b630e),
	.w7(32'hbb23acd8),
	.w8(32'hbb95531a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d220),
	.w1(32'h3a5a2b1a),
	.w2(32'h3bc7fa28),
	.w3(32'h3b3721c9),
	.w4(32'hba65f578),
	.w5(32'hb94d9cbe),
	.w6(32'h3b96bf9f),
	.w7(32'h3b8a69a7),
	.w8(32'hb92b36e1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e67f4a),
	.w1(32'h3a44fd0a),
	.w2(32'hba1463a9),
	.w3(32'h3aa4f6ae),
	.w4(32'h38ed5058),
	.w5(32'hbb74df23),
	.w6(32'hb7953a9f),
	.w7(32'h3a90c217),
	.w8(32'hbb56c638),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb914da32),
	.w1(32'h3a9301d1),
	.w2(32'h3b3d4236),
	.w3(32'hbaf61982),
	.w4(32'hbb4bf722),
	.w5(32'hbb0bb6f2),
	.w6(32'hbb33a736),
	.w7(32'hbb0d686c),
	.w8(32'hbb9a43d0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7968fb),
	.w1(32'hba065ec3),
	.w2(32'hbbc7811e),
	.w3(32'hbb108651),
	.w4(32'hbbc49890),
	.w5(32'hbaec6437),
	.w6(32'h3b3ccb3c),
	.w7(32'hbb94d731),
	.w8(32'hbb1950ea),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f13f2),
	.w1(32'h3bc8003b),
	.w2(32'h3a8829c9),
	.w3(32'h3a6066d1),
	.w4(32'h3add2b1a),
	.w5(32'hbb8b39c5),
	.w6(32'h3be2e43b),
	.w7(32'h3ba39708),
	.w8(32'hbbfc51b2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44d1bf),
	.w1(32'hbb023c86),
	.w2(32'hbaaca2a8),
	.w3(32'hbaed7c64),
	.w4(32'hbac91f4a),
	.w5(32'h38d79cb9),
	.w6(32'hbc04f82b),
	.w7(32'hbae02fa1),
	.w8(32'hbae9a2c6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a23b3),
	.w1(32'hbb83a6eb),
	.w2(32'hbc50a0a1),
	.w3(32'h3c418fef),
	.w4(32'hbc2a2f56),
	.w5(32'hbc8fa080),
	.w6(32'h3c9c1d4f),
	.w7(32'hbbf261e9),
	.w8(32'hbc926871),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08806e),
	.w1(32'hbc1c84af),
	.w2(32'hbc0f06d8),
	.w3(32'hbc242bd3),
	.w4(32'hbc8803c1),
	.w5(32'h3ac6dcd2),
	.w6(32'hbc904aa1),
	.w7(32'hbc362398),
	.w8(32'h3a326213),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f9c8a),
	.w1(32'h3a7f681d),
	.w2(32'h3a9a559d),
	.w3(32'hba3594a3),
	.w4(32'hbb25fd37),
	.w5(32'h3b79f0c8),
	.w6(32'hbaae53ba),
	.w7(32'h3b0b7593),
	.w8(32'hbb4bf3f1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa38ebe),
	.w1(32'hbb0d2ec5),
	.w2(32'hba9e7c9b),
	.w3(32'h3adb6e0f),
	.w4(32'hb80b827a),
	.w5(32'h37ca57ac),
	.w6(32'hbb814af7),
	.w7(32'hbb7dd766),
	.w8(32'hbb08ff50),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9570fd),
	.w1(32'h39fa26d6),
	.w2(32'h3ae378fb),
	.w3(32'hbb176381),
	.w4(32'hbb48c77b),
	.w5(32'h3b733bd6),
	.w6(32'hbb347c29),
	.w7(32'hbaf0b99f),
	.w8(32'h3b1b89ea),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61eb8a),
	.w1(32'h39f3e7f2),
	.w2(32'hb999036e),
	.w3(32'h3af1db83),
	.w4(32'h3a299a53),
	.w5(32'h3999ac58),
	.w6(32'hbb9b777d),
	.w7(32'h3addc647),
	.w8(32'hbacfb717),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27f3eb),
	.w1(32'hbaff7d52),
	.w2(32'hbb18d917),
	.w3(32'h3a31e9a3),
	.w4(32'hb9f3cb2f),
	.w5(32'hbb27c5d2),
	.w6(32'h3b2e95e7),
	.w7(32'h3a240e41),
	.w8(32'hbb832fb9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea78e9),
	.w1(32'hbad06415),
	.w2(32'h3ba5b4eb),
	.w3(32'h3a790f6d),
	.w4(32'h3ad916b1),
	.w5(32'h3bec25cc),
	.w6(32'h3bad725e),
	.w7(32'h3bffdf25),
	.w8(32'h3c0c30ba),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2965bb),
	.w1(32'hbb8229cc),
	.w2(32'hb97dae1a),
	.w3(32'h3bbfe6cf),
	.w4(32'h3a88c4dc),
	.w5(32'hb9b5f2ac),
	.w6(32'h3b8ec84b),
	.w7(32'h3b4f4111),
	.w8(32'hb819465c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e189),
	.w1(32'hb8b4bd77),
	.w2(32'hbb59f53a),
	.w3(32'h3b1a951d),
	.w4(32'hbb501176),
	.w5(32'hbb240d59),
	.w6(32'hb920aca4),
	.w7(32'hbaae0139),
	.w8(32'h3a6ca3fd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7859d8),
	.w1(32'hbb53d112),
	.w2(32'hbbad3ecd),
	.w3(32'h3ac791e2),
	.w4(32'hb97d63d8),
	.w5(32'hbb9e57ee),
	.w6(32'h3c461662),
	.w7(32'h3b8f1694),
	.w8(32'hbaba9928),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5311),
	.w1(32'hbb628548),
	.w2(32'hba99c8e0),
	.w3(32'hbaa1aab4),
	.w4(32'h37be6b29),
	.w5(32'h3a9b39bc),
	.w6(32'hba3bbd4a),
	.w7(32'hb92c707b),
	.w8(32'h3aae4fd2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231fc9),
	.w1(32'h3b8073e7),
	.w2(32'h3b6193a2),
	.w3(32'h3bac9e7e),
	.w4(32'hbaa5f96b),
	.w5(32'h3b928d52),
	.w6(32'h3b0b37e1),
	.w7(32'h3bd72cc3),
	.w8(32'h3c185003),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd8ee0),
	.w1(32'h3c537ce6),
	.w2(32'h3b3fcd06),
	.w3(32'h3bd34c24),
	.w4(32'h3b34d02d),
	.w5(32'h3b80296f),
	.w6(32'h3c639a62),
	.w7(32'h3c47b533),
	.w8(32'h3afa4c8b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b490),
	.w1(32'h3b92db8d),
	.w2(32'h3aa56c47),
	.w3(32'h3a89ff30),
	.w4(32'h3b2ba365),
	.w5(32'h398b514c),
	.w6(32'hb94ce68f),
	.w7(32'hb9ebc943),
	.w8(32'hbab9f6d2),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b798ce4),
	.w1(32'h3a719210),
	.w2(32'h3b6187b8),
	.w3(32'h3b4932b3),
	.w4(32'h3a9d830b),
	.w5(32'hbab0074c),
	.w6(32'h3bfa9d19),
	.w7(32'h3c429115),
	.w8(32'h3b98acd4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb592b7),
	.w1(32'h3ac725b3),
	.w2(32'hbb1a2d6d),
	.w3(32'h3aa8eeda),
	.w4(32'h391bf1fc),
	.w5(32'hb9ae9cc5),
	.w6(32'h3b80fdce),
	.w7(32'h3a9a6b09),
	.w8(32'h3ac3387a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9262717),
	.w1(32'hbaf973bc),
	.w2(32'hbabc65e0),
	.w3(32'hb96dfcdc),
	.w4(32'hbb6877b1),
	.w5(32'hbc18850f),
	.w6(32'h3a6dc45c),
	.w7(32'hbac60e7f),
	.w8(32'hbbfac0b9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f9395),
	.w1(32'hbb8d643b),
	.w2(32'hbb168a32),
	.w3(32'hbbf99c54),
	.w4(32'hbb0c1cc0),
	.w5(32'hbb1d408f),
	.w6(32'hbb9ced1b),
	.w7(32'hbb44f4d8),
	.w8(32'hba9d9b7c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de0282),
	.w1(32'hbb4e838c),
	.w2(32'hbb90cbaa),
	.w3(32'h3904c85b),
	.w4(32'hbb81f9af),
	.w5(32'hbad38c62),
	.w6(32'h3b7a8b4e),
	.w7(32'hbb50768b),
	.w8(32'hba95d1a9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3562f6fe),
	.w1(32'h3bac01a5),
	.w2(32'h3b857bc4),
	.w3(32'h3ba72925),
	.w4(32'hbb83616a),
	.w5(32'hbba61ebf),
	.w6(32'h3c48f74c),
	.w7(32'h3b9a7433),
	.w8(32'h3afe0351),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d08f3),
	.w1(32'hbc3a74eb),
	.w2(32'hbc62944e),
	.w3(32'hbb16a313),
	.w4(32'hbbd30c11),
	.w5(32'hbc1cd5da),
	.w6(32'h397950a5),
	.w7(32'hbbcbebc2),
	.w8(32'h3a0ef195),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96d09b),
	.w1(32'h3aff02f9),
	.w2(32'h37a404a7),
	.w3(32'h3b076770),
	.w4(32'h3b793bb3),
	.w5(32'h3b68755e),
	.w6(32'h3b79390a),
	.w7(32'h3a7e1844),
	.w8(32'h3b8fc360),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedcbce),
	.w1(32'hbb5e1dc1),
	.w2(32'hba9a8d21),
	.w3(32'hbb8bd9df),
	.w4(32'hbb6bb575),
	.w5(32'hba76dea2),
	.w6(32'hbaed7c1f),
	.w7(32'hba2113f3),
	.w8(32'hbb16caea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6143bf),
	.w1(32'hbb4c7f77),
	.w2(32'hb9f63d2d),
	.w3(32'h3b22ba55),
	.w4(32'h388d876f),
	.w5(32'hbb44a388),
	.w6(32'h3b2d53a6),
	.w7(32'h3b0c713a),
	.w8(32'h3a3a9000),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25f9e8),
	.w1(32'hbaf159d2),
	.w2(32'hbb45dce5),
	.w3(32'h3bc1cb9c),
	.w4(32'h39b71b3d),
	.w5(32'h3ba0c49a),
	.w6(32'h3c34bb99),
	.w7(32'h3b5f8044),
	.w8(32'h3c2cf920),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5ddb8),
	.w1(32'hbbfe1aef),
	.w2(32'hbbd6efe7),
	.w3(32'h3b7436bc),
	.w4(32'hbb96dd77),
	.w5(32'hbbde6da6),
	.w6(32'h3ba01acd),
	.w7(32'hb99d1e52),
	.w8(32'hbba3f33d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9127c97),
	.w1(32'h3aba55d0),
	.w2(32'hba953869),
	.w3(32'h3a172c12),
	.w4(32'hbb0c70e9),
	.w5(32'hbb25e25e),
	.w6(32'hb8ab1107),
	.w7(32'hbb877927),
	.w8(32'hbc1b5c52),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c5509),
	.w1(32'hb9d9860a),
	.w2(32'hba1ba0cf),
	.w3(32'hbabcf6c7),
	.w4(32'h37ad1d83),
	.w5(32'hbb066bcf),
	.w6(32'hbb84ece0),
	.w7(32'hbaa9ffd1),
	.w8(32'hbb7187d3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaf837),
	.w1(32'h3a4d50f6),
	.w2(32'h3b38db0a),
	.w3(32'hbb87e3df),
	.w4(32'hbafe265f),
	.w5(32'h3b6b61d0),
	.w6(32'hbb4cfdca),
	.w7(32'h3aec6ed8),
	.w8(32'h3b95d524),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ca1b4),
	.w1(32'hb990e5c2),
	.w2(32'h3b37dbe7),
	.w3(32'h3aa89ba4),
	.w4(32'h3b143bd6),
	.w5(32'hbbacbacd),
	.w6(32'h3c0e3fa3),
	.w7(32'h3c22faa3),
	.w8(32'hbb2f4069),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57d1fe),
	.w1(32'hbc26059a),
	.w2(32'hbb89901d),
	.w3(32'h3acf412d),
	.w4(32'hbb8bccc6),
	.w5(32'hbaff6b95),
	.w6(32'h3ae938be),
	.w7(32'hba7783d6),
	.w8(32'h3b0f7a60),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aa7e2),
	.w1(32'hb967d5a8),
	.w2(32'h3af01b1d),
	.w3(32'h3bb7900a),
	.w4(32'h3bab8f11),
	.w5(32'hba9f5578),
	.w6(32'h3c448cca),
	.w7(32'h3c3df423),
	.w8(32'h3a826adf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb945d237),
	.w1(32'hbac8494c),
	.w2(32'h3b86eedf),
	.w3(32'hb91006fe),
	.w4(32'h3b6b9b51),
	.w5(32'h3b3aa119),
	.w6(32'hbb683e61),
	.w7(32'h38d80dd3),
	.w8(32'h3b6a7607),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc2ccd),
	.w1(32'h3b97463f),
	.w2(32'hbb4b9dbd),
	.w3(32'h3c2a04e3),
	.w4(32'hbb07f104),
	.w5(32'h3be4d777),
	.w6(32'h3bf6ad25),
	.w7(32'hbb4d0c8f),
	.w8(32'h3c19d688),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3364da),
	.w1(32'h3ad35dc5),
	.w2(32'h3ba13d12),
	.w3(32'h3b0c4ad1),
	.w4(32'h3c2ec687),
	.w5(32'h3a93a344),
	.w6(32'hbb3319bc),
	.w7(32'h3c13460a),
	.w8(32'hbb9357e9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996970b),
	.w1(32'hbac858e2),
	.w2(32'hbb462f50),
	.w3(32'hbb3a01d2),
	.w4(32'hb93cabc2),
	.w5(32'hba286e57),
	.w6(32'hbb68ed73),
	.w7(32'h3b355880),
	.w8(32'h3b0a6713),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a909ab2),
	.w1(32'h3b7e8fda),
	.w2(32'hba8ab72a),
	.w3(32'h3b85b563),
	.w4(32'h3b0e5b32),
	.w5(32'hba5bb78f),
	.w6(32'h3c0f48e8),
	.w7(32'h3b52e685),
	.w8(32'hb995fb2e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4d243),
	.w1(32'h3a0a960f),
	.w2(32'h39bac77f),
	.w3(32'h3a14bd83),
	.w4(32'hbb249411),
	.w5(32'hb825feee),
	.w6(32'hbaa428af),
	.w7(32'hbb5199a1),
	.w8(32'hb92e94b6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa63dc3),
	.w1(32'hbba06952),
	.w2(32'h3a0039bf),
	.w3(32'hbaac7318),
	.w4(32'h3abc966c),
	.w5(32'h3c08c05b),
	.w6(32'h3b6b1a05),
	.w7(32'h3b3dc7c1),
	.w8(32'h3b77b508),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c984d),
	.w1(32'hbc527526),
	.w2(32'h3b9ea6aa),
	.w3(32'h3bdedb3f),
	.w4(32'h3af18a43),
	.w5(32'hb90a8489),
	.w6(32'h3c2926ea),
	.w7(32'h3b9ce41a),
	.w8(32'h3bc1d860),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9685fa),
	.w1(32'hbc680d9f),
	.w2(32'hbc389da1),
	.w3(32'hb8dcbf13),
	.w4(32'h39f0fe4b),
	.w5(32'hbbebf978),
	.w6(32'h3bb72e62),
	.w7(32'h3b0c6442),
	.w8(32'hbbc84df9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a9485),
	.w1(32'h3ca81c7b),
	.w2(32'h3c73c6f4),
	.w3(32'h3a5412bf),
	.w4(32'hbbab241c),
	.w5(32'h3abaed1a),
	.w6(32'hbc64b720),
	.w7(32'hbbef30d7),
	.w8(32'h3b890b42),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eb0d8),
	.w1(32'h3bae9a74),
	.w2(32'h3a4d488a),
	.w3(32'hbacad4c8),
	.w4(32'h3b26d69b),
	.w5(32'h38a31a71),
	.w6(32'h3c4441a8),
	.w7(32'h3c396ae2),
	.w8(32'h3b2d401d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52462),
	.w1(32'h3b40dad3),
	.w2(32'h3b57dcbe),
	.w3(32'h3b65bc45),
	.w4(32'h3b9c4562),
	.w5(32'hbc038e19),
	.w6(32'h3b5164bb),
	.w7(32'h3bcdd2de),
	.w8(32'hbc4ed612),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29f4c1),
	.w1(32'h3b9fe590),
	.w2(32'hbb99ccc1),
	.w3(32'h3c00b1b3),
	.w4(32'hbbd11079),
	.w5(32'hba43e711),
	.w6(32'h3bbbabe4),
	.w7(32'hbb123f2a),
	.w8(32'h3ad54244),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7f7df),
	.w1(32'hbbbfcd34),
	.w2(32'h3c0237d1),
	.w3(32'h3b3d2b15),
	.w4(32'h3b02d2a9),
	.w5(32'hbc29f3ef),
	.w6(32'h3b03a278),
	.w7(32'h3bc7c04d),
	.w8(32'hbbaf01b5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7fb7),
	.w1(32'hba2de014),
	.w2(32'h3c078215),
	.w3(32'hbb603902),
	.w4(32'h3a5e2ac9),
	.w5(32'hba9819b8),
	.w6(32'h3bafb7ff),
	.w7(32'hbb40e7d3),
	.w8(32'h3ad80ff2),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd75abb),
	.w1(32'hbbc7aaab),
	.w2(32'hbbfbb53c),
	.w3(32'hbaf4bbd3),
	.w4(32'hbb8b3271),
	.w5(32'h3b08f95a),
	.w6(32'h3b356c55),
	.w7(32'hbb67ab3a),
	.w8(32'h3a90a933),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6bbdd),
	.w1(32'hbb8649ce),
	.w2(32'h39b4f117),
	.w3(32'hba8ccf4b),
	.w4(32'h3b1024a1),
	.w5(32'h39a9d4e0),
	.w6(32'h3abd0d2d),
	.w7(32'hb9b6f1e4),
	.w8(32'hbb8a5fdc),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa4bbe),
	.w1(32'hbbaa4b26),
	.w2(32'hbb439356),
	.w3(32'h3a3b3f37),
	.w4(32'hb9cf834d),
	.w5(32'h3bee0bae),
	.w6(32'hba654384),
	.w7(32'h3a9234b9),
	.w8(32'h3bc94198),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9777eb),
	.w1(32'hbb0722dc),
	.w2(32'h3bc387b4),
	.w3(32'h3b169b84),
	.w4(32'h3993780e),
	.w5(32'hbb992f1a),
	.w6(32'h3c720cac),
	.w7(32'h3b49d806),
	.w8(32'hbc1c373c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07b485),
	.w1(32'hbaf0325a),
	.w2(32'h39386059),
	.w3(32'hba7c8797),
	.w4(32'hbb85f295),
	.w5(32'hbb1fdb30),
	.w6(32'hba8a3ee2),
	.w7(32'h3c0ae81d),
	.w8(32'hbbc432b2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39804161),
	.w1(32'hbbae25c0),
	.w2(32'h3bbd3b81),
	.w3(32'h3b45e0d5),
	.w4(32'h3b8692d7),
	.w5(32'hbbf3ae73),
	.w6(32'h3c2decd7),
	.w7(32'h3c23bdeb),
	.w8(32'hbbdfedbf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcf743),
	.w1(32'h3b53825a),
	.w2(32'h3a69b281),
	.w3(32'hbad32327),
	.w4(32'hbc2daf9a),
	.w5(32'hbbc22285),
	.w6(32'hbbf8cd07),
	.w7(32'hbbc357d6),
	.w8(32'hbb968ec8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ebaa5),
	.w1(32'hbc6a5950),
	.w2(32'hbc86336b),
	.w3(32'h3bd89bbd),
	.w4(32'h3b9010ae),
	.w5(32'hbbd98d93),
	.w6(32'h3bfc2726),
	.w7(32'h3b18cccc),
	.w8(32'hbbc3001a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca56e1),
	.w1(32'h3c07a6e9),
	.w2(32'h3b9dab17),
	.w3(32'hbb88b89d),
	.w4(32'hbb5c80fc),
	.w5(32'h3abd2fcf),
	.w6(32'hbc37e01e),
	.w7(32'hbaf7cdeb),
	.w8(32'h3abac594),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0975),
	.w1(32'h39ebe140),
	.w2(32'hb9b419ae),
	.w3(32'hbb7354fc),
	.w4(32'hbb2a76de),
	.w5(32'hbb4b9b80),
	.w6(32'h3a51927e),
	.w7(32'hbb2f4a2b),
	.w8(32'hbb73f508),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34a932),
	.w1(32'h3c9e5b6e),
	.w2(32'h3c537838),
	.w3(32'h3bfe2cc4),
	.w4(32'h3b559b54),
	.w5(32'h3b605773),
	.w6(32'hbc851821),
	.w7(32'h3be2af1c),
	.w8(32'h3b22fc66),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cab60),
	.w1(32'hbc6d8c7a),
	.w2(32'hbc250938),
	.w3(32'hba285792),
	.w4(32'hbb8dfa5e),
	.w5(32'hbb74dc0d),
	.w6(32'h39f50b27),
	.w7(32'hbb3a2a14),
	.w8(32'h3b3e1f6a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63efe9),
	.w1(32'hbc3c601e),
	.w2(32'h3bde49eb),
	.w3(32'hbc1a04d3),
	.w4(32'hbb6496ab),
	.w5(32'h3b1531c5),
	.w6(32'hbbf5fed3),
	.w7(32'hba7c95d1),
	.w8(32'hbbc1aa82),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3757a),
	.w1(32'h3ce5210b),
	.w2(32'h3cf07de8),
	.w3(32'h3b0152b4),
	.w4(32'h3c1320b1),
	.w5(32'hbb391d84),
	.w6(32'hbc94f675),
	.w7(32'h3c68ddc4),
	.w8(32'hba5ce20b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbb09d),
	.w1(32'hbb00732a),
	.w2(32'h3a7082f1),
	.w3(32'h3af96616),
	.w4(32'h3b116e1a),
	.w5(32'h3a88bc0f),
	.w6(32'hbb258721),
	.w7(32'h3b454c4c),
	.w8(32'hbb2cb125),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6fef),
	.w1(32'h3c57593f),
	.w2(32'h3c26fbfe),
	.w3(32'hbb205c16),
	.w4(32'hbb4e2abd),
	.w5(32'hbb57ed2a),
	.w6(32'hbb85f79a),
	.w7(32'hbb978981),
	.w8(32'hbb26a207),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaa0ad),
	.w1(32'hba8a51b0),
	.w2(32'hbb8022f5),
	.w3(32'h3ad5b524),
	.w4(32'h3a0d88ce),
	.w5(32'hba76232a),
	.w6(32'hbb277274),
	.w7(32'h3b80d769),
	.w8(32'h3b778df5),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa72ed6),
	.w1(32'hba507671),
	.w2(32'h3b70c89f),
	.w3(32'h3b760f93),
	.w4(32'h3a6512f3),
	.w5(32'hbb8a4587),
	.w6(32'h3a6626a2),
	.w7(32'h3b947f42),
	.w8(32'hbab2b596),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb5324),
	.w1(32'h3bd241c5),
	.w2(32'h3ad9c8b4),
	.w3(32'h3abfb64b),
	.w4(32'hbbfa8a06),
	.w5(32'h3bbc6495),
	.w6(32'h3af29218),
	.w7(32'hba8538a7),
	.w8(32'h3b73b0bd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718231),
	.w1(32'hbb8b9e24),
	.w2(32'hbbd99457),
	.w3(32'h3b8ef89c),
	.w4(32'h3ac13aec),
	.w5(32'h3b98301c),
	.w6(32'h3b41e3ea),
	.w7(32'h3a29a8a0),
	.w8(32'h3a78a72f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d77e0),
	.w1(32'hbac85f44),
	.w2(32'hbbc5e597),
	.w3(32'h3a28a13f),
	.w4(32'hbbb357c0),
	.w5(32'h3b0089f5),
	.w6(32'h3a7941e1),
	.w7(32'hbada63a2),
	.w8(32'h39340a6c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule