module layer_6_featuremap_99(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a3035c),
	.w1(32'hbbc53ad2),
	.w2(32'hbba605fa),
	.w3(32'hba92d035),
	.w4(32'hbb380b55),
	.w5(32'h39be39c9),
	.w6(32'hbb259600),
	.w7(32'hbb21778f),
	.w8(32'hbb68eb30),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb412110),
	.w1(32'h3abb3b81),
	.w2(32'h3b1378eb),
	.w3(32'hbaaf25df),
	.w4(32'hbb6beaf8),
	.w5(32'hbbc67d3c),
	.w6(32'h3a4ec3a4),
	.w7(32'h3b84718e),
	.w8(32'hba7f3cf3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad868e0),
	.w1(32'hbbfa3557),
	.w2(32'h3c0e8d99),
	.w3(32'h3bda9143),
	.w4(32'hbc1005e7),
	.w5(32'h3a29e7e4),
	.w6(32'hbb782efa),
	.w7(32'hbb20956a),
	.w8(32'hbbd16fe3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6267ce),
	.w1(32'hb984e80f),
	.w2(32'h3b7e2054),
	.w3(32'hb9e9ccb3),
	.w4(32'h3b437f12),
	.w5(32'h3b1d5616),
	.w6(32'hb972c9a8),
	.w7(32'h3a04805b),
	.w8(32'h3b8b431a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42e84a),
	.w1(32'hbc995295),
	.w2(32'h3c0745b8),
	.w3(32'h3cc35bff),
	.w4(32'hbbb1973f),
	.w5(32'hbc17cc5b),
	.w6(32'hbadb3b37),
	.w7(32'h3d3a2823),
	.w8(32'hbd038cc9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d589449),
	.w1(32'hbbddfa0b),
	.w2(32'hbbb4f017),
	.w3(32'hbabfa198),
	.w4(32'hb9b9b9dd),
	.w5(32'h3baa80ac),
	.w6(32'hbb84422c),
	.w7(32'hbba3a884),
	.w8(32'hbb8b95b8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ec5f),
	.w1(32'h3bbd5b46),
	.w2(32'h3b20ccdb),
	.w3(32'hbbf288ce),
	.w4(32'hbb20c9a0),
	.w5(32'hbbcc4689),
	.w6(32'h3a91750a),
	.w7(32'hba6b17d3),
	.w8(32'h3ab05262),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93311),
	.w1(32'hbcd951dd),
	.w2(32'h3d0ccbcf),
	.w3(32'h3bdf9fb8),
	.w4(32'hbc4e27c7),
	.w5(32'h3c144e86),
	.w6(32'h3cb2bcc5),
	.w7(32'h3a6af3e4),
	.w8(32'hbd08877e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ef322),
	.w1(32'h3b01c48a),
	.w2(32'hbd89b657),
	.w3(32'hbc26b524),
	.w4(32'h3cc59c29),
	.w5(32'hbcbb9695),
	.w6(32'hbd4b5775),
	.w7(32'h3d1b88be),
	.w8(32'h3c734db0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d93ecf8),
	.w1(32'hbbadc400),
	.w2(32'hbb8abb3d),
	.w3(32'hba90ca43),
	.w4(32'h3ababcca),
	.w5(32'h3ad0995f),
	.w6(32'hbb791fdf),
	.w7(32'hba2154ea),
	.w8(32'hba2ef16e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fcc45),
	.w1(32'hbba728a8),
	.w2(32'hbc26f7ba),
	.w3(32'h3bd4b66d),
	.w4(32'h3c3bd5c0),
	.w5(32'hbc079054),
	.w6(32'h397a6e4a),
	.w7(32'hbc172181),
	.w8(32'h3c1482a9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9914a),
	.w1(32'h3a77d923),
	.w2(32'hbb6fbdd9),
	.w3(32'h3929eb0a),
	.w4(32'h3aedcc96),
	.w5(32'h3b624384),
	.w6(32'hbb21c0dc),
	.w7(32'h3b4fcd1a),
	.w8(32'h3a957b01),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ed374),
	.w1(32'hbb028686),
	.w2(32'h3b8d37c7),
	.w3(32'hbbf9abf0),
	.w4(32'h3c0177f1),
	.w5(32'hbb83e053),
	.w6(32'hbb264549),
	.w7(32'h3bd73638),
	.w8(32'hbac32886),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049e01),
	.w1(32'hbb8f1c0d),
	.w2(32'h3adb74de),
	.w3(32'hbb8fe93b),
	.w4(32'hbc9e55df),
	.w5(32'h3c72cebf),
	.w6(32'h3b8c6f11),
	.w7(32'hbca13c2c),
	.w8(32'hbbbd5b51),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccceab),
	.w1(32'h3b69ec83),
	.w2(32'h3be1dde9),
	.w3(32'h3b864d4c),
	.w4(32'h3c3bc9b5),
	.w5(32'h3bff712e),
	.w6(32'h3b9560b7),
	.w7(32'h3b8cfadf),
	.w8(32'h3c345f56),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfd8c1),
	.w1(32'hbb51dd2d),
	.w2(32'hba51899e),
	.w3(32'h3a9be132),
	.w4(32'h3b5ac22e),
	.w5(32'h3b16c6cd),
	.w6(32'hba82b86d),
	.w7(32'hbb75ec3f),
	.w8(32'h3a957e99),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2338b),
	.w1(32'h3b7300e3),
	.w2(32'hbc03a6bb),
	.w3(32'h3c2e3931),
	.w4(32'hbc156388),
	.w5(32'h3c1445fd),
	.w6(32'hbb1ec698),
	.w7(32'hbbcc6c7c),
	.w8(32'h3b8b6876),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5d14e),
	.w1(32'h3b11654e),
	.w2(32'h3b4d1551),
	.w3(32'h3a767732),
	.w4(32'h3b8fc733),
	.w5(32'hb9b1a84c),
	.w6(32'hb9dd6236),
	.w7(32'hbb26605a),
	.w8(32'h3ab04519),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499efb),
	.w1(32'hbb7b0287),
	.w2(32'hbb32b482),
	.w3(32'h39fe82c0),
	.w4(32'h3b1f64b0),
	.w5(32'h3baac59a),
	.w6(32'hbad727be),
	.w7(32'hba9a251f),
	.w8(32'h396834ba),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24908c),
	.w1(32'h3cad7ae8),
	.w2(32'hbcbfd687),
	.w3(32'h3bde1307),
	.w4(32'h3aeb8680),
	.w5(32'h3b5d7b88),
	.w6(32'hbc98dccf),
	.w7(32'h3ca8fd16),
	.w8(32'h3bcdffd2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c993eff),
	.w1(32'hba878293),
	.w2(32'h3ad3d3f2),
	.w3(32'h3ad662a9),
	.w4(32'hbb33f3f8),
	.w5(32'hbb477d12),
	.w6(32'hba442d78),
	.w7(32'hbb193431),
	.w8(32'hba1facc5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb311dee),
	.w1(32'hbbb08c98),
	.w2(32'hbb569c0d),
	.w3(32'h3ac0373f),
	.w4(32'h3b9772b0),
	.w5(32'hb9fbf56d),
	.w6(32'hba72a2f6),
	.w7(32'h39bd090d),
	.w8(32'h3b91bd75),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e60b74),
	.w1(32'hbc5cc9e4),
	.w2(32'h3cb4c7b6),
	.w3(32'hbc549fb8),
	.w4(32'h398d9331),
	.w5(32'h3c943a30),
	.w6(32'h3c4e9069),
	.w7(32'h3b7438cf),
	.w8(32'hbca50aa2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba576b9),
	.w1(32'h3c4cab1a),
	.w2(32'hbd000f95),
	.w3(32'hbcfb2390),
	.w4(32'h3c8cd3f5),
	.w5(32'hba9b4cd8),
	.w6(32'hbc9524a3),
	.w7(32'hbcd7d5e5),
	.w8(32'h3d16744e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8548d0),
	.w1(32'hbc192c84),
	.w2(32'hbc2b2b78),
	.w3(32'h39a90405),
	.w4(32'hbc1bf26f),
	.w5(32'hbbffae8e),
	.w6(32'hbc0a44e2),
	.w7(32'hbc885321),
	.w8(32'hbbbbb18e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e6055),
	.w1(32'hbbfa5e7e),
	.w2(32'hbc28c69e),
	.w3(32'hbc0e797f),
	.w4(32'hbbfcabd4),
	.w5(32'h3b2ef912),
	.w6(32'hbc5c9ae4),
	.w7(32'hbbfa661d),
	.w8(32'hbbb0911e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe10ead),
	.w1(32'hbb29b87a),
	.w2(32'h3bb5a709),
	.w3(32'h3be1b3a4),
	.w4(32'h3ad55da2),
	.w5(32'h3bd9bb06),
	.w6(32'h3c2e7fb5),
	.w7(32'hbb8787cf),
	.w8(32'h3846d4ca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09d589),
	.w1(32'h3adc9eb3),
	.w2(32'h3ab3e232),
	.w3(32'hba77d874),
	.w4(32'h3b51504d),
	.w5(32'h3a77c5a1),
	.w6(32'hba1d6dcb),
	.w7(32'h3b01f7bf),
	.w8(32'h3b1091cb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a8069),
	.w1(32'hbae67250),
	.w2(32'hba96e866),
	.w3(32'h3b17f1cd),
	.w4(32'h3a5e20a7),
	.w5(32'hbb386f4c),
	.w6(32'h3a1a9df7),
	.w7(32'h3a2582ce),
	.w8(32'hba240f81),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59265e),
	.w1(32'h3ca94f27),
	.w2(32'h3ce9c4a4),
	.w3(32'hbbed2c14),
	.w4(32'h3cb8e93b),
	.w5(32'hbc139961),
	.w6(32'h3c78ccc5),
	.w7(32'h3ce4d5bd),
	.w8(32'h3c99f224),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d07f6cb),
	.w1(32'hbc6b4b3a),
	.w2(32'h3c984b7a),
	.w3(32'h3c45ef6c),
	.w4(32'hbc8ca514),
	.w5(32'hbbbf0e4c),
	.w6(32'h3c4c6751),
	.w7(32'h3cd8c49c),
	.w8(32'hbcafca38),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e2098),
	.w1(32'hbbb2da5f),
	.w2(32'h3b59ea29),
	.w3(32'h3b83ae31),
	.w4(32'h3a547d59),
	.w5(32'hbb11060b),
	.w6(32'hbc834e4c),
	.w7(32'h3c17741b),
	.w8(32'hbadbdda5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2dccd),
	.w1(32'h3c3e54ee),
	.w2(32'hbc663eef),
	.w3(32'hbc50c063),
	.w4(32'h3c6da577),
	.w5(32'h3b232c77),
	.w6(32'hbba31efc),
	.w7(32'hbd15c5c1),
	.w8(32'h3ca73213),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd2793),
	.w1(32'h3b1058a0),
	.w2(32'h3d097f39),
	.w3(32'h3b94e08c),
	.w4(32'hbba1b506),
	.w5(32'h3c96b27f),
	.w6(32'h3c453623),
	.w7(32'h3d2214b8),
	.w8(32'h3c72bcaf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f5772),
	.w1(32'hbb80e822),
	.w2(32'hbaef248a),
	.w3(32'hba6ee1ae),
	.w4(32'hbaccfad4),
	.w5(32'hb8721e73),
	.w6(32'hbb10d601),
	.w7(32'hba470648),
	.w8(32'hbb6f0057),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24fba),
	.w1(32'hbb0989e0),
	.w2(32'h3c1883c9),
	.w3(32'hbb6d04a2),
	.w4(32'hbbe10057),
	.w5(32'hbb694533),
	.w6(32'h3b4fb0b8),
	.w7(32'h37e4b7a1),
	.w8(32'hbbc7a2ab),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825963),
	.w1(32'hba08a945),
	.w2(32'hbb848efc),
	.w3(32'h3ac2e879),
	.w4(32'hbaa2701a),
	.w5(32'h3c288951),
	.w6(32'hbac04a06),
	.w7(32'hbb3d2df9),
	.w8(32'hbbd19185),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394806a2),
	.w1(32'hbaac8e39),
	.w2(32'h3a948dfe),
	.w3(32'h3a68166c),
	.w4(32'hb9be857d),
	.w5(32'hba1295eb),
	.w6(32'hbaab7297),
	.w7(32'h3a8cfcf6),
	.w8(32'hbb10e415),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b363260),
	.w1(32'hbb739287),
	.w2(32'hbc5f0b13),
	.w3(32'h3ba42265),
	.w4(32'h3c4c56fa),
	.w5(32'h3baa3990),
	.w6(32'hbc00739f),
	.w7(32'h39572e9c),
	.w8(32'hbbc50de1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50ec8a),
	.w1(32'h3c77a241),
	.w2(32'hbda7d461),
	.w3(32'h3933145c),
	.w4(32'h3d3d3dec),
	.w5(32'hbd13845f),
	.w6(32'hbd5a2478),
	.w7(32'h3d302130),
	.w8(32'h3c976b36),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d546bb7),
	.w1(32'hbcabcc8a),
	.w2(32'h3ca5ad12),
	.w3(32'h3cfbacb9),
	.w4(32'hbc0e6fd4),
	.w5(32'hbc20ce7e),
	.w6(32'h3c44823c),
	.w7(32'h3d0c4e0c),
	.w8(32'hbce974f9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d12cfbc),
	.w1(32'hbace5f07),
	.w2(32'h3b47da97),
	.w3(32'hbab18ee7),
	.w4(32'h3b33cfd3),
	.w5(32'h3a28e10c),
	.w6(32'hba32ea6d),
	.w7(32'h38db8aed),
	.w8(32'h3b3609d8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46a2b2),
	.w1(32'hbb303f94),
	.w2(32'hbb03969c),
	.w3(32'h3c018633),
	.w4(32'h3b837a2e),
	.w5(32'h3c1ec8cb),
	.w6(32'hba5cf4b3),
	.w7(32'h3bdaa2c0),
	.w8(32'hbb42bb9a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d268d),
	.w1(32'hbbadeeda),
	.w2(32'hba499342),
	.w3(32'hbb725675),
	.w4(32'hbab1af74),
	.w5(32'h3b1db720),
	.w6(32'hbba32d52),
	.w7(32'hba8319ad),
	.w8(32'hbae0020f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd7a0e),
	.w1(32'hbb913ce9),
	.w2(32'hbb05ef94),
	.w3(32'hbb154646),
	.w4(32'h3a84f78f),
	.w5(32'h3a19ba66),
	.w6(32'hbb52631d),
	.w7(32'hbb1a8330),
	.w8(32'hba7e247d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f56f0),
	.w1(32'hbcc6a3b1),
	.w2(32'h3c5b6a6c),
	.w3(32'h3c325948),
	.w4(32'hbb44ecb2),
	.w5(32'hbc67412e),
	.w6(32'h3b9d11d1),
	.w7(32'hbbeb5268),
	.w8(32'hbb7a4343),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc912a17),
	.w1(32'h3b9869a1),
	.w2(32'h3c4fd5d7),
	.w3(32'hbb98d16a),
	.w4(32'hbad01433),
	.w5(32'hbbbee309),
	.w6(32'hbba83db2),
	.w7(32'h39b98526),
	.w8(32'h3c6efa59),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde8e25),
	.w1(32'hbb7674ad),
	.w2(32'hbc877b1e),
	.w3(32'hbbc54c09),
	.w4(32'hbba51a0f),
	.w5(32'hbb3c0b04),
	.w6(32'hbc861c01),
	.w7(32'hbcde232a),
	.w8(32'h3c52bd83),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd08cc0),
	.w1(32'hb9c84a60),
	.w2(32'hbb1698fe),
	.w3(32'hbad22b1e),
	.w4(32'h3aeb11b1),
	.w5(32'h3bd32367),
	.w6(32'hbb41d559),
	.w7(32'hbad2a0d8),
	.w8(32'h3adcbb06),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3972b7),
	.w1(32'h3aa45d9c),
	.w2(32'h3d811708),
	.w3(32'hbb8ddc1c),
	.w4(32'hbd1180ad),
	.w5(32'h3cc77771),
	.w6(32'h3d1b3c8b),
	.w7(32'hbd3cda26),
	.w8(32'hbc309572),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdac742e),
	.w1(32'hbaf49617),
	.w2(32'h3be39bfb),
	.w3(32'hbb97f0a5),
	.w4(32'h3a2338bd),
	.w5(32'hbb39bf0a),
	.w6(32'hbb2415b5),
	.w7(32'hbaabdaf5),
	.w8(32'hbb16d628),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc173f3a),
	.w1(32'h3ba97606),
	.w2(32'h39393fc9),
	.w3(32'hbb8f540c),
	.w4(32'hbad55e8f),
	.w5(32'h39666e82),
	.w6(32'h39bcd7b4),
	.w7(32'hbb7b6637),
	.w8(32'h3af539dc),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6e968),
	.w1(32'h39320ba8),
	.w2(32'hb9e79ea7),
	.w3(32'hbaa8d9b8),
	.w4(32'hb99ecf73),
	.w5(32'h3b58a8c6),
	.w6(32'hba1a404f),
	.w7(32'hbb985836),
	.w8(32'h3b96993f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa51236),
	.w1(32'hba0ac49b),
	.w2(32'h3b97fcfa),
	.w3(32'hbabc7205),
	.w4(32'h3ad2cdf8),
	.w5(32'hbb5ef6d9),
	.w6(32'h3ac47e96),
	.w7(32'hbab81412),
	.w8(32'h3ba01af9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b628188),
	.w1(32'hb94ff1d6),
	.w2(32'h399c2c51),
	.w3(32'hbac09951),
	.w4(32'h3ab50e86),
	.w5(32'hb99442d2),
	.w6(32'hbb9ee9f5),
	.w7(32'hbbac02eb),
	.w8(32'h3b7771f0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc2f0d),
	.w1(32'h3ae25a5c),
	.w2(32'h3c025307),
	.w3(32'hbc070306),
	.w4(32'h3bc078ac),
	.w5(32'h3c443831),
	.w6(32'h3c6edbef),
	.w7(32'h3d06aa1a),
	.w8(32'h3cbcba4b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379fbdd1),
	.w1(32'h3a2a8057),
	.w2(32'h3bb562a1),
	.w3(32'h3a8f30c9),
	.w4(32'hbc0017a1),
	.w5(32'hbbc8f68d),
	.w6(32'hbb8a7cdd),
	.w7(32'hbbe36d47),
	.w8(32'h3ae7edda),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e31e8),
	.w1(32'h3b60db93),
	.w2(32'h3bbc86b4),
	.w3(32'h39fb9bb6),
	.w4(32'h3ba3a25f),
	.w5(32'h3b90297f),
	.w6(32'hbb729c48),
	.w7(32'h3c241fbc),
	.w8(32'hbb2da8c2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf81a9),
	.w1(32'hba9f93ed),
	.w2(32'hbb1605e0),
	.w3(32'hbb019d84),
	.w4(32'hbb4f40ad),
	.w5(32'hbb94cfc6),
	.w6(32'hba696539),
	.w7(32'hba3b5618),
	.w8(32'hbb7d28a2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf405e8),
	.w1(32'hbcba0bcb),
	.w2(32'hbd02f0bd),
	.w3(32'hbb05c2b4),
	.w4(32'hbbdb516d),
	.w5(32'hbd1028f3),
	.w6(32'hbc9193ca),
	.w7(32'hbd65efca),
	.w8(32'hbd76a9e7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3da4a),
	.w1(32'hbb4e6ad3),
	.w2(32'hbc0f8168),
	.w3(32'hbb13c05c),
	.w4(32'hbb4b5cb4),
	.w5(32'hbb5c6ae5),
	.w6(32'h3a89d759),
	.w7(32'hba177589),
	.w8(32'hbc36ffb8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc817b49),
	.w1(32'hbcbb6711),
	.w2(32'hbcfa650d),
	.w3(32'hbc941acb),
	.w4(32'hbcb8363f),
	.w5(32'hbc40642c),
	.w6(32'hbc8340fd),
	.w7(32'hbc8b35c3),
	.w8(32'hbcc27a9a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61d7cf),
	.w1(32'hbc8bdfdb),
	.w2(32'hbb8f82cf),
	.w3(32'hbd1522e4),
	.w4(32'hbd37fc6f),
	.w5(32'hbc8b9231),
	.w6(32'hbd061f0d),
	.w7(32'hbc3d7a8a),
	.w8(32'h3c6e6df7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca92a2c),
	.w1(32'h3b6403f4),
	.w2(32'hbc117093),
	.w3(32'hbc074093),
	.w4(32'h3bb2decf),
	.w5(32'h3c0a6afd),
	.w6(32'h3c1e28e0),
	.w7(32'h3c4e0fcf),
	.w8(32'hbac283d7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule