module layer_8_featuremap_243(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfedf5d),
	.w1(32'hbb445b40),
	.w2(32'h3b8be796),
	.w3(32'hbbaa232b),
	.w4(32'h36f5c57c),
	.w5(32'hbb3818d1),
	.w6(32'h3b045833),
	.w7(32'h39d1143f),
	.w8(32'hbb7eaf14),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0e68a),
	.w1(32'hb9dbc5a6),
	.w2(32'hbb0c49a1),
	.w3(32'hbba6b25f),
	.w4(32'hbb3beebb),
	.w5(32'hbb68bc10),
	.w6(32'h38945466),
	.w7(32'hb9282655),
	.w8(32'h3ad9fd30),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad208f1),
	.w1(32'hbb65a28c),
	.w2(32'h3adadbfe),
	.w3(32'hbacdf458),
	.w4(32'h3a8d957c),
	.w5(32'h3ad5e913),
	.w6(32'h3a873cbb),
	.w7(32'h3b2d65a1),
	.w8(32'h3bd0ffca),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b343),
	.w1(32'hbab77b22),
	.w2(32'h3b37396a),
	.w3(32'h3ba6f2d9),
	.w4(32'h39eb7f2b),
	.w5(32'h3b7afb3d),
	.w6(32'hbbb1589b),
	.w7(32'h3af4f4a8),
	.w8(32'hbac48c90),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49005e),
	.w1(32'hbbd12e36),
	.w2(32'hbbf15abc),
	.w3(32'hb93eabeb),
	.w4(32'hbbd39d82),
	.w5(32'hbbfeed40),
	.w6(32'hbbba2610),
	.w7(32'hbbdc1175),
	.w8(32'hbb92e744),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47fc3),
	.w1(32'hba806174),
	.w2(32'h3be1c599),
	.w3(32'hbbb2654d),
	.w4(32'hbc04329e),
	.w5(32'hbb55f8a1),
	.w6(32'hbb56351f),
	.w7(32'h3c0344f1),
	.w8(32'h3b99436b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb63811),
	.w1(32'h3a5312d1),
	.w2(32'h3af0aa98),
	.w3(32'hbbe8f7e8),
	.w4(32'h3b17feaf),
	.w5(32'h3b88a0c7),
	.w6(32'h3af258af),
	.w7(32'hb86fb8af),
	.w8(32'hbb0ff129),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60c1f9),
	.w1(32'hbaf94573),
	.w2(32'hbbd359b4),
	.w3(32'h3b06a071),
	.w4(32'hb984d7e1),
	.w5(32'h3aa13445),
	.w6(32'hbb1f5837),
	.w7(32'hbc0471c9),
	.w8(32'hbc0283b4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0c943),
	.w1(32'hb9067f7d),
	.w2(32'hbb34b382),
	.w3(32'h3bb4da66),
	.w4(32'hbb39f176),
	.w5(32'hbbaf1f0b),
	.w6(32'h3b45a6e9),
	.w7(32'h39c4b2e8),
	.w8(32'hba761e6f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f6478),
	.w1(32'h3b9575d9),
	.w2(32'hbbc48c0c),
	.w3(32'hbb64b894),
	.w4(32'hbbca32c1),
	.w5(32'hbbb49493),
	.w6(32'h3acd6c68),
	.w7(32'h3819229e),
	.w8(32'hbc292fd3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04d8b1),
	.w1(32'hbba7e01b),
	.w2(32'hbc4ad2ac),
	.w3(32'hbc1c97f6),
	.w4(32'h3ab01df8),
	.w5(32'hbbc0d9a5),
	.w6(32'hbb6f49e2),
	.w7(32'hbb377006),
	.w8(32'h3c01d2ca),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989d126),
	.w1(32'h3be7a1de),
	.w2(32'h3c0aab73),
	.w3(32'h39ddb92e),
	.w4(32'h3c016fe8),
	.w5(32'h3c0270d5),
	.w6(32'h3bf60dd3),
	.w7(32'h3c0912a6),
	.w8(32'h3abde1dc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4267f3),
	.w1(32'hbb9e6d38),
	.w2(32'hbbcb22ad),
	.w3(32'hbb99ac5f),
	.w4(32'hbba8b4c0),
	.w5(32'hbbb42157),
	.w6(32'hbba612a1),
	.w7(32'hbb84fcf6),
	.w8(32'h3a51321b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3bf1e),
	.w1(32'h3ac7bdf4),
	.w2(32'hbb03b90d),
	.w3(32'hb9bc9677),
	.w4(32'h3b0db221),
	.w5(32'h3a79c934),
	.w6(32'hbb8c96b2),
	.w7(32'h3b94e174),
	.w8(32'hbab0048c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e571),
	.w1(32'hbbcbc96e),
	.w2(32'hbc048015),
	.w3(32'h3b9e792f),
	.w4(32'hbb9eea6b),
	.w5(32'hbbe9ebd5),
	.w6(32'hbb8426b0),
	.w7(32'hbbe22307),
	.w8(32'hbbf419de),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf3b77),
	.w1(32'h3bf63d91),
	.w2(32'h3addad74),
	.w3(32'hbbe43ec6),
	.w4(32'h3b56ad1d),
	.w5(32'hbb9c6243),
	.w6(32'h3be5502f),
	.w7(32'hbb880239),
	.w8(32'hbba3f167),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb489a8),
	.w1(32'hbae89dbe),
	.w2(32'h39d0ca7e),
	.w3(32'hbb826d95),
	.w4(32'hbbb4b21c),
	.w5(32'hbadad1fb),
	.w6(32'hbb3ec9ef),
	.w7(32'hbb333dec),
	.w8(32'hbbb9b10a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8163c),
	.w1(32'h3af14d7c),
	.w2(32'h3b42274f),
	.w3(32'hbb296c58),
	.w4(32'h3af71ed0),
	.w5(32'h3ba30575),
	.w6(32'hbab3cd74),
	.w7(32'h3bdbc863),
	.w8(32'h3beb6f6a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bce4a),
	.w1(32'hbb308255),
	.w2(32'h3a9b37f3),
	.w3(32'h3b4ab202),
	.w4(32'hba03dd91),
	.w5(32'hbb5278c1),
	.w6(32'hbb8f9c78),
	.w7(32'hbbf9340d),
	.w8(32'hbbe851af),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea5bde),
	.w1(32'hbb66e14e),
	.w2(32'hbbb0696d),
	.w3(32'hbb94e2d5),
	.w4(32'hbb958fd2),
	.w5(32'hbb518453),
	.w6(32'hbbf50e50),
	.w7(32'hbc0791d3),
	.w8(32'hbc1c077e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb324d7),
	.w1(32'hbbb3ea32),
	.w2(32'hbc141af2),
	.w3(32'hbbbf1a97),
	.w4(32'hb9962531),
	.w5(32'hbb2dadd0),
	.w6(32'hba9971a7),
	.w7(32'hbb53a4f3),
	.w8(32'h3c21ae4f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7f36),
	.w1(32'h3b639b79),
	.w2(32'h3c25391f),
	.w3(32'h3b8639cd),
	.w4(32'h3b4ec611),
	.w5(32'h3a6be2a3),
	.w6(32'hbb9b69f8),
	.w7(32'h3b73be04),
	.w8(32'h3b1482fc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35ccd0),
	.w1(32'hbb9cc98d),
	.w2(32'hbbee43ab),
	.w3(32'h3b93e72c),
	.w4(32'h3b5a90be),
	.w5(32'hbba7b1fe),
	.w6(32'hbb62b599),
	.w7(32'hbb9b39ec),
	.w8(32'hb768891c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8f27),
	.w1(32'h3b983ef4),
	.w2(32'h3b7f60b4),
	.w3(32'h3bd9bdb0),
	.w4(32'h3b910c5f),
	.w5(32'h3ba7d1c7),
	.w6(32'h3bcdadec),
	.w7(32'h3b5412c2),
	.w8(32'hbafae8ca),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ad3af),
	.w1(32'hbb070c5c),
	.w2(32'h39a6ed15),
	.w3(32'h3b9b02d0),
	.w4(32'hbc2920da),
	.w5(32'hbbd425a2),
	.w6(32'hba821e27),
	.w7(32'h3aafdf36),
	.w8(32'h38851cad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43819a),
	.w1(32'hbb028f26),
	.w2(32'hba1078f4),
	.w3(32'hbb5d0b82),
	.w4(32'h3c5785fd),
	.w5(32'h3ba26660),
	.w6(32'hbb745bd1),
	.w7(32'hbbbd24fe),
	.w8(32'h3b107ae7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a980a91),
	.w1(32'h3b0086ea),
	.w2(32'h3a54b3dc),
	.w3(32'h3b5128a5),
	.w4(32'hbb5b6032),
	.w5(32'h3aa3a398),
	.w6(32'h3a2cb3ed),
	.w7(32'h39d5c209),
	.w8(32'hbbbdd492),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaedcc6),
	.w1(32'hbc2a0697),
	.w2(32'hbbfcfbd5),
	.w3(32'hbaf1f520),
	.w4(32'hba0bbd1c),
	.w5(32'hbc0a4dd9),
	.w6(32'hbb924df2),
	.w7(32'hbade1396),
	.w8(32'h3b9bc680),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8ac5),
	.w1(32'hba764704),
	.w2(32'h3adc0b86),
	.w3(32'h3aa9cbf6),
	.w4(32'hba026222),
	.w5(32'h3b091e92),
	.w6(32'h3b0fcd62),
	.w7(32'h3b885ac1),
	.w8(32'h3ba49b85),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02bf1b),
	.w1(32'hb889a5eb),
	.w2(32'h3a3356f9),
	.w3(32'h3b826cfd),
	.w4(32'hbb2c3639),
	.w5(32'hbb87e71d),
	.w6(32'h39e30d2a),
	.w7(32'h3a45788a),
	.w8(32'hbbfa2e5e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc064c23),
	.w1(32'h3b43c75c),
	.w2(32'h3a95a60b),
	.w3(32'hbc4a6ec8),
	.w4(32'h3c06640d),
	.w5(32'h3bc60fa8),
	.w6(32'hbb70af6f),
	.w7(32'hba7e6a4d),
	.w8(32'hbb838dfc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba468980),
	.w1(32'h3bb68501),
	.w2(32'h3abd8c95),
	.w3(32'h3bf3ce02),
	.w4(32'h3c3dbb6a),
	.w5(32'h3b9ebc88),
	.w6(32'h3bb8d419),
	.w7(32'h3a729818),
	.w8(32'h3bb4d319),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61d353),
	.w1(32'h3b67cc36),
	.w2(32'h3b31b5b6),
	.w3(32'h3bcf65d6),
	.w4(32'h3989e878),
	.w5(32'hbb4e6212),
	.w6(32'h3b458e86),
	.w7(32'h3a2e6c7a),
	.w8(32'hbb3502bd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a4a7e),
	.w1(32'h3a8d44cf),
	.w2(32'h397412e9),
	.w3(32'hbbcf339e),
	.w4(32'hbb1a9b84),
	.w5(32'h3ae7266e),
	.w6(32'h3b5eb8a5),
	.w7(32'hba12c761),
	.w8(32'h39a937ff),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890aedb),
	.w1(32'hbabe0636),
	.w2(32'h3b9c9c71),
	.w3(32'h3ad1e4c3),
	.w4(32'hbb6136c5),
	.w5(32'hba71b8b2),
	.w6(32'hbc1c93a8),
	.w7(32'hbadb7f3d),
	.w8(32'hbbb8c393),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecebd2),
	.w1(32'hbb683c3e),
	.w2(32'hb9e806fd),
	.w3(32'hbc13b946),
	.w4(32'h3a8dfcfb),
	.w5(32'h3b904ae3),
	.w6(32'hba47cfe4),
	.w7(32'h3b8035fd),
	.w8(32'h3abb87a6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ea13c),
	.w1(32'h3b27f275),
	.w2(32'hbaad8c2b),
	.w3(32'h3a44e8e9),
	.w4(32'h3c06f30c),
	.w5(32'h3b40ea84),
	.w6(32'hbaa7dfb8),
	.w7(32'hbb6e1127),
	.w8(32'hbbbe16f2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63c680),
	.w1(32'h39d9d696),
	.w2(32'hbba31fbd),
	.w3(32'hbb10cc3e),
	.w4(32'hba0d2917),
	.w5(32'hbbb2163f),
	.w6(32'h3baa4bcf),
	.w7(32'hbaa25aa2),
	.w8(32'h3ab541c7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d6f3b),
	.w1(32'h3a4f04dd),
	.w2(32'h37e16603),
	.w3(32'hbabf6835),
	.w4(32'hb95a8fc4),
	.w5(32'h3b18bd94),
	.w6(32'h3b23fe41),
	.w7(32'h3b992e02),
	.w8(32'hb9e62e41),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade2cb5),
	.w1(32'h3b5c82ae),
	.w2(32'h3b08bfe8),
	.w3(32'hb98d4506),
	.w4(32'h3b969b46),
	.w5(32'h3bc75ace),
	.w6(32'hb94ddf95),
	.w7(32'hba7628b0),
	.w8(32'h3b30e3c2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c3107),
	.w1(32'h3caab09e),
	.w2(32'h3ca9ee38),
	.w3(32'h3ba66ed9),
	.w4(32'h3ccb229e),
	.w5(32'h3cb4143a),
	.w6(32'h3ca6dc5b),
	.w7(32'h3ca90751),
	.w8(32'h3cd941ab),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd0541),
	.w1(32'h3b33869b),
	.w2(32'hbaa15c1e),
	.w3(32'h3ccd9a49),
	.w4(32'h3b558b97),
	.w5(32'h39a5a5fb),
	.w6(32'h3b83b2d9),
	.w7(32'hbb8f6dc9),
	.w8(32'hbc6eeb47),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f41d6),
	.w1(32'hbae6c388),
	.w2(32'hbb32e369),
	.w3(32'hbc2334e6),
	.w4(32'hbc027f11),
	.w5(32'hbbf93bcf),
	.w6(32'hbb889212),
	.w7(32'hbb1c9456),
	.w8(32'hba7d5017),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75908c),
	.w1(32'h3a7cab2a),
	.w2(32'h3bf02cc5),
	.w3(32'hbbc41735),
	.w4(32'h3b56312e),
	.w5(32'h3ab6382e),
	.w6(32'hbb5c557c),
	.w7(32'h3afe33c0),
	.w8(32'h3b2dc8f8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2f9aa),
	.w1(32'h3b1574bb),
	.w2(32'hbab4d3e4),
	.w3(32'h3b2323d0),
	.w4(32'h3b25f7c2),
	.w5(32'hbbbe4c06),
	.w6(32'h3b62cda2),
	.w7(32'hbb1b6219),
	.w8(32'hba1641e7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd21ea7),
	.w1(32'hbb22504e),
	.w2(32'hbb0de957),
	.w3(32'hbbbc5b30),
	.w4(32'hbb1aab2b),
	.w5(32'hbb76eec0),
	.w6(32'hbba4c617),
	.w7(32'hbbc554e0),
	.w8(32'hbbc5cb95),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77dbac),
	.w1(32'hbbdc4b60),
	.w2(32'hbb8ebdb2),
	.w3(32'hbb7ccb01),
	.w4(32'hbbcbce0f),
	.w5(32'hbb9e9db0),
	.w6(32'hbbb64d5e),
	.w7(32'hbba850b8),
	.w8(32'hbb4cbe8d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb588248),
	.w1(32'h3ac498e6),
	.w2(32'hbaa0c65d),
	.w3(32'hbb384673),
	.w4(32'h3bbb9da0),
	.w5(32'hba642fc4),
	.w6(32'h3b96160c),
	.w7(32'h3b699580),
	.w8(32'h3a5378ed),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89f5f0),
	.w1(32'h3be20d46),
	.w2(32'h3a833fe9),
	.w3(32'h39da8d91),
	.w4(32'hbba4f5b1),
	.w5(32'hbac4d773),
	.w6(32'h3ab23cfb),
	.w7(32'h3bd15d0c),
	.w8(32'h3baf100e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c110605),
	.w1(32'hbb03f894),
	.w2(32'hba34d4ea),
	.w3(32'hbae28921),
	.w4(32'hbab73904),
	.w5(32'hbb19deca),
	.w6(32'hbc57b35d),
	.w7(32'hbbe329d3),
	.w8(32'h3b8a363b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac84f9a),
	.w1(32'hbc14b92e),
	.w2(32'hbc1696b5),
	.w3(32'hbb554fa8),
	.w4(32'hb90e07a9),
	.w5(32'hb98d98db),
	.w6(32'h39d9e671),
	.w7(32'hbacf19f2),
	.w8(32'h3a9d2ec1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588bcc),
	.w1(32'hbbb22051),
	.w2(32'hbb718bc1),
	.w3(32'hba932610),
	.w4(32'hbb507f95),
	.w5(32'hbbc25e17),
	.w6(32'hbbc1d8d3),
	.w7(32'hbbb5bfb6),
	.w8(32'hbb9fda67),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34fbb2),
	.w1(32'hbc08c7ed),
	.w2(32'hbc605fb2),
	.w3(32'hbb377c7b),
	.w4(32'hbbf80464),
	.w5(32'hbc486724),
	.w6(32'hbb9b4676),
	.w7(32'hbc087c8c),
	.w8(32'hbafca14a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9acb2f),
	.w1(32'h3bd5ae49),
	.w2(32'h3b66f865),
	.w3(32'hbb938ee0),
	.w4(32'h397d7c1d),
	.w5(32'h3ab633d2),
	.w6(32'h3bcad915),
	.w7(32'h3c13936e),
	.w8(32'h3b803110),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18fedd),
	.w1(32'h3b7a0cf6),
	.w2(32'h3ba8488f),
	.w3(32'h3b73ee1f),
	.w4(32'h397a2a37),
	.w5(32'h399b7e14),
	.w6(32'h3a82e445),
	.w7(32'h3bf24e92),
	.w8(32'h3b03d182),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924492),
	.w1(32'h38b0d9ea),
	.w2(32'h3c246e4e),
	.w3(32'h3b32e8b2),
	.w4(32'h3c518b77),
	.w5(32'h3bb0e6c4),
	.w6(32'h3b507aff),
	.w7(32'h3c0f092b),
	.w8(32'h3bfa95f2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce2dff),
	.w1(32'h3b6a6455),
	.w2(32'h398dec85),
	.w3(32'h3b675d8d),
	.w4(32'h3b36ef61),
	.w5(32'h3aba5c89),
	.w6(32'h3b1b5ae0),
	.w7(32'h3ac65b1b),
	.w8(32'hbb577235),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0439),
	.w1(32'hbad1e17d),
	.w2(32'h39e34fa9),
	.w3(32'hbaedf2ed),
	.w4(32'h3b51a377),
	.w5(32'hb9543368),
	.w6(32'hbab7bd1f),
	.w7(32'h3b15031d),
	.w8(32'hbb6a98e9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae181d),
	.w1(32'hb9f4cc05),
	.w2(32'h3b331b51),
	.w3(32'hbb9dad6b),
	.w4(32'hbbb2be51),
	.w5(32'hbad8b5ed),
	.w6(32'hb903118b),
	.w7(32'h3af451c4),
	.w8(32'h3a1d6939),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a75bb6),
	.w1(32'h3b827a21),
	.w2(32'h3aa9014f),
	.w3(32'hbb296e57),
	.w4(32'hbbc56f19),
	.w5(32'h3a2a7f33),
	.w6(32'hbba2070c),
	.w7(32'hbb9ee65c),
	.w8(32'h3a84fd15),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ce27),
	.w1(32'hbbf150fb),
	.w2(32'hbaa621a1),
	.w3(32'h3badeafc),
	.w4(32'hbab044a9),
	.w5(32'hbac4a918),
	.w6(32'hba6ed582),
	.w7(32'hbbadd387),
	.w8(32'hbb922d03),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993738),
	.w1(32'h3c273b16),
	.w2(32'h3bd4dfc2),
	.w3(32'h3b373af3),
	.w4(32'h3c770e4e),
	.w5(32'h3c67bd6b),
	.w6(32'hbb9913bd),
	.w7(32'hbc7c6b18),
	.w8(32'hbc54a05b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0df93),
	.w1(32'h3b730445),
	.w2(32'hbb2b05bb),
	.w3(32'h3c512ba9),
	.w4(32'h3bc9f025),
	.w5(32'hba0d9e58),
	.w6(32'h3b8e0c02),
	.w7(32'hb9096d41),
	.w8(32'hbaf43d64),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4f7ae),
	.w1(32'h3cd0b083),
	.w2(32'h3ce4e10b),
	.w3(32'hbb68e36f),
	.w4(32'h3ca0e24e),
	.w5(32'h3cc3c907),
	.w6(32'h3cdd135f),
	.w7(32'h3cfa49ec),
	.w8(32'h3c72f96b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51e31c),
	.w1(32'h3bc662cb),
	.w2(32'h3bd43982),
	.w3(32'h3c59203d),
	.w4(32'h3b913d45),
	.w5(32'h3b9c0339),
	.w6(32'h3c0b48f4),
	.w7(32'h3c0bd98e),
	.w8(32'h3bcece69),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568692),
	.w1(32'h3a98e849),
	.w2(32'h3b489107),
	.w3(32'h3b699b02),
	.w4(32'h3a51ce73),
	.w5(32'h3bc8cf98),
	.w6(32'h3bbe796a),
	.w7(32'h3b63fe2a),
	.w8(32'h3b72b75a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb07d0),
	.w1(32'h3bcc45c8),
	.w2(32'h3b3e84ff),
	.w3(32'h3b9a1ce3),
	.w4(32'hbc15fcab),
	.w5(32'hbbc5c74f),
	.w6(32'h3c01ee05),
	.w7(32'hbb11c6db),
	.w8(32'h39a9de4a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26094c),
	.w1(32'hbba2e65c),
	.w2(32'hbac841cc),
	.w3(32'hbbc60532),
	.w4(32'h3a6f860b),
	.w5(32'h3a897662),
	.w6(32'hbb894e84),
	.w7(32'h3a9031ba),
	.w8(32'h3ba31d94),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7c902),
	.w1(32'hb96ba502),
	.w2(32'hb9464044),
	.w3(32'h3ba645ac),
	.w4(32'hb7e6d7c6),
	.w5(32'hbb02ce37),
	.w6(32'h39338dfc),
	.w7(32'hbab370d6),
	.w8(32'hb9c87864),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabce9b0),
	.w1(32'hbb9c2f77),
	.w2(32'hba123d2b),
	.w3(32'hb98d5ee6),
	.w4(32'h3bb585c7),
	.w5(32'hbb55c331),
	.w6(32'hba7c8886),
	.w7(32'hbba275a3),
	.w8(32'h3af5f151),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf083),
	.w1(32'hbbc6d09c),
	.w2(32'h3c9133fd),
	.w3(32'h3b1401d6),
	.w4(32'hbc86957e),
	.w5(32'h3bd7d3cf),
	.w6(32'h3b11d8be),
	.w7(32'h3cb3c597),
	.w8(32'h3cdec848),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdaee53),
	.w1(32'h3a51d029),
	.w2(32'h3bdedeed),
	.w3(32'h3c9d563e),
	.w4(32'hbae6a05e),
	.w5(32'h3b3ffd7a),
	.w6(32'h3a145775),
	.w7(32'hba51fff6),
	.w8(32'h3aafbf69),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd81fa),
	.w1(32'h3ba889b9),
	.w2(32'h3ba039fd),
	.w3(32'hbadbb3e7),
	.w4(32'hbb751740),
	.w5(32'h3989f2bc),
	.w6(32'h3aa1c997),
	.w7(32'hbadb1a35),
	.w8(32'hbafed7d9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2279fb),
	.w1(32'hb81f6f89),
	.w2(32'hba4c81a1),
	.w3(32'hbabde495),
	.w4(32'h3b907b4e),
	.w5(32'h3b90dd8e),
	.w6(32'hbafdc762),
	.w7(32'h3b1536d6),
	.w8(32'h3b530e93),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f15ab),
	.w1(32'h3b9c8157),
	.w2(32'h3c41e000),
	.w3(32'h3c05b08d),
	.w4(32'h3ad5c5e2),
	.w5(32'h3c231d77),
	.w6(32'hbb2ed85d),
	.w7(32'h3b7bfdb1),
	.w8(32'h3b9bcac5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57cb55),
	.w1(32'h3bb3ff21),
	.w2(32'h3bb90dbd),
	.w3(32'h3c7a9f00),
	.w4(32'h3b962c0b),
	.w5(32'h3bb00732),
	.w6(32'h3bec0252),
	.w7(32'h3bbcacec),
	.w8(32'h3ba4e74c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8547c7),
	.w1(32'hba7f3cdf),
	.w2(32'h3b8014fd),
	.w3(32'h3c185563),
	.w4(32'h3b36eb82),
	.w5(32'h3b776666),
	.w6(32'hba01e550),
	.w7(32'h3a637bce),
	.w8(32'h3b6cd7a0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59d22c),
	.w1(32'hbaacf4bf),
	.w2(32'hbb334aa4),
	.w3(32'h3c0265b2),
	.w4(32'h39ba8d52),
	.w5(32'hbb36a4d2),
	.w6(32'h39bc17af),
	.w7(32'h381c2f74),
	.w8(32'hbb142e1e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83fc63),
	.w1(32'h3b9811d9),
	.w2(32'h3c4b0042),
	.w3(32'hbb2e299d),
	.w4(32'h3b0ff309),
	.w5(32'h3b4f9f6f),
	.w6(32'h3b1f719f),
	.w7(32'h3bee0508),
	.w8(32'h3c3202e9),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c1416),
	.w1(32'h3bc60ee1),
	.w2(32'h3bc0d562),
	.w3(32'h3ba6b000),
	.w4(32'h3b43418a),
	.w5(32'h3ba9173e),
	.w6(32'h3bd5464f),
	.w7(32'h3ba31ea2),
	.w8(32'h3a2fb31a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e98cb),
	.w1(32'h3b7397b0),
	.w2(32'h3b5169c9),
	.w3(32'h3aee2509),
	.w4(32'h3a56d3aa),
	.w5(32'h3a655577),
	.w6(32'h3b18aef0),
	.w7(32'h3ae81fb6),
	.w8(32'h3b64f25f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba832ef),
	.w1(32'h3b7afe27),
	.w2(32'h3b1bc17d),
	.w3(32'h3b564b5f),
	.w4(32'h3ac08c64),
	.w5(32'hb610bfd8),
	.w6(32'h3a5330f6),
	.w7(32'hba57d873),
	.w8(32'h3bcd445c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaace2c3),
	.w1(32'h3b9a3754),
	.w2(32'h3bd22042),
	.w3(32'hb930bc62),
	.w4(32'hb828df75),
	.w5(32'hba867a14),
	.w6(32'h3bf045f6),
	.w7(32'h3bd35813),
	.w8(32'hba574358),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb899e25),
	.w1(32'h3b7f6d63),
	.w2(32'h3b9257a1),
	.w3(32'h3b6e2208),
	.w4(32'hbaeebe69),
	.w5(32'h3b2ad80b),
	.w6(32'hbabec56d),
	.w7(32'h3b0e14c5),
	.w8(32'hba4ece46),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd8369),
	.w1(32'hba285732),
	.w2(32'h3babc00c),
	.w3(32'hbbb1b457),
	.w4(32'h3b3e4484),
	.w5(32'h3b561ab7),
	.w6(32'h3acac34b),
	.w7(32'h3c06762b),
	.w8(32'h3bbb4859),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d163),
	.w1(32'h3b021201),
	.w2(32'h3af81779),
	.w3(32'h3b3b6932),
	.w4(32'hbb0667d8),
	.w5(32'hbb7d9474),
	.w6(32'h3b29a4f8),
	.w7(32'h3b9b7520),
	.w8(32'h3b81122b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cdc5c),
	.w1(32'h3a3bb1f0),
	.w2(32'h3b612e12),
	.w3(32'h3a837de7),
	.w4(32'hbc217b3b),
	.w5(32'hbc2a5df1),
	.w6(32'h3c10d838),
	.w7(32'h3c673de2),
	.w8(32'h3c861757),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb772c6),
	.w1(32'h3acda139),
	.w2(32'h3b53342a),
	.w3(32'hbbd8056a),
	.w4(32'hbbfeb7e3),
	.w5(32'hbbc4e1ee),
	.w6(32'h3ba16331),
	.w7(32'h3b9e70ba),
	.w8(32'h3b8fa620),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1733f2),
	.w1(32'h3b8c1888),
	.w2(32'h3b9affca),
	.w3(32'hbb25fada),
	.w4(32'hbc01f316),
	.w5(32'hbc0a0940),
	.w6(32'h3b86454d),
	.w7(32'h3bd88c6b),
	.w8(32'h3b9bd86e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34fb14),
	.w1(32'h3b857ed5),
	.w2(32'h3bde32f1),
	.w3(32'hbc31823b),
	.w4(32'hb9f4a922),
	.w5(32'h3a4b7c6e),
	.w6(32'hbbc9796b),
	.w7(32'hbb81f23b),
	.w8(32'hbb626ac9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac99e93),
	.w1(32'hbb213df6),
	.w2(32'h3b9704b5),
	.w3(32'h39336e12),
	.w4(32'h3a13a075),
	.w5(32'h3c12e4e8),
	.w6(32'hb9986ec0),
	.w7(32'h3b9d3824),
	.w8(32'h3b6ad480),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0d3f),
	.w1(32'hbaf714ce),
	.w2(32'h3bd52ac9),
	.w3(32'h3bd025a6),
	.w4(32'h3bbf8b13),
	.w5(32'h3ba4a188),
	.w6(32'h3a43f751),
	.w7(32'h3bd75c14),
	.w8(32'h3b70def2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb13bfe),
	.w1(32'h3bfc3447),
	.w2(32'h3bf0b220),
	.w3(32'h3b7c8715),
	.w4(32'h3af394e8),
	.w5(32'h3badb767),
	.w6(32'h3bd37970),
	.w7(32'h3bca9bfd),
	.w8(32'h3b75bd35),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaaf04),
	.w1(32'h3a834fe2),
	.w2(32'h3b22a0e6),
	.w3(32'h3b86eba8),
	.w4(32'hba0faa49),
	.w5(32'h3a3bfc24),
	.w6(32'h3ac091f2),
	.w7(32'h3b49d232),
	.w8(32'h3b5b4bd5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291c40),
	.w1(32'hb9ac7d34),
	.w2(32'hbc0e6229),
	.w3(32'h3b4a3f28),
	.w4(32'h3bd6ff12),
	.w5(32'hbaa394a6),
	.w6(32'hbb4ad8d5),
	.w7(32'h3b75216c),
	.w8(32'hbb254793),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81413c),
	.w1(32'h3b0dfeb7),
	.w2(32'hbb30b678),
	.w3(32'h3b09eeca),
	.w4(32'hba181e62),
	.w5(32'hbb89eab3),
	.w6(32'h3ba227b7),
	.w7(32'h3aac7485),
	.w8(32'hbaf662c3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0666a),
	.w1(32'hbb34f5f1),
	.w2(32'h3a5adee9),
	.w3(32'hbbe27aee),
	.w4(32'hbac8abed),
	.w5(32'hbb6fc63c),
	.w6(32'hbb10a24d),
	.w7(32'hb9c254b4),
	.w8(32'h3a7c4bd2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151087),
	.w1(32'h3b890feb),
	.w2(32'h3bc30e59),
	.w3(32'h3b0a4382),
	.w4(32'hbb1a0107),
	.w5(32'h3b897d8e),
	.w6(32'h3a4699a6),
	.w7(32'h3b8166f3),
	.w8(32'h3b87d1ce),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c254b),
	.w1(32'h3b000973),
	.w2(32'h3b85df60),
	.w3(32'h3bbc7d73),
	.w4(32'h3b2da45d),
	.w5(32'hba384e05),
	.w6(32'h3b6cc189),
	.w7(32'hb98adab0),
	.w8(32'h3c0b9049),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b927ac2),
	.w1(32'h3a87fe30),
	.w2(32'hbba01e0c),
	.w3(32'h3c01851d),
	.w4(32'hbbd2182e),
	.w5(32'hbb89c509),
	.w6(32'hbbccfadc),
	.w7(32'hbae7eefb),
	.w8(32'hbbdffcb9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f4ea6),
	.w1(32'h39f8819d),
	.w2(32'hbafd9829),
	.w3(32'hbba1413f),
	.w4(32'hbba1b1e0),
	.w5(32'hbb54b3e1),
	.w6(32'h3b5daf92),
	.w7(32'h3986faaf),
	.w8(32'h3bc523e0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e96b7),
	.w1(32'h3ae077e3),
	.w2(32'hbbdfba50),
	.w3(32'hb9213955),
	.w4(32'h3bb19f3c),
	.w5(32'hbab71ed8),
	.w6(32'hbb9a44ef),
	.w7(32'h3b1c9629),
	.w8(32'hba6673e3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeee3cc),
	.w1(32'h3b72b461),
	.w2(32'h3b56bf18),
	.w3(32'hb972d604),
	.w4(32'hb985aae7),
	.w5(32'h3be7666b),
	.w6(32'hbaeab3bc),
	.w7(32'h3bc14206),
	.w8(32'h3b936792),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94456e),
	.w1(32'hbb816caa),
	.w2(32'h3a00b7ca),
	.w3(32'h3b542e98),
	.w4(32'hbbabc87e),
	.w5(32'hbb5ea509),
	.w6(32'h3b0b9da7),
	.w7(32'hba0300ae),
	.w8(32'h3b8c14fd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa2252),
	.w1(32'hbb98c879),
	.w2(32'hbb816c6e),
	.w3(32'hbb48b81f),
	.w4(32'hbc1900c2),
	.w5(32'hbb95c431),
	.w6(32'hbb63b47d),
	.w7(32'hba9fd166),
	.w8(32'h3a587646),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f3e4),
	.w1(32'hba81a5a0),
	.w2(32'hbb8534e7),
	.w3(32'h3abade72),
	.w4(32'hb91c1ec5),
	.w5(32'hbb9a0f10),
	.w6(32'hba1740eb),
	.w7(32'hbb893c5d),
	.w8(32'h398f1ecc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70bfd5),
	.w1(32'h39d0cc26),
	.w2(32'hba22cf83),
	.w3(32'h3ab9feaf),
	.w4(32'hbbbd088d),
	.w5(32'hbbd55a51),
	.w6(32'hb8dbd695),
	.w7(32'h3b493d87),
	.w8(32'hbae52a43),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa70529),
	.w1(32'h3c14bf2c),
	.w2(32'h3be94820),
	.w3(32'hbb894bbf),
	.w4(32'h3bd1046c),
	.w5(32'h3bb2b360),
	.w6(32'hbb582c0b),
	.w7(32'hbb85966b),
	.w8(32'hbba9d93d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b764b53),
	.w1(32'h3b9b8af5),
	.w2(32'h3bbe568c),
	.w3(32'h39f7e30b),
	.w4(32'h3b70f78f),
	.w5(32'h3bf0333a),
	.w6(32'h3c0aab5a),
	.w7(32'h3bc0a139),
	.w8(32'h3bdaac72),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d9ab),
	.w1(32'hbaadd799),
	.w2(32'hbb37badf),
	.w3(32'h3bed9df4),
	.w4(32'hbafade98),
	.w5(32'hbb33b48d),
	.w6(32'h3a9acc0b),
	.w7(32'hb9abbd6e),
	.w8(32'h3b2e86c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab58865),
	.w1(32'h3974f807),
	.w2(32'h3980c9d8),
	.w3(32'hb9761a54),
	.w4(32'h3abaf589),
	.w5(32'hba2cc5b7),
	.w6(32'h3ab14b03),
	.w7(32'hbb823523),
	.w8(32'h3b2aa9e7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e809e4),
	.w1(32'h3c79efda),
	.w2(32'h3c8ea132),
	.w3(32'hbaeee0e6),
	.w4(32'h3c672d9c),
	.w5(32'h3c8ae539),
	.w6(32'h3c5fffd0),
	.w7(32'h3c8a5097),
	.w8(32'h3c5ea719),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c782fd0),
	.w1(32'hbba1c9f9),
	.w2(32'hbb5584ff),
	.w3(32'h3c60b3eb),
	.w4(32'h3900bad3),
	.w5(32'h3a83960b),
	.w6(32'hbab3e56b),
	.w7(32'hbb068b0e),
	.w8(32'hba96e480),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eb5b2),
	.w1(32'hbb44857c),
	.w2(32'h3a27d286),
	.w3(32'h3bb5fb32),
	.w4(32'h3bc6ffd2),
	.w5(32'h3bfa9f81),
	.w6(32'hbbbe57eb),
	.w7(32'h3b5049da),
	.w8(32'hbaa4d8ce),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815063f),
	.w1(32'h3a8481b9),
	.w2(32'h3a383c4d),
	.w3(32'h3c0b682f),
	.w4(32'h3940d682),
	.w5(32'hbb908f5f),
	.w6(32'hba4f0a6b),
	.w7(32'hbb3fe34a),
	.w8(32'hbba0517f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc053b13),
	.w1(32'hba90922e),
	.w2(32'hbb343c15),
	.w3(32'hbc184ae9),
	.w4(32'hba0274f4),
	.w5(32'hbb298146),
	.w6(32'h3b01bee9),
	.w7(32'h3a929348),
	.w8(32'h3b3c222d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad23d10),
	.w1(32'hbb4d3f9d),
	.w2(32'hbbf2a1b6),
	.w3(32'hb953784d),
	.w4(32'h3aa5b696),
	.w5(32'hbb15ea8d),
	.w6(32'hbb1aa21c),
	.w7(32'hbbf36589),
	.w8(32'hba8bada8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255bab),
	.w1(32'hb913e590),
	.w2(32'hbbcb78f7),
	.w3(32'h3bf5f75a),
	.w4(32'h3ab19bc9),
	.w5(32'hbb3212b5),
	.w6(32'h3aa62fba),
	.w7(32'hbb2141dc),
	.w8(32'h3937a6b8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb942ebf),
	.w1(32'h39697815),
	.w2(32'h3c2395bb),
	.w3(32'hbb0f9e58),
	.w4(32'h3b2f46ec),
	.w5(32'h3b981401),
	.w6(32'h3b3efad2),
	.w7(32'h3ad56702),
	.w8(32'h3b5069eb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcfdd7),
	.w1(32'h3b411fdd),
	.w2(32'h3b9a5535),
	.w3(32'h3b99f980),
	.w4(32'hbbc699ee),
	.w5(32'hbbd5c8b5),
	.w6(32'h3b71d4ce),
	.w7(32'h3b63449d),
	.w8(32'hbab6269b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dee1d),
	.w1(32'h3b8fb230),
	.w2(32'h3b4eacd0),
	.w3(32'hbc02b6e5),
	.w4(32'h3b0bbc0a),
	.w5(32'h3aafa5e4),
	.w6(32'hb99395e3),
	.w7(32'h3b144b48),
	.w8(32'h3b9c8ffc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ae129),
	.w1(32'h3b8161e4),
	.w2(32'h3aed86bc),
	.w3(32'h38e2c4db),
	.w4(32'hbae679dc),
	.w5(32'h3a2eb967),
	.w6(32'hbb3951b5),
	.w7(32'hbb2ea86d),
	.w8(32'hbbe3b262),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1e69),
	.w1(32'h3b489003),
	.w2(32'h3b9edfba),
	.w3(32'hbbca20f7),
	.w4(32'h3a1cf86a),
	.w5(32'h3b336d68),
	.w6(32'h3a11f4ba),
	.w7(32'h3b40b437),
	.w8(32'h38b898f4),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b8dfd),
	.w1(32'hb9deefe0),
	.w2(32'hbbc646c7),
	.w3(32'hb7a1fcb3),
	.w4(32'hba7e3d62),
	.w5(32'hba1ca391),
	.w6(32'hba67d79d),
	.w7(32'hbb318c06),
	.w8(32'hbaa620cb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3e349),
	.w1(32'h3bb25d1e),
	.w2(32'h3b0912b5),
	.w3(32'h3b68235b),
	.w4(32'hbacd69b9),
	.w5(32'hbb114fe9),
	.w6(32'h3c072b3c),
	.w7(32'h3a92983d),
	.w8(32'hba5969b1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb283d84),
	.w1(32'h399efb22),
	.w2(32'h3bc51adc),
	.w3(32'h3b80bb58),
	.w4(32'h39ac0a35),
	.w5(32'h3bd32ee5),
	.w6(32'h3aacd243),
	.w7(32'hbb2ee6d3),
	.w8(32'h3affd29e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5b34d),
	.w1(32'hb860d7e6),
	.w2(32'hb9b2ddc4),
	.w3(32'h3ba1cb34),
	.w4(32'h3a772e40),
	.w5(32'hba1eb97f),
	.w6(32'h39f2ffe3),
	.w7(32'h398ee75e),
	.w8(32'h3997d642),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba958602),
	.w1(32'hbbce4e50),
	.w2(32'hbad422dc),
	.w3(32'hb992ce67),
	.w4(32'hbb3b522d),
	.w5(32'h3bf824bb),
	.w6(32'hbb88cf57),
	.w7(32'h3a735a3f),
	.w8(32'hbaa27a55),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule