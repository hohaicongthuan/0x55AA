module layer_10_featuremap_40(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a0d2),
	.w1(32'hbba917c6),
	.w2(32'hbade6145),
	.w3(32'hbcabdf0f),
	.w4(32'hbc9fcbfb),
	.w5(32'hbbaa26fc),
	.w6(32'hbc107994),
	.w7(32'hbc3d4354),
	.w8(32'h3b6a8138),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a1dec),
	.w1(32'hbb7f7043),
	.w2(32'h3c5628d5),
	.w3(32'h3cd4dc7d),
	.w4(32'h3aa5bdc3),
	.w5(32'h3c9fb4db),
	.w6(32'h3c33e05f),
	.w7(32'hbbb0f5bc),
	.w8(32'h3b9b11fc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85280d),
	.w1(32'hbbb0f10d),
	.w2(32'hbb71ca3d),
	.w3(32'hbabbf56e),
	.w4(32'h3b9c6708),
	.w5(32'hbb9106dd),
	.w6(32'hbc1a7f4c),
	.w7(32'h3c155ae9),
	.w8(32'hbb9c531a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11d840),
	.w1(32'h3977c27f),
	.w2(32'h3b28de7c),
	.w3(32'hbbeb7d07),
	.w4(32'hbbd32344),
	.w5(32'hbbf73e65),
	.w6(32'h3bb7a791),
	.w7(32'h3bd1172a),
	.w8(32'hbb12758d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13155a),
	.w1(32'h3b47160b),
	.w2(32'h3ae2ea41),
	.w3(32'h3b4fd8e8),
	.w4(32'h3b72ab5b),
	.w5(32'h3c4a0471),
	.w6(32'h3c756c0a),
	.w7(32'hbbef8cc8),
	.w8(32'h3c5d6cb1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b2ff),
	.w1(32'h3b1e88b2),
	.w2(32'hbc80bce7),
	.w3(32'h3cacab36),
	.w4(32'h3c035155),
	.w5(32'hbc6877e5),
	.w6(32'h3cbde028),
	.w7(32'h3bf6046e),
	.w8(32'hbc0140b7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51d240),
	.w1(32'h3b7a9e68),
	.w2(32'h3aebead5),
	.w3(32'h3c35a56e),
	.w4(32'h3c37da84),
	.w5(32'h3b4023b6),
	.w6(32'h3c414102),
	.w7(32'h3c440234),
	.w8(32'h3bbf887f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c973ea5),
	.w1(32'h3a76dd38),
	.w2(32'hbb1c005b),
	.w3(32'h3c8312e6),
	.w4(32'h398e2b89),
	.w5(32'hbb5efc7e),
	.w6(32'h3c1becce),
	.w7(32'h3b272a57),
	.w8(32'h3c055164),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d509),
	.w1(32'hbc51bda2),
	.w2(32'h3bd27fd1),
	.w3(32'h3a89deab),
	.w4(32'hbc1a27bd),
	.w5(32'h3b1acd52),
	.w6(32'h3b20aac0),
	.w7(32'hbbbec604),
	.w8(32'h3b8c53b7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1df64f),
	.w1(32'h3c936f71),
	.w2(32'h3b825520),
	.w3(32'h3ac3ed2e),
	.w4(32'h3c47b697),
	.w5(32'h3b986ec7),
	.w6(32'h3b43a0ec),
	.w7(32'h3c6e2119),
	.w8(32'h3be71cbd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38b5af),
	.w1(32'hbb0db819),
	.w2(32'h3b9dddd4),
	.w3(32'hbb748c8d),
	.w4(32'hbb3daaf4),
	.w5(32'hbae90699),
	.w6(32'hba9ea3be),
	.w7(32'hb90833f9),
	.w8(32'hbb9ec2b9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba634e59),
	.w1(32'h3a231d87),
	.w2(32'hbb2513f4),
	.w3(32'h3bf3f63d),
	.w4(32'h3bcc3522),
	.w5(32'hbbc305f7),
	.w6(32'h3c09b7d3),
	.w7(32'h3c2dd3cf),
	.w8(32'hbb3c27ad),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515749),
	.w1(32'hbad5b0ba),
	.w2(32'h3c99a816),
	.w3(32'hba2a650e),
	.w4(32'h3b284ee9),
	.w5(32'h3c0a3a0d),
	.w6(32'hbaf1aae2),
	.w7(32'h3b41302d),
	.w8(32'h3c908404),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e6ea6),
	.w1(32'h3c4a15e8),
	.w2(32'hbc4569af),
	.w3(32'h3c543656),
	.w4(32'h3c5e679b),
	.w5(32'hbbd1cdfc),
	.w6(32'h3ca50bdf),
	.w7(32'h3c65e35c),
	.w8(32'h3bb98b91),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b863575),
	.w1(32'h3bdb80f9),
	.w2(32'h3a830674),
	.w3(32'h3c978e11),
	.w4(32'hbb914c81),
	.w5(32'hbbc6565b),
	.w6(32'h3addbb02),
	.w7(32'hbba28c07),
	.w8(32'hbb0c63fa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52ccfb),
	.w1(32'h3c27eef0),
	.w2(32'h3c1acce7),
	.w3(32'h3bcd08e7),
	.w4(32'h3b172efd),
	.w5(32'h3bc7f27d),
	.w6(32'h39c870a3),
	.w7(32'h3aea6dc8),
	.w8(32'h3c1b9058),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96587d9),
	.w1(32'hbab9ba43),
	.w2(32'h3aa7e7c6),
	.w3(32'hb9e1f139),
	.w4(32'h3968413f),
	.w5(32'h3b9e36e4),
	.w6(32'h3b44db9d),
	.w7(32'h3b556b13),
	.w8(32'h3bc9d96e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86cf23),
	.w1(32'h3c1d2e0f),
	.w2(32'h3c99e43f),
	.w3(32'h3c19b5b0),
	.w4(32'h3c3c6742),
	.w5(32'h3c8ff904),
	.w6(32'h3bbbb30b),
	.w7(32'h3bc38735),
	.w8(32'h3c90283c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73fe5),
	.w1(32'h3c6b5944),
	.w2(32'hbb13e410),
	.w3(32'h3c2bb639),
	.w4(32'h3c80412e),
	.w5(32'hbc012228),
	.w6(32'h3bd6620c),
	.w7(32'h3c2848f3),
	.w8(32'h3b5ee004),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96a290),
	.w1(32'hbb97d2cb),
	.w2(32'hbb1b51c6),
	.w3(32'hbc8d2390),
	.w4(32'hbc991b53),
	.w5(32'hbb339048),
	.w6(32'hbc4b25ac),
	.w7(32'hbca89f1b),
	.w8(32'hbaa15853),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85e374),
	.w1(32'h3a7d3b24),
	.w2(32'hbbd70c5c),
	.w3(32'hbb0837d0),
	.w4(32'hbb6f0020),
	.w5(32'hbb3a883c),
	.w6(32'hbbcb6a27),
	.w7(32'hbb48fc6d),
	.w8(32'hbb3f5adb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c98a6),
	.w1(32'h3af2298b),
	.w2(32'hbc1ca88b),
	.w3(32'hbb477278),
	.w4(32'hbbc80fb7),
	.w5(32'hbc9c1d73),
	.w6(32'h3be20c85),
	.w7(32'hbba1d709),
	.w8(32'hbc8dcfdb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96c4bc),
	.w1(32'hbc22228d),
	.w2(32'h3b1f93ba),
	.w3(32'hbcc534bd),
	.w4(32'hbcad3302),
	.w5(32'h38f8d486),
	.w6(32'hbca2d627),
	.w7(32'hbc949bef),
	.w8(32'h3b39e304),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb713e1b),
	.w1(32'h3ab4570e),
	.w2(32'h3c19981c),
	.w3(32'hbab30b12),
	.w4(32'h3af911ef),
	.w5(32'h3bed2bc3),
	.w6(32'h38e53426),
	.w7(32'h3b96540f),
	.w8(32'h3b84f904),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20224e),
	.w1(32'h3a303f14),
	.w2(32'hbcaf9971),
	.w3(32'h3ba6f165),
	.w4(32'h3ae53bfd),
	.w5(32'hbca21a97),
	.w6(32'h3c39bb92),
	.w7(32'h3b480623),
	.w8(32'hbc8ee736),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69fb77),
	.w1(32'h3ae90006),
	.w2(32'h3b925111),
	.w3(32'hbca9a8f5),
	.w4(32'hbb8cf395),
	.w5(32'hb8c3e2dd),
	.w6(32'hbc530bba),
	.w7(32'hbbf8f12f),
	.w8(32'hba20b999),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae55645),
	.w1(32'hbb85a6d5),
	.w2(32'h3a805c47),
	.w3(32'hbb839dbb),
	.w4(32'hbb8c9370),
	.w5(32'h39b405ff),
	.w6(32'hbb95f8a3),
	.w7(32'h3aa27763),
	.w8(32'h39d1ce9e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f8b04),
	.w1(32'hbae7ab84),
	.w2(32'h3bde90a9),
	.w3(32'h3ba922d3),
	.w4(32'hbb9b0f25),
	.w5(32'h3c053214),
	.w6(32'h3a7b31f6),
	.w7(32'h38c059ab),
	.w8(32'h3c7ab624),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd69a21),
	.w1(32'hbac4f894),
	.w2(32'hba704c99),
	.w3(32'h3c8f1614),
	.w4(32'h3b379aeb),
	.w5(32'h3a8a36e5),
	.w6(32'h3ca05190),
	.w7(32'h3bc0b0c4),
	.w8(32'h3c5ac21b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28a3e2),
	.w1(32'hbb6bc7de),
	.w2(32'hbc0299d0),
	.w3(32'h3c20080f),
	.w4(32'hbbbe648c),
	.w5(32'hbca5cc52),
	.w6(32'h3caaf3a6),
	.w7(32'hbaace92c),
	.w8(32'hbc86a86e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede903),
	.w1(32'h3ae474d7),
	.w2(32'h3bf34e40),
	.w3(32'hbb90f22b),
	.w4(32'hba096832),
	.w5(32'h3b7e0969),
	.w6(32'hbb7ad0d5),
	.w7(32'h398cf76f),
	.w8(32'hbb0b0582),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb159f0a),
	.w1(32'hbae295f8),
	.w2(32'h3c31de58),
	.w3(32'h3a01f364),
	.w4(32'hbba130aa),
	.w5(32'h3aefaba0),
	.w6(32'hbb20fea5),
	.w7(32'hbbb65ac0),
	.w8(32'hbc0235f2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed144),
	.w1(32'hbb9803eb),
	.w2(32'h3b8a0f83),
	.w3(32'h3aab2b76),
	.w4(32'h3aeb2088),
	.w5(32'h3b7267a5),
	.w6(32'hbb854511),
	.w7(32'hbb83091f),
	.w8(32'h3bc36b5a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42dae),
	.w1(32'h3b5c70a8),
	.w2(32'h3b2e14c3),
	.w3(32'h39e0e583),
	.w4(32'hbb1fe432),
	.w5(32'hbb6a544e),
	.w6(32'h3b948116),
	.w7(32'h3aa93a8a),
	.w8(32'hbc6be054),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47e8eb),
	.w1(32'h3c09f365),
	.w2(32'hbac3ae30),
	.w3(32'h3b8a90ed),
	.w4(32'h3c47fc3b),
	.w5(32'hbb96479d),
	.w6(32'h3a9c8d1f),
	.w7(32'h3c28d86d),
	.w8(32'hbb16b0e0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d60c2),
	.w1(32'hbb1933b8),
	.w2(32'h39528844),
	.w3(32'hbbd0bc35),
	.w4(32'hbbe6d3a9),
	.w5(32'h3b9c8670),
	.w6(32'hbc09526b),
	.w7(32'hbbce1c83),
	.w8(32'h3b221fb2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d6276),
	.w1(32'h3b5ea954),
	.w2(32'h3b1221cd),
	.w3(32'h3b3d841d),
	.w4(32'hbb981660),
	.w5(32'h3c0e3b30),
	.w6(32'h3ba41fd0),
	.w7(32'hb9da90d5),
	.w8(32'hbacac2bc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5b39),
	.w1(32'hbcbed82c),
	.w2(32'hbc9fac8b),
	.w3(32'hbc577dfc),
	.w4(32'hbd0fc745),
	.w5(32'hbcbc35e1),
	.w6(32'hbbb377ec),
	.w7(32'hbcf000c5),
	.w8(32'hbc91837d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c812773),
	.w1(32'h3b05190f),
	.w2(32'h39f19d5b),
	.w3(32'h3c26774c),
	.w4(32'h3b870f40),
	.w5(32'hbc8e096d),
	.w6(32'h3c47a078),
	.w7(32'hbac7e979),
	.w8(32'hbd023ab1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58c439),
	.w1(32'h3c3fd386),
	.w2(32'hbb8708d6),
	.w3(32'h3c58056a),
	.w4(32'h3c9030d3),
	.w5(32'hbc1ac9a9),
	.w6(32'hbba993ec),
	.w7(32'h3bf43345),
	.w8(32'hbbce2c37),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb85836),
	.w1(32'h3be6da47),
	.w2(32'h3baa13d8),
	.w3(32'hbc045993),
	.w4(32'h3bea3837),
	.w5(32'h3af492fa),
	.w6(32'hbb52e75e),
	.w7(32'h3c21828c),
	.w8(32'h3b488b2d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb742f),
	.w1(32'h3b8a36c1),
	.w2(32'hbbbe8f5a),
	.w3(32'h399019c9),
	.w4(32'h3a71c81e),
	.w5(32'hbba3b1c9),
	.w6(32'h3b881a4a),
	.w7(32'h37ed850e),
	.w8(32'hbb454fb8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc062eb4),
	.w1(32'hba2e1b48),
	.w2(32'hbb4abec5),
	.w3(32'h3b284fcb),
	.w4(32'hba645d89),
	.w5(32'h3b1bfc14),
	.w6(32'h39a491a5),
	.w7(32'hb9ac6d60),
	.w8(32'h3b67ea68),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbc62),
	.w1(32'hbbae8ac8),
	.w2(32'h3c8730c3),
	.w3(32'hb98d53cc),
	.w4(32'hbb88ffe9),
	.w5(32'h3c660f9e),
	.w6(32'h3a83ab74),
	.w7(32'hbb115a26),
	.w8(32'h3cb77ac0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24d5c),
	.w1(32'hbb7da1a1),
	.w2(32'h3bde93df),
	.w3(32'h3ba01733),
	.w4(32'h3b2cf8b3),
	.w5(32'h3c0f622e),
	.w6(32'h3c1c1f27),
	.w7(32'hb9db0e25),
	.w8(32'h3c2acf6c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f558b),
	.w1(32'h3c63e260),
	.w2(32'hbc408166),
	.w3(32'h3c986a23),
	.w4(32'h3c37d8c6),
	.w5(32'hbc22cbb2),
	.w6(32'h3c902d57),
	.w7(32'h3c2e5a81),
	.w8(32'hbc8aeac5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc810835),
	.w1(32'hbc409170),
	.w2(32'h3bf71422),
	.w3(32'hbc8f27eb),
	.w4(32'hbc3a1da3),
	.w5(32'h3a96bb9b),
	.w6(32'hbc99dde1),
	.w7(32'hbc82a202),
	.w8(32'h3b6f824f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7186b),
	.w1(32'h3c998ae4),
	.w2(32'h3c51861a),
	.w3(32'h3c03bd4d),
	.w4(32'h3c8f8a57),
	.w5(32'h3c446fd0),
	.w6(32'hba5f2b19),
	.w7(32'h3c31e2e4),
	.w8(32'h3c67b569),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35afbe),
	.w1(32'hbbe85b02),
	.w2(32'h3b828af7),
	.w3(32'h3a2d01a5),
	.w4(32'hbbec4c09),
	.w5(32'h3ba2dad9),
	.w6(32'h3a99c960),
	.w7(32'hbbf75236),
	.w8(32'hbb09ad53),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287a4a),
	.w1(32'h3b1cb730),
	.w2(32'hbbbcc6bb),
	.w3(32'h3b1909c2),
	.w4(32'h3aba3704),
	.w5(32'hbc31a4fc),
	.w6(32'hbb2fd7c4),
	.w7(32'hbb52293c),
	.w8(32'hbc3b73f6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5524a),
	.w1(32'hbc526694),
	.w2(32'hbbe3fa5b),
	.w3(32'hbcc23a63),
	.w4(32'hbc27f02d),
	.w5(32'h3c54c018),
	.w6(32'hbc3076ed),
	.w7(32'h39507515),
	.w8(32'h3c1c2bf0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63d0fe),
	.w1(32'h3c061e1e),
	.w2(32'hbac01eaa),
	.w3(32'h3cc8a5b7),
	.w4(32'h3cba5f3d),
	.w5(32'hbc8c561a),
	.w6(32'h3c862501),
	.w7(32'h3c95598d),
	.w8(32'hbcb20518),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4cb8),
	.w1(32'hbc06668b),
	.w2(32'hb96e5bd1),
	.w3(32'hbce7376c),
	.w4(32'hbc28c02f),
	.w5(32'h3b69f119),
	.w6(32'hbcd3e2bd),
	.w7(32'hbc0f463f),
	.w8(32'h3b91b083),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad37a6),
	.w1(32'h3b789bc4),
	.w2(32'h3c05c55e),
	.w3(32'h3befcdf9),
	.w4(32'h3c1625f1),
	.w5(32'h3be0b36d),
	.w6(32'h3c5d491e),
	.w7(32'h3c9184bd),
	.w8(32'h3c91644b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bc83a),
	.w1(32'hbbeca000),
	.w2(32'h3c90ce02),
	.w3(32'hbaaa2783),
	.w4(32'hbba7564f),
	.w5(32'h3bf2577b),
	.w6(32'h3be63602),
	.w7(32'hbb7a3810),
	.w8(32'h3c43c75c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c412ac7),
	.w1(32'h3bb45827),
	.w2(32'hbc84dcc7),
	.w3(32'h3c3950d9),
	.w4(32'h3bbcad86),
	.w5(32'hbbbaec1c),
	.w6(32'h3c4f074a),
	.w7(32'h3c3cbdb6),
	.w8(32'hbc510f67),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc776d3b),
	.w1(32'hbc586c09),
	.w2(32'h3c4f878e),
	.w3(32'hbca3eb82),
	.w4(32'hbc8a6a86),
	.w5(32'h3c819093),
	.w6(32'hbc6fdadf),
	.w7(32'hbc8a403d),
	.w8(32'h3c5eec6a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71ffd0),
	.w1(32'h395883ad),
	.w2(32'hbb875d8d),
	.w3(32'h3ccc57ed),
	.w4(32'h3bc0455c),
	.w5(32'hbb951547),
	.w6(32'h3ca4f002),
	.w7(32'h3b7d651c),
	.w8(32'h3beda85d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55c5b6),
	.w1(32'hbb3f2118),
	.w2(32'h3b4b88c4),
	.w3(32'hbb16d4fe),
	.w4(32'hbba42dd7),
	.w5(32'h3b9ec06e),
	.w6(32'h3c47e9b7),
	.w7(32'h3c17425a),
	.w8(32'h3ae361de),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49a206),
	.w1(32'h3becfce1),
	.w2(32'hbb0b6a4c),
	.w3(32'h3c439b1d),
	.w4(32'h3c095cc5),
	.w5(32'hbc8768f7),
	.w6(32'h3b8dd4e5),
	.w7(32'h3a9653e7),
	.w8(32'hbc62ecaf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c08ec),
	.w1(32'h3c12a725),
	.w2(32'h3cbf46cd),
	.w3(32'hbbcf5cb7),
	.w4(32'h3b3636ac),
	.w5(32'h3cf0a3c8),
	.w6(32'hbc4c8d80),
	.w7(32'h38f7f2d9),
	.w8(32'h3c9eb399),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a2e2c),
	.w1(32'hbba6edea),
	.w2(32'h3b83e2f3),
	.w3(32'h3d170cbc),
	.w4(32'h3b413549),
	.w5(32'h3bc6f1ce),
	.w6(32'h3ce0ba83),
	.w7(32'h3c28dc96),
	.w8(32'h3c084f87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab578bd),
	.w1(32'h3c003eab),
	.w2(32'h3a492543),
	.w3(32'hbbf9057a),
	.w4(32'h3b3c7d26),
	.w5(32'h3c0fe292),
	.w6(32'hbaec7227),
	.w7(32'h3c258e99),
	.w8(32'h3c07087c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42b68),
	.w1(32'h39826b13),
	.w2(32'h3b5c2566),
	.w3(32'h3b7c4273),
	.w4(32'hba74d844),
	.w5(32'h3b5b0a45),
	.w6(32'h3c5e765b),
	.w7(32'h3c3cf553),
	.w8(32'hba2189f4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad075ce),
	.w1(32'h3a6ce74b),
	.w2(32'h3bf502bb),
	.w3(32'hbba34363),
	.w4(32'hbb336e7f),
	.w5(32'h3c034a93),
	.w6(32'h3b43d2c6),
	.w7(32'h3a58acf6),
	.w8(32'h3abf04a4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03a5ce),
	.w1(32'hb937ea5f),
	.w2(32'hbbaa0e7c),
	.w3(32'h3c5219e8),
	.w4(32'h3b388636),
	.w5(32'h3b3e9f66),
	.w6(32'h3be6cc20),
	.w7(32'h3b12a6ff),
	.w8(32'h3b6135d1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2931d),
	.w1(32'hbc1a133c),
	.w2(32'h3c12049a),
	.w3(32'hbba6e21a),
	.w4(32'hbb954768),
	.w5(32'hbc149e92),
	.w6(32'h398ba172),
	.w7(32'hbbec9b80),
	.w8(32'hbc2a6310),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb5f95),
	.w1(32'hbc908272),
	.w2(32'h3c01b119),
	.w3(32'hbd1306b6),
	.w4(32'hbc8f4dc6),
	.w5(32'h3b9bd0a2),
	.w6(32'hbd2067e5),
	.w7(32'hbc1e3b90),
	.w8(32'h3abe9e8c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c70c1),
	.w1(32'h3c1e2531),
	.w2(32'h3c0fbdbe),
	.w3(32'hba9d130e),
	.w4(32'h3c062b2d),
	.w5(32'h3c2bce79),
	.w6(32'hbbbb47b0),
	.w7(32'h3bf26f5e),
	.w8(32'h3c825c2a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c399774),
	.w1(32'h39f82b4f),
	.w2(32'hbcb5421d),
	.w3(32'h3c4ef41f),
	.w4(32'hbaab0098),
	.w5(32'hbd0edd5b),
	.w6(32'h3c815e5b),
	.w7(32'h3aab101d),
	.w8(32'hbd0e1d56),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9eebc),
	.w1(32'h3c06030c),
	.w2(32'h3c2fe57a),
	.w3(32'hbcee6ca5),
	.w4(32'h3bbd11f3),
	.w5(32'h3c5b736c),
	.w6(32'hbce8f866),
	.w7(32'h3b8f6eb5),
	.w8(32'h3c0e624e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ac99),
	.w1(32'hbb4d50ca),
	.w2(32'hbc55c81a),
	.w3(32'h3c6054a1),
	.w4(32'h3b38ff60),
	.w5(32'hbc58999b),
	.w6(32'h3c2fc038),
	.w7(32'h3bf0dbad),
	.w8(32'hbc58c306),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e01b6),
	.w1(32'hbb9b21f8),
	.w2(32'hbae5f8d1),
	.w3(32'hbce941a6),
	.w4(32'hbc75463e),
	.w5(32'h3c2b81be),
	.w6(32'hbcf5fa5a),
	.w7(32'hbc8c5d68),
	.w8(32'h3c292ec6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed5321),
	.w1(32'hbc0e9744),
	.w2(32'h3b66d632),
	.w3(32'h3ca6afd8),
	.w4(32'h3a14741c),
	.w5(32'hbb391ec5),
	.w6(32'h3ca6540f),
	.w7(32'h3b8a423d),
	.w8(32'hb916e659),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfb754),
	.w1(32'h3b8b07b6),
	.w2(32'hbc34cec7),
	.w3(32'hbc08b387),
	.w4(32'hbb82bc10),
	.w5(32'hbc4e58cb),
	.w6(32'hbc01e567),
	.w7(32'hbb4f708a),
	.w8(32'hbc70f395),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88d33c),
	.w1(32'hbc22ebee),
	.w2(32'h3c22e7c9),
	.w3(32'hbcd394f2),
	.w4(32'hbc62af2c),
	.w5(32'h3ad8c273),
	.w6(32'hbc984222),
	.w7(32'hbc67ea4f),
	.w8(32'h3b6fa2d6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55adf4),
	.w1(32'hbb9627d0),
	.w2(32'h3c2ade8a),
	.w3(32'hbb83a7e7),
	.w4(32'hba51b438),
	.w5(32'h3b9a9119),
	.w6(32'hbbaf0e29),
	.w7(32'h3aae14b6),
	.w8(32'h39043f4f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10e579),
	.w1(32'hbc31683a),
	.w2(32'hbc04304c),
	.w3(32'hbbba40ee),
	.w4(32'hbb54ad66),
	.w5(32'hbc8e6bc0),
	.w6(32'h3ba4a70c),
	.w7(32'hb97fb642),
	.w8(32'hbc710943),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373746),
	.w1(32'h3c19b6b6),
	.w2(32'h3b9e8412),
	.w3(32'hbbfceeb2),
	.w4(32'h3b83e8d4),
	.w5(32'hb9ea33c9),
	.w6(32'hbc0d31a0),
	.w7(32'hbb6906fd),
	.w8(32'h3bb909dc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f828),
	.w1(32'h3aeaebf5),
	.w2(32'hbab9e535),
	.w3(32'hbbdfbf82),
	.w4(32'h3ba81efc),
	.w5(32'hbbd0ba4b),
	.w6(32'h3a33b020),
	.w7(32'h3b813587),
	.w8(32'hba788d70),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f643e),
	.w1(32'hbad445a4),
	.w2(32'h3bbc96f1),
	.w3(32'hbc49ed5d),
	.w4(32'hbbf2d4b8),
	.w5(32'hba315c6b),
	.w6(32'hbc09bd75),
	.w7(32'hbbbc7d89),
	.w8(32'h3a9fdab8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a0dc1),
	.w1(32'h3c1f62cc),
	.w2(32'h3c1e61ca),
	.w3(32'hb9d5f36f),
	.w4(32'h3be731ec),
	.w5(32'h3c828b1d),
	.w6(32'hb9709904),
	.w7(32'h3c094f6f),
	.w8(32'h3c4d52ec),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7a12),
	.w1(32'h3b58850a),
	.w2(32'h3c089ae4),
	.w3(32'h3c453fd2),
	.w4(32'h3bcaa0bf),
	.w5(32'h3cd7044d),
	.w6(32'h3c022380),
	.w7(32'h3c445414),
	.w8(32'h3c96d71c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b441a2d),
	.w1(32'hbc24b1f1),
	.w2(32'hbc97bf6c),
	.w3(32'h3bca04dc),
	.w4(32'hbbaddbfe),
	.w5(32'hbc7bd2c5),
	.w6(32'h3b4e18de),
	.w7(32'hbb3f8290),
	.w8(32'hbcae1d06),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4be57f),
	.w1(32'hbc4bef99),
	.w2(32'h3a8715c2),
	.w3(32'hbcc2f2d9),
	.w4(32'hbca9a022),
	.w5(32'h3c076c30),
	.w6(32'hbcd5d5f1),
	.w7(32'hbca33137),
	.w8(32'h3b0ba624),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befc216),
	.w1(32'hb81bac29),
	.w2(32'h3b9ab8e6),
	.w3(32'h3c78811a),
	.w4(32'h3b935125),
	.w5(32'h3b86ada7),
	.w6(32'h3c1f1ff5),
	.w7(32'h3c0afa17),
	.w8(32'h3bdf979d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f04f6),
	.w1(32'h3bb2cde1),
	.w2(32'hbb2abafa),
	.w3(32'h3c9e6742),
	.w4(32'h3c09a8b6),
	.w5(32'hbbb7676b),
	.w6(32'h3c96e42e),
	.w7(32'h3c136454),
	.w8(32'hbb9c382d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe3b4d),
	.w1(32'h3a8851be),
	.w2(32'hbbdc858d),
	.w3(32'hba0890fe),
	.w4(32'h3a61a66b),
	.w5(32'hbc8004ae),
	.w6(32'h3aa6980c),
	.w7(32'h3b117d3a),
	.w8(32'hbc8c871b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7634ae),
	.w1(32'hbc401625),
	.w2(32'h3b8088fc),
	.w3(32'hbcbc532f),
	.w4(32'hbca32ef5),
	.w5(32'hbb4f14f3),
	.w6(32'hbc96ebd1),
	.w7(32'hbc5f9ff0),
	.w8(32'hbc3a748d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b358047),
	.w1(32'h3c1b676a),
	.w2(32'h3c2de9d6),
	.w3(32'h39de7e9c),
	.w4(32'h3c164f52),
	.w5(32'h3bb6a33b),
	.w6(32'hbbec0056),
	.w7(32'h3a925693),
	.w8(32'hbc4ab0a8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c715dd3),
	.w1(32'hbabb3309),
	.w2(32'hbc667bc8),
	.w3(32'h3a2a291c),
	.w4(32'hbc1bfb44),
	.w5(32'hbc8ad557),
	.w6(32'hbc2c24f9),
	.w7(32'hbc55479e),
	.w8(32'hbc7f7447),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d9113),
	.w1(32'hbae9852f),
	.w2(32'h3ba7bfd1),
	.w3(32'hbbe6b624),
	.w4(32'h3952ebcc),
	.w5(32'h3b426f3d),
	.w6(32'hbb49ef94),
	.w7(32'h39d64254),
	.w8(32'h3921635f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad351a),
	.w1(32'hbb68fff0),
	.w2(32'hbc06b41a),
	.w3(32'h3b5868dd),
	.w4(32'hbbd3747f),
	.w5(32'hbc4f9fc1),
	.w6(32'h3bd4a534),
	.w7(32'hbb940ab6),
	.w8(32'hbc6387d8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb417500),
	.w1(32'h3b534210),
	.w2(32'h3c99773b),
	.w3(32'hbaf791e8),
	.w4(32'h3b903698),
	.w5(32'h3b6e21db),
	.w6(32'hba1bb9f7),
	.w7(32'h3b05f332),
	.w8(32'h3b91fd77),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb321114),
	.w1(32'h3c10e5d3),
	.w2(32'h3c0c829b),
	.w3(32'hbc68aa64),
	.w4(32'h3a4b6163),
	.w5(32'h3c8adb58),
	.w6(32'hbb9fa4ff),
	.w7(32'hba897a63),
	.w8(32'hba1b9af1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5613c0),
	.w1(32'hb97e20b8),
	.w2(32'hbc97b7fa),
	.w3(32'h3c936aab),
	.w4(32'h3bafa271),
	.w5(32'hbc84e0b7),
	.w6(32'h3ba0d3b9),
	.w7(32'hbadd7015),
	.w8(32'hbc343e0e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9704b2),
	.w1(32'hbc0c418a),
	.w2(32'hbc93a35d),
	.w3(32'hbc9152df),
	.w4(32'hbc2abb1d),
	.w5(32'hbc808aaa),
	.w6(32'hbbf26d45),
	.w7(32'hbb314fa8),
	.w8(32'hbc336b7b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6423a8),
	.w1(32'h3ac17d21),
	.w2(32'h3c43f7d5),
	.w3(32'hbcbfa671),
	.w4(32'hbc4e924d),
	.w5(32'h3c9c9eb5),
	.w6(32'hbcb88bd6),
	.w7(32'hbc7345d3),
	.w8(32'h3c89a35c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3b226),
	.w1(32'h3c078331),
	.w2(32'hbb58d900),
	.w3(32'h3bde0b81),
	.w4(32'h3b3565c6),
	.w5(32'hbbfe03fe),
	.w6(32'h3c22cfa5),
	.w7(32'hbb6f2669),
	.w8(32'h3b32eeac),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceadd47),
	.w1(32'h3b26e698),
	.w2(32'h3c3d08f2),
	.w3(32'hbcf62609),
	.w4(32'hbc90d79d),
	.w5(32'h3bf424ac),
	.w6(32'hbd173a1c),
	.w7(32'hbc89851f),
	.w8(32'h3b1ae393),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d15c4),
	.w1(32'hbc3424f7),
	.w2(32'hbc07f5b2),
	.w3(32'h3a19cc55),
	.w4(32'hbc66a759),
	.w5(32'hbc930e3e),
	.w6(32'h3b4aa25a),
	.w7(32'hbc5654e3),
	.w8(32'hbc8c24ba),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4b06c),
	.w1(32'h3b6222e0),
	.w2(32'hbb2742d4),
	.w3(32'h39c0cdd9),
	.w4(32'hbc27f781),
	.w5(32'h3b87713d),
	.w6(32'h3b46932c),
	.w7(32'hbbd8afc0),
	.w8(32'hbb859a93),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba431f5c),
	.w1(32'h3bc38cc0),
	.w2(32'h3aaebed0),
	.w3(32'h3c8aa59a),
	.w4(32'h3c49a81e),
	.w5(32'hbac91258),
	.w6(32'h3be0a2c4),
	.w7(32'h3bdce44c),
	.w8(32'hba683c7a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d3070),
	.w1(32'h3bc8ca0f),
	.w2(32'hbae353a6),
	.w3(32'hbc930ea9),
	.w4(32'h3aa969d9),
	.w5(32'hbb2f1c15),
	.w6(32'hbc416142),
	.w7(32'h3b1a22a1),
	.w8(32'hbb2b51ea),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2573a7),
	.w1(32'h3b69710e),
	.w2(32'h3c28c783),
	.w3(32'h3c652ec1),
	.w4(32'h3bd3ec97),
	.w5(32'h3c3bd766),
	.w6(32'h3c25cd39),
	.w7(32'hbc14c7cc),
	.w8(32'h3bd7204c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdab73b),
	.w1(32'h3bc4eb46),
	.w2(32'h3c45fdea),
	.w3(32'h3c14a39f),
	.w4(32'h3c0ec2b8),
	.w5(32'h3c291bee),
	.w6(32'h3bdb841f),
	.w7(32'h3c3a2a73),
	.w8(32'h3c5639b2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d91f8),
	.w1(32'h3c122e7d),
	.w2(32'hbbcceef8),
	.w3(32'h3c583128),
	.w4(32'h3c14821b),
	.w5(32'hbc0d2e10),
	.w6(32'h3c3a2d7f),
	.w7(32'h3c497079),
	.w8(32'hbb694d24),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54b1ca),
	.w1(32'hbb189010),
	.w2(32'hbb533cbf),
	.w3(32'hbccac8f5),
	.w4(32'hbc38c368),
	.w5(32'hbc961a72),
	.w6(32'hbc63bde4),
	.w7(32'hbba96cc7),
	.w8(32'hbc2b645c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac44c73),
	.w1(32'h3bc0a2d3),
	.w2(32'h3c689eef),
	.w3(32'hbbfeeb91),
	.w4(32'h3bc24bf0),
	.w5(32'h3c2b4f21),
	.w6(32'hbc9f4193),
	.w7(32'h3ae43109),
	.w8(32'h3c203984),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad43f8e),
	.w1(32'hbc28b65d),
	.w2(32'hbbedd7c5),
	.w3(32'h3be8eb6f),
	.w4(32'hbc14d7cc),
	.w5(32'hbbb33ca0),
	.w6(32'h3922c6f0),
	.w7(32'hbc0078be),
	.w8(32'hbbef7c9e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3041c),
	.w1(32'hbbb55f21),
	.w2(32'hbc2fb9e9),
	.w3(32'hbb8d4b14),
	.w4(32'hbb905416),
	.w5(32'hbc7ad443),
	.w6(32'h3a598678),
	.w7(32'hbc299966),
	.w8(32'hbc4f2cb9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ab6b5),
	.w1(32'hbb6f470f),
	.w2(32'h3ca84285),
	.w3(32'hbc1dfaee),
	.w4(32'hb9f93833),
	.w5(32'h3ccfd5b3),
	.w6(32'hbbb7ec3d),
	.w7(32'h3b31821d),
	.w8(32'h3c4fc254),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3516f),
	.w1(32'h3aed4987),
	.w2(32'h395ad9ec),
	.w3(32'h3bc99621),
	.w4(32'h3b870f99),
	.w5(32'h3be79e43),
	.w6(32'hbbabb228),
	.w7(32'hbb981828),
	.w8(32'h3b7fcf9c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfa6f3),
	.w1(32'hbb0af0df),
	.w2(32'h3bfb2be7),
	.w3(32'h3ae51eab),
	.w4(32'hbc08b14d),
	.w5(32'h3c42f0b9),
	.w6(32'hbbe9cfc6),
	.w7(32'hb92f98ad),
	.w8(32'h3a90bc14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cdb8c),
	.w1(32'hbbeff0ac),
	.w2(32'hbc17a6ec),
	.w3(32'h3bb50288),
	.w4(32'hbbc712af),
	.w5(32'hbc3ce0be),
	.w6(32'hbab71849),
	.w7(32'hbb899fcf),
	.w8(32'hbb6a6a49),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16faf),
	.w1(32'hbb3b0423),
	.w2(32'hbaa2c2f0),
	.w3(32'hbc113046),
	.w4(32'hbb9ff71d),
	.w5(32'hb9bda5b0),
	.w6(32'hba8ec624),
	.w7(32'hbb4ed509),
	.w8(32'hbaa34e8c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176c5c),
	.w1(32'hbae1fa0d),
	.w2(32'hb9f439ac),
	.w3(32'h3b295b56),
	.w4(32'hb822e411),
	.w5(32'hb98c8160),
	.w6(32'h3bca663f),
	.w7(32'h3c2fcb24),
	.w8(32'h3b4bbd57),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92daeb),
	.w1(32'hbb4a26e5),
	.w2(32'h3b1810f7),
	.w3(32'hbb6d46ae),
	.w4(32'hbba8246b),
	.w5(32'hbba9efc9),
	.w6(32'h3c05af57),
	.w7(32'h3b559eec),
	.w8(32'h3b9a8c28),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836fa1),
	.w1(32'h3bca1a97),
	.w2(32'h3ad2840f),
	.w3(32'h3b90a6fd),
	.w4(32'h3c43ea0e),
	.w5(32'hbba5822f),
	.w6(32'h3ac1d99f),
	.w7(32'h3b000908),
	.w8(32'h3b6c9c5f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a343c94),
	.w1(32'hbacac8c4),
	.w2(32'h3b660b6c),
	.w3(32'hbb228d21),
	.w4(32'hb92e55fe),
	.w5(32'hbb955524),
	.w6(32'h3b8bc78c),
	.w7(32'h3a92e708),
	.w8(32'hbb70aa1d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aaa79),
	.w1(32'h3b91d87c),
	.w2(32'hbb78d479),
	.w3(32'hbc16241e),
	.w4(32'h3b2a732b),
	.w5(32'hbbf19ab1),
	.w6(32'hbbaac170),
	.w7(32'hbb3a0807),
	.w8(32'hbbbb76c5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9346f07),
	.w1(32'h3ab44e48),
	.w2(32'hb908313a),
	.w3(32'hbb99390c),
	.w4(32'hbb507cb3),
	.w5(32'hbbff3464),
	.w6(32'hbb7ee6ab),
	.w7(32'hbaea90fb),
	.w8(32'hbbdc56c3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8a30d),
	.w1(32'hbb9c5774),
	.w2(32'h3b3753b4),
	.w3(32'hbc2ef93d),
	.w4(32'hbc213d76),
	.w5(32'hbb6d460d),
	.w6(32'hbbf32ff0),
	.w7(32'hbc1a973f),
	.w8(32'hbaeaf2b3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895427),
	.w1(32'h3bc6744b),
	.w2(32'h3b762799),
	.w3(32'h3bf7d8c6),
	.w4(32'h3c4077f6),
	.w5(32'h3c2acd7d),
	.w6(32'h3bcd054a),
	.w7(32'h3c340952),
	.w8(32'h3c4b4c83),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac167b),
	.w1(32'h3a8fd5e3),
	.w2(32'h3b6341f4),
	.w3(32'h3c575958),
	.w4(32'h3bc8dd49),
	.w5(32'h3bdcadff),
	.w6(32'h3c47ea29),
	.w7(32'h3b9d0663),
	.w8(32'h3c642949),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6006),
	.w1(32'h3a5b7ece),
	.w2(32'hbb4aa1fd),
	.w3(32'h3c46ed1f),
	.w4(32'hbb8c0f77),
	.w5(32'hbbdd7141),
	.w6(32'hbbbcd033),
	.w7(32'hbbc80d6f),
	.w8(32'hbc160e0e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c2ea9),
	.w1(32'hbbbd8001),
	.w2(32'hbc975e1c),
	.w3(32'hbca059f7),
	.w4(32'hbc075e2c),
	.w5(32'hbcf2d69a),
	.w6(32'hbca470e8),
	.w7(32'hbb78ca3b),
	.w8(32'hbcd891d8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06bf5d),
	.w1(32'hbb627980),
	.w2(32'h3c349e86),
	.w3(32'hbd159dda),
	.w4(32'hbc63ef03),
	.w5(32'h3ca90fdd),
	.w6(32'hbd1d4555),
	.w7(32'hbc077edf),
	.w8(32'h3c9d6097),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d6b29),
	.w1(32'h3c45175a),
	.w2(32'h3bf8432a),
	.w3(32'h3cf8893c),
	.w4(32'h3c8677b7),
	.w5(32'h3c3a9163),
	.w6(32'h3ccff207),
	.w7(32'h3c884bbb),
	.w8(32'h3c69c795),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4f5a9),
	.w1(32'h3b6714d0),
	.w2(32'h3b317b83),
	.w3(32'h3c2b1ccb),
	.w4(32'h3c2fefda),
	.w5(32'h3c4e148f),
	.w6(32'hbb895a09),
	.w7(32'hb9ddae63),
	.w8(32'h3c8c27e2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef30f6),
	.w1(32'hb9f4387c),
	.w2(32'hbb2053aa),
	.w3(32'h3c50617a),
	.w4(32'h3b350e05),
	.w5(32'hba2b72bd),
	.w6(32'h3c5f12de),
	.w7(32'h3ac400b0),
	.w8(32'h3c56e221),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22b21),
	.w1(32'h39ae2faf),
	.w2(32'hbbfc9e41),
	.w3(32'hb89d1f8f),
	.w4(32'hba60d572),
	.w5(32'hbc9a31b3),
	.w6(32'h3b9b7838),
	.w7(32'h3a8e1f74),
	.w8(32'hbc01e1dc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b685),
	.w1(32'h3bc5eeb2),
	.w2(32'h3b828941),
	.w3(32'hbc144982),
	.w4(32'hbbef39e0),
	.w5(32'hbba6704d),
	.w6(32'hbb1bc5c0),
	.w7(32'hbb57a858),
	.w8(32'hb9a69f00),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d812),
	.w1(32'h3b571c15),
	.w2(32'h3a8fbcfd),
	.w3(32'h3bf78e9e),
	.w4(32'h3c40f2e8),
	.w5(32'hbc317b1e),
	.w6(32'h3bec4479),
	.w7(32'h3c3640cc),
	.w8(32'hbb8c9ef7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe673a4),
	.w1(32'h3c2486d3),
	.w2(32'h3c5a1ce3),
	.w3(32'hbc75fa74),
	.w4(32'h3b75f027),
	.w5(32'h3c6963de),
	.w6(32'hbc67e51a),
	.w7(32'h3b7a0e0c),
	.w8(32'h3c9bf466),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74c40b),
	.w1(32'hbb61afdc),
	.w2(32'h3bd1cace),
	.w3(32'h3b719c9b),
	.w4(32'hbb3854fe),
	.w5(32'h3c43e6ff),
	.w6(32'h3c5c5277),
	.w7(32'hbac66dc1),
	.w8(32'hbb6e5aec),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfac78a),
	.w1(32'hb90de8eb),
	.w2(32'hbb76fbd1),
	.w3(32'h3c4883dc),
	.w4(32'h3b2e763f),
	.w5(32'hbc1a224c),
	.w6(32'hba23b000),
	.w7(32'hbaf9208d),
	.w8(32'hbba94a7b),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb5228),
	.w1(32'h3b1e8e0a),
	.w2(32'hba25332b),
	.w3(32'hbc1cf23e),
	.w4(32'hba7465c6),
	.w5(32'hbbbf0cc0),
	.w6(32'hbbea5daf),
	.w7(32'h3a9c5bce),
	.w8(32'hbb407840),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe586a6),
	.w1(32'h3b0f94d6),
	.w2(32'hb9854def),
	.w3(32'hbc154ef1),
	.w4(32'hbaa4e21d),
	.w5(32'hbb8607a5),
	.w6(32'hbc3f1b1c),
	.w7(32'hbac73133),
	.w8(32'h3983f041),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d5f70),
	.w1(32'hb9e4e145),
	.w2(32'hb8b279b3),
	.w3(32'h39fea358),
	.w4(32'h3b64d269),
	.w5(32'hbbf6236f),
	.w6(32'hbaf44b03),
	.w7(32'hba95d588),
	.w8(32'hbba28715),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4073f2),
	.w1(32'h3a3879d5),
	.w2(32'h3c1c0738),
	.w3(32'hbbc67419),
	.w4(32'hbb28153e),
	.w5(32'h3c433a37),
	.w6(32'hbbc73e8c),
	.w7(32'hbb7f167f),
	.w8(32'h3ba9824e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c872021),
	.w1(32'hbaa81135),
	.w2(32'hba9f6252),
	.w3(32'h3c87cf88),
	.w4(32'h3aa45489),
	.w5(32'hbaf799b6),
	.w6(32'h3c96eab4),
	.w7(32'hb979dc53),
	.w8(32'hbc29d7e9),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce0818),
	.w1(32'hbb1e719e),
	.w2(32'hbbdecbbc),
	.w3(32'h3c2f1e70),
	.w4(32'hbaa9fb17),
	.w5(32'hbc56b80a),
	.w6(32'h3ab29469),
	.w7(32'hbb01f0dc),
	.w8(32'hbbe74b7c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f160),
	.w1(32'hbb43fe7a),
	.w2(32'hbb924a65),
	.w3(32'hbccc2bc1),
	.w4(32'hbc3e42b2),
	.w5(32'hbbd7d67e),
	.w6(32'hbc5c0394),
	.w7(32'hbbc9bee1),
	.w8(32'hbb9b3fda),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4abcfb),
	.w1(32'h3b777bd9),
	.w2(32'hbb3d7686),
	.w3(32'h3aacb514),
	.w4(32'h3bc5aff7),
	.w5(32'hba85c8da),
	.w6(32'h3a8c5ef3),
	.w7(32'h3bcdac5a),
	.w8(32'h3b929712),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade87fb),
	.w1(32'hb968edc6),
	.w2(32'h3b65e54a),
	.w3(32'h3b653805),
	.w4(32'h3ac5d408),
	.w5(32'h3ad15469),
	.w6(32'h3b877794),
	.w7(32'h3b3e56ec),
	.w8(32'h3bc85756),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3925a),
	.w1(32'h38a577d8),
	.w2(32'h3b7bb15d),
	.w3(32'h3bdb67a1),
	.w4(32'h3b91e2bf),
	.w5(32'hbb9a1abb),
	.w6(32'h3bfb92f3),
	.w7(32'h3bbf4ed1),
	.w8(32'hbc3931d8),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8aadfb),
	.w1(32'h3bb57d18),
	.w2(32'hb90762ad),
	.w3(32'h3c9eb83d),
	.w4(32'h3c0b98c5),
	.w5(32'hbbca60d1),
	.w6(32'h3b12818f),
	.w7(32'h3b9b1cd3),
	.w8(32'hba037d9d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d1351),
	.w1(32'hbb0fafce),
	.w2(32'hbc5a0618),
	.w3(32'hbc9de208),
	.w4(32'hbc18839b),
	.w5(32'hbc35cb90),
	.w6(32'hbc50d649),
	.w7(32'hbbc18006),
	.w8(32'hbbeb0222),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0777ad),
	.w1(32'h3baf410b),
	.w2(32'h3c18cb7e),
	.w3(32'hbc76f3ca),
	.w4(32'hbb9d6be8),
	.w5(32'h3b8e297a),
	.w6(32'hbc882016),
	.w7(32'hbc291298),
	.w8(32'h3c00eb79),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4830e9),
	.w1(32'hba2f1e02),
	.w2(32'hbbf545e6),
	.w3(32'h3c08ea85),
	.w4(32'h3ba8dc28),
	.w5(32'hbc72a884),
	.w6(32'h3915a362),
	.w7(32'hba3542b2),
	.w8(32'hbc284566),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf80c40),
	.w1(32'h3b2e3960),
	.w2(32'h3c8c8725),
	.w3(32'hbc65d845),
	.w4(32'hbba207bb),
	.w5(32'h3c29e707),
	.w6(32'hbc06221d),
	.w7(32'hbb9f90f5),
	.w8(32'h3bf655b9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41f013),
	.w1(32'hbb7fc6bd),
	.w2(32'h3c1d784b),
	.w3(32'h3c1c94e0),
	.w4(32'hbbab9ed8),
	.w5(32'h3b59629f),
	.w6(32'h3c2b570a),
	.w7(32'h3b85d778),
	.w8(32'h3a457fea),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d86ad),
	.w1(32'hbab6b98f),
	.w2(32'h3c3c8ae7),
	.w3(32'h3c10677e),
	.w4(32'hba9dd269),
	.w5(32'h3bb742ac),
	.w6(32'h3beb2f8e),
	.w7(32'hbab9e9ab),
	.w8(32'hbb0379e6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c860b),
	.w1(32'h3c07c539),
	.w2(32'h3ba727ba),
	.w3(32'h39e3aebf),
	.w4(32'h3b1a6b26),
	.w5(32'h3b623c3e),
	.w6(32'hba038337),
	.w7(32'h38c326c7),
	.w8(32'h3b65256c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b237160),
	.w1(32'h3a444b7a),
	.w2(32'hbc141010),
	.w3(32'hbb36d577),
	.w4(32'hbaecf4ca),
	.w5(32'hbbdd474d),
	.w6(32'h3a3cedaf),
	.w7(32'hbaa0d980),
	.w8(32'hbb94539e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437324),
	.w1(32'h3b81cb47),
	.w2(32'h3976378d),
	.w3(32'h3c18c8b0),
	.w4(32'h3c1f9834),
	.w5(32'hbb509ca6),
	.w6(32'h3c30851a),
	.w7(32'h3c64d63a),
	.w8(32'hbb0cbf66),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58920b),
	.w1(32'hbb2aad7c),
	.w2(32'hbcc11e9a),
	.w3(32'h3b170147),
	.w4(32'h391fb0ea),
	.w5(32'hbd437c27),
	.w6(32'h3ad291fb),
	.w7(32'hbb180314),
	.w8(32'hbd076602),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd26ed4c),
	.w1(32'hbcd7a7f5),
	.w2(32'h3b359c5a),
	.w3(32'hbd9777ea),
	.w4(32'hbd6ea2f3),
	.w5(32'h3b8428dc),
	.w6(32'hbd5b6009),
	.w7(32'hbd1db59c),
	.w8(32'h3bcc9e99),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7dfe4),
	.w1(32'h3b8e34d9),
	.w2(32'hb9f54736),
	.w3(32'h3bbb49ae),
	.w4(32'h3ba74b65),
	.w5(32'h3c219198),
	.w6(32'h3bcae374),
	.w7(32'h3be89f54),
	.w8(32'h3aad1408),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37ea5),
	.w1(32'h3bf98fae),
	.w2(32'h3ccc5350),
	.w3(32'h3bcd0d78),
	.w4(32'h3c00367b),
	.w5(32'h3bc97d6b),
	.w6(32'hbb50bcaa),
	.w7(32'h3b0bb95d),
	.w8(32'h3cac079f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29ff92),
	.w1(32'h3c6415d7),
	.w2(32'h3a68451a),
	.w3(32'hbcb1bfd2),
	.w4(32'hbbcd068c),
	.w5(32'hbb88b3aa),
	.w6(32'hbb6baed3),
	.w7(32'h3c222f9b),
	.w8(32'hbac5e059),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971006),
	.w1(32'h3b97f9a6),
	.w2(32'h3bdb6de0),
	.w3(32'hbb8fb1d6),
	.w4(32'h3b845107),
	.w5(32'h3cb53648),
	.w6(32'hbb1f46b8),
	.w7(32'h3c220474),
	.w8(32'h3c433f8d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd03f0f),
	.w1(32'h3c502409),
	.w2(32'hbc3e905e),
	.w3(32'h3d59c412),
	.w4(32'h3d24d00d),
	.w5(32'hbbb5549f),
	.w6(32'h3d1a94d5),
	.w7(32'h3cd35b0d),
	.w8(32'hbc06fc5a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6d48),
	.w1(32'h3919f7bd),
	.w2(32'h3c265d7c),
	.w3(32'hbb5e8e33),
	.w4(32'h3aeaf818),
	.w5(32'h3b6f8962),
	.w6(32'hbb7e5183),
	.w7(32'h3c0364f3),
	.w8(32'h3c849782),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2be94),
	.w1(32'h3c9e1977),
	.w2(32'hba917473),
	.w3(32'hbb3016f2),
	.w4(32'h3c3278a5),
	.w5(32'h378875c9),
	.w6(32'h3c66f821),
	.w7(32'h3ccc80e6),
	.w8(32'hbb9975b9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bc484),
	.w1(32'hbad29587),
	.w2(32'hbbcbc609),
	.w3(32'h3b3f48ed),
	.w4(32'h3b5ba10d),
	.w5(32'hbaf824c0),
	.w6(32'h3b9a38a7),
	.w7(32'h3a4408d2),
	.w8(32'h3bb30aae),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e3235),
	.w1(32'hbbd17a9c),
	.w2(32'h39ef2352),
	.w3(32'hbab007f3),
	.w4(32'hbbaecf01),
	.w5(32'hbbe4b4ab),
	.w6(32'h3bd6f315),
	.w7(32'hbaa129b0),
	.w8(32'hbbfb4ae6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab37eb5),
	.w1(32'h3a732be3),
	.w2(32'h3a7d8b19),
	.w3(32'hbb25c0da),
	.w4(32'hbbee1776),
	.w5(32'h3c014cd6),
	.w6(32'hbc63ccbd),
	.w7(32'hbc170b37),
	.w8(32'h383d70f5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964680e),
	.w1(32'h39fd385e),
	.w2(32'h3bc4e1dc),
	.w3(32'h3c24245f),
	.w4(32'h3c366cfc),
	.w5(32'h3b630efe),
	.w6(32'h3b4fe776),
	.w7(32'h3b6ad540),
	.w8(32'h3bb83418),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ad62),
	.w1(32'h3b4fcca3),
	.w2(32'hbbea4392),
	.w3(32'h3c15518c),
	.w4(32'h3b6de0c9),
	.w5(32'h3c665739),
	.w6(32'h3babae02),
	.w7(32'h3bb9f04c),
	.w8(32'hba88c86d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9dfb3c),
	.w1(32'h3b4c7258),
	.w2(32'hb9f93b30),
	.w3(32'h3d46d812),
	.w4(32'h3d060d84),
	.w5(32'hbbf9bed2),
	.w6(32'h3cea2eff),
	.w7(32'h3c58b8db),
	.w8(32'hbb8e2b09),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108114),
	.w1(32'h3bd928b6),
	.w2(32'h3c3e44b2),
	.w3(32'h3ba147ac),
	.w4(32'h3b87fc6f),
	.w5(32'h3af08881),
	.w6(32'h3b7f92ca),
	.w7(32'h3c2ac1cd),
	.w8(32'h3c39538e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba719e14),
	.w1(32'h3a80d337),
	.w2(32'h3bae5106),
	.w3(32'h3bf723f1),
	.w4(32'hbb1c616d),
	.w5(32'h3baa1c2a),
	.w6(32'h3b17a7f7),
	.w7(32'h3b9641a7),
	.w8(32'h3c02246e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48114),
	.w1(32'h3c5122ea),
	.w2(32'h3b73cb5e),
	.w3(32'h3c3ee60b),
	.w4(32'h3c1c85f3),
	.w5(32'h3b0bbd19),
	.w6(32'h3bbee5b0),
	.w7(32'h3b9bdbc9),
	.w8(32'h3bb5f486),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30bf41),
	.w1(32'hba477f05),
	.w2(32'h3be414c4),
	.w3(32'hbc6d7274),
	.w4(32'hb916df27),
	.w5(32'h3d25c969),
	.w6(32'hbb80c0a3),
	.w7(32'h38a3658c),
	.w8(32'h3cb4d434),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d269530),
	.w1(32'h3ccea3b6),
	.w2(32'h3bd87e23),
	.w3(32'h3db92b19),
	.w4(32'h3d8c4635),
	.w5(32'h3c2c674f),
	.w6(32'h3d868a62),
	.w7(32'h3d3e39de),
	.w8(32'h3c24282c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91bf45),
	.w1(32'h3b48a0a1),
	.w2(32'h3b18e1ec),
	.w3(32'h3c1f2f81),
	.w4(32'h3baf6784),
	.w5(32'hbb746b96),
	.w6(32'h3c1ec935),
	.w7(32'h3c0c8d53),
	.w8(32'hb9d4afc2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb863f9f),
	.w1(32'hba80a4d7),
	.w2(32'h3b52ecbf),
	.w3(32'hbb38683f),
	.w4(32'h3b4bab23),
	.w5(32'h3b54bb18),
	.w6(32'hb9d0913e),
	.w7(32'h3a25d98e),
	.w8(32'h3a2cfc88),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99265f),
	.w1(32'hbadd3b36),
	.w2(32'h3b0b5889),
	.w3(32'hbb7ebd38),
	.w4(32'hbb460296),
	.w5(32'hb9b7afef),
	.w6(32'h3b9219ad),
	.w7(32'hbb3a8587),
	.w8(32'h3a5da27e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba407588),
	.w1(32'h3b0db229),
	.w2(32'h3c35887d),
	.w3(32'hbb024ce3),
	.w4(32'h3b59da05),
	.w5(32'h3bfe7c70),
	.w6(32'hbab0d2c2),
	.w7(32'h3b18aacb),
	.w8(32'h3b012233),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be64ef8),
	.w1(32'h3c04f6c4),
	.w2(32'h3b28b3df),
	.w3(32'h3b735eb7),
	.w4(32'h3bf9f2c0),
	.w5(32'h3b726d07),
	.w6(32'h3b0a11da),
	.w7(32'h3ae22fca),
	.w8(32'hba346f2e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebee2a),
	.w1(32'h3c2c5131),
	.w2(32'h38abc8f6),
	.w3(32'h3c4121cd),
	.w4(32'h3be8ec44),
	.w5(32'h3a1151ec),
	.w6(32'h3b220555),
	.w7(32'hbb1d05d1),
	.w8(32'hbb47daa9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb024517),
	.w1(32'hbb8d8b50),
	.w2(32'h398f5759),
	.w3(32'hbb9ecd95),
	.w4(32'h3a7c2cf9),
	.w5(32'hbb5644f0),
	.w6(32'h3ba0b88a),
	.w7(32'hb9e9d3df),
	.w8(32'hbb72bd0b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84f06),
	.w1(32'h3b3d451b),
	.w2(32'hbc4e2e09),
	.w3(32'h3c240bd8),
	.w4(32'h3c20ac45),
	.w5(32'hbcb41d72),
	.w6(32'h3b66cdc2),
	.w7(32'h3bf42fff),
	.w8(32'hbc497383),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14dcf5),
	.w1(32'h3a21b7cb),
	.w2(32'h3be2d808),
	.w3(32'hbc212f79),
	.w4(32'h3a2c1ea0),
	.w5(32'h3bf69401),
	.w6(32'hbbb70fc1),
	.w7(32'h3bc483f9),
	.w8(32'h3b2dc782),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0488),
	.w1(32'h3c4e9b0a),
	.w2(32'hbb54f222),
	.w3(32'h3bad7963),
	.w4(32'h3c5a4761),
	.w5(32'hbc05d497),
	.w6(32'h3b307354),
	.w7(32'h3c1e2765),
	.w8(32'h38f5b525),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98375a),
	.w1(32'h3ba8e4d1),
	.w2(32'h3a3b2b04),
	.w3(32'hbbef6a09),
	.w4(32'hbb5db1c0),
	.w5(32'hbb9634e2),
	.w6(32'h39c0bd81),
	.w7(32'h3c52b239),
	.w8(32'h3bc2949d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d6b7),
	.w1(32'hbae4767c),
	.w2(32'h3b21563f),
	.w3(32'h3a0fef9f),
	.w4(32'hbbad7661),
	.w5(32'h3b7f5ca2),
	.w6(32'h3ab3f176),
	.w7(32'h3b8147ca),
	.w8(32'hbad4fa92),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa2958),
	.w1(32'h3b9a6702),
	.w2(32'h3ae8b31d),
	.w3(32'h3bd2c01a),
	.w4(32'h3bd7416e),
	.w5(32'h3b4a6548),
	.w6(32'h3c3d3782),
	.w7(32'hb8c86659),
	.w8(32'hb97c2f1c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce8370),
	.w1(32'h3b00338f),
	.w2(32'hba9230f9),
	.w3(32'h3baf31f8),
	.w4(32'h3b9cc7ff),
	.w5(32'h3ca480fc),
	.w6(32'h3b816ef0),
	.w7(32'h3b9d19b5),
	.w8(32'h399a5e89),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50d975),
	.w1(32'hbabc4bdc),
	.w2(32'hbaaa2b3d),
	.w3(32'h3cebf812),
	.w4(32'h3cb6e5d2),
	.w5(32'hbb99afc8),
	.w6(32'h3b4b1043),
	.w7(32'hba8c6d71),
	.w8(32'h3afad2a7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a962ef1),
	.w1(32'h3afa0ab1),
	.w2(32'hbb6deba3),
	.w3(32'hba1174c3),
	.w4(32'hbb87f281),
	.w5(32'hbbba3faf),
	.w6(32'hbab48f83),
	.w7(32'hba9104dd),
	.w8(32'hbc0b774a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b222414),
	.w1(32'h3ba1b372),
	.w2(32'h3c505839),
	.w3(32'h3ae26f16),
	.w4(32'h3bdce753),
	.w5(32'h3c2168aa),
	.w6(32'hbb30b846),
	.w7(32'h3b0e3122),
	.w8(32'h3c3b8657),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205e5b),
	.w1(32'h3bf939f3),
	.w2(32'h3b214b70),
	.w3(32'h3abd6ae8),
	.w4(32'h3b5bbed5),
	.w5(32'h3ad2d77a),
	.w6(32'h3bdc80b9),
	.w7(32'h3bbf538c),
	.w8(32'h3b118dbd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90458e9),
	.w1(32'h3989399e),
	.w2(32'h3bcf3ff0),
	.w3(32'h3a95224d),
	.w4(32'h3915962b),
	.w5(32'h3bc2c640),
	.w6(32'h3b8b319b),
	.w7(32'h3a750172),
	.w8(32'h3bb55350),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c422561),
	.w1(32'h3c069beb),
	.w2(32'hbba18cde),
	.w3(32'h3c34b200),
	.w4(32'h3c22affe),
	.w5(32'hbbdd55f7),
	.w6(32'h3c06ed80),
	.w7(32'h3c085be1),
	.w8(32'hbbed7da3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2a66),
	.w1(32'hbaea803f),
	.w2(32'h3b3640be),
	.w3(32'h3b6c7698),
	.w4(32'hbba23184),
	.w5(32'h3b877233),
	.w6(32'h3b03287e),
	.w7(32'hbb9524c1),
	.w8(32'h3c0014c7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d7c2f),
	.w1(32'hbc08cca1),
	.w2(32'h3c1efc96),
	.w3(32'h3b247192),
	.w4(32'hbc5634c7),
	.w5(32'h3be83a88),
	.w6(32'h3bdcd4e4),
	.w7(32'hbc3753ca),
	.w8(32'h3b290839),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf13f2a),
	.w1(32'h3ba2ab9d),
	.w2(32'h3b97cc55),
	.w3(32'hbbf2d7dc),
	.w4(32'h3bbda7c1),
	.w5(32'hba1a6856),
	.w6(32'hbc03e6c3),
	.w7(32'h3bcaad90),
	.w8(32'h38826a8a),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9bc6),
	.w1(32'h3bbef22c),
	.w2(32'h3abf3634),
	.w3(32'h3c191e1f),
	.w4(32'h3ba6a424),
	.w5(32'h3b150b3c),
	.w6(32'h3bf6c23e),
	.w7(32'h3b1fffb4),
	.w8(32'hbba4e94c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c3d6b),
	.w1(32'hbb562179),
	.w2(32'hbc2d4863),
	.w3(32'hb8402229),
	.w4(32'h3a1e0bc8),
	.w5(32'h3c2517b8),
	.w6(32'hbbae6f1a),
	.w7(32'hbb0dee6f),
	.w8(32'hbb8a20ec),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af189),
	.w1(32'h3aa98366),
	.w2(32'h3ba29606),
	.w3(32'h3d22b3de),
	.w4(32'h3ce15dc3),
	.w5(32'h3baa7018),
	.w6(32'h3c9304a4),
	.w7(32'h3c1b83f2),
	.w8(32'h3b4c75f2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad0b9),
	.w1(32'h3a3c1f27),
	.w2(32'h3b884a51),
	.w3(32'h3c0e07ac),
	.w4(32'h3af97667),
	.w5(32'h39bc41ed),
	.w6(32'h3b8e5f87),
	.w7(32'h3a02e4f8),
	.w8(32'hbb6246fc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc5de5),
	.w1(32'hbb16ef88),
	.w2(32'hbba14a4f),
	.w3(32'h3c03f643),
	.w4(32'h3a445726),
	.w5(32'h3b93f35d),
	.w6(32'h3af80431),
	.w7(32'h3ba5c045),
	.w8(32'hbaffe558),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d2b58),
	.w1(32'h3b86af93),
	.w2(32'h3a2ccc1f),
	.w3(32'h3bd6c1c7),
	.w4(32'h3aab44e3),
	.w5(32'hbafde822),
	.w6(32'h3a36cd6e),
	.w7(32'h3c085fa6),
	.w8(32'h3b9e50d4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b911fc8),
	.w1(32'hbb48552d),
	.w2(32'h3bcd6164),
	.w3(32'h3be8cd83),
	.w4(32'h3b272358),
	.w5(32'hbb8e3dc5),
	.w6(32'h3beafb6c),
	.w7(32'h3b8965cd),
	.w8(32'h3b5a97fe),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf33ec5),
	.w1(32'h3b908fe5),
	.w2(32'h3c4e246e),
	.w3(32'hbb03c485),
	.w4(32'hbb939e2e),
	.w5(32'h3c3f1ab6),
	.w6(32'h3be06735),
	.w7(32'h3abca346),
	.w8(32'h3c2860f4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c50c6),
	.w1(32'hbb050d74),
	.w2(32'h3b072f3f),
	.w3(32'h3bf57579),
	.w4(32'hbbe2e3bb),
	.w5(32'hbc7168a6),
	.w6(32'h3c220424),
	.w7(32'hbb49a8ad),
	.w8(32'hbbca703c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a34d9),
	.w1(32'hbbccb9d9),
	.w2(32'h3ace9fdd),
	.w3(32'hbd25821a),
	.w4(32'hbce09979),
	.w5(32'h3b54d234),
	.w6(32'hbcd5975c),
	.w7(32'hbc811cc8),
	.w8(32'h392a849d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba094e6),
	.w1(32'h3c063ada),
	.w2(32'h3bc12c98),
	.w3(32'h3b20ab19),
	.w4(32'h3b6dbea0),
	.w5(32'h3c20169d),
	.w6(32'h3c04c78d),
	.w7(32'h3c0441c4),
	.w8(32'h3be21e4f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7dd1c),
	.w1(32'h3c5aa22e),
	.w2(32'h39e350bf),
	.w3(32'h3c8bd9cc),
	.w4(32'h3bedb365),
	.w5(32'h3b59dcc9),
	.w6(32'h3c71e411),
	.w7(32'h3b964923),
	.w8(32'hba2dd5a2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb69db),
	.w1(32'h3bbbcf33),
	.w2(32'h3ba32bc5),
	.w3(32'h3a55fb06),
	.w4(32'h39b68367),
	.w5(32'hba8ab32c),
	.w6(32'hbb84bd06),
	.w7(32'h3b669101),
	.w8(32'hb9366937),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38fe43),
	.w1(32'hb9ef59bd),
	.w2(32'h39d9d4bf),
	.w3(32'hb9fcaef8),
	.w4(32'h3b58648d),
	.w5(32'hbb3437bb),
	.w6(32'h3b9095eb),
	.w7(32'h3b50c45f),
	.w8(32'hbb89df17),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcc277),
	.w1(32'hb927acdb),
	.w2(32'hbbc21919),
	.w3(32'h3c3fb9aa),
	.w4(32'h3ba5e654),
	.w5(32'hbc1d7f9f),
	.w6(32'h3c889442),
	.w7(32'h39d6704c),
	.w8(32'hbbfa1159),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e684),
	.w1(32'hbc2e2f52),
	.w2(32'hb9858bf0),
	.w3(32'hbc2b19b5),
	.w4(32'hbc440cde),
	.w5(32'hbad8d51a),
	.w6(32'hbc240bde),
	.w7(32'hbc28b038),
	.w8(32'hbb47449a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a560fce),
	.w1(32'hbb26aefb),
	.w2(32'h3a89a428),
	.w3(32'h38f3d68c),
	.w4(32'h3c093f86),
	.w5(32'hbad4bd6c),
	.w6(32'h395ed9a8),
	.w7(32'hba90e7ab),
	.w8(32'hbb8fd390),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc048b08),
	.w1(32'h3c1bfa42),
	.w2(32'h3b6f087a),
	.w3(32'hbba75f1e),
	.w4(32'h3b22d2f2),
	.w5(32'h3b28e5fb),
	.w6(32'hbb837232),
	.w7(32'h3bc4553b),
	.w8(32'hbc06f6f0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52a882),
	.w1(32'h3c8f85c2),
	.w2(32'hbc7be303),
	.w3(32'h3c63f9ad),
	.w4(32'h3cc42a5d),
	.w5(32'hbc2e1834),
	.w6(32'h3b231c67),
	.w7(32'h3c4dce57),
	.w8(32'hbc282ecc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc300b67),
	.w1(32'hbb9e0fee),
	.w2(32'hba959727),
	.w3(32'hbb96b2da),
	.w4(32'hbba53357),
	.w5(32'hbaee9c4d),
	.w6(32'hbc4b5386),
	.w7(32'hbc220e73),
	.w8(32'hbb9ba829),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baab3b4),
	.w1(32'hbb82690d),
	.w2(32'hbc93189a),
	.w3(32'h3b816951),
	.w4(32'hbc07a514),
	.w5(32'hbcb2c6fe),
	.w6(32'h3b8ade67),
	.w7(32'hbbc42a9b),
	.w8(32'hbcb61cfe),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d5df5),
	.w1(32'hbc4d9245),
	.w2(32'h3b5c1a03),
	.w3(32'hbc14e9a7),
	.w4(32'hbc8ea7c2),
	.w5(32'h3a32aa7d),
	.w6(32'hbbe404a4),
	.w7(32'hbc6d13e2),
	.w8(32'hbb590470),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8227d),
	.w1(32'h3b64d7a3),
	.w2(32'h3a842212),
	.w3(32'h3c28e30b),
	.w4(32'h3bda653a),
	.w5(32'h3ba54f8b),
	.w6(32'h3ba2f3e0),
	.w7(32'h3b30780a),
	.w8(32'hbb2710fe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66df5a),
	.w1(32'h3b75c643),
	.w2(32'h3bc4bc10),
	.w3(32'h3c1e71a4),
	.w4(32'h3b9f1ccf),
	.w5(32'h3c07ad9e),
	.w6(32'h3a30721f),
	.w7(32'h3a7eef99),
	.w8(32'h3bf52716),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b937569),
	.w1(32'h3bbca7e0),
	.w2(32'hbb331ba0),
	.w3(32'h3c46dca0),
	.w4(32'h3c3fccdb),
	.w5(32'h3b4cfa26),
	.w6(32'h3c10edc4),
	.w7(32'h3c14c8e5),
	.w8(32'h3b8981aa),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4baf9),
	.w1(32'h3ab8b26b),
	.w2(32'h3c31e4ac),
	.w3(32'h39b1af28),
	.w4(32'h3bbf47b4),
	.w5(32'h3c157b76),
	.w6(32'h3b065211),
	.w7(32'h391986ce),
	.w8(32'h3b2a27bf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14ca1e),
	.w1(32'h3aec4462),
	.w2(32'h363cf0a0),
	.w3(32'h3c4967a9),
	.w4(32'h3bf85ac6),
	.w5(32'h3bdd808b),
	.w6(32'h3c128c45),
	.w7(32'h3bddf5db),
	.w8(32'h3c065304),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332509),
	.w1(32'h3b9f5058),
	.w2(32'hba539705),
	.w3(32'h3bf53ce6),
	.w4(32'h3c525bff),
	.w5(32'h3a376f22),
	.w6(32'h3c0e4cdf),
	.w7(32'h3c6ce1e4),
	.w8(32'h3b18cbd2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b6cbd),
	.w1(32'h3b0993e0),
	.w2(32'h3b60e98c),
	.w3(32'hba006f49),
	.w4(32'h3b1468e3),
	.w5(32'h3ae36e96),
	.w6(32'hbb7bf1f8),
	.w7(32'h3c1a7233),
	.w8(32'h3bbb6e73),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b701e8c),
	.w1(32'h3a151764),
	.w2(32'h3978709c),
	.w3(32'h3b314f92),
	.w4(32'hba08fc42),
	.w5(32'h3aecb2e2),
	.w6(32'h3ba14dba),
	.w7(32'h3be89cc0),
	.w8(32'h3a354d86),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f118),
	.w1(32'h3adf2092),
	.w2(32'h3c847f7a),
	.w3(32'h3bb34b06),
	.w4(32'h3b3a5b1d),
	.w5(32'h3c24c391),
	.w6(32'h3b4c7366),
	.w7(32'h3b50202b),
	.w8(32'h3bfe1037),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72fcb6),
	.w1(32'h3ad2b554),
	.w2(32'h3c044585),
	.w3(32'h3a9cdaf6),
	.w4(32'hb9d05d1a),
	.w5(32'h3b60c01b),
	.w6(32'hb4b0b614),
	.w7(32'h3aa3c7de),
	.w8(32'h3bf78d3f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d3644),
	.w1(32'h3afbfffa),
	.w2(32'h3c2a6133),
	.w3(32'hb8171124),
	.w4(32'h3b35682e),
	.w5(32'h3bd1924e),
	.w6(32'hba8f5ceb),
	.w7(32'h3bd24b56),
	.w8(32'h3bcfaf0b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b924195),
	.w1(32'h3c03164e),
	.w2(32'h3c374c1b),
	.w3(32'h3ab8b618),
	.w4(32'h3baf1633),
	.w5(32'h3c284968),
	.w6(32'hbb01c15d),
	.w7(32'h3c124950),
	.w8(32'h3c3f5981),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29346d),
	.w1(32'h3c1b858d),
	.w2(32'h3c0e3605),
	.w3(32'h3c49c588),
	.w4(32'h3c6a9242),
	.w5(32'h3c14715f),
	.w6(32'h3c4d526b),
	.w7(32'h3c73958d),
	.w8(32'h3c5a3eef),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9211d),
	.w1(32'h3b3747eb),
	.w2(32'h3b8a597b),
	.w3(32'h3c1cbd26),
	.w4(32'h3c0f4ef1),
	.w5(32'h3b6e6723),
	.w6(32'h3c52e940),
	.w7(32'h3c2d594a),
	.w8(32'h3b923b18),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08ed64),
	.w1(32'h3bc8791f),
	.w2(32'h3a45caaa),
	.w3(32'h3af64c44),
	.w4(32'h3c310295),
	.w5(32'h3a9a162e),
	.w6(32'hbb92ca0f),
	.w7(32'h3bb244ee),
	.w8(32'h3b9d482f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835e59),
	.w1(32'h3a0d58fb),
	.w2(32'h39ddc121),
	.w3(32'h3c08c52e),
	.w4(32'h3b9ceecd),
	.w5(32'h3a90f2ab),
	.w6(32'h3bebb55e),
	.w7(32'h3b6e01d5),
	.w8(32'hbb0c33a4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38909b4c),
	.w1(32'hbb2f4fa3),
	.w2(32'hbbec7b2e),
	.w3(32'h3ac968b0),
	.w4(32'hbaac714d),
	.w5(32'hbbf8a65a),
	.w6(32'h3b22946f),
	.w7(32'h39930e35),
	.w8(32'hbc127841),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4922d3),
	.w1(32'hba742926),
	.w2(32'h3c80fab7),
	.w3(32'h3a95dc92),
	.w4(32'h3c0734dd),
	.w5(32'h3c3ec11a),
	.w6(32'h3b225fa0),
	.w7(32'h3ad565a1),
	.w8(32'h3c100828),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd6fb5),
	.w1(32'h3bf7f052),
	.w2(32'h3bc3b628),
	.w3(32'h3b75e255),
	.w4(32'h3b86e920),
	.w5(32'h3bae9d3e),
	.w6(32'hbaeb0559),
	.w7(32'h3b4fbe9a),
	.w8(32'h3c038770),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf78aaf),
	.w1(32'h3c1e960f),
	.w2(32'h3bcc4bcf),
	.w3(32'h3c61d546),
	.w4(32'h3c353671),
	.w5(32'h3bace25b),
	.w6(32'h3bd783c8),
	.w7(32'h3c1b5520),
	.w8(32'h3bfd99c6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c43d8),
	.w1(32'h3bdbb163),
	.w2(32'hbbd83d75),
	.w3(32'h3ba25bcb),
	.w4(32'h3a7cb996),
	.w5(32'hbb8fb055),
	.w6(32'h3bc9e93b),
	.w7(32'h3c13c7c6),
	.w8(32'h3ad13799),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b3db0),
	.w1(32'hbbe05a44),
	.w2(32'hbc074ed6),
	.w3(32'hbbf24b27),
	.w4(32'hbba39587),
	.w5(32'hbbf1b1e5),
	.w6(32'h3b805615),
	.w7(32'h3b941290),
	.w8(32'hbc862e18),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b254c72),
	.w1(32'h3b0d7a36),
	.w2(32'hbba73fed),
	.w3(32'h3b6d1d6c),
	.w4(32'h3ae2cdb6),
	.w5(32'h3bfa4a92),
	.w6(32'hbc4e3482),
	.w7(32'hbc16b56e),
	.w8(32'hbb953198),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcce79e),
	.w1(32'hbbe3caa1),
	.w2(32'h3b8a0a09),
	.w3(32'h3bf929dc),
	.w4(32'h3c171ead),
	.w5(32'h3bac0432),
	.w6(32'hba69e6de),
	.w7(32'hba032f4d),
	.w8(32'h3ad9a530),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3971),
	.w1(32'h3ba359b5),
	.w2(32'h3c119c68),
	.w3(32'h3bfb7760),
	.w4(32'h3b558cdb),
	.w5(32'h3ba8b69e),
	.w6(32'h3bea873f),
	.w7(32'h3ba68414),
	.w8(32'h3a9716cf),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105656),
	.w1(32'hbb35792b),
	.w2(32'h3b1fc7b7),
	.w3(32'hb8cfced9),
	.w4(32'h3aaa6c1a),
	.w5(32'hbb4c4c5d),
	.w6(32'h3b508452),
	.w7(32'h3b6fd057),
	.w8(32'h3bcf08c9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb260bd),
	.w1(32'h3bb6a946),
	.w2(32'hbb2248f6),
	.w3(32'h3bfe0fcc),
	.w4(32'h3b1e1172),
	.w5(32'hbb17fa95),
	.w6(32'h3c4dafa4),
	.w7(32'h3b3537ed),
	.w8(32'hbb05f7b0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba16974),
	.w1(32'hba8b32bf),
	.w2(32'hbc2dd60e),
	.w3(32'hbb219024),
	.w4(32'hba18c528),
	.w5(32'hbcb90d4d),
	.w6(32'hbb1284d0),
	.w7(32'h398ba854),
	.w8(32'hbc3ef54e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca47b10),
	.w1(32'hbc454c7e),
	.w2(32'hbaeca2db),
	.w3(32'hbd13e00a),
	.w4(32'hbcd80625),
	.w5(32'h3b068330),
	.w6(32'hbccfe0bf),
	.w7(32'hbc74fe97),
	.w8(32'hbb4edfb1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b003f),
	.w1(32'h3bdd053b),
	.w2(32'hbbc8d0a2),
	.w3(32'h3bcf2ce7),
	.w4(32'h3c066b7b),
	.w5(32'hbbda27df),
	.w6(32'h3b17c6b6),
	.w7(32'h3bf45d90),
	.w8(32'hbbb11740),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12b26),
	.w1(32'hba934613),
	.w2(32'h3c0a5e63),
	.w3(32'h3a001474),
	.w4(32'h3a8d02cb),
	.w5(32'h3c4b61d5),
	.w6(32'h3b71e752),
	.w7(32'h3ba872ee),
	.w8(32'h3bd7d754),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f86d2),
	.w1(32'h3c1b543e),
	.w2(32'h3c311d9f),
	.w3(32'h3c9b947c),
	.w4(32'h3c49a4be),
	.w5(32'h3b48c41a),
	.w6(32'h3ca3e4a4),
	.w7(32'h3c38e513),
	.w8(32'h3bed23d3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54becd),
	.w1(32'h3b872fc3),
	.w2(32'h3b2a040f),
	.w3(32'hbb8a6994),
	.w4(32'h3bb013e2),
	.w5(32'hbb82e8a0),
	.w6(32'hba8ce726),
	.w7(32'h3be50b35),
	.w8(32'hbbd3da13),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d0a73),
	.w1(32'h3b6467d2),
	.w2(32'hbc0334f9),
	.w3(32'h3adc5dd1),
	.w4(32'h3a4e4576),
	.w5(32'hbbe124ad),
	.w6(32'hbb01d02f),
	.w7(32'hb98856a4),
	.w8(32'hbb9960d3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule