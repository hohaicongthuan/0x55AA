module layer_10_featuremap_496(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34b97864),
	.w1(32'h350f1526),
	.w2(32'h3572978b),
	.w3(32'h34fc27e9),
	.w4(32'h355a692b),
	.w5(32'h3583e840),
	.w6(32'hb2927d68),
	.w7(32'h35779421),
	.w8(32'h358ba09b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978c5e4),
	.w1(32'hb8a9163f),
	.w2(32'hb834188c),
	.w3(32'hb950005f),
	.w4(32'hb900be1b),
	.w5(32'hb89e0bc7),
	.w6(32'hb98683a4),
	.w7(32'hb8699fa0),
	.w8(32'h37c8fff6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33675f43),
	.w1(32'h350ea0ac),
	.w2(32'h354f7648),
	.w3(32'h34abd2e7),
	.w4(32'h34ee6aa5),
	.w5(32'h35397cbc),
	.w6(32'hb3095bdd),
	.w7(32'h352e6a09),
	.w8(32'h35590006),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d8bd7),
	.w1(32'h393919aa),
	.w2(32'h38883cb6),
	.w3(32'h391e67d4),
	.w4(32'h39690e4a),
	.w5(32'h38d743d6),
	.w6(32'h394418fa),
	.w7(32'h3941180f),
	.w8(32'hb4dfda3b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354bfbfd),
	.w1(32'hb58f1c49),
	.w2(32'hb4e64411),
	.w3(32'h358dc238),
	.w4(32'hb408614f),
	.w5(32'h359019b5),
	.w6(32'h3653feab),
	.w7(32'h35db8daa),
	.w8(32'h359e5c79),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3392ce2d),
	.w1(32'hb4e7263e),
	.w2(32'h33d2dc8e),
	.w3(32'h35828ad8),
	.w4(32'h3359aa46),
	.w5(32'h35a8e68e),
	.w6(32'h3573a290),
	.w7(32'h350304d9),
	.w8(32'h3580d9e6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d67221),
	.w1(32'h38930b1f),
	.w2(32'h382f863f),
	.w3(32'h38ffb80c),
	.w4(32'h38b9e72a),
	.w5(32'h38b4249d),
	.w6(32'h3901d39c),
	.w7(32'h38c00152),
	.w8(32'h387993cd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ea396),
	.w1(32'h39bc6809),
	.w2(32'hb8889395),
	.w3(32'h3a50b0ec),
	.w4(32'h39d108e3),
	.w5(32'hb8ab1de7),
	.w6(32'h3a11fa3f),
	.w7(32'h391c3a41),
	.w8(32'hb940ebd8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3757fb9e),
	.w1(32'h37ac31ee),
	.w2(32'h381b3623),
	.w3(32'hb75976c3),
	.w4(32'hb67cb688),
	.w5(32'h376f5fba),
	.w6(32'hb802b47d),
	.w7(32'hb7bf790a),
	.w8(32'h374b20cc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971d0a2),
	.w1(32'hb7aa3d30),
	.w2(32'hb8fe6bb0),
	.w3(32'hb9d27d60),
	.w4(32'hb9626caa),
	.w5(32'hb9666885),
	.w6(32'hba017bce),
	.w7(32'hb9ac5e11),
	.w8(32'hb96af10d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6429bcd),
	.w1(32'h35bc45c4),
	.w2(32'h36202091),
	.w3(32'hb754bcf9),
	.w4(32'hb64d07a4),
	.w5(32'h36b8223f),
	.w6(32'hb670a9b7),
	.w7(32'hb5a794bf),
	.w8(32'h36dbc4b6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09744a),
	.w1(32'h39bc6238),
	.w2(32'h394cc7e1),
	.w3(32'h39f8cceb),
	.w4(32'h39c3575a),
	.w5(32'h39863453),
	.w6(32'h3a015775),
	.w7(32'h39d46180),
	.w8(32'h38aba8cc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8007c8c),
	.w1(32'h38920746),
	.w2(32'h37b3a1fd),
	.w3(32'hb6fc7571),
	.w4(32'h388274fa),
	.w5(32'hb8409cbf),
	.w6(32'hb8d8e9cf),
	.w7(32'hb7d98f68),
	.w8(32'hb8ec2397),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb736d134),
	.w1(32'h3445f7a1),
	.w2(32'h36ed3263),
	.w3(32'hb7d4b5f0),
	.w4(32'hb6fd7dab),
	.w5(32'hb5ac6712),
	.w6(32'hb6e28ff1),
	.w7(32'hb60986e0),
	.w8(32'hb6d19587),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939311e),
	.w1(32'hb9084037),
	.w2(32'hb8c4f035),
	.w3(32'hb88b2958),
	.w4(32'hb8e72ad0),
	.w5(32'hb8e68724),
	.w6(32'hb98321bd),
	.w7(32'hb929689e),
	.w8(32'hb89f3be6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d51ec),
	.w1(32'h38492ca8),
	.w2(32'hb91830fc),
	.w3(32'hb848131c),
	.w4(32'h38084fb4),
	.w5(32'hb9002498),
	.w6(32'hb8aa55db),
	.w7(32'hb803db13),
	.w8(32'hb9155bbd),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b79662),
	.w1(32'h3540fc55),
	.w2(32'h353c5c5a),
	.w3(32'hb61726a7),
	.w4(32'hb5d98857),
	.w5(32'h354000f0),
	.w6(32'h35f863b0),
	.w7(32'h35cddbb9),
	.w8(32'h362f4eb5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a932e86),
	.w1(32'h395958de),
	.w2(32'hb9a3697b),
	.w3(32'h3ad1f18d),
	.w4(32'h3a6907bd),
	.w5(32'h39edd4a0),
	.w6(32'h3ac0b5f4),
	.w7(32'h3a6a94e6),
	.w8(32'hb8f3c674),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebdfae),
	.w1(32'h396ea89b),
	.w2(32'h379e4f07),
	.w3(32'h3a100293),
	.w4(32'h39b162fc),
	.w5(32'h3915fc4b),
	.w6(32'h3a02fa3d),
	.w7(32'h39ced6bc),
	.w8(32'h3749090f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59dfd02),
	.w1(32'hb5a853bb),
	.w2(32'hb47ea8fd),
	.w3(32'h33ad90bc),
	.w4(32'hb51bb95b),
	.w5(32'hb571ada8),
	.w6(32'h331bae96),
	.w7(32'h342281cc),
	.w8(32'h3563bf08),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367974b1),
	.w1(32'h3548fc7e),
	.w2(32'h339e8d01),
	.w3(32'h360c7030),
	.w4(32'h360bc5fb),
	.w5(32'h35df5c9a),
	.w6(32'h36128c52),
	.w7(32'h3611f5c1),
	.w8(32'h3513af08),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881b622),
	.w1(32'h38980216),
	.w2(32'hb68b7f7b),
	.w3(32'h3816fa2b),
	.w4(32'h3860e26f),
	.w5(32'h377e144b),
	.w6(32'h36f7a98f),
	.w7(32'h38348381),
	.w8(32'h37db82ab),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5a8ff),
	.w1(32'h39e7b695),
	.w2(32'hb9225917),
	.w3(32'h3ac88e5f),
	.w4(32'h3a7a819e),
	.w5(32'h3924970d),
	.w6(32'h3ae3302a),
	.w7(32'h3a675a10),
	.w8(32'hba0a5715),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff5b45),
	.w1(32'h383f116b),
	.w2(32'hb8388423),
	.w3(32'hb9b3d451),
	.w4(32'hb8723b35),
	.w5(32'hb96ec472),
	.w6(32'hb9fb58c6),
	.w7(32'hb99e27d8),
	.w8(32'hb984f7c0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b762a9),
	.w1(32'hb8e663de),
	.w2(32'hb940e498),
	.w3(32'hb9f84144),
	.w4(32'hb95eada4),
	.w5(32'hb9a84a16),
	.w6(32'hba1b8a0f),
	.w7(32'hb9a597e7),
	.w8(32'hb96bb757),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357ce778),
	.w1(32'hb6a4d1bf),
	.w2(32'hb624c1ae),
	.w3(32'h34f1006a),
	.w4(32'hb738a84b),
	.w5(32'hb7963b4e),
	.w6(32'h3508951c),
	.w7(32'hb78c08cb),
	.w8(32'hb7ead200),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb645fe23),
	.w1(32'hb64beda9),
	.w2(32'h36225dfe),
	.w3(32'hb5a9ed64),
	.w4(32'hb601ee0a),
	.w5(32'h366f8461),
	.w6(32'hb3a8da7a),
	.w7(32'h359b6763),
	.w8(32'h36db4a08),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d3e807),
	.w1(32'h383275ac),
	.w2(32'hb6b01433),
	.w3(32'hb7ca3e9d),
	.w4(32'h37b47590),
	.w5(32'hb7856874),
	.w6(32'h368ae59b),
	.w7(32'h3709943a),
	.w8(32'h38406952),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e0b1b8),
	.w1(32'h37ef9fbd),
	.w2(32'h372ba968),
	.w3(32'h37896f98),
	.w4(32'h37e8d299),
	.w5(32'h36c31b8a),
	.w6(32'h3763f69e),
	.w7(32'h37f0b758),
	.w8(32'h373522c4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c22cf4),
	.w1(32'hb922e1b1),
	.w2(32'hb9374b99),
	.w3(32'hb9e15565),
	.w4(32'hb952f4b4),
	.w5(32'hb9786744),
	.w6(32'hba0b5469),
	.w7(32'hb997c347),
	.w8(32'hb909f391),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb464d25d),
	.w1(32'h33989967),
	.w2(32'h34a46ee3),
	.w3(32'hb48d3a3d),
	.w4(32'hb51adb5e),
	.w5(32'hb477c1a2),
	.w6(32'h3506c763),
	.w7(32'h35242d4b),
	.w8(32'h352a23d4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34eddf7c),
	.w1(32'hb511cf53),
	.w2(32'h34c725d9),
	.w3(32'hb4ae5dac),
	.w4(32'hb5563d7a),
	.w5(32'h3480e371),
	.w6(32'h3560d0d4),
	.w7(32'h34d79870),
	.w8(32'h3514b9d5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8956a40),
	.w1(32'h36e36499),
	.w2(32'hb7ccf4b9),
	.w3(32'hb8a0cc88),
	.w4(32'hb7859281),
	.w5(32'hb8645ba1),
	.w6(32'hb8e9ca56),
	.w7(32'hb86fc942),
	.w8(32'hb890eadf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9037c01),
	.w1(32'hb7d5e463),
	.w2(32'hb7ee0b78),
	.w3(32'hb903d91b),
	.w4(32'hb821a55c),
	.w5(32'hb819d08b),
	.w6(32'hb91aa778),
	.w7(32'hb815d864),
	.w8(32'h36fb21ae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c05b2f),
	.w1(32'h37060004),
	.w2(32'h36355fcb),
	.w3(32'h35c0c3ee),
	.w4(32'h3442296c),
	.w5(32'hb69e4424),
	.w6(32'h36bd2244),
	.w7(32'h36d2abdf),
	.w8(32'h36c4faf2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ba530),
	.w1(32'h3922086b),
	.w2(32'hb81f71d2),
	.w3(32'h39b7072b),
	.w4(32'h39be8dc3),
	.w5(32'h38a2a08f),
	.w6(32'h397c5ad4),
	.w7(32'h389b8f15),
	.w8(32'hb8bb3b2f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39deaebf),
	.w1(32'h39902158),
	.w2(32'hb8b1b636),
	.w3(32'h3a29b88e),
	.w4(32'h39c2b52c),
	.w5(32'h3966542e),
	.w6(32'h3a005946),
	.w7(32'h3a037d5e),
	.w8(32'h38934403),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bccc8),
	.w1(32'hb9140866),
	.w2(32'hb974dc63),
	.w3(32'hb9e014ce),
	.w4(32'hb8abce19),
	.w5(32'hb9262f93),
	.w6(32'hba121904),
	.w7(32'hb8121d0a),
	.w8(32'h38bdfe2a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a1496),
	.w1(32'hb7ac3e36),
	.w2(32'hb8d18561),
	.w3(32'hb9750bbe),
	.w4(32'hb818db70),
	.w5(32'hb8cd0eae),
	.w6(32'hb98485f8),
	.w7(32'hb79406e2),
	.w8(32'h38a108ee),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b38b15),
	.w1(32'hb7b027c1),
	.w2(32'hb7421e81),
	.w3(32'hb8af46d0),
	.w4(32'hb78903db),
	.w5(32'hb7aab446),
	.w6(32'hb8c28c35),
	.w7(32'hb81bdfa9),
	.w8(32'h37153a4e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e43093),
	.w1(32'h34921d96),
	.w2(32'h360f7042),
	.w3(32'h35e1e046),
	.w4(32'hb3de6a08),
	.w5(32'h361852f4),
	.w6(32'h36214442),
	.w7(32'h348c79ab),
	.w8(32'h362512e7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a117fd),
	.w1(32'hb671bd5b),
	.w2(32'h36219ff5),
	.w3(32'hb6a2264d),
	.w4(32'hb6870479),
	.w5(32'h35f7e783),
	.w6(32'hb6a8037a),
	.w7(32'hb4e46710),
	.w8(32'h372a3969),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825d116),
	.w1(32'h37c4eb37),
	.w2(32'h3717bddc),
	.w3(32'h3808ae85),
	.w4(32'h373d13d0),
	.w5(32'hb7273027),
	.w6(32'h37f7cb78),
	.w7(32'h3754f44e),
	.w8(32'hb6893b26),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7699c77),
	.w1(32'h3852c4a4),
	.w2(32'hb8bef4ee),
	.w3(32'hb79dd5fb),
	.w4(32'h3757ef65),
	.w5(32'hb8d74fe5),
	.w6(32'hb8d72a1e),
	.w7(32'hb8d0edee),
	.w8(32'hb973bf4c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b50ec),
	.w1(32'hb879e414),
	.w2(32'hb8d9a0e9),
	.w3(32'hb9b24efd),
	.w4(32'hb936e1ba),
	.w5(32'hb932fce0),
	.w6(32'hb9dff0cd),
	.w7(32'hb96bd1ab),
	.w8(32'hb906d15c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b0bb6),
	.w1(32'h38a66cfa),
	.w2(32'hb8eedb5c),
	.w3(32'hb9ca08c0),
	.w4(32'hb8a29139),
	.w5(32'hb95c2820),
	.w6(32'hba02a852),
	.w7(32'hb9995196),
	.w8(32'hb99c9190),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ce469),
	.w1(32'h39677a54),
	.w2(32'hb90436a7),
	.w3(32'h38fae1d3),
	.w4(32'h395480b5),
	.w5(32'hb89ecc5d),
	.w6(32'h38c88d29),
	.w7(32'h38a9384e),
	.w8(32'hb97c1371),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e275),
	.w1(32'h3a2c99b7),
	.w2(32'hb9224398),
	.w3(32'h3ac0e995),
	.w4(32'h3a74bff7),
	.w5(32'h39934015),
	.w6(32'h3ac2602b),
	.w7(32'h3a9bb485),
	.w8(32'hb8e09841),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59ddb20),
	.w1(32'hb5b3c1d2),
	.w2(32'hb499ec0b),
	.w3(32'hb47637f6),
	.w4(32'hb530d9a0),
	.w5(32'h33bc0f41),
	.w6(32'hb50ee5ce),
	.w7(32'hb472219b),
	.w8(32'h353db4c3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37162af4),
	.w1(32'h3568387a),
	.w2(32'h372f3ce8),
	.w3(32'hb7627fc4),
	.w4(32'hb7965570),
	.w5(32'h371d25ca),
	.w6(32'hb6db5316),
	.w7(32'hb73757e7),
	.w8(32'h370c8a49),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb632e39b),
	.w1(32'hb5da810b),
	.w2(32'h3678b003),
	.w3(32'hb677d3ad),
	.w4(32'hb6a3971a),
	.w5(32'hb685916d),
	.w6(32'hb6d711d3),
	.w7(32'hb6d11fad),
	.w8(32'hb6b708a5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e4dbb8),
	.w1(32'hb70a3e0e),
	.w2(32'hb8a8cf97),
	.w3(32'hb83aab10),
	.w4(32'h36827a6d),
	.w5(32'hb899279a),
	.w6(32'hb8840c95),
	.w7(32'hb84cc2f8),
	.w8(32'hb9130773),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948329b),
	.w1(32'h38dc9f24),
	.w2(32'hb710a167),
	.w3(32'h391a1638),
	.w4(32'h38d4b877),
	.w5(32'hb5fa1db4),
	.w6(32'h39291a2b),
	.w7(32'h38d955e3),
	.w8(32'hb8292e57),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80bf15),
	.w1(32'h39bfcb8e),
	.w2(32'hb968ab96),
	.w3(32'h3a8568c0),
	.w4(32'h3a3ac180),
	.w5(32'h39992dce),
	.w6(32'h3a85d138),
	.w7(32'h3a499f87),
	.w8(32'hb91c5c76),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dfc17),
	.w1(32'h3811c608),
	.w2(32'hb810ed74),
	.w3(32'h38f15f5e),
	.w4(32'h38c3def6),
	.w5(32'h35af0d1a),
	.w6(32'h388ca65e),
	.w7(32'h378adf91),
	.w8(32'hb816d851),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb637e942),
	.w1(32'hb54cf520),
	.w2(32'hb54eb47c),
	.w3(32'hb608b026),
	.w4(32'hb635b43b),
	.w5(32'hb62c10e4),
	.w6(32'hb57e091f),
	.w7(32'hb640440c),
	.w8(32'hb6afd174),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5368e56),
	.w1(32'hb4ed5015),
	.w2(32'h350be0f3),
	.w3(32'hb50f89f8),
	.w4(32'hb52f38c1),
	.w5(32'h34c45a34),
	.w6(32'h30f12d56),
	.w7(32'hb47852e8),
	.w8(32'h357423df),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37170222),
	.w1(32'h3723bcca),
	.w2(32'h344ab121),
	.w3(32'h3653e72b),
	.w4(32'h36a5b510),
	.w5(32'hb50e1d56),
	.w6(32'h36993cdf),
	.w7(32'h36c839b1),
	.w8(32'hb5027781),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37543e7c),
	.w1(32'h373f14a0),
	.w2(32'h34ac074e),
	.w3(32'h373b1766),
	.w4(32'h37697807),
	.w5(32'h35e60b54),
	.w6(32'h36fa6f77),
	.w7(32'h3751d58f),
	.w8(32'h36b8f770),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f58cb0),
	.w1(32'h35ec015b),
	.w2(32'hb67ee160),
	.w3(32'h36d72af5),
	.w4(32'h3586324f),
	.w5(32'hb69b4f0f),
	.w6(32'h366bd19c),
	.w7(32'hb516ad98),
	.w8(32'hb5c701fb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9fad8),
	.w1(32'h398420bf),
	.w2(32'h386fea05),
	.w3(32'h39dc3ed4),
	.w4(32'h39c2f274),
	.w5(32'h3960837e),
	.w6(32'h39dcdf55),
	.w7(32'h399e4a4b),
	.w8(32'hb8949d98),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980c50c),
	.w1(32'hb8b7a80c),
	.w2(32'hb907dc7d),
	.w3(32'h392bf70d),
	.w4(32'h383ebf81),
	.w5(32'hb9011f88),
	.w6(32'h394d148e),
	.w7(32'hb7d62121),
	.w8(32'hb968716f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3595667c),
	.w1(32'h351bfaa6),
	.w2(32'h35da42b2),
	.w3(32'hb4a63d9d),
	.w4(32'hb4f40a1f),
	.w5(32'h352beeb7),
	.w6(32'h32c76386),
	.w7(32'h3449c102),
	.w8(32'h3603b39b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb48acd5f),
	.w1(32'hb4b25f34),
	.w2(32'h356aae46),
	.w3(32'hb5075b21),
	.w4(32'hb5ab0acd),
	.w5(32'hb47dd31b),
	.w6(32'hb512f23c),
	.w7(32'hb55e028a),
	.w8(32'h355be5ba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f6a387),
	.w1(32'hb5b94a81),
	.w2(32'hb538e2f7),
	.w3(32'hb50ee2fd),
	.w4(32'hb5ad77cc),
	.w5(32'hb519b07b),
	.w6(32'h359beb68),
	.w7(32'hb59c1b6d),
	.w8(32'hb48211e4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h340906b2),
	.w1(32'h35937ee0),
	.w2(32'h35af4c5e),
	.w3(32'h345e6dff),
	.w4(32'h36064824),
	.w5(32'h362e290e),
	.w6(32'h35b3a4e2),
	.w7(32'h362b843b),
	.w8(32'h3671afd1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930a1fd),
	.w1(32'h38205b6e),
	.w2(32'hb8dc1569),
	.w3(32'h398edd37),
	.w4(32'h395158c6),
	.w5(32'h373a6902),
	.w6(32'h39915573),
	.w7(32'h3936273b),
	.w8(32'hb914dc02),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ca2fd3),
	.w1(32'h391f0a4c),
	.w2(32'hb926f0bc),
	.w3(32'hb935979b),
	.w4(32'h373ebd55),
	.w5(32'hb9760293),
	.w6(32'hb96e197b),
	.w7(32'hb9125186),
	.w8(32'hb96b133d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f3b6),
	.w1(32'h3914183a),
	.w2(32'hb973aae8),
	.w3(32'h39d53fd2),
	.w4(32'h39ea24d8),
	.w5(32'hb872474c),
	.w6(32'h396dd27e),
	.w7(32'hb8ee9c6f),
	.w8(32'hba210a1c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c972ab),
	.w1(32'h3b88deec),
	.w2(32'hbb5291f6),
	.w3(32'hba26587d),
	.w4(32'hbb495950),
	.w5(32'hbc3b02f2),
	.w6(32'hba41de6e),
	.w7(32'h3bca3eac),
	.w8(32'hbb851725),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27c10c),
	.w1(32'hbb721522),
	.w2(32'h3b1f60f0),
	.w3(32'h3b5ee09d),
	.w4(32'hb9f9fe42),
	.w5(32'hbbb5d7ac),
	.w6(32'h38dfccae),
	.w7(32'hbb0f6995),
	.w8(32'hbad3f969),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd4243),
	.w1(32'hbaf4124e),
	.w2(32'hbb0a2364),
	.w3(32'hbbb43949),
	.w4(32'hbbf7180f),
	.w5(32'h3ad3060d),
	.w6(32'hba8b3770),
	.w7(32'hbb85f824),
	.w8(32'hbaac0847),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe200a),
	.w1(32'hbbce1a58),
	.w2(32'hbc3a8a37),
	.w3(32'hbb6e59e2),
	.w4(32'hbb669573),
	.w5(32'hb9818622),
	.w6(32'h3a74cff2),
	.w7(32'hba88c91e),
	.w8(32'h3a1f6461),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3cdee),
	.w1(32'hbbd794ab),
	.w2(32'hbb7c1c92),
	.w3(32'h3b17926f),
	.w4(32'hbb211a08),
	.w5(32'h3bf11491),
	.w6(32'h3b8b96dd),
	.w7(32'h3a8616da),
	.w8(32'h3be32e39),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8baead),
	.w1(32'hbbf0ea43),
	.w2(32'hbc2a2eef),
	.w3(32'h3a5be80b),
	.w4(32'hbb1f72ee),
	.w5(32'h3ab584b0),
	.w6(32'hba7cc549),
	.w7(32'h3b330739),
	.w8(32'h3b79af92),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c19f),
	.w1(32'h3bf0865e),
	.w2(32'hbb02be00),
	.w3(32'hbc26e342),
	.w4(32'h3a82bd05),
	.w5(32'h3bdccc79),
	.w6(32'h3b24b4df),
	.w7(32'h39fc02df),
	.w8(32'h3897fc1b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a751),
	.w1(32'hbc102607),
	.w2(32'hbb4172f2),
	.w3(32'h3b0a2f25),
	.w4(32'hbbcbc6e3),
	.w5(32'hb8927c17),
	.w6(32'h3bc8d98b),
	.w7(32'h3b58c2e3),
	.w8(32'h3c1e2aa5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296843),
	.w1(32'hbc14b9ae),
	.w2(32'hbb9ecb88),
	.w3(32'h3bef039b),
	.w4(32'hbc5e0df4),
	.w5(32'h3b5b9032),
	.w6(32'h3b99c52f),
	.w7(32'hbc543609),
	.w8(32'h3b1daf77),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2539c),
	.w1(32'hbba3d8c0),
	.w2(32'h3b3e1113),
	.w3(32'hbb9c9ad6),
	.w4(32'h39ba196f),
	.w5(32'h3c102763),
	.w6(32'h3b308492),
	.w7(32'hb94ba1d9),
	.w8(32'h3a55b064),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7832dc),
	.w1(32'hbc34c1aa),
	.w2(32'hbc53c488),
	.w3(32'hbb24fa4b),
	.w4(32'hbc85b6e6),
	.w5(32'hbc6c2922),
	.w6(32'hbbdd8f4e),
	.w7(32'hbc0d1003),
	.w8(32'hbbe0ad86),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a6363),
	.w1(32'h3c4369a4),
	.w2(32'h3c40a8aa),
	.w3(32'hbc4a516b),
	.w4(32'hba8df100),
	.w5(32'h3b8b73a2),
	.w6(32'hbb285be0),
	.w7(32'hb9bba882),
	.w8(32'h3b87545d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e2d0e),
	.w1(32'h3b047716),
	.w2(32'h3b01f86e),
	.w3(32'h3a33a534),
	.w4(32'h3b8e7632),
	.w5(32'hba124c56),
	.w6(32'h3b2b2a74),
	.w7(32'h3a78ad7c),
	.w8(32'h3b44d158),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a59761e),
	.w1(32'hbb546f46),
	.w2(32'h3b8a5dc0),
	.w3(32'h39d1bd1e),
	.w4(32'h3b38c5d7),
	.w5(32'h3c1139ee),
	.w6(32'hbb8a6931),
	.w7(32'h3c154c7b),
	.w8(32'h3bf46a5a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99aa8e5),
	.w1(32'hbbf90573),
	.w2(32'hbac2aa45),
	.w3(32'hbb423b97),
	.w4(32'hbba64af4),
	.w5(32'h3ca99245),
	.w6(32'hb9125565),
	.w7(32'h3b66abbf),
	.w8(32'hba3a365c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fa391),
	.w1(32'hbb992eb0),
	.w2(32'hbaf37f7a),
	.w3(32'h39f0dfaf),
	.w4(32'hbbc881f2),
	.w5(32'hbaa3dca3),
	.w6(32'hbb061808),
	.w7(32'hbba11f75),
	.w8(32'h3b04f082),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1c00c),
	.w1(32'h39d616b2),
	.w2(32'h3cc7a44f),
	.w3(32'hbaebcdb3),
	.w4(32'h3d178df1),
	.w5(32'h3c83c80d),
	.w6(32'h3a007dae),
	.w7(32'h3c8882b1),
	.w8(32'h3be52573),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35d55e),
	.w1(32'hbb8ca318),
	.w2(32'hb9e68039),
	.w3(32'h3c17cbfb),
	.w4(32'hbad826a9),
	.w5(32'hbc0c5f21),
	.w6(32'h3b6fde34),
	.w7(32'hbb4182f5),
	.w8(32'hbb421cb3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a34ff),
	.w1(32'hb9aed1a9),
	.w2(32'h3c2933bc),
	.w3(32'hbb21c9c4),
	.w4(32'h3c0f24b9),
	.w5(32'h3c226010),
	.w6(32'hbbf3a189),
	.w7(32'h3bf00b94),
	.w8(32'hba3835ac),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25b41),
	.w1(32'hbb709f86),
	.w2(32'hbbfba039),
	.w3(32'hbab9ddc5),
	.w4(32'hbb9c656b),
	.w5(32'h3b8a65a8),
	.w6(32'hbc025323),
	.w7(32'h3988f6a5),
	.w8(32'h3b63d73d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073402),
	.w1(32'h3b60a658),
	.w2(32'hbb26ac9f),
	.w3(32'hbb686ecc),
	.w4(32'h3bfdc9ba),
	.w5(32'hbbcb428d),
	.w6(32'hbbb4e967),
	.w7(32'h39bbc552),
	.w8(32'h3ac5e450),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b053994),
	.w1(32'hbb05d7cc),
	.w2(32'hba95e12f),
	.w3(32'hbb733e1d),
	.w4(32'hbb0dfa56),
	.w5(32'hbbbc74fd),
	.w6(32'hbb62d4a6),
	.w7(32'hbb86d52d),
	.w8(32'hbbfffee2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba217),
	.w1(32'hbb9b126f),
	.w2(32'h3c073ba5),
	.w3(32'h3c0389d1),
	.w4(32'h3cbf0f57),
	.w5(32'h3c1758ab),
	.w6(32'h3bd9c1f1),
	.w7(32'hbbf49a36),
	.w8(32'hbbe7170b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c172b75),
	.w1(32'h3b7be38a),
	.w2(32'h39bdffd4),
	.w3(32'h3b215d26),
	.w4(32'h3ad64973),
	.w5(32'hb9e33bb0),
	.w6(32'hbb1647ec),
	.w7(32'hb9c56564),
	.w8(32'hba902e57),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c383d9),
	.w1(32'h3b449e87),
	.w2(32'h3c234b5f),
	.w3(32'h3b6cd946),
	.w4(32'h3bbedc76),
	.w5(32'h3b79a888),
	.w6(32'hbab44922),
	.w7(32'h39941b2d),
	.w8(32'h3af270a1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf668da),
	.w1(32'hbbccdfab),
	.w2(32'hbc6f1708),
	.w3(32'h3b378510),
	.w4(32'hbbbc81e6),
	.w5(32'hbbe23dc8),
	.w6(32'h3a32a8a1),
	.w7(32'hbc5304d5),
	.w8(32'hbc25a371),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105226),
	.w1(32'hba233613),
	.w2(32'hbaa2a4c2),
	.w3(32'hbb19d9d0),
	.w4(32'hbc0569f7),
	.w5(32'hbaeace58),
	.w6(32'hb919c3d0),
	.w7(32'hb99a33bd),
	.w8(32'h3a8cc056),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6018),
	.w1(32'h39422250),
	.w2(32'h3c340248),
	.w3(32'h3c08ab34),
	.w4(32'h3bd1bcac),
	.w5(32'h3c6dad63),
	.w6(32'h395839f7),
	.w7(32'h3bfbbbfe),
	.w8(32'h3c566a98),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c02d),
	.w1(32'h3b5a4d6b),
	.w2(32'hb9ba84c6),
	.w3(32'h3bdb4e2c),
	.w4(32'h3bbec98a),
	.w5(32'h3ba7318d),
	.w6(32'hbbc19777),
	.w7(32'hbb6c3b91),
	.w8(32'h3be5ed34),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabed539),
	.w1(32'hbc28ab3c),
	.w2(32'hbbb993ec),
	.w3(32'h3bf05233),
	.w4(32'h3b001860),
	.w5(32'hbc46d3c9),
	.w6(32'h3c3f0b7e),
	.w7(32'hbb52903e),
	.w8(32'h3b6705b0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51c6d4),
	.w1(32'h3b8cfcfb),
	.w2(32'hbc0060e7),
	.w3(32'h3b077591),
	.w4(32'hbbcc3bb4),
	.w5(32'hbade4286),
	.w6(32'h3b356a17),
	.w7(32'hbb7f65fa),
	.w8(32'hbbb316cb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d0c4),
	.w1(32'hbbdb8dc6),
	.w2(32'h3a932ee3),
	.w3(32'hbc23e645),
	.w4(32'hbbe96d00),
	.w5(32'h3b1cdeff),
	.w6(32'h3b519d15),
	.w7(32'hbb884413),
	.w8(32'h3b08f515),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab838ce),
	.w1(32'hbb341be6),
	.w2(32'h3a8bb26d),
	.w3(32'hb9a0f80a),
	.w4(32'hbaf2ea8f),
	.w5(32'h3b12c0bb),
	.w6(32'hbb46c4a0),
	.w7(32'hbbda3407),
	.w8(32'hbbb17487),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c58f0),
	.w1(32'hbb303740),
	.w2(32'h3c182103),
	.w3(32'h3a38a5f3),
	.w4(32'hba369b0b),
	.w5(32'h3c574f36),
	.w6(32'hbb8bc1cf),
	.w7(32'hbb0037a0),
	.w8(32'h3c31dc9e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba77cc4),
	.w1(32'h3bcd7e78),
	.w2(32'h3b92f5b2),
	.w3(32'h3baad641),
	.w4(32'h3b0db3b9),
	.w5(32'h3b86effb),
	.w6(32'h3c3e2be7),
	.w7(32'h3b0bf606),
	.w8(32'hba081c14),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee5ebd),
	.w1(32'hbbbc6353),
	.w2(32'h3bca05d4),
	.w3(32'h3b9ecbe3),
	.w4(32'h3aba8100),
	.w5(32'h3c18ff5f),
	.w6(32'h3b4f5bba),
	.w7(32'h3a05f0d9),
	.w8(32'hbbe5d1de),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ad64c),
	.w1(32'hba2ba673),
	.w2(32'h3c0eb332),
	.w3(32'h3aac2624),
	.w4(32'h3b9d42c9),
	.w5(32'h3bd68c60),
	.w6(32'hbb70b472),
	.w7(32'h3b776574),
	.w8(32'h3b4c50a4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d072d),
	.w1(32'h3b26848f),
	.w2(32'h3b608d28),
	.w3(32'h3b011d74),
	.w4(32'h3b81f817),
	.w5(32'hbb3af807),
	.w6(32'hbb707bb3),
	.w7(32'h3b4e0e17),
	.w8(32'h3ba7a005),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070108),
	.w1(32'hbaa08b6b),
	.w2(32'h387e9f22),
	.w3(32'hbbb92bf6),
	.w4(32'h3a1cc543),
	.w5(32'hbade611e),
	.w6(32'hbb9ac831),
	.w7(32'hbbd744c7),
	.w8(32'hbab9aab4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223192),
	.w1(32'h3c4a307f),
	.w2(32'hbb94b26d),
	.w3(32'h3a60c177),
	.w4(32'h3b81887a),
	.w5(32'hb9a17013),
	.w6(32'h3a8ac71a),
	.w7(32'h3b926ade),
	.w8(32'h361be597),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd6ac),
	.w1(32'hbafda5bf),
	.w2(32'hbb797390),
	.w3(32'hbb7e2fd4),
	.w4(32'hbb990180),
	.w5(32'h38a2c84b),
	.w6(32'h3b15dba4),
	.w7(32'hbc35717f),
	.w8(32'hbc1d8dd0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd887f9),
	.w1(32'h3ca73c27),
	.w2(32'h3c8abe94),
	.w3(32'h3afa54ee),
	.w4(32'h3caa4ae5),
	.w5(32'h3b20073a),
	.w6(32'hbbcb9114),
	.w7(32'h3b8b9995),
	.w8(32'hb88db8e2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9baf80),
	.w1(32'h3bcc813e),
	.w2(32'h3b743619),
	.w3(32'h3c26654f),
	.w4(32'h3c564a42),
	.w5(32'h3b079a09),
	.w6(32'h3bbb4e70),
	.w7(32'h3c2d5528),
	.w8(32'h3c6f299a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7653b),
	.w1(32'hbb752938),
	.w2(32'h3b6bf3c5),
	.w3(32'h3c27d9ec),
	.w4(32'h3ba50934),
	.w5(32'h3c099db7),
	.w6(32'h3c275fec),
	.w7(32'h3b29e469),
	.w8(32'h3c1bc057),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb185de),
	.w1(32'h3c12ba60),
	.w2(32'hbba5d007),
	.w3(32'h3b342025),
	.w4(32'hbbc618cc),
	.w5(32'h3c702267),
	.w6(32'h3b1a7bc1),
	.w7(32'h3c043a5f),
	.w8(32'hbb3f4baa),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56fabb),
	.w1(32'hbc18d2d3),
	.w2(32'hb9fe6487),
	.w3(32'hbb5eadb4),
	.w4(32'hbc1d040a),
	.w5(32'h3b5aef3a),
	.w6(32'hbc19bb21),
	.w7(32'hbb99b445),
	.w8(32'h3b911e36),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c1212),
	.w1(32'h3afc0741),
	.w2(32'hbc0e5dcc),
	.w3(32'h3c3a04bd),
	.w4(32'hbbf3756c),
	.w5(32'hbbcd65f1),
	.w6(32'h39e3c921),
	.w7(32'hbc0f5cea),
	.w8(32'hb9feb9fc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06ecc8),
	.w1(32'h3aedbb0a),
	.w2(32'hb8f75886),
	.w3(32'h3a88e901),
	.w4(32'hbb060a81),
	.w5(32'h3bc93ede),
	.w6(32'h3b29db4e),
	.w7(32'h3ac26c3e),
	.w8(32'h3b4f82d2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8713f),
	.w1(32'hbb836589),
	.w2(32'hbafe288e),
	.w3(32'h3c6d05b7),
	.w4(32'h3a9bf9a3),
	.w5(32'h3b14d5ca),
	.w6(32'h3c0b1234),
	.w7(32'h3b545aec),
	.w8(32'h3bd157ea),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a365),
	.w1(32'hbb6fa30f),
	.w2(32'hbbae91f4),
	.w3(32'hbb3d2a2c),
	.w4(32'hba5c41ec),
	.w5(32'h3af88e71),
	.w6(32'h3b02ad5c),
	.w7(32'hbbe91fc3),
	.w8(32'hbbcfed68),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb508a13),
	.w1(32'h3babeaa4),
	.w2(32'h3acc3f88),
	.w3(32'h3ac2c604),
	.w4(32'hbbb352e7),
	.w5(32'hbb62271c),
	.w6(32'hbb56b44f),
	.w7(32'hbc164068),
	.w8(32'hbb93bc34),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3a0db),
	.w1(32'hbbd5512e),
	.w2(32'hbad42541),
	.w3(32'hbaaa543f),
	.w4(32'hbbfb05b3),
	.w5(32'h3a1dd2bb),
	.w6(32'h3bf8a078),
	.w7(32'hbbcfa071),
	.w8(32'h3a20c924),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9efd0),
	.w1(32'h3c3b45f1),
	.w2(32'h3b54ba46),
	.w3(32'h3b148f97),
	.w4(32'h3bec52e5),
	.w5(32'hbc863e0e),
	.w6(32'hb95f2a1f),
	.w7(32'h3bb9ccb1),
	.w8(32'hbba858f5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8994a2),
	.w1(32'h3adf2a67),
	.w2(32'h3c42e39c),
	.w3(32'hbabcbc54),
	.w4(32'h3bdca23b),
	.w5(32'h3c1447df),
	.w6(32'h3ba0ad11),
	.w7(32'h3b83e4c9),
	.w8(32'h3bb8ec2a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7efc80),
	.w1(32'h3aed1ba8),
	.w2(32'h3c41172e),
	.w3(32'h3b895b20),
	.w4(32'h3bb0e802),
	.w5(32'h3b57cf52),
	.w6(32'hb9dd6d26),
	.w7(32'h3b2af845),
	.w8(32'hba93b6c1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e4756),
	.w1(32'h3a79d6f2),
	.w2(32'hbaeda95f),
	.w3(32'hbb4a441c),
	.w4(32'hbbbaf927),
	.w5(32'h3b10ec7d),
	.w6(32'hbbfc4d7e),
	.w7(32'hbaa0d749),
	.w8(32'hbaa7008a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dbe42),
	.w1(32'hbbbb325b),
	.w2(32'hbb91398e),
	.w3(32'hbb96790b),
	.w4(32'hbb2f1b89),
	.w5(32'h3c037431),
	.w6(32'hbb0f6423),
	.w7(32'hbb55e15c),
	.w8(32'hbb98e0e3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9cee7),
	.w1(32'h3b234dfa),
	.w2(32'h3c6c8957),
	.w3(32'hbb6eba19),
	.w4(32'h3b4a4e87),
	.w5(32'h3c542c3a),
	.w6(32'hbbc55bea),
	.w7(32'h3acd89cf),
	.w8(32'h3b7a77c9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8812ecc),
	.w1(32'hbba4054e),
	.w2(32'h3c7068f2),
	.w3(32'h3c116eb0),
	.w4(32'h3baa23ae),
	.w5(32'h3c23b3c0),
	.w6(32'h3b70d04a),
	.w7(32'h3c6a50db),
	.w8(32'h3b7b4e42),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9688),
	.w1(32'hbb87c470),
	.w2(32'hbc0e9ff5),
	.w3(32'h3ba7278c),
	.w4(32'hbc1a4f2a),
	.w5(32'hbbbf8806),
	.w6(32'h39e1b8d6),
	.w7(32'hbbb8f0c0),
	.w8(32'hbb6a1d31),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89d553),
	.w1(32'hbc164d49),
	.w2(32'h3bb8b496),
	.w3(32'hbb2d3074),
	.w4(32'hbbcdfc0c),
	.w5(32'h3bfc0a7d),
	.w6(32'hba6c1e0c),
	.w7(32'hba99d6fb),
	.w8(32'h3b0325f3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab05193),
	.w1(32'h3b80aa31),
	.w2(32'hba92c4f6),
	.w3(32'h3b77ef7c),
	.w4(32'h3afc65d6),
	.w5(32'h3b8c1c7e),
	.w6(32'h3b465401),
	.w7(32'hbb0d4d94),
	.w8(32'hbaf8161e),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59da68),
	.w1(32'h3bf4ba30),
	.w2(32'hbb9e01e4),
	.w3(32'h3be40c0f),
	.w4(32'hbb2521d1),
	.w5(32'h3abeca51),
	.w6(32'hbb7888dd),
	.w7(32'h3c06e64b),
	.w8(32'h3a070614),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20c1f1),
	.w1(32'h3b0eada9),
	.w2(32'hba837ea8),
	.w3(32'h3ba84bfc),
	.w4(32'hba6fd92d),
	.w5(32'hbbd34848),
	.w6(32'h3be23af6),
	.w7(32'hbae404db),
	.w8(32'hbbf66de8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ea784),
	.w1(32'hb92ed647),
	.w2(32'hbb5b5ba5),
	.w3(32'hbb6b2ae9),
	.w4(32'h3a0409c1),
	.w5(32'h3c8f4549),
	.w6(32'hbb9d5365),
	.w7(32'h3bcd924e),
	.w8(32'h3c272b03),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dce03),
	.w1(32'h386da695),
	.w2(32'hbbc042ef),
	.w3(32'h3bb39593),
	.w4(32'hbac9f19b),
	.w5(32'h3b6377ce),
	.w6(32'hb9266b3f),
	.w7(32'h3afe3fab),
	.w8(32'h3ad02f69),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88d3a0),
	.w1(32'h3bf9b16d),
	.w2(32'h3ba22131),
	.w3(32'h3b5591d3),
	.w4(32'h3c25ba06),
	.w5(32'hbb98f721),
	.w6(32'h3b7f4e15),
	.w7(32'h3b2f8be7),
	.w8(32'h3be7a7f8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbca96),
	.w1(32'h3ae40881),
	.w2(32'h3b009cab),
	.w3(32'h3a07c0d4),
	.w4(32'h394e7a18),
	.w5(32'h3a8b3b21),
	.w6(32'hbb1565b6),
	.w7(32'h3aad471d),
	.w8(32'h3a40fdd2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce6f05),
	.w1(32'h3b0328be),
	.w2(32'hbb188724),
	.w3(32'h3c288579),
	.w4(32'hbb9dc4b4),
	.w5(32'hbc2cfa18),
	.w6(32'h3c0458b3),
	.w7(32'h3bc65606),
	.w8(32'hbb875beb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f09a1),
	.w1(32'hbbf29126),
	.w2(32'hbb17fc6b),
	.w3(32'hbbf453ae),
	.w4(32'hbbe785a3),
	.w5(32'hbae88d11),
	.w6(32'h39f5674a),
	.w7(32'hbb9d28e3),
	.w8(32'h3aa209e6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3eb6),
	.w1(32'hbb68de99),
	.w2(32'h3bae7901),
	.w3(32'hbb874039),
	.w4(32'hbaa7fa55),
	.w5(32'hbb6d836f),
	.w6(32'h3c1a0118),
	.w7(32'hbab4b5f8),
	.w8(32'h3b2fbc0a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56251),
	.w1(32'hbc419327),
	.w2(32'h3c9239db),
	.w3(32'hbbc0af51),
	.w4(32'hbba9565e),
	.w5(32'h3c77cc0a),
	.w6(32'hbc15a298),
	.w7(32'h3b631e2e),
	.w8(32'h3c3e8106),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31ef9a),
	.w1(32'h3b379a08),
	.w2(32'h3ba8ab29),
	.w3(32'hb97d758b),
	.w4(32'h3b869262),
	.w5(32'h3aa8811b),
	.w6(32'hbbb29fa1),
	.w7(32'h3bbf9dbe),
	.w8(32'hbbe56d3e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39230ba8),
	.w1(32'hba005ce0),
	.w2(32'hbb0ab9c7),
	.w3(32'h3bf94c1e),
	.w4(32'hbb88e3b9),
	.w5(32'hba40dfed),
	.w6(32'h3b4083a0),
	.w7(32'hbc04682c),
	.w8(32'h3afadb28),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8f138),
	.w1(32'hbb63830c),
	.w2(32'hbaf3ad3d),
	.w3(32'h3ae69107),
	.w4(32'hbb2d53bf),
	.w5(32'hbb2614da),
	.w6(32'h38b4e953),
	.w7(32'hbbca1f9b),
	.w8(32'hb976cebd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d51b),
	.w1(32'hbc2048b2),
	.w2(32'hbba19e25),
	.w3(32'hbaa755a3),
	.w4(32'hbc204f2e),
	.w5(32'hbbf30ad0),
	.w6(32'hbb82faa4),
	.w7(32'hbc1de8ce),
	.w8(32'hbc56ff7b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a79b),
	.w1(32'hbb55590b),
	.w2(32'hbc437a0b),
	.w3(32'hbac5f9fe),
	.w4(32'hbbae1b32),
	.w5(32'hbc1fa242),
	.w6(32'h3aae61d5),
	.w7(32'hbc0146c7),
	.w8(32'hbc0f31cf),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3876d5),
	.w1(32'h3ad5b5b0),
	.w2(32'h3b4957c2),
	.w3(32'h3b158f09),
	.w4(32'hba4eafb6),
	.w5(32'h39c079ea),
	.w6(32'hba3e711d),
	.w7(32'hb9b82073),
	.w8(32'h3ad52b33),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913933d),
	.w1(32'hbbed6c14),
	.w2(32'hbbec5d73),
	.w3(32'h3b86b1f4),
	.w4(32'hbc05a038),
	.w5(32'hbbdf5d6c),
	.w6(32'hba83a080),
	.w7(32'hbc34aead),
	.w8(32'hba4856fc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd473c3),
	.w1(32'hbbfe8ddc),
	.w2(32'h3c5a3592),
	.w3(32'hbc5723ec),
	.w4(32'hbad40183),
	.w5(32'h3b529946),
	.w6(32'hba99fc48),
	.w7(32'h3a32fb95),
	.w8(32'h3b679cf7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d1710),
	.w1(32'h3a73f206),
	.w2(32'h3cbd9f30),
	.w3(32'hbb24c8d1),
	.w4(32'hbc755d00),
	.w5(32'h3cfa1329),
	.w6(32'hbbc7d2ff),
	.w7(32'hbbfb81a0),
	.w8(32'h3c9dc210),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc347b66),
	.w1(32'h3c3f4f06),
	.w2(32'hbb86e631),
	.w3(32'h3bb9682b),
	.w4(32'hbbc42b68),
	.w5(32'hbbc0bbda),
	.w6(32'h3b44d4c2),
	.w7(32'h3c6f113e),
	.w8(32'h3bb28e4a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292f6d),
	.w1(32'hbb14281b),
	.w2(32'hb9345ad8),
	.w3(32'h3be65969),
	.w4(32'hbb8198bc),
	.w5(32'hbbdcc033),
	.w6(32'h3afd719c),
	.w7(32'hbbfa3685),
	.w8(32'hbc1ddaf9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0e83d),
	.w1(32'h3bce85e0),
	.w2(32'hbba7048a),
	.w3(32'hbc05c63a),
	.w4(32'h3bff6050),
	.w5(32'hba1ec2f9),
	.w6(32'hbb914bd0),
	.w7(32'h3c8bbe5f),
	.w8(32'h3c133790),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e66d0),
	.w1(32'hbb932e5c),
	.w2(32'h3c231b2d),
	.w3(32'h3ca5c1fa),
	.w4(32'h3b4c4c49),
	.w5(32'h3c165b3c),
	.w6(32'h3c4371dd),
	.w7(32'hba3ca033),
	.w8(32'h3c2cda5d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cc224),
	.w1(32'hbc13d854),
	.w2(32'h3c71722f),
	.w3(32'h3bbd72f1),
	.w4(32'hbb0c719f),
	.w5(32'h3c8b396b),
	.w6(32'h3b034d76),
	.w7(32'h3b990d4e),
	.w8(32'h3bf75159),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c60c5),
	.w1(32'h3c140315),
	.w2(32'hbb303802),
	.w3(32'h3bbc6c7f),
	.w4(32'h3b8ef8d4),
	.w5(32'hbc25f89c),
	.w6(32'h3b3f4df3),
	.w7(32'h3c050b67),
	.w8(32'h3a58a317),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20157e),
	.w1(32'hbbcd478e),
	.w2(32'hbbc87924),
	.w3(32'h3c35cd61),
	.w4(32'hbbba0e2f),
	.w5(32'h3c30364a),
	.w6(32'h3c39f592),
	.w7(32'h3b283587),
	.w8(32'h3b8b4353),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f11bb),
	.w1(32'hbadea10b),
	.w2(32'h3a9b92fb),
	.w3(32'h3bfd86e3),
	.w4(32'hba557dcd),
	.w5(32'hbb14007a),
	.w6(32'h3b3ae029),
	.w7(32'h3acaa696),
	.w8(32'h3aa8878d),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17cd5f),
	.w1(32'hbbe87766),
	.w2(32'hbc3652c7),
	.w3(32'hbc14df82),
	.w4(32'hbbd88639),
	.w5(32'hbb0b036c),
	.w6(32'hbc1da743),
	.w7(32'hbb667873),
	.w8(32'hbac3a02b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2116),
	.w1(32'h3b94c38d),
	.w2(32'h3b096ae3),
	.w3(32'hbb4311d3),
	.w4(32'h3b3e8af8),
	.w5(32'h3b081980),
	.w6(32'hbad648eb),
	.w7(32'h3aaab6be),
	.w8(32'h3ab3358e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39271c6d),
	.w1(32'h3b762b26),
	.w2(32'h3a90a997),
	.w3(32'h39cd12a1),
	.w4(32'h3b5b9755),
	.w5(32'h3b362511),
	.w6(32'hb7b89665),
	.w7(32'h3ac28e25),
	.w8(32'h3ac1be86),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a45707),
	.w1(32'h3b0e3a5d),
	.w2(32'hba19f680),
	.w3(32'hbb6a2a08),
	.w4(32'h39fb9238),
	.w5(32'hba8ed9b6),
	.w6(32'hba9d4319),
	.w7(32'h395909a4),
	.w8(32'h3c019165),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1f39a),
	.w1(32'h3a4617f3),
	.w2(32'h3abdad1c),
	.w3(32'h3b1dc5d0),
	.w4(32'h3b9ef11d),
	.w5(32'hbbb424a1),
	.w6(32'h3c217354),
	.w7(32'h3b4829db),
	.w8(32'h3ade5089),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa66bb),
	.w1(32'hbb94d64c),
	.w2(32'hbbd92e26),
	.w3(32'hbb837dbc),
	.w4(32'hbc1a5a8e),
	.w5(32'hbc0829a7),
	.w6(32'h3ba3ec45),
	.w7(32'hbbd53fca),
	.w8(32'hbb35b1fe),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae21f2b),
	.w1(32'h3af3e57c),
	.w2(32'h3b4a17a6),
	.w3(32'hbb99585d),
	.w4(32'h3b74670b),
	.w5(32'h3c8f358b),
	.w6(32'hbb1de49e),
	.w7(32'h3c381f05),
	.w8(32'hba91a309),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9874820),
	.w1(32'hbad2b03e),
	.w2(32'h3a3f9283),
	.w3(32'hbb46073f),
	.w4(32'hba558442),
	.w5(32'h3c1393c5),
	.w6(32'hba9b1677),
	.w7(32'hbb81c73b),
	.w8(32'h3b12147f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b01be),
	.w1(32'hbb7fac78),
	.w2(32'hbb839ac4),
	.w3(32'h3b56cfd6),
	.w4(32'hbc3b5246),
	.w5(32'hbc114fc7),
	.w6(32'h3ba2dc66),
	.w7(32'hbc03d272),
	.w8(32'hbb4ce622),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90def5),
	.w1(32'h3aff563d),
	.w2(32'h3a0ec5d2),
	.w3(32'h3c012b65),
	.w4(32'h3b25d6a0),
	.w5(32'hbb901b3d),
	.w6(32'h3b1cd55f),
	.w7(32'h3af730d5),
	.w8(32'h39d16d4e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9564c8),
	.w1(32'h3b793fbe),
	.w2(32'h3b9f3893),
	.w3(32'h39a6f242),
	.w4(32'hba2a0740),
	.w5(32'h3c8c7de0),
	.w6(32'h3b85e6d8),
	.w7(32'h3bcb2eb5),
	.w8(32'h3a3e9118),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61e6e2),
	.w1(32'hba54f46a),
	.w2(32'h3bd8e925),
	.w3(32'h3bdd3836),
	.w4(32'h3a3620f9),
	.w5(32'h3c656dbf),
	.w6(32'h3c59204a),
	.w7(32'hbb4041f1),
	.w8(32'h3b983423),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf67b28),
	.w1(32'h3b75d667),
	.w2(32'hbbf8b3d3),
	.w3(32'hbb1649f4),
	.w4(32'hbbba0e0b),
	.w5(32'h3b1405b1),
	.w6(32'hbb99c56a),
	.w7(32'h3bb39345),
	.w8(32'h3a291440),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb8b9),
	.w1(32'h3b54cb49),
	.w2(32'hbc0ffc4f),
	.w3(32'h3b194787),
	.w4(32'h3b1252c4),
	.w5(32'hbbca44ed),
	.w6(32'hba94ac71),
	.w7(32'h3ab7aa2d),
	.w8(32'hbbdef648),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff075e),
	.w1(32'hbb41e705),
	.w2(32'hbb097435),
	.w3(32'h3c0745aa),
	.w4(32'hbaaf7ef3),
	.w5(32'h3bb7e8ca),
	.w6(32'h3c4b1419),
	.w7(32'h3b1c72c7),
	.w8(32'hba5a2de3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd44c3),
	.w1(32'hbb82b378),
	.w2(32'hbbbaa685),
	.w3(32'h3b6c4d0c),
	.w4(32'hba6a97bc),
	.w5(32'hbc1b7183),
	.w6(32'h3b19e940),
	.w7(32'hbbcb3f90),
	.w8(32'hbbbaf7fa),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb192dd6),
	.w1(32'hb9bbd1b9),
	.w2(32'h3c4d6b48),
	.w3(32'hbaf33e75),
	.w4(32'h3b8d4b0c),
	.w5(32'h3b592384),
	.w6(32'h3b0a170b),
	.w7(32'h3b9fa2fd),
	.w8(32'h3a92c1c5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc3f1a),
	.w1(32'hbb9bdeac),
	.w2(32'h3b2243a6),
	.w3(32'h3bfd9795),
	.w4(32'hbbd34561),
	.w5(32'hbb02090f),
	.w6(32'h3b217d6b),
	.w7(32'hbc04ef61),
	.w8(32'hbaf1a427),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac44042),
	.w1(32'h3b653a95),
	.w2(32'hba952863),
	.w3(32'hbb06065b),
	.w4(32'hbba0d422),
	.w5(32'hbc1080dd),
	.w6(32'h3b519403),
	.w7(32'hbb11b51a),
	.w8(32'hbb9881f5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5198ad),
	.w1(32'hba72552b),
	.w2(32'h3b4f8641),
	.w3(32'h3bbc7206),
	.w4(32'hbb8465d8),
	.w5(32'hbbbc5ac5),
	.w6(32'h3b2af5b5),
	.w7(32'hbbc43558),
	.w8(32'h37c3d842),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8664a7),
	.w1(32'h3981baa6),
	.w2(32'h3b260092),
	.w3(32'hba9109c5),
	.w4(32'hbaff17e6),
	.w5(32'h3a67a4f6),
	.w6(32'hbb03040d),
	.w7(32'hba5f4398),
	.w8(32'hbb56e7de),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02c1cb),
	.w1(32'hbb546517),
	.w2(32'h3ba02602),
	.w3(32'h3b56906b),
	.w4(32'hbc345347),
	.w5(32'h3c4a82d2),
	.w6(32'h3c3572fb),
	.w7(32'hbb24220e),
	.w8(32'h3c2dfa8e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ffb18),
	.w1(32'hbb8a1a81),
	.w2(32'hbbe586cb),
	.w3(32'h3b4b4aa4),
	.w4(32'hbb7eb3f5),
	.w5(32'h370c20ed),
	.w6(32'h3c27564d),
	.w7(32'hbb4fe8da),
	.w8(32'h3b51f52f),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6e89),
	.w1(32'h3bbd9136),
	.w2(32'h3b980b73),
	.w3(32'h3aa43685),
	.w4(32'h3bcd75bb),
	.w5(32'hbaddb382),
	.w6(32'hbba8d9a0),
	.w7(32'h3b9dc1fa),
	.w8(32'h3bee2d07),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb516ac),
	.w1(32'hbc0911c8),
	.w2(32'hbba5e212),
	.w3(32'hba8bbe2b),
	.w4(32'hb8383fb0),
	.w5(32'hbb9f9cc8),
	.w6(32'hbaffa493),
	.w7(32'hbbeda057),
	.w8(32'hbb579bf2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2071c8),
	.w1(32'hba746df3),
	.w2(32'h38c8df80),
	.w3(32'hba957c1f),
	.w4(32'hbbaba9c1),
	.w5(32'h3a079593),
	.w6(32'h3b3a0510),
	.w7(32'hbaa8ce4d),
	.w8(32'hbba4f314),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3df38a),
	.w1(32'h3c13475c),
	.w2(32'h3b89a8b4),
	.w3(32'hbb2b81e3),
	.w4(32'h3c38bed2),
	.w5(32'hbb232344),
	.w6(32'hba77355b),
	.w7(32'h3ab3c2a3),
	.w8(32'h3bad95b4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6274b1),
	.w1(32'h39e63f19),
	.w2(32'hba16db9b),
	.w3(32'h3bfc69dd),
	.w4(32'h3c0deb22),
	.w5(32'h3bac84c8),
	.w6(32'h3ba68f41),
	.w7(32'h3b59a63c),
	.w8(32'h3c3a2742),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c4fdb),
	.w1(32'h39f2549a),
	.w2(32'hbc18506b),
	.w3(32'h3bf2167c),
	.w4(32'hbb7a042e),
	.w5(32'h3b0a97fd),
	.w6(32'h39c79353),
	.w7(32'h3aa02b7c),
	.w8(32'hbb8a8fe1),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be26bd5),
	.w1(32'hba6dbfc6),
	.w2(32'hbb1a6554),
	.w3(32'h3bedae74),
	.w4(32'h3af30240),
	.w5(32'hbbe07213),
	.w6(32'h3bda6b87),
	.w7(32'h3adfba0d),
	.w8(32'h3b8bd841),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d4b6),
	.w1(32'hbc9fd762),
	.w2(32'h3c2e7842),
	.w3(32'h3aefcf87),
	.w4(32'h3b6ecf68),
	.w5(32'hbba695af),
	.w6(32'h3a92cd3b),
	.w7(32'hbbdf220b),
	.w8(32'h3be4b88b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa01f6),
	.w1(32'h3b0b84ab),
	.w2(32'h3be50584),
	.w3(32'hbb5317ba),
	.w4(32'h3b267078),
	.w5(32'h3b1d6407),
	.w6(32'h3a0cd6a9),
	.w7(32'hbb817ec0),
	.w8(32'hbb5ae27b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab7c5a),
	.w1(32'h3bafc3c4),
	.w2(32'h3b0fbfaf),
	.w3(32'h3b17bca5),
	.w4(32'hba89322b),
	.w5(32'hbb0f08d9),
	.w6(32'hbacffcbe),
	.w7(32'h3ba26df9),
	.w8(32'h3b05157b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c577e),
	.w1(32'h3b648fb8),
	.w2(32'h3a0e8ff5),
	.w3(32'hbbb4e294),
	.w4(32'hbaf827eb),
	.w5(32'h3ad232e3),
	.w6(32'h39db59d8),
	.w7(32'hbba05ecd),
	.w8(32'h3bd46553),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a229c3b),
	.w1(32'h3bb250a3),
	.w2(32'h3bb765d8),
	.w3(32'h3c10e73e),
	.w4(32'h3aad6961),
	.w5(32'hb9b8b8a0),
	.w6(32'h3b296feb),
	.w7(32'h3af73a5b),
	.w8(32'h3be2f33f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0331a),
	.w1(32'hbb759b75),
	.w2(32'h39270907),
	.w3(32'h3b0cb52c),
	.w4(32'hbc29c03d),
	.w5(32'h3b18a977),
	.w6(32'h3c1141b6),
	.w7(32'hbbf74847),
	.w8(32'hbbc6fe37),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa090b),
	.w1(32'hb903a0ec),
	.w2(32'h3ba8cd40),
	.w3(32'hbc1019dc),
	.w4(32'hbb1569c9),
	.w5(32'h3ba54c98),
	.w6(32'hbc5334f8),
	.w7(32'hbb0cbfda),
	.w8(32'h3b7ed466),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8de97),
	.w1(32'hb991f1dd),
	.w2(32'h3b20c268),
	.w3(32'h3c70bde2),
	.w4(32'hb9cbba71),
	.w5(32'hbbe2288d),
	.w6(32'h3c0208dc),
	.w7(32'hbb066882),
	.w8(32'hbae4d2bf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d9e4d),
	.w1(32'hbb6c9685),
	.w2(32'h3a41390b),
	.w3(32'h391672c0),
	.w4(32'hbc018c49),
	.w5(32'h3a81db5c),
	.w6(32'h3ac9af16),
	.w7(32'hba8108a5),
	.w8(32'hbbd92d17),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9863351),
	.w1(32'h3b98eedc),
	.w2(32'h3c1cd9ef),
	.w3(32'hb9e42596),
	.w4(32'h3a892cf1),
	.w5(32'h3c70005a),
	.w6(32'h3ba39ceb),
	.w7(32'hbb9ecb3a),
	.w8(32'h3c828fe3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923fa80),
	.w1(32'h3cbb1ccd),
	.w2(32'h3c01c327),
	.w3(32'h3bbf63d4),
	.w4(32'h3c84b906),
	.w5(32'hbbdad9a7),
	.w6(32'h3b5135a1),
	.w7(32'h3b9608d6),
	.w8(32'h39f334ef),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80443c),
	.w1(32'hbb88a230),
	.w2(32'h3bab3d7f),
	.w3(32'h3afb00e7),
	.w4(32'hbae686c5),
	.w5(32'h3c8fafdc),
	.w6(32'h3c95670c),
	.w7(32'hba6eb996),
	.w8(32'hb9e52a68),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07d47b),
	.w1(32'hbb41254a),
	.w2(32'hbb91a4b3),
	.w3(32'h3b78994c),
	.w4(32'hbb914de8),
	.w5(32'hbb5cbc58),
	.w6(32'hbc3dd373),
	.w7(32'hbb3d4cb9),
	.w8(32'h39f2ff27),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80c134),
	.w1(32'hbb836acf),
	.w2(32'hbb11b001),
	.w3(32'h39538a2a),
	.w4(32'hb83203e5),
	.w5(32'h3c77b9e4),
	.w6(32'hbc256e12),
	.w7(32'hbac2369e),
	.w8(32'h3abd4ad9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb481d31),
	.w1(32'hbbe6a68d),
	.w2(32'hbbded979),
	.w3(32'hbbc2a608),
	.w4(32'h3adc98fe),
	.w5(32'h3ca13593),
	.w6(32'hbc2cd598),
	.w7(32'h3b2db52d),
	.w8(32'hbace4d00),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c3ced),
	.w1(32'hbb114773),
	.w2(32'hbb00cc1f),
	.w3(32'hb9e7c062),
	.w4(32'h3bd27a1d),
	.w5(32'h3cc237e0),
	.w6(32'hbc3e1900),
	.w7(32'h38479233),
	.w8(32'hbb9a6b45),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ec94e),
	.w1(32'h3b8c5a92),
	.w2(32'h3c0e3a23),
	.w3(32'h3c0ccf06),
	.w4(32'h3b8e5a60),
	.w5(32'hba25fa26),
	.w6(32'hbbae3c27),
	.w7(32'h3bb9defe),
	.w8(32'h3a2db8f1),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d475),
	.w1(32'hbb4a87db),
	.w2(32'hbc8f48fd),
	.w3(32'hbc795616),
	.w4(32'hb9a155db),
	.w5(32'hbbdf7913),
	.w6(32'hbc7b9352),
	.w7(32'hbb490594),
	.w8(32'hbc798dbf),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c422f),
	.w1(32'hbae77650),
	.w2(32'hbb42a141),
	.w3(32'h3b942fef),
	.w4(32'hbb91080c),
	.w5(32'h3bd6bf4b),
	.w6(32'hbb92659c),
	.w7(32'hbb9fb52b),
	.w8(32'hbb9e6cd1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379fe9c3),
	.w1(32'hbbfcab9e),
	.w2(32'hbbd08aee),
	.w3(32'h39e3e14b),
	.w4(32'hbbbb5351),
	.w5(32'hbc1a1172),
	.w6(32'h3b2dabda),
	.w7(32'hbb3e0334),
	.w8(32'hbb92ef9d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05328d),
	.w1(32'h3c733b37),
	.w2(32'hba94b361),
	.w3(32'hbc2dbf25),
	.w4(32'hba20e00b),
	.w5(32'hbc85171a),
	.w6(32'hbc0a64a0),
	.w7(32'h3bba1750),
	.w8(32'h3a69267e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12ca61),
	.w1(32'h3b29688c),
	.w2(32'hbabf70f7),
	.w3(32'hbb19fa17),
	.w4(32'h39053cfa),
	.w5(32'hb9ea227a),
	.w6(32'h3bcc6329),
	.w7(32'hbab485ee),
	.w8(32'hbb2d6b49),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c898),
	.w1(32'hbb18484e),
	.w2(32'hbb13549d),
	.w3(32'h3b00917f),
	.w4(32'h39c18290),
	.w5(32'hbb73fd4f),
	.w6(32'hbb178188),
	.w7(32'h3bb1753d),
	.w8(32'hbb435b1e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b385),
	.w1(32'hb957affd),
	.w2(32'hbbb27b28),
	.w3(32'hba701c8c),
	.w4(32'h3bda285a),
	.w5(32'hbbc40c72),
	.w6(32'hba0b7da2),
	.w7(32'h3bb07c9a),
	.w8(32'hbc22302c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7a52),
	.w1(32'h3b85cef3),
	.w2(32'hbb408019),
	.w3(32'hbc2c5b4a),
	.w4(32'h3b60071f),
	.w5(32'hbbf2baf7),
	.w6(32'hbae9c14b),
	.w7(32'hbb395cbb),
	.w8(32'hbc554f03),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489839),
	.w1(32'hbb9f3e0d),
	.w2(32'hbbfd7c46),
	.w3(32'hbb5359f8),
	.w4(32'hbc36b049),
	.w5(32'h3b21c06c),
	.w6(32'hbc0420c8),
	.w7(32'hbbcd9ec1),
	.w8(32'hbb26997c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee03b0),
	.w1(32'hbc359341),
	.w2(32'h3a3ac137),
	.w3(32'h3c09c7c2),
	.w4(32'hbbe8617b),
	.w5(32'h3acc3e45),
	.w6(32'h3c200b1c),
	.w7(32'hba2cce3b),
	.w8(32'h3bc55642),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbffa96),
	.w1(32'hbaf3bbbc),
	.w2(32'hbc4cad14),
	.w3(32'hbc132f0e),
	.w4(32'hba828c5c),
	.w5(32'h3c5c16d9),
	.w6(32'hbbb49d03),
	.w7(32'h3b86cee3),
	.w8(32'h3c025e99),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9586a),
	.w1(32'h3b0528ed),
	.w2(32'h3bee29f7),
	.w3(32'hbb94a49f),
	.w4(32'h3b67b5e0),
	.w5(32'hbc11ee4f),
	.w6(32'hbb21f19c),
	.w7(32'hbae91f42),
	.w8(32'hbc6cfc02),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0875b7),
	.w1(32'hbbf585f9),
	.w2(32'hbc20dcee),
	.w3(32'hbc20001e),
	.w4(32'hba924c42),
	.w5(32'hbba15fad),
	.w6(32'hbc297edb),
	.w7(32'h3b34e2ce),
	.w8(32'hbb03d461),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd943bf),
	.w1(32'hbbd0eed4),
	.w2(32'h3ab4b249),
	.w3(32'hbbde4b1e),
	.w4(32'hbc15c720),
	.w5(32'h3b262012),
	.w6(32'hba580f6d),
	.w7(32'hbc1d3e9e),
	.w8(32'hbbd9c483),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba311ee),
	.w1(32'h3b278e7f),
	.w2(32'hbbf791fd),
	.w3(32'h3b5bf3b8),
	.w4(32'hbc20191f),
	.w5(32'hbc63db2e),
	.w6(32'h3b59c538),
	.w7(32'h3a169371),
	.w8(32'hba01cc42),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad1c6),
	.w1(32'hbbac8ffd),
	.w2(32'hbb6b63b0),
	.w3(32'hbc392d47),
	.w4(32'hbbc1cb8b),
	.w5(32'h3c04c415),
	.w6(32'h3b58ac6c),
	.w7(32'hbba887a4),
	.w8(32'hbb488010),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b907752),
	.w1(32'hbacb976f),
	.w2(32'hbbed0d00),
	.w3(32'hba93d2ca),
	.w4(32'h3bb98bf1),
	.w5(32'h3a2eaa5d),
	.w6(32'hbb986521),
	.w7(32'h3b34c1bf),
	.w8(32'hbb486d09),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d6d6c),
	.w1(32'h3adf944e),
	.w2(32'hbc0da57c),
	.w3(32'h3ba39577),
	.w4(32'hbbf242ee),
	.w5(32'hbc3e12af),
	.w6(32'h3ba0315f),
	.w7(32'hbbfd3971),
	.w8(32'hbc698e23),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849643),
	.w1(32'hbb7b730e),
	.w2(32'h3c988ad7),
	.w3(32'hbc95e15c),
	.w4(32'h3bffc7ba),
	.w5(32'h3cb334f5),
	.w6(32'hbc6408c0),
	.w7(32'h3bc65e95),
	.w8(32'h3c92f44d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18ab16),
	.w1(32'h3bb6bec9),
	.w2(32'hbba3c2d7),
	.w3(32'h3b942a4a),
	.w4(32'h3b67f9b9),
	.w5(32'h3c105156),
	.w6(32'hbb590363),
	.w7(32'h3b266aec),
	.w8(32'hbb4cce25),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59c2a9),
	.w1(32'hbbdd606c),
	.w2(32'hba3028bb),
	.w3(32'hba46889b),
	.w4(32'hbc345cf5),
	.w5(32'hbb229c53),
	.w6(32'h3b29a818),
	.w7(32'hbb106558),
	.w8(32'h3b261505),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1db57),
	.w1(32'hbb830b7d),
	.w2(32'hbaa4c9d5),
	.w3(32'hbbbf5ab7),
	.w4(32'hbb97a9db),
	.w5(32'hbb731fd7),
	.w6(32'hbb648f39),
	.w7(32'hbb7965c9),
	.w8(32'h3a1a8095),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3e082),
	.w1(32'hbb3b2def),
	.w2(32'hbc11bd35),
	.w3(32'hbad5420f),
	.w4(32'h3caf50bb),
	.w5(32'h3c3782e0),
	.w6(32'h3bbdeb8b),
	.w7(32'h3b75ac42),
	.w8(32'h3adbf753),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a14fa),
	.w1(32'h3bc7ae15),
	.w2(32'hbae7338a),
	.w3(32'h3c6cfec7),
	.w4(32'h3ba3ae5f),
	.w5(32'h3ba0c3c0),
	.w6(32'h3c02b24e),
	.w7(32'h3b591f24),
	.w8(32'hbb9b54af),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50eaba),
	.w1(32'hbc1f85f3),
	.w2(32'hbc0ffb71),
	.w3(32'hbc01e12f),
	.w4(32'hbc1d9fa7),
	.w5(32'h3ad12d43),
	.w6(32'hbc1f24e6),
	.w7(32'hbc0c9f5d),
	.w8(32'h3a93168f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd167a5),
	.w1(32'h39e2d0b3),
	.w2(32'hbb942bf3),
	.w3(32'hbb4fffff),
	.w4(32'hbbafea5b),
	.w5(32'h3c6c02b4),
	.w6(32'h39f28c9b),
	.w7(32'hba97ff9d),
	.w8(32'hbbc211ad),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb557aa),
	.w1(32'h3b222e65),
	.w2(32'h3b88cdd3),
	.w3(32'h3b816049),
	.w4(32'hbc00dcac),
	.w5(32'h3b06cd15),
	.w6(32'hbc15ebdf),
	.w7(32'hba7b6ca0),
	.w8(32'hbac49667),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932987b),
	.w1(32'h3c26f69c),
	.w2(32'hbbcd0088),
	.w3(32'h3a89c4ce),
	.w4(32'hba97efdd),
	.w5(32'hbb7fb6e6),
	.w6(32'hbae2cab3),
	.w7(32'h3bef1139),
	.w8(32'hb993b6f4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba861769),
	.w1(32'hba19bec0),
	.w2(32'hbab56658),
	.w3(32'hbbcdb0e6),
	.w4(32'hbb027abd),
	.w5(32'hbb1244f0),
	.w6(32'h3b5890fe),
	.w7(32'h3b2995a5),
	.w8(32'h3a3c3410),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7b1f),
	.w1(32'h3c3a260c),
	.w2(32'hbb5563dd),
	.w3(32'h3b57e84a),
	.w4(32'h3b935e56),
	.w5(32'hbb8cbe07),
	.w6(32'h3bbf3285),
	.w7(32'hba15f1a8),
	.w8(32'hbaf0a6cb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128bfd),
	.w1(32'h3a957b87),
	.w2(32'hbbd57327),
	.w3(32'h3bf258e9),
	.w4(32'hbb0b1a97),
	.w5(32'hbb9dadc2),
	.w6(32'h3c6b1879),
	.w7(32'hbc2ffbf8),
	.w8(32'hbc2ed478),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a6ae3),
	.w1(32'hba47f8e1),
	.w2(32'hba6016d0),
	.w3(32'h3c32ddc7),
	.w4(32'h3828ff0d),
	.w5(32'h3b8de1bc),
	.w6(32'h3b0d1dbb),
	.w7(32'h3b03fe07),
	.w8(32'h3b52721e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8869cc),
	.w1(32'hbb2bdc79),
	.w2(32'hbba7ee97),
	.w3(32'h39f263c9),
	.w4(32'h39381548),
	.w5(32'h3b2e509d),
	.w6(32'hbb46912b),
	.w7(32'h3b7d5729),
	.w8(32'hbb483084),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac993a0),
	.w1(32'hbbd9deea),
	.w2(32'hbbbe27e5),
	.w3(32'hbc8d0bd0),
	.w4(32'hbbb2aa8a),
	.w5(32'h3b7d4793),
	.w6(32'hbb857abd),
	.w7(32'hba6a786c),
	.w8(32'hbac381e1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4686b),
	.w1(32'h398ce350),
	.w2(32'hba86021b),
	.w3(32'h39f00a4e),
	.w4(32'hbb98c3e4),
	.w5(32'hbc05b798),
	.w6(32'h3b9c157e),
	.w7(32'hb940d6ed),
	.w8(32'h37428a0f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5d17),
	.w1(32'hb9f3fac7),
	.w2(32'hbba8179a),
	.w3(32'h3b8d8ab9),
	.w4(32'hbae8e855),
	.w5(32'h3be5fd32),
	.w6(32'h3afdfbd8),
	.w7(32'hbb33a317),
	.w8(32'hbb919d60),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89158c),
	.w1(32'h3bed9ff0),
	.w2(32'hbba0eba8),
	.w3(32'hbbd5ab6f),
	.w4(32'hbb859746),
	.w5(32'h3c0575f5),
	.w6(32'hbb76205f),
	.w7(32'hbc116015),
	.w8(32'h3b29bed6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc184421),
	.w1(32'hbb3a8b5f),
	.w2(32'h3a25e6ad),
	.w3(32'hbb59839a),
	.w4(32'hbc001147),
	.w5(32'hbc1e5ffa),
	.w6(32'hbb5ae6f7),
	.w7(32'hbb9f48f1),
	.w8(32'hbb898e0e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852bc5),
	.w1(32'h391598b7),
	.w2(32'hbb276e49),
	.w3(32'hbbc6e291),
	.w4(32'h3b8aa3bc),
	.w5(32'h3bc17f78),
	.w6(32'h39cdd8cc),
	.w7(32'hbb1013d4),
	.w8(32'hbba9134a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaa9f7),
	.w1(32'hbae324cf),
	.w2(32'h3b79a86a),
	.w3(32'h3b906257),
	.w4(32'h3af2d6a5),
	.w5(32'h3c0fb9e6),
	.w6(32'hb96f0eac),
	.w7(32'hba2eeb0a),
	.w8(32'h3bf6f75c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79a0a4),
	.w1(32'h3ac0a7c9),
	.w2(32'hbc1d8214),
	.w3(32'hbb87598e),
	.w4(32'hba886588),
	.w5(32'hbc816462),
	.w6(32'hbae3c54b),
	.w7(32'hbaaaa77e),
	.w8(32'hbc6c2d47),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18865d),
	.w1(32'hbc5c0b57),
	.w2(32'hbb2c7ca6),
	.w3(32'hbbe07f81),
	.w4(32'hbb334d7b),
	.w5(32'h3c93d274),
	.w6(32'hbb043bf2),
	.w7(32'hbbe8c4dc),
	.w8(32'hb9db588b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0451c),
	.w1(32'hbaa28dcb),
	.w2(32'hba97cae2),
	.w3(32'hbb7cbb46),
	.w4(32'hbb52c6d0),
	.w5(32'h3c6e1b86),
	.w6(32'hbc846711),
	.w7(32'hbb567541),
	.w8(32'h3c1338ee),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b026d77),
	.w1(32'h3c14f78c),
	.w2(32'h3b6b0438),
	.w3(32'hbc01183b),
	.w4(32'h3c134565),
	.w5(32'h3bc60d40),
	.w6(32'hbc0211db),
	.w7(32'h3a807612),
	.w8(32'h3b3fed24),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de2c7),
	.w1(32'hbb1dbff8),
	.w2(32'hbb102468),
	.w3(32'hbc777b51),
	.w4(32'hbb81a4bb),
	.w5(32'h3c79fb51),
	.w6(32'hbc0fb0e3),
	.w7(32'h3c7e8d9c),
	.w8(32'h3c92e4b4),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a7ea9),
	.w1(32'h3c60789d),
	.w2(32'h3b3e53a6),
	.w3(32'h3ca04293),
	.w4(32'h3c186507),
	.w5(32'h3a98456a),
	.w6(32'h3cd310d6),
	.w7(32'h3c100eda),
	.w8(32'hbb10eb65),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f69a5),
	.w1(32'h3a9fcb39),
	.w2(32'hba063c33),
	.w3(32'hbc12c3f9),
	.w4(32'hbb997281),
	.w5(32'h3b692c3c),
	.w6(32'h3c0b6507),
	.w7(32'hba98f2b4),
	.w8(32'h3b91567b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c36f4),
	.w1(32'hbc1d32bc),
	.w2(32'hbb8f950e),
	.w3(32'h3c55ff74),
	.w4(32'hbb151cef),
	.w5(32'hbb8bc7c0),
	.w6(32'h3be3e32a),
	.w7(32'hbc083e04),
	.w8(32'hbbd907d6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba86c16),
	.w1(32'h3bdaedf8),
	.w2(32'hba3bc2b2),
	.w3(32'h3bc4006b),
	.w4(32'hb8bdcdf0),
	.w5(32'h3c33472f),
	.w6(32'hbb0886ec),
	.w7(32'hb8829a9a),
	.w8(32'hb9aa39c1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e289c),
	.w1(32'hbbf31f07),
	.w2(32'h3b027415),
	.w3(32'hbbfa42b9),
	.w4(32'h3bcf5362),
	.w5(32'hbc0f250a),
	.w6(32'hbbc02d7c),
	.w7(32'hbc15a3ab),
	.w8(32'hbba7dad1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0a22),
	.w1(32'h3b93ff96),
	.w2(32'hbb4321fc),
	.w3(32'hbacb01ad),
	.w4(32'hbb951da6),
	.w5(32'h3bfbaa09),
	.w6(32'h3c37d843),
	.w7(32'hbafec3df),
	.w8(32'hbb75ac8f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule