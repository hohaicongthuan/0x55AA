module layer_10_featuremap_88(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacf733),
	.w1(32'hbab51ef0),
	.w2(32'h3b095374),
	.w3(32'hbaf811f3),
	.w4(32'h3b9609b8),
	.w5(32'h3c88e9c0),
	.w6(32'h3bb35f19),
	.w7(32'hba8430e6),
	.w8(32'h39e0750b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68f6b3),
	.w1(32'h3b457750),
	.w2(32'hba08286e),
	.w3(32'h3b978f4d),
	.w4(32'hba4d7e97),
	.w5(32'hba6731dc),
	.w6(32'hbafa83bc),
	.w7(32'hb98d1290),
	.w8(32'hbae86883),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7e30a),
	.w1(32'hba933288),
	.w2(32'hbb986c34),
	.w3(32'h3bb8e83c),
	.w4(32'hbbcb4f5e),
	.w5(32'hbb73df46),
	.w6(32'h3b45894d),
	.w7(32'h3b75bdb6),
	.w8(32'hbbfbb524),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38bb9f),
	.w1(32'h3ac2e0ab),
	.w2(32'h3a82698a),
	.w3(32'hbbbd084f),
	.w4(32'hbbd96de4),
	.w5(32'hbac094d5),
	.w6(32'hbb94ee44),
	.w7(32'hbb04a257),
	.w8(32'h3b6ddedf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae20a9c),
	.w1(32'h3c07b125),
	.w2(32'hba0cc682),
	.w3(32'hbbaa392f),
	.w4(32'hbb31c7e9),
	.w5(32'hbaff6ded),
	.w6(32'hbb25b060),
	.w7(32'h3bbcd599),
	.w8(32'h3c060f76),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba169b10),
	.w1(32'hb9420b1b),
	.w2(32'h3ae55564),
	.w3(32'h39962ec2),
	.w4(32'hba123439),
	.w5(32'h3aaeeaff),
	.w6(32'hbca83ecd),
	.w7(32'hba805738),
	.w8(32'hbb73b395),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba147ba1),
	.w1(32'h3b23de6f),
	.w2(32'hbc1cd4e9),
	.w3(32'h3be8f20e),
	.w4(32'hba34ad72),
	.w5(32'hbc8e80ad),
	.w6(32'h3bc48f37),
	.w7(32'h3b9dc043),
	.w8(32'h3c260dca),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db856),
	.w1(32'h3bbebc44),
	.w2(32'hbbd8699e),
	.w3(32'hbc40ac40),
	.w4(32'h3ae04184),
	.w5(32'hb9e172e9),
	.w6(32'h3acbb176),
	.w7(32'hbc008fc6),
	.w8(32'hbbe466fa),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2783a2),
	.w1(32'hb96d477d),
	.w2(32'hb9f30b0a),
	.w3(32'h3bb45593),
	.w4(32'h3b179440),
	.w5(32'hbaad2db4),
	.w6(32'hbc16bbc2),
	.w7(32'h39fe9706),
	.w8(32'h3811d80e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2f641),
	.w1(32'hbbb456e0),
	.w2(32'hbc509ccd),
	.w3(32'h3c2ecfc2),
	.w4(32'h3bce9e8f),
	.w5(32'hbc434692),
	.w6(32'hbbe8b68f),
	.w7(32'h3cdb843f),
	.w8(32'h3b5743d1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabca1c),
	.w1(32'hba60c642),
	.w2(32'h3a67c217),
	.w3(32'h3c53b01a),
	.w4(32'hbb41d3dd),
	.w5(32'hbbcfba96),
	.w6(32'h3ab7c7c0),
	.w7(32'h3b176ffe),
	.w8(32'hbafb9561),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba617e6),
	.w1(32'hba4d7f11),
	.w2(32'hbc3f4dae),
	.w3(32'h3c246a9a),
	.w4(32'h3c405cab),
	.w5(32'hbba2c577),
	.w6(32'h3a0240d0),
	.w7(32'h3a8b354d),
	.w8(32'hbc2d67f9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f6d4),
	.w1(32'hbb9463e6),
	.w2(32'hbc178bc0),
	.w3(32'h3b496042),
	.w4(32'h3a18f161),
	.w5(32'hbbaccbf0),
	.w6(32'h3bb79e11),
	.w7(32'hbae7f4b9),
	.w8(32'hbb5e5676),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a0d9b),
	.w1(32'hba6e7ca4),
	.w2(32'hbbbdbc2a),
	.w3(32'hbbf79ef6),
	.w4(32'h3c167f6e),
	.w5(32'hbb9d514c),
	.w6(32'h3b8b2aeb),
	.w7(32'hbb9cf51e),
	.w8(32'h3b968787),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcec44),
	.w1(32'h3bb6c892),
	.w2(32'h3aa4f974),
	.w3(32'hbb94b3de),
	.w4(32'h3ae70ad9),
	.w5(32'h3afba360),
	.w6(32'h3b432f0e),
	.w7(32'h3bd3d1b4),
	.w8(32'hba84a3f9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba701fc4),
	.w1(32'hbbad6188),
	.w2(32'hbb890ae3),
	.w3(32'hbc5e05f1),
	.w4(32'hbb4a0715),
	.w5(32'hbb340ccd),
	.w6(32'hba8c14ec),
	.w7(32'hbb1f3037),
	.w8(32'hbc21c8e5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f076c),
	.w1(32'h3bced286),
	.w2(32'h3ae93be1),
	.w3(32'h3bad08d1),
	.w4(32'h387c8f1c),
	.w5(32'h3b8e9721),
	.w6(32'h3a95a6f7),
	.w7(32'h3b896b03),
	.w8(32'hbaeab7ac),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8eefda),
	.w1(32'hbaebe8de),
	.w2(32'hbb5b566d),
	.w3(32'h3b05f296),
	.w4(32'h3b0f7f11),
	.w5(32'hbc1df98f),
	.w6(32'hbb7b08d0),
	.w7(32'h3b79fda7),
	.w8(32'hbb4275b4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f510e),
	.w1(32'hbc3f49db),
	.w2(32'hbc217ff8),
	.w3(32'h3b778f98),
	.w4(32'h3b46c867),
	.w5(32'hbbb9d779),
	.w6(32'hbbbe02c7),
	.w7(32'hbbf71d77),
	.w8(32'hbb04b385),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34d87d),
	.w1(32'h3a1aa8da),
	.w2(32'hbb5a5830),
	.w3(32'h3a31eb45),
	.w4(32'h3b9c8edd),
	.w5(32'h3aed48bb),
	.w6(32'hbbe7c587),
	.w7(32'hbacd2f9e),
	.w8(32'hbaf50310),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab82b1a),
	.w1(32'hba6ed3d7),
	.w2(32'hbc200891),
	.w3(32'hbba9f271),
	.w4(32'hb8a0b7cd),
	.w5(32'h3a2cf1e9),
	.w6(32'hbbd353eb),
	.w7(32'hbb8cc4f7),
	.w8(32'hbba352e7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa7fe7),
	.w1(32'h3b721bd2),
	.w2(32'h3b4e6eef),
	.w3(32'hb9b49e58),
	.w4(32'h3b0b9bb8),
	.w5(32'hba116304),
	.w6(32'hb9af5d9a),
	.w7(32'h3a08c5a5),
	.w8(32'h3b9b4414),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd871),
	.w1(32'hbb95b96f),
	.w2(32'hbc8b1e79),
	.w3(32'h3c0957ef),
	.w4(32'h3b69d1e7),
	.w5(32'hbb63f2a9),
	.w6(32'h3a690a17),
	.w7(32'h3bf04346),
	.w8(32'hbc2d5a63),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae38059),
	.w1(32'hbb8ea3b3),
	.w2(32'hbba1719c),
	.w3(32'h3b5b1528),
	.w4(32'hbab56818),
	.w5(32'h3b3b8975),
	.w6(32'h3a35ccdc),
	.w7(32'h3a344eda),
	.w8(32'h3b4f269e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdff48e),
	.w1(32'h3c235774),
	.w2(32'h3c75ca2c),
	.w3(32'h3bef7090),
	.w4(32'h3b4c644c),
	.w5(32'h3bddef1e),
	.w6(32'h3af9ab2f),
	.w7(32'h3a88ffff),
	.w8(32'hbb6f29db),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12599),
	.w1(32'hbb0a3285),
	.w2(32'h3c728ff1),
	.w3(32'hbb6375df),
	.w4(32'hba4212fa),
	.w5(32'h3ad9a5f5),
	.w6(32'h3b8f8924),
	.w7(32'h3b80a4fe),
	.w8(32'hbaa99b25),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a565f03),
	.w1(32'hb9e18ce8),
	.w2(32'h3bf12ef1),
	.w3(32'hba0eb543),
	.w4(32'hbb3a35a8),
	.w5(32'hba883b26),
	.w6(32'h3b88c769),
	.w7(32'h3be3e089),
	.w8(32'hbb9b8141),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a650d88),
	.w1(32'h3b1051a0),
	.w2(32'hbc8feb64),
	.w3(32'hbb3187d5),
	.w4(32'hbb8f008e),
	.w5(32'h3c1ada0f),
	.w6(32'hba83df4f),
	.w7(32'h3d354d2e),
	.w8(32'h3bb8ef75),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306bf5),
	.w1(32'hbac0275d),
	.w2(32'hbc1c5d7e),
	.w3(32'h3a729170),
	.w4(32'hba8dc3af),
	.w5(32'hbc0ed94f),
	.w6(32'h3bf5ccca),
	.w7(32'hba5c8bc1),
	.w8(32'h3b82840f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f8eda),
	.w1(32'h3a79ed57),
	.w2(32'h3c29be8f),
	.w3(32'hbbb74e56),
	.w4(32'hbc96e1e8),
	.w5(32'h3c06342c),
	.w6(32'h3c3f8ab2),
	.w7(32'h3abdaf07),
	.w8(32'hb891a6db),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b939b35),
	.w1(32'hbb816840),
	.w2(32'h3a194813),
	.w3(32'hbace6c6f),
	.w4(32'hbc1173cc),
	.w5(32'hbb00fe4c),
	.w6(32'h3c188103),
	.w7(32'h3ac32471),
	.w8(32'hbc3d9b24),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a2ffd),
	.w1(32'h3afdb3ff),
	.w2(32'h3b9c24c3),
	.w3(32'hbb200494),
	.w4(32'h3b5e2f07),
	.w5(32'h3ca1d047),
	.w6(32'h392690be),
	.w7(32'h3b7ae679),
	.w8(32'hbbb7e8be),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcbfc5),
	.w1(32'hbb0d9a42),
	.w2(32'hbbb2eca6),
	.w3(32'h3c293abb),
	.w4(32'h3c415728),
	.w5(32'h3c20f19e),
	.w6(32'h3b2b8577),
	.w7(32'h3ae73c89),
	.w8(32'hbbd3cfdd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde5b14),
	.w1(32'h3d428a9c),
	.w2(32'h3aa1d7d7),
	.w3(32'hb8b901ea),
	.w4(32'hbb9138ce),
	.w5(32'h3a10e864),
	.w6(32'h3a9bbf5a),
	.w7(32'hbac0402e),
	.w8(32'hbb2ee6d3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdd804),
	.w1(32'h3b46f28e),
	.w2(32'hbc040524),
	.w3(32'h3bc3717f),
	.w4(32'h3b4d1be3),
	.w5(32'hbb69f090),
	.w6(32'hba014a06),
	.w7(32'hbc1b98f7),
	.w8(32'hbce884fe),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5849),
	.w1(32'h3cd9966b),
	.w2(32'hbbf9777e),
	.w3(32'h3c872df5),
	.w4(32'hbb20196b),
	.w5(32'hbbeb7d45),
	.w6(32'hbd1d7636),
	.w7(32'h3bc2157f),
	.w8(32'hba9e3119),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca65dca),
	.w1(32'h3c12a170),
	.w2(32'hbc4d8506),
	.w3(32'hbc8ef021),
	.w4(32'h3befc368),
	.w5(32'hbc9c4cbe),
	.w6(32'hbbff13a9),
	.w7(32'hbb5d1b76),
	.w8(32'hbc108613),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b4aff),
	.w1(32'h3c403327),
	.w2(32'h3cab832b),
	.w3(32'h3c2c2035),
	.w4(32'h3bdf2e3e),
	.w5(32'h3c39cc3f),
	.w6(32'h3c4cb7c6),
	.w7(32'h39db95a1),
	.w8(32'h3b110ff7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d642a),
	.w1(32'hba995de6),
	.w2(32'h3c10b97f),
	.w3(32'hbbd8cb8d),
	.w4(32'hbc44d2a6),
	.w5(32'h3ba4d7b0),
	.w6(32'h3ba4ee6e),
	.w7(32'h3ba2b454),
	.w8(32'h3d0ff69a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba900289),
	.w1(32'h3b642143),
	.w2(32'h3c30ba62),
	.w3(32'hba27d911),
	.w4(32'h3c07ff2e),
	.w5(32'h3bd38561),
	.w6(32'h3c1d520d),
	.w7(32'h3b1ff980),
	.w8(32'h3c759423),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c4254),
	.w1(32'h3b3c0612),
	.w2(32'hbc27cda8),
	.w3(32'h3c1b46d1),
	.w4(32'h3b8ae05d),
	.w5(32'hbb369d85),
	.w6(32'hb97f646c),
	.w7(32'hbb09eef6),
	.w8(32'h3b81f87e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0ac9c),
	.w1(32'h3b23cb65),
	.w2(32'hbbc713b4),
	.w3(32'hba6fa171),
	.w4(32'hbbdec559),
	.w5(32'h3bbe33c2),
	.w6(32'hbbc10d3d),
	.w7(32'h3aa6cf92),
	.w8(32'hbca26771),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea1623),
	.w1(32'h3b808101),
	.w2(32'h3acac607),
	.w3(32'h3afea3e2),
	.w4(32'h3a9c5563),
	.w5(32'h393869f6),
	.w6(32'h3ba4a4c9),
	.w7(32'hbb63ba93),
	.w8(32'hba3667e0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb38cc),
	.w1(32'hbc87c213),
	.w2(32'hbca75d63),
	.w3(32'hbbcbc60f),
	.w4(32'h3a93f423),
	.w5(32'hbc092edd),
	.w6(32'hbbed8f62),
	.w7(32'hbca25e40),
	.w8(32'hbbae7a44),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a546107),
	.w1(32'hbcd4a039),
	.w2(32'h3b018b54),
	.w3(32'hbbf2749a),
	.w4(32'hbb6081f8),
	.w5(32'h3a0fcf1f),
	.w6(32'h3c05bbdf),
	.w7(32'h3bb86260),
	.w8(32'h3b3c8323),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4184c5),
	.w1(32'h3a6289f7),
	.w2(32'hb93a9f00),
	.w3(32'hba1acd58),
	.w4(32'hbb2522f1),
	.w5(32'h3c151663),
	.w6(32'h3c8f38b2),
	.w7(32'hbb890ae5),
	.w8(32'h3ae5a9b4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32a1ec),
	.w1(32'hbb2d7b05),
	.w2(32'hbba3075a),
	.w3(32'h3c0ab25d),
	.w4(32'h3914055c),
	.w5(32'hbc99a181),
	.w6(32'h38234bdf),
	.w7(32'h3a38c071),
	.w8(32'hbb947923),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4469),
	.w1(32'hbc014ffe),
	.w2(32'hbc78e70a),
	.w3(32'h3bb9fb45),
	.w4(32'h3afb50a9),
	.w5(32'hbb972063),
	.w6(32'h3c7429b5),
	.w7(32'h3ba376eb),
	.w8(32'hbc1e158e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af85a43),
	.w1(32'hbbe7c920),
	.w2(32'hbcb4300f),
	.w3(32'hba8f777c),
	.w4(32'h3b6b1d1e),
	.w5(32'hbba86608),
	.w6(32'hbbc45104),
	.w7(32'hbbb651d2),
	.w8(32'h39728872),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28eefa),
	.w1(32'hbaa162fa),
	.w2(32'hbb23851a),
	.w3(32'hbc7f4d0a),
	.w4(32'h3c34ae43),
	.w5(32'hbb780e58),
	.w6(32'h3c0d096b),
	.w7(32'hbb03b270),
	.w8(32'hb99e1515),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919c2b1),
	.w1(32'hbb7e3734),
	.w2(32'hbaad3569),
	.w3(32'hbbd55c2b),
	.w4(32'h3915976c),
	.w5(32'h3a2b9fc5),
	.w6(32'hba66e058),
	.w7(32'hbb947bf4),
	.w8(32'hbacce47a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc254318),
	.w1(32'hbb224142),
	.w2(32'h3aa7b39b),
	.w3(32'hbcef7f95),
	.w4(32'hbb6655a9),
	.w5(32'hbbc13222),
	.w6(32'hbc889c7d),
	.w7(32'h3b6224a7),
	.w8(32'hba05cd73),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128fcc),
	.w1(32'hbb02e5bb),
	.w2(32'hbb308ca1),
	.w3(32'hbbef7a71),
	.w4(32'hbb234971),
	.w5(32'h3bf1ad3b),
	.w6(32'h3b8dd6e9),
	.w7(32'hba46d150),
	.w8(32'hbc16b657),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fb392),
	.w1(32'hbd091f48),
	.w2(32'hbc03bd16),
	.w3(32'h3c424b8c),
	.w4(32'h3c8df639),
	.w5(32'hbb291904),
	.w6(32'hbbba2653),
	.w7(32'hbc2bbc77),
	.w8(32'hbb8678b3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba940fa2),
	.w1(32'h3909eb66),
	.w2(32'hbb057103),
	.w3(32'h3b9968e7),
	.w4(32'h3c0ecf93),
	.w5(32'hbb1cfdbc),
	.w6(32'hba96129e),
	.w7(32'hbb2036cc),
	.w8(32'hbbb32dc3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ec352),
	.w1(32'h3a34ada5),
	.w2(32'hbaa1f666),
	.w3(32'hbb5a9181),
	.w4(32'hbae37e9c),
	.w5(32'hb9c27806),
	.w6(32'h3b144bef),
	.w7(32'hba13c3bc),
	.w8(32'h3aa6b7e3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05f88a),
	.w1(32'hbada5021),
	.w2(32'hbb89ac51),
	.w3(32'hbb093ce8),
	.w4(32'h3b095a76),
	.w5(32'h3a437b34),
	.w6(32'h3c725a37),
	.w7(32'hba85281e),
	.w8(32'hb989972f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8541682),
	.w1(32'h3b0b369a),
	.w2(32'h3b357266),
	.w3(32'hbb74bb1f),
	.w4(32'hba4afb1b),
	.w5(32'h39207af0),
	.w6(32'hb94867d6),
	.w7(32'h3add979c),
	.w8(32'hbbda3c0e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aedaf),
	.w1(32'h3981d860),
	.w2(32'h3b54ab2d),
	.w3(32'hbac348cd),
	.w4(32'h3a6177ca),
	.w5(32'hba77dc06),
	.w6(32'hba9742d4),
	.w7(32'h3a9b0bbe),
	.w8(32'hba7e690f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab44aef),
	.w1(32'h3c2646d6),
	.w2(32'h3a569a83),
	.w3(32'hbb36a095),
	.w4(32'h3a74d15c),
	.w5(32'hbad020cf),
	.w6(32'h3a43daaa),
	.w7(32'hbafbb305),
	.w8(32'hbae4660c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac06953),
	.w1(32'hbbaf9da8),
	.w2(32'hbbe29b6e),
	.w3(32'hb8f3ba7a),
	.w4(32'h3a90a55d),
	.w5(32'hbba47dc0),
	.w6(32'hbb25005e),
	.w7(32'h39fc59c8),
	.w8(32'hbb86aa20),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53d88a),
	.w1(32'hbb4179a2),
	.w2(32'hbc02bf1b),
	.w3(32'hbbc8fccb),
	.w4(32'hbaffa79d),
	.w5(32'hbb87b376),
	.w6(32'hbb89d9ef),
	.w7(32'h3a993800),
	.w8(32'hbb51d300),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d65b3),
	.w1(32'h384881a3),
	.w2(32'h3a8d39dc),
	.w3(32'hbc02e05c),
	.w4(32'hbb1546b3),
	.w5(32'h39fe546b),
	.w6(32'h39dee4eb),
	.w7(32'hb9b08bee),
	.w8(32'h38ec467b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03fe04),
	.w1(32'hbb0097b9),
	.w2(32'h3c63b947),
	.w3(32'h3ac636cd),
	.w4(32'h390eba47),
	.w5(32'h3bffd4b2),
	.w6(32'hba3ac5bc),
	.w7(32'hba107af4),
	.w8(32'h3b1235b1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef2304),
	.w1(32'h394ab2ba),
	.w2(32'h3a551809),
	.w3(32'hbb21b946),
	.w4(32'h3bc24216),
	.w5(32'hb92c812b),
	.w6(32'h3b6058c7),
	.w7(32'hbb7ddd3a),
	.w8(32'hbb256e1f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967f6c9),
	.w1(32'hba186b4d),
	.w2(32'h3a6965b2),
	.w3(32'hbb0ccb5c),
	.w4(32'hbb10cef0),
	.w5(32'h37d605ac),
	.w6(32'h3bf4f06f),
	.w7(32'hbb773f71),
	.w8(32'hba959003),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897c40c),
	.w1(32'hbc5326ef),
	.w2(32'hbcc4c79c),
	.w3(32'h3c901fd7),
	.w4(32'h3c2dcc0d),
	.w5(32'hbbf4bd5e),
	.w6(32'h3b963bf7),
	.w7(32'hb98610e4),
	.w8(32'hbbe17ee5),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79a9db),
	.w1(32'h3c0dfa40),
	.w2(32'hbc316d82),
	.w3(32'h3bd047cb),
	.w4(32'h3abdd81e),
	.w5(32'hbacfc1e9),
	.w6(32'h3ac43340),
	.w7(32'h3a592227),
	.w8(32'hbc06632a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397776),
	.w1(32'hbb4a8ddf),
	.w2(32'hbbc3cc19),
	.w3(32'h3b125f34),
	.w4(32'hbab0ab29),
	.w5(32'hbbc65406),
	.w6(32'hb94f758c),
	.w7(32'h3b0310c3),
	.w8(32'hb9b99e36),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c765fb4),
	.w1(32'h3c3245a9),
	.w2(32'h3c69464f),
	.w3(32'h3b8fab1b),
	.w4(32'hba89e069),
	.w5(32'h3c1f3bd3),
	.w6(32'h3ba90e25),
	.w7(32'h3bb62bef),
	.w8(32'h3d013047),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb261a),
	.w1(32'hbbd1d71b),
	.w2(32'h39bd02f8),
	.w3(32'hba314480),
	.w4(32'h3c0d7023),
	.w5(32'h3afb5597),
	.w6(32'hbae8f7cc),
	.w7(32'hbb852f27),
	.w8(32'h3b585972),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dbae8),
	.w1(32'hba93d042),
	.w2(32'h3a8575b7),
	.w3(32'hbb00ec9f),
	.w4(32'h3aab7293),
	.w5(32'hbaac2d3d),
	.w6(32'h3b0d2945),
	.w7(32'hbb076a20),
	.w8(32'h3aae5fc1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7167a8),
	.w1(32'h392a5e2c),
	.w2(32'hba2c382a),
	.w3(32'hba6fb4a6),
	.w4(32'hbabbba94),
	.w5(32'h3c5f69ef),
	.w6(32'hb9ea40fb),
	.w7(32'hba29651a),
	.w8(32'h3af00d96),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395590a7),
	.w1(32'hb9863a56),
	.w2(32'hbc1ec69d),
	.w3(32'h3a94852c),
	.w4(32'h3a7f3ddd),
	.w5(32'hbb60211b),
	.w6(32'h3c7814f1),
	.w7(32'hb9077e32),
	.w8(32'hbb380a05),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7dae54),
	.w1(32'hba84b6b9),
	.w2(32'h38c95fd3),
	.w3(32'hba4a31e9),
	.w4(32'h3b84f797),
	.w5(32'h3af0485c),
	.w6(32'hbc02cbb7),
	.w7(32'hb8f9bbac),
	.w8(32'h3c5e9f7e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb1bb),
	.w1(32'hbba33db6),
	.w2(32'hbc164b17),
	.w3(32'h3b98e9eb),
	.w4(32'h3ba5eceb),
	.w5(32'hba899979),
	.w6(32'hbafc92b2),
	.w7(32'hbaaf7a3a),
	.w8(32'hbb06fb06),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae08848),
	.w1(32'h3aa519b9),
	.w2(32'hbc0863a1),
	.w3(32'h3b66719f),
	.w4(32'h3b90b558),
	.w5(32'hbb1da452),
	.w6(32'h3ac2f8af),
	.w7(32'hbaa52ea9),
	.w8(32'hb9855f58),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895987),
	.w1(32'h3b7ed610),
	.w2(32'h3bb981ea),
	.w3(32'hbb6a4355),
	.w4(32'hba879e6f),
	.w5(32'hba55cb8c),
	.w6(32'h3a0c6e55),
	.w7(32'hbb4968a4),
	.w8(32'h3bc752ce),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cb728),
	.w1(32'hba9de490),
	.w2(32'hbb9f3e0a),
	.w3(32'hb909cb6c),
	.w4(32'h3aec31eb),
	.w5(32'hbb0422f7),
	.w6(32'h3b534271),
	.w7(32'h39b33c0e),
	.w8(32'hbb6ace73),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82becc),
	.w1(32'hba7e35e7),
	.w2(32'hbc6adde7),
	.w3(32'h3c175b4b),
	.w4(32'h3be195c2),
	.w5(32'hbb9bec0a),
	.w6(32'h3a999e3f),
	.w7(32'hbbff8782),
	.w8(32'hbaacd4a4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953adef),
	.w1(32'hbb2f7417),
	.w2(32'hba82dd52),
	.w3(32'hba848d2c),
	.w4(32'hbb3205d6),
	.w5(32'hba224177),
	.w6(32'hbb1bf256),
	.w7(32'h3abeb614),
	.w8(32'hb92b9d77),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15d5b6),
	.w1(32'hbb3f6101),
	.w2(32'hbba074dd),
	.w3(32'h3b0d45fd),
	.w4(32'h3a8a4994),
	.w5(32'hbbd4d4b2),
	.w6(32'h3b1371f8),
	.w7(32'h3be97beb),
	.w8(32'hbb3fdc22),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99f18f),
	.w1(32'h3b4efdc8),
	.w2(32'hbb4ab357),
	.w3(32'hba0c31bf),
	.w4(32'h3a741348),
	.w5(32'h3ad24f85),
	.w6(32'h39cf2a7e),
	.w7(32'h3b481f5f),
	.w8(32'h392932e0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952b89c),
	.w1(32'h395f9a7a),
	.w2(32'h3a7bcef6),
	.w3(32'h3a22d55d),
	.w4(32'h3a06299e),
	.w5(32'hbb322515),
	.w6(32'hb9679a1a),
	.w7(32'h3b56892a),
	.w8(32'hbbcd0fae),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f55c5),
	.w1(32'h3ab8b8d2),
	.w2(32'h3a62b7fa),
	.w3(32'hbab946fc),
	.w4(32'hbc2c3650),
	.w5(32'h399fa78f),
	.w6(32'h3b6d48e2),
	.w7(32'hbc2db911),
	.w8(32'h3b3a9343),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab749df),
	.w1(32'h39109b9c),
	.w2(32'h3ad19877),
	.w3(32'h3b10b7a2),
	.w4(32'h398f0957),
	.w5(32'h3ab77e95),
	.w6(32'h3a476e6f),
	.w7(32'h3c832d5b),
	.w8(32'hbad11989),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b591f),
	.w1(32'h3c641107),
	.w2(32'hba23f12c),
	.w3(32'hbac9488b),
	.w4(32'h3b0f23cf),
	.w5(32'hba75669e),
	.w6(32'h3c02337c),
	.w7(32'h3a05d5ac),
	.w8(32'hbafeb77b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b025f),
	.w1(32'hbb7f117a),
	.w2(32'h3ab9a72c),
	.w3(32'hba489f34),
	.w4(32'hbaf3b4e3),
	.w5(32'h3b8fe1b9),
	.w6(32'hbae8192b),
	.w7(32'hbc245924),
	.w8(32'hbb416998),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2771d1),
	.w1(32'h3bfb3061),
	.w2(32'h3b4ef56f),
	.w3(32'h3b756386),
	.w4(32'h3b5a074a),
	.w5(32'h3a9a2584),
	.w6(32'h3940ca37),
	.w7(32'h3b0796e6),
	.w8(32'h39a4c8ee),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba651ccb),
	.w1(32'hbb3e6779),
	.w2(32'hbbd2cf46),
	.w3(32'h3b88312e),
	.w4(32'h3b361e5c),
	.w5(32'hbba72659),
	.w6(32'h3b6a6d87),
	.w7(32'h3a92f8b9),
	.w8(32'hbb67f148),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70f3cc),
	.w1(32'hbbb0bb98),
	.w2(32'h3bd9e842),
	.w3(32'hbac57db1),
	.w4(32'hbb87b432),
	.w5(32'hba5152de),
	.w6(32'hbbd44f84),
	.w7(32'h3cf14d5a),
	.w8(32'h3be95ab8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14d434),
	.w1(32'hbb76e25f),
	.w2(32'hbc9c3bc2),
	.w3(32'h3c8e37c2),
	.w4(32'h3bf332ed),
	.w5(32'h3b5f6cd0),
	.w6(32'h3ab048c6),
	.w7(32'h3b88450c),
	.w8(32'hbb0b2de2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad244a),
	.w1(32'hba9c3941),
	.w2(32'h3bfe4461),
	.w3(32'h3a527f0a),
	.w4(32'h3a2e9b10),
	.w5(32'h3b88b858),
	.w6(32'hbb4257c4),
	.w7(32'hb97133f2),
	.w8(32'h3b8b8a46),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a1390),
	.w1(32'h3a3f43b0),
	.w2(32'hbbc19b9f),
	.w3(32'h3bf72484),
	.w4(32'h3a9c26b5),
	.w5(32'hbc4159fa),
	.w6(32'h3b252eda),
	.w7(32'hbbe0ff9a),
	.w8(32'hbb652c06),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced045c),
	.w1(32'h3b15a670),
	.w2(32'hbb002497),
	.w3(32'h3b317b87),
	.w4(32'h3b87b8b8),
	.w5(32'hbabda436),
	.w6(32'h38f6caf4),
	.w7(32'hbb863cfd),
	.w8(32'hbac975e0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0d9e9),
	.w1(32'h3ba65b1d),
	.w2(32'h3c2e53b1),
	.w3(32'h3a61c6cf),
	.w4(32'hba99bee8),
	.w5(32'hbbc7627f),
	.w6(32'h3af5e0a4),
	.w7(32'h3bbbee17),
	.w8(32'h3b55c126),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0bde4),
	.w1(32'h3c2b698e),
	.w2(32'hbb417351),
	.w3(32'h3c04b862),
	.w4(32'h3aa63e7a),
	.w5(32'hbb1b76cf),
	.w6(32'h3995a1e5),
	.w7(32'hb9793e77),
	.w8(32'h379cf67f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54725),
	.w1(32'hbacbe603),
	.w2(32'hbbf3c017),
	.w3(32'h3b49c1bb),
	.w4(32'hba8fe2e4),
	.w5(32'hbb34011a),
	.w6(32'h3bcdbba9),
	.w7(32'hbaac56f6),
	.w8(32'hbb1b28c3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959463c),
	.w1(32'hbb956e53),
	.w2(32'hbc713d74),
	.w3(32'h3c49cf70),
	.w4(32'h3b804e85),
	.w5(32'h3ab5cf5b),
	.w6(32'h39f21d26),
	.w7(32'hbc1f5911),
	.w8(32'hbc929993),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890f883),
	.w1(32'h3bbbe95d),
	.w2(32'hbacbeb89),
	.w3(32'hbaf85ead),
	.w4(32'h3bf133f9),
	.w5(32'h3b16292b),
	.w6(32'hbc1b29a5),
	.w7(32'h3c6ef587),
	.w8(32'hbb5d9983),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73c710),
	.w1(32'h3c331a9c),
	.w2(32'h3c4979df),
	.w3(32'h3b85e5b8),
	.w4(32'h3b3c4097),
	.w5(32'h3c1206ed),
	.w6(32'h3b62626a),
	.w7(32'h3c4a0479),
	.w8(32'h3c4b44db),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874e3b),
	.w1(32'h3b9ebf6d),
	.w2(32'hbaf02d96),
	.w3(32'hba279acd),
	.w4(32'h3a965314),
	.w5(32'h3b5a33f1),
	.w6(32'h39d90858),
	.w7(32'h3b091361),
	.w8(32'h3ac0ac68),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d14aa),
	.w1(32'hbbb4b433),
	.w2(32'h3b83f399),
	.w3(32'h3c642b90),
	.w4(32'h3b97f678),
	.w5(32'h3acaa8b1),
	.w6(32'hbb875d96),
	.w7(32'h3b8964ef),
	.w8(32'h3b1cd453),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba23ae),
	.w1(32'hbb0a08df),
	.w2(32'h3c9295b9),
	.w3(32'h38c3fd43),
	.w4(32'hbb8cbcd6),
	.w5(32'h3a024806),
	.w6(32'h3a0b7064),
	.w7(32'hbbaff8d0),
	.w8(32'hbb1fd99c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc672128),
	.w1(32'h3c862716),
	.w2(32'hbc07868d),
	.w3(32'hbc227b50),
	.w4(32'h3b8e29bb),
	.w5(32'hbba9630b),
	.w6(32'hbc51c4ed),
	.w7(32'hbc098ae4),
	.w8(32'hbba272a8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1afb0a),
	.w1(32'h3beeda1c),
	.w2(32'hba565dc3),
	.w3(32'h3a21a0f5),
	.w4(32'h3ab58d7d),
	.w5(32'hbb73d821),
	.w6(32'hb88a92b2),
	.w7(32'h3c738352),
	.w8(32'hbb78e02f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6a6cb),
	.w1(32'hbb52cad7),
	.w2(32'h3bb4a942),
	.w3(32'hbaf07a41),
	.w4(32'hb7caac27),
	.w5(32'hba241c8b),
	.w6(32'hbb52b9ec),
	.w7(32'h3a8a0a1f),
	.w8(32'h39751247),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e45b2),
	.w1(32'hbadb26b8),
	.w2(32'hba01b809),
	.w3(32'h3a8f0291),
	.w4(32'hbb917908),
	.w5(32'hbacb3285),
	.w6(32'hba092eb9),
	.w7(32'h3a8a8c79),
	.w8(32'hbbdb80ad),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bb31),
	.w1(32'h3b01816a),
	.w2(32'hbc0fa764),
	.w3(32'h3a67ed56),
	.w4(32'h3b6e7109),
	.w5(32'hbb6ceb75),
	.w6(32'hbb0fc462),
	.w7(32'h3a118108),
	.w8(32'hbb1737dd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad9a44),
	.w1(32'h3bc6525b),
	.w2(32'h3c11e6f1),
	.w3(32'hbb12995f),
	.w4(32'hbab3bb12),
	.w5(32'hb8dbe999),
	.w6(32'h3bdd3707),
	.w7(32'h3ad1f690),
	.w8(32'hba82767f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f7603),
	.w1(32'h3bead143),
	.w2(32'h3b05c756),
	.w3(32'hbb38525f),
	.w4(32'hbb7214f9),
	.w5(32'h3b35feb2),
	.w6(32'hbb1c4e86),
	.w7(32'hbc7c1463),
	.w8(32'h3ac93be0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338b0e),
	.w1(32'hba62ab63),
	.w2(32'h3a734ae3),
	.w3(32'hbae07fec),
	.w4(32'hb9aa4c17),
	.w5(32'hb9b43f63),
	.w6(32'h3b41afc5),
	.w7(32'h3aab5bd6),
	.w8(32'h3ace651d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b953ac0),
	.w1(32'h3c5102cc),
	.w2(32'h3b005e47),
	.w3(32'h3c18ff5f),
	.w4(32'h3c02c603),
	.w5(32'hba147ffa),
	.w6(32'hbac28fd1),
	.w7(32'h3b8ab7db),
	.w8(32'h3afb6dfd),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aad6b),
	.w1(32'hb9ca1017),
	.w2(32'hbbedb240),
	.w3(32'h3cc06567),
	.w4(32'hbb0f2c7d),
	.w5(32'hbbb8cc0c),
	.w6(32'hbac2664f),
	.w7(32'hbb9829c4),
	.w8(32'hbb88526d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847f75),
	.w1(32'hbae647e6),
	.w2(32'h3a1020a4),
	.w3(32'h3a3486cb),
	.w4(32'h3b25d8a2),
	.w5(32'hbbf10df6),
	.w6(32'h3b407859),
	.w7(32'h3b7d6a72),
	.w8(32'h3b0bdc82),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaa4ae),
	.w1(32'hbaf1b352),
	.w2(32'hbaf5d38c),
	.w3(32'h3ad4799f),
	.w4(32'h3a795e2c),
	.w5(32'h3a3c28a0),
	.w6(32'hbb4e2b78),
	.w7(32'h3bb17bb7),
	.w8(32'hba167afb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59fa64),
	.w1(32'hbb0fa3a7),
	.w2(32'hbb1886f5),
	.w3(32'h3b06b61b),
	.w4(32'hba66e099),
	.w5(32'hbb3eff88),
	.w6(32'h3c806183),
	.w7(32'hbac7f15f),
	.w8(32'hbbf1f792),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cde697),
	.w1(32'h39381baf),
	.w2(32'hb7939bab),
	.w3(32'h3b36c6af),
	.w4(32'h3aec3ad9),
	.w5(32'hbae0f728),
	.w6(32'hbb64873e),
	.w7(32'h3b42356c),
	.w8(32'hbadb5bf3),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b610),
	.w1(32'hba9bbe67),
	.w2(32'hba8265ff),
	.w3(32'hbaaf1e0f),
	.w4(32'h3b6cd171),
	.w5(32'hba2fbdd4),
	.w6(32'hba0ee043),
	.w7(32'h389e5047),
	.w8(32'h39d191c7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1ab36),
	.w1(32'hba1e95eb),
	.w2(32'h3b55c010),
	.w3(32'hba55e750),
	.w4(32'hbb2d9aff),
	.w5(32'h3a90b7b4),
	.w6(32'h3af4bdb7),
	.w7(32'h3b883a82),
	.w8(32'h398e511c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e32bdb),
	.w1(32'hbbba29e2),
	.w2(32'h3ca468a2),
	.w3(32'hbbf15987),
	.w4(32'hba89ea9d),
	.w5(32'hbb2801ea),
	.w6(32'h3947a24f),
	.w7(32'h3c3a0183),
	.w8(32'h3a696721),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7db5b8),
	.w1(32'h3bf42441),
	.w2(32'hbbae7e0e),
	.w3(32'h3b81fbf8),
	.w4(32'hba9592d6),
	.w5(32'hbbaa09c5),
	.w6(32'h3a25dedd),
	.w7(32'h3b05f728),
	.w8(32'hbb9a764a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d339),
	.w1(32'h3b43d50c),
	.w2(32'h3bf52752),
	.w3(32'h3c445682),
	.w4(32'hbba0d511),
	.w5(32'h3b29ea93),
	.w6(32'hbac520b0),
	.w7(32'h3ae9d962),
	.w8(32'h3bb6a239),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb274c25),
	.w1(32'hbbdc8b30),
	.w2(32'h3a385947),
	.w3(32'hb604c3ce),
	.w4(32'h398c867f),
	.w5(32'h3a1ae7ea),
	.w6(32'hbab82b12),
	.w7(32'hbb3b4ac2),
	.w8(32'hbb6b7754),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b529e19),
	.w1(32'hb9b8128a),
	.w2(32'hb9aa31e0),
	.w3(32'hb9b36215),
	.w4(32'h3b883bbc),
	.w5(32'hbb0a6063),
	.w6(32'h3beef878),
	.w7(32'hbc5b0340),
	.w8(32'h39d8269c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ac588),
	.w1(32'h367b849f),
	.w2(32'hb95c8cd1),
	.w3(32'h3b07972f),
	.w4(32'h38d9cc36),
	.w5(32'hbacc4518),
	.w6(32'h3b579778),
	.w7(32'hb95f229e),
	.w8(32'hbb5b5485),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b289c),
	.w1(32'hba584482),
	.w2(32'h3a234a49),
	.w3(32'hbaa5b8ce),
	.w4(32'h3a4ea364),
	.w5(32'h3d04c48f),
	.w6(32'h3a91f3ca),
	.w7(32'h3ba3e905),
	.w8(32'h3a8b130a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4c7fa),
	.w1(32'h3c9ec02d),
	.w2(32'hbc25e0f2),
	.w3(32'h3c049ac0),
	.w4(32'hbb103416),
	.w5(32'hbb938763),
	.w6(32'hbbcdd54d),
	.w7(32'h3a9352ae),
	.w8(32'h3b03b5a5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad95279),
	.w1(32'hbc00455b),
	.w2(32'hbc495ec1),
	.w3(32'h3be96c01),
	.w4(32'h3a9cb795),
	.w5(32'hbb7b9006),
	.w6(32'h3b3d050e),
	.w7(32'h3b129b2c),
	.w8(32'hba99cfac),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba0f3),
	.w1(32'hba772d9d),
	.w2(32'h3cae4f46),
	.w3(32'h3b35dda0),
	.w4(32'h3b2b7686),
	.w5(32'h3bfc360e),
	.w6(32'h3a989392),
	.w7(32'h39af1fc6),
	.w8(32'hba924f00),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9926315),
	.w1(32'hb9d00a19),
	.w2(32'hbb9483f2),
	.w3(32'h3c968d1c),
	.w4(32'hb999215d),
	.w5(32'hbb913643),
	.w6(32'h3b0be42c),
	.w7(32'hbc026bb9),
	.w8(32'h39bcb0dd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1761a),
	.w1(32'hba847d19),
	.w2(32'h3a4d894f),
	.w3(32'hbc851e29),
	.w4(32'h3a3fed4a),
	.w5(32'h3c74e29e),
	.w6(32'h39b6ec48),
	.w7(32'h3a10fcb0),
	.w8(32'h3ad41e2f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba625fc8),
	.w1(32'hbb85e755),
	.w2(32'hbb889b5f),
	.w3(32'hbc127f28),
	.w4(32'hbae5e922),
	.w5(32'hbb912186),
	.w6(32'hba9a3f56),
	.w7(32'h3ad68e1d),
	.w8(32'hbb8b03c8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00edd2),
	.w1(32'hbb2e4485),
	.w2(32'hbb9fbe02),
	.w3(32'hbad1824c),
	.w4(32'hbb7474ff),
	.w5(32'h3b2489e3),
	.w6(32'h3c045fd9),
	.w7(32'hba2f24cd),
	.w8(32'h3a8fad75),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ae620),
	.w1(32'hbbe52281),
	.w2(32'hbc4aabc5),
	.w3(32'h3c04f824),
	.w4(32'h3c06d1f3),
	.w5(32'hbba100f1),
	.w6(32'h3b036989),
	.w7(32'h3bca52f4),
	.w8(32'hbb74310a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af30f4c),
	.w1(32'h3b8b8acf),
	.w2(32'h3bd5daf3),
	.w3(32'h3a00663a),
	.w4(32'h3924beaa),
	.w5(32'h3b1bd86a),
	.w6(32'h3af74ada),
	.w7(32'h3a965b1c),
	.w8(32'h3b76d042),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34308d),
	.w1(32'hb9b51a46),
	.w2(32'hbba60b43),
	.w3(32'h3b6c1e4c),
	.w4(32'hbba77765),
	.w5(32'hb9c6fc00),
	.w6(32'h3a202a2b),
	.w7(32'hbc7c71da),
	.w8(32'h3ac07e8e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab603b3),
	.w1(32'hbbfb412f),
	.w2(32'hbbeca6af),
	.w3(32'h3b3e3a31),
	.w4(32'h3b0b233f),
	.w5(32'hbba9999a),
	.w6(32'hba935ac7),
	.w7(32'h3b884f77),
	.w8(32'hbaca5cb6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb258ef),
	.w1(32'h3bad8194),
	.w2(32'h3b692c05),
	.w3(32'h3ab63d29),
	.w4(32'h3c4fc7a4),
	.w5(32'h3bb5d27a),
	.w6(32'h3b84f8b4),
	.w7(32'h3bb217e7),
	.w8(32'hb89df0f6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed6771),
	.w1(32'hbae8323e),
	.w2(32'hbb87e718),
	.w3(32'h3b4db436),
	.w4(32'h3aa3c00e),
	.w5(32'hbbde3557),
	.w6(32'h3ba7fe9d),
	.w7(32'hbb0e5a39),
	.w8(32'hbb7efe80),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac51b1f),
	.w1(32'hba30c901),
	.w2(32'h3b02a368),
	.w3(32'hb9f09db4),
	.w4(32'hba8bfc0c),
	.w5(32'hbbcf6c63),
	.w6(32'hbaf16938),
	.w7(32'h3b1883c9),
	.w8(32'h38d6a073),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c625643),
	.w1(32'h3c3bdb8b),
	.w2(32'h3c3e41ed),
	.w3(32'h3aeb8e4e),
	.w4(32'hbb3a3756),
	.w5(32'h3b91ed3f),
	.w6(32'h3c7d3b1c),
	.w7(32'h3c7391f3),
	.w8(32'h3bdf616f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77b566),
	.w1(32'hbaaf8c56),
	.w2(32'hbab1aab0),
	.w3(32'hb7e3381c),
	.w4(32'hbb18ea52),
	.w5(32'h39b8e474),
	.w6(32'h3b1ceb4a),
	.w7(32'hbac5b2d3),
	.w8(32'h3a82300f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5746ea),
	.w1(32'hbbb3bb39),
	.w2(32'hbb7a5432),
	.w3(32'hbaa52c05),
	.w4(32'hbb0ca138),
	.w5(32'hbba9a0d4),
	.w6(32'hbc06631e),
	.w7(32'hbab00b43),
	.w8(32'h3a107b5e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a615984),
	.w1(32'h3a55c8e4),
	.w2(32'h3b967a05),
	.w3(32'hbad5fde4),
	.w4(32'h38a48381),
	.w5(32'hbacb111f),
	.w6(32'hbab7e6d1),
	.w7(32'h3ab04e53),
	.w8(32'h3bc3cacb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08c87d),
	.w1(32'h3c207590),
	.w2(32'hbac709bd),
	.w3(32'h3b15cecc),
	.w4(32'hbab7ec0d),
	.w5(32'h3b446675),
	.w6(32'h3a4f34de),
	.w7(32'hba821ace),
	.w8(32'hbabb16b2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63f811),
	.w1(32'h3ae70cbe),
	.w2(32'h3bd44b8d),
	.w3(32'hbb500f9e),
	.w4(32'h3bdd63dd),
	.w5(32'h3b2759c2),
	.w6(32'h3b954cfe),
	.w7(32'hba461255),
	.w8(32'h3b23299a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5a9cd),
	.w1(32'h3a27a880),
	.w2(32'hbb300fad),
	.w3(32'h3ba4b81f),
	.w4(32'hbb800671),
	.w5(32'hb986c21b),
	.w6(32'hba8d82c2),
	.w7(32'h3a080450),
	.w8(32'h3aed63b3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad082fa),
	.w1(32'h3b4a42ab),
	.w2(32'hbbc6a79c),
	.w3(32'hbb3f53ec),
	.w4(32'hbb2ad23b),
	.w5(32'h3ab5cc33),
	.w6(32'h3b1d3810),
	.w7(32'hbb1c9cfe),
	.w8(32'hbb0e5816),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dd295),
	.w1(32'hbb7ca678),
	.w2(32'hbc0d1dae),
	.w3(32'h3c4ed817),
	.w4(32'h3b41fc3a),
	.w5(32'hbb26689e),
	.w6(32'h3b32708e),
	.w7(32'h3b3f3605),
	.w8(32'hbb649fe2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39fe3e),
	.w1(32'h3b34b398),
	.w2(32'hbb09eb7d),
	.w3(32'h3af129e8),
	.w4(32'hbb486640),
	.w5(32'hbb5a3603),
	.w6(32'hbb1a2d87),
	.w7(32'h3c23f61d),
	.w8(32'hbb4963dc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f2d56),
	.w1(32'h39a1f499),
	.w2(32'hbc0a0f1a),
	.w3(32'h3bf6dd58),
	.w4(32'h3b1a9afe),
	.w5(32'hbc35670f),
	.w6(32'hbc0938ad),
	.w7(32'h3aeb3bf5),
	.w8(32'h3b2900c6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dbc4e),
	.w1(32'h3c0763d5),
	.w2(32'h3bcc3801),
	.w3(32'hbb8361ef),
	.w4(32'hbb088170),
	.w5(32'hba5356e1),
	.w6(32'h3b847bde),
	.w7(32'hbabd83d9),
	.w8(32'h3a9de50e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802361d),
	.w1(32'h3b4fc4d2),
	.w2(32'hbbb59b6b),
	.w3(32'h3a544bcc),
	.w4(32'h3b6ffc83),
	.w5(32'hbac008e8),
	.w6(32'h3ad817e7),
	.w7(32'h3a93059e),
	.w8(32'hbbd76610),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398df86b),
	.w1(32'h3ba3ad03),
	.w2(32'h39f4f6b0),
	.w3(32'hbb7e6d80),
	.w4(32'hbb1c3c12),
	.w5(32'h39993543),
	.w6(32'hbb2317c8),
	.w7(32'h3ae65b3e),
	.w8(32'hbae14dc7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e17bf),
	.w1(32'h3b847c70),
	.w2(32'h3c3498a4),
	.w3(32'h3b06a37b),
	.w4(32'hbb3c9992),
	.w5(32'h3c013329),
	.w6(32'h3d02065c),
	.w7(32'hbb8e42ad),
	.w8(32'h392ec9ae),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a9d4),
	.w1(32'h3ad91afa),
	.w2(32'h3b3d3e66),
	.w3(32'h3babe075),
	.w4(32'hbaf39ea1),
	.w5(32'h3b97f348),
	.w6(32'h3c3e4538),
	.w7(32'h3a4486fc),
	.w8(32'h3b5627c6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90be15),
	.w1(32'h3c27e87c),
	.w2(32'h3b548398),
	.w3(32'h3a0dafbd),
	.w4(32'hbb6bd09a),
	.w5(32'h3af7a6ce),
	.w6(32'hb9982f2a),
	.w7(32'h3b3bbea0),
	.w8(32'h3af30af4),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a23fa),
	.w1(32'hbb5abb1e),
	.w2(32'hbb1e8ff7),
	.w3(32'h3c1abf8c),
	.w4(32'h3b0407df),
	.w5(32'hbb9adb16),
	.w6(32'hbaf9cba8),
	.w7(32'h3c46c934),
	.w8(32'hbaf0b2f3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc88d),
	.w1(32'h39abe416),
	.w2(32'hbae19660),
	.w3(32'hba9e0bdd),
	.w4(32'h3b3af43d),
	.w5(32'h398baea3),
	.w6(32'h3a18063e),
	.w7(32'hbb8f11eb),
	.w8(32'h3aa043f6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f673d),
	.w1(32'hb797fbab),
	.w2(32'hbbb14d52),
	.w3(32'h3bbc5b1a),
	.w4(32'h3b06aafa),
	.w5(32'hbb9e8017),
	.w6(32'h3c46cbde),
	.w7(32'hba811c0e),
	.w8(32'hbaab52c1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc723f1),
	.w1(32'hba86b77f),
	.w2(32'hba94b59a),
	.w3(32'h3b074442),
	.w4(32'h3b2364cf),
	.w5(32'h3a3e585f),
	.w6(32'h3c12e947),
	.w7(32'hbb50d420),
	.w8(32'hba9034f3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdef5b5),
	.w1(32'h3b862e0e),
	.w2(32'h3c1c9519),
	.w3(32'hbb293b0e),
	.w4(32'h3b0171a4),
	.w5(32'h3b1533a8),
	.w6(32'h3b2a8d59),
	.w7(32'hbadd426c),
	.w8(32'hbb171462),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b921bb7),
	.w1(32'hb81232fe),
	.w2(32'h3a88ff1a),
	.w3(32'h3b245370),
	.w4(32'hba682133),
	.w5(32'hb8547d84),
	.w6(32'h3b85356c),
	.w7(32'hbabe56d6),
	.w8(32'hbaed5d8e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0630d5),
	.w1(32'h3b056863),
	.w2(32'hbad8037c),
	.w3(32'h3b8e2058),
	.w4(32'h39d4d56c),
	.w5(32'hbb7e738a),
	.w6(32'h3b4f9bf9),
	.w7(32'h3a1cf835),
	.w8(32'hbc715ea8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20326a),
	.w1(32'hbacc54ef),
	.w2(32'h3a1d91b2),
	.w3(32'hbb4d4cfe),
	.w4(32'h3a0fc9b3),
	.w5(32'h3ae3a38f),
	.w6(32'h38f37b5f),
	.w7(32'h3b86f5c9),
	.w8(32'hbab0bb77),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfc82),
	.w1(32'hbb28b37f),
	.w2(32'h3a762fda),
	.w3(32'hbb05ec1b),
	.w4(32'h3a0b9333),
	.w5(32'hbb3e1f71),
	.w6(32'hba6e264c),
	.w7(32'hbab48020),
	.w8(32'h3bfae910),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a304883),
	.w1(32'hba82104b),
	.w2(32'h3b21f6c6),
	.w3(32'hbbf69f6a),
	.w4(32'hbaeca389),
	.w5(32'h3a8f9c66),
	.w6(32'hbaf3efe7),
	.w7(32'hbb36fc1c),
	.w8(32'h3a74d249),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92399cc),
	.w1(32'h3ba6b2ce),
	.w2(32'hbb56d5fb),
	.w3(32'h3bb4f69b),
	.w4(32'h3bd1e5d1),
	.w5(32'hb9159e29),
	.w6(32'h3913a210),
	.w7(32'h3a933c8e),
	.w8(32'hba9ebd63),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6b15),
	.w1(32'h3b6ee6e5),
	.w2(32'h3b845791),
	.w3(32'h3b4fd9ae),
	.w4(32'hb99f20ab),
	.w5(32'h3d282cac),
	.w6(32'hbb8b38aa),
	.w7(32'h3b67452b),
	.w8(32'hbb68cb2e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb91af1),
	.w1(32'h3be31481),
	.w2(32'h3bab463e),
	.w3(32'hbb157d46),
	.w4(32'hbbe6fe7b),
	.w5(32'hbb70ede4),
	.w6(32'hbb1cf38b),
	.w7(32'hba9588ab),
	.w8(32'h3d040c61),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1904b9),
	.w1(32'hb8ae79d7),
	.w2(32'h3ca5c3f9),
	.w3(32'h39933cf6),
	.w4(32'h3c0d380e),
	.w5(32'hbb60c281),
	.w6(32'hbae3263f),
	.w7(32'hbafcd0dd),
	.w8(32'hbb94a438),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac9e0c),
	.w1(32'hbc1451a2),
	.w2(32'hbbe95476),
	.w3(32'hbc17e5d6),
	.w4(32'hbb3abe72),
	.w5(32'h3a8ee916),
	.w6(32'hbc0bb3ca),
	.w7(32'hbb1e6b70),
	.w8(32'hbc30f844),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93370f),
	.w1(32'hbb9e5dd9),
	.w2(32'hba8b2c6c),
	.w3(32'h3c647007),
	.w4(32'h3c35fa12),
	.w5(32'hb9b438f1),
	.w6(32'h3b5c5cfc),
	.w7(32'hbb7b23da),
	.w8(32'hbb7127c5),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde3409),
	.w1(32'hbc151920),
	.w2(32'hbbb06e07),
	.w3(32'hbb5d5d24),
	.w4(32'hbb2a3130),
	.w5(32'hbc0a1092),
	.w6(32'hbb6d3b64),
	.w7(32'h3bd6034d),
	.w8(32'h3a0ac405),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80401e),
	.w1(32'hba2ef872),
	.w2(32'h3ba7ccfb),
	.w3(32'h39828882),
	.w4(32'h3a5a75ec),
	.w5(32'hba8fd06a),
	.w6(32'hbb9d1a59),
	.w7(32'hbcbace6c),
	.w8(32'hbc24c190),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad06372),
	.w1(32'h3a392ef0),
	.w2(32'hbaeda85b),
	.w3(32'hb9937b38),
	.w4(32'hb886d3da),
	.w5(32'hbb233ca7),
	.w6(32'h3b4efa40),
	.w7(32'hbb96ba56),
	.w8(32'h3b576c77),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fd0bc),
	.w1(32'hbba3fea4),
	.w2(32'h3c00ab03),
	.w3(32'h3c0e8b1d),
	.w4(32'hbd207b19),
	.w5(32'hbbdc42e1),
	.w6(32'h3b8f9981),
	.w7(32'h3c4d90b3),
	.w8(32'hbc4a0816),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd30fb),
	.w1(32'h3c71d3f0),
	.w2(32'h3c0d7da9),
	.w3(32'h38021256),
	.w4(32'hba3aa46d),
	.w5(32'h3be4ca84),
	.w6(32'h3a114b8d),
	.w7(32'hba1af0c5),
	.w8(32'hbb8bfee3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc94d9e),
	.w1(32'h3c6d6823),
	.w2(32'h3ab910bf),
	.w3(32'hb8a8d063),
	.w4(32'hbba03e3e),
	.w5(32'h3b9e0435),
	.w6(32'h3ab648f6),
	.w7(32'hb82fd92e),
	.w8(32'hbb37a494),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b38f62),
	.w1(32'hbb9b3a00),
	.w2(32'hbba0eaec),
	.w3(32'h3b205f9f),
	.w4(32'hbc10199d),
	.w5(32'h3b0aede7),
	.w6(32'h3d0d9e1c),
	.w7(32'h3bffcc78),
	.w8(32'h3b336761),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db6d2),
	.w1(32'hbadd580f),
	.w2(32'h3c9c15ef),
	.w3(32'hb85dfcf6),
	.w4(32'h3c8f2a47),
	.w5(32'h3b764ddc),
	.w6(32'hbac73e65),
	.w7(32'hbb9d97a2),
	.w8(32'h3a168244),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aee372),
	.w1(32'hbbfbc5e2),
	.w2(32'hbb5060e9),
	.w3(32'h3c26b8f4),
	.w4(32'hb98e0e15),
	.w5(32'hba8649b9),
	.w6(32'hb6fe38ba),
	.w7(32'h3aff96c2),
	.w8(32'h3aefa3ea),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4147c0),
	.w1(32'hba282c9a),
	.w2(32'hbd124803),
	.w3(32'hbb835cb5),
	.w4(32'hb9e4a828),
	.w5(32'hbbac3074),
	.w6(32'h3b1cd2df),
	.w7(32'hba8102a5),
	.w8(32'h3c2a0375),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c5076),
	.w1(32'hbb0d105a),
	.w2(32'hbb3fc426),
	.w3(32'h3c1cd112),
	.w4(32'hba4087b4),
	.w5(32'hbc05dfe9),
	.w6(32'hbc8e4e7d),
	.w7(32'hbb82e566),
	.w8(32'h39f0b8bb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23bca2),
	.w1(32'h3ade70ea),
	.w2(32'hbbf9c082),
	.w3(32'hbbb16a9f),
	.w4(32'h391f35d4),
	.w5(32'hbd347b1b),
	.w6(32'hbad84568),
	.w7(32'hbc5bcdfd),
	.w8(32'hbbd7fca1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fca4c),
	.w1(32'h3b0575fc),
	.w2(32'hb8e7dcec),
	.w3(32'hba0b4186),
	.w4(32'hb9c64370),
	.w5(32'h3baa1fd7),
	.w6(32'h3a8a7735),
	.w7(32'hbca2c580),
	.w8(32'hba9b98a9),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc67ffd),
	.w1(32'hbbeb8e62),
	.w2(32'hbc77d806),
	.w3(32'h3b87e8e7),
	.w4(32'h3cb885d9),
	.w5(32'hbc36960d),
	.w6(32'hbb50ce68),
	.w7(32'hbb040fdc),
	.w8(32'hbbac865d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cabd6cb),
	.w1(32'h3c82dced),
	.w2(32'h3c1c9aea),
	.w3(32'h3bbd7128),
	.w4(32'h3b96f293),
	.w5(32'hbac7d355),
	.w6(32'hbbd0b64b),
	.w7(32'hbb8dcb46),
	.w8(32'hbaf2d113),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd89d45),
	.w1(32'hbb9fc97d),
	.w2(32'h3c0d50f0),
	.w3(32'h3b73fce5),
	.w4(32'hbbe3f8dc),
	.w5(32'hb9370d80),
	.w6(32'hbb00dc81),
	.w7(32'hbb330df5),
	.w8(32'hbb5cbe21),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab540c1),
	.w1(32'h3b87baab),
	.w2(32'h3ad33fc3),
	.w3(32'h3bfae814),
	.w4(32'h3b8980d3),
	.w5(32'hbbd29fd2),
	.w6(32'hbb438f37),
	.w7(32'hbb9bf2f4),
	.w8(32'hbd04c3ac),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba859e46),
	.w1(32'h3b1fb473),
	.w2(32'h3ced2ed0),
	.w3(32'h3b00d2ba),
	.w4(32'h3965ce37),
	.w5(32'h38802db6),
	.w6(32'hbba69e44),
	.w7(32'hbb1d3b99),
	.w8(32'hba140c89),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc69238),
	.w1(32'h3afc62eb),
	.w2(32'hbb24d012),
	.w3(32'h3b32e75f),
	.w4(32'hbaabc064),
	.w5(32'h3b410a52),
	.w6(32'h39b03c16),
	.w7(32'hbb74ef43),
	.w8(32'h3aea4256),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a358b),
	.w1(32'h3c7471d6),
	.w2(32'hba03b26c),
	.w3(32'h3acdc28f),
	.w4(32'hbcbfd9a5),
	.w5(32'hbbffe2ca),
	.w6(32'h3b87223a),
	.w7(32'h391e149b),
	.w8(32'hbbe5b7cd),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b3ef),
	.w1(32'h3b96b43b),
	.w2(32'hbb022475),
	.w3(32'hba7354ff),
	.w4(32'hbac5e85c),
	.w5(32'hb9da4657),
	.w6(32'hb96ab1b0),
	.w7(32'hba5d6e1e),
	.w8(32'hbb429de8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d54e4),
	.w1(32'h3c437b38),
	.w2(32'h3c85316d),
	.w3(32'hbb9a6e71),
	.w4(32'hbb3959e9),
	.w5(32'hbba6b6f3),
	.w6(32'h3b89ad01),
	.w7(32'hbc1a8f99),
	.w8(32'h3b74254e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0b225),
	.w1(32'h3b57a6a2),
	.w2(32'h3a3ee31b),
	.w3(32'h3b09505e),
	.w4(32'h3b313c73),
	.w5(32'hbc04b576),
	.w6(32'h3b86d7c3),
	.w7(32'hbb73b69a),
	.w8(32'h3b08d5d5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134de0),
	.w1(32'h3af5be95),
	.w2(32'hbc1078e3),
	.w3(32'h3ab6e267),
	.w4(32'h3be1df92),
	.w5(32'hbb2e31a7),
	.w6(32'h39783922),
	.w7(32'hba8f6b34),
	.w8(32'hbb4cafeb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed000e),
	.w1(32'hbb10dbfa),
	.w2(32'h3a90c1a0),
	.w3(32'hbb80afb8),
	.w4(32'hbc886794),
	.w5(32'hba71c2b1),
	.w6(32'hbc989138),
	.w7(32'h3a6dabf9),
	.w8(32'hbb57e4ed),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24054d),
	.w1(32'h3ced8166),
	.w2(32'hbac1d6c8),
	.w3(32'hbb218ccd),
	.w4(32'hbb7729b3),
	.w5(32'hbb30ba69),
	.w6(32'hbac952b8),
	.w7(32'hb9a07ce9),
	.w8(32'h3b54d358),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0702),
	.w1(32'hbc0928ee),
	.w2(32'hbacbe5b8),
	.w3(32'h3cb6286b),
	.w4(32'h3a3d2436),
	.w5(32'hb9ba125c),
	.w6(32'h3b28fdba),
	.w7(32'hbb03de68),
	.w8(32'h3a430936),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fa7438),
	.w1(32'hbb50f54d),
	.w2(32'h3a94a2ef),
	.w3(32'h3b9c58c2),
	.w4(32'h39fff6c5),
	.w5(32'hbbc49cd6),
	.w6(32'hbaa84bdc),
	.w7(32'h3a4d3719),
	.w8(32'hbb4f14a5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace27b3),
	.w1(32'h3a80c77f),
	.w2(32'hbb903a37),
	.w3(32'h3bf948e7),
	.w4(32'hbb318dd2),
	.w5(32'hbb2f2b61),
	.w6(32'h3b9dd9b1),
	.w7(32'h3ac073e5),
	.w8(32'hb9f33208),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f00f3),
	.w1(32'h3a4e533c),
	.w2(32'h3b665bc3),
	.w3(32'h3b4e4b96),
	.w4(32'h3b61e30e),
	.w5(32'h3a8fc571),
	.w6(32'h399a21a2),
	.w7(32'hba8d1e94),
	.w8(32'h3a61b2b3),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf4676),
	.w1(32'h3c8ca956),
	.w2(32'hbac752ee),
	.w3(32'hb9968bd8),
	.w4(32'hba4cfb79),
	.w5(32'h3b6b739a),
	.w6(32'h3a53d43e),
	.w7(32'h3ba74901),
	.w8(32'hbb73d17f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b853),
	.w1(32'h3aa0cf48),
	.w2(32'hba437bbd),
	.w3(32'hbaae6636),
	.w4(32'h3bd7a632),
	.w5(32'h3b48fb9e),
	.w6(32'hba1f2c75),
	.w7(32'hbc241d5b),
	.w8(32'h3cb1d1d4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b7c6b),
	.w1(32'hbb04a6f8),
	.w2(32'hbb50ee88),
	.w3(32'hbb2464f3),
	.w4(32'h3bbba284),
	.w5(32'h3c294c14),
	.w6(32'hbb067e6d),
	.w7(32'hbb10e4f8),
	.w8(32'h3b8ef2cf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f81e67),
	.w1(32'hbafca150),
	.w2(32'hbb8beac9),
	.w3(32'h3c091746),
	.w4(32'hbad7de4a),
	.w5(32'h3c903ea0),
	.w6(32'h3b8641d3),
	.w7(32'hb8fc6843),
	.w8(32'h3b08ac97),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac62148),
	.w1(32'hbb1d6dc1),
	.w2(32'hbc53c000),
	.w3(32'hbc09ccfa),
	.w4(32'h3a566e8b),
	.w5(32'hbb9a0304),
	.w6(32'h39f071ee),
	.w7(32'hb835f489),
	.w8(32'h3af18a89),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8792a5),
	.w1(32'hb8d309e4),
	.w2(32'h39e32e49),
	.w3(32'hbbd782b0),
	.w4(32'hb9a2c6c2),
	.w5(32'h3a5180f3),
	.w6(32'h3bd64ea7),
	.w7(32'hbcabcab0),
	.w8(32'h3c9ff37e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e74ec),
	.w1(32'h39fc94ee),
	.w2(32'h38284608),
	.w3(32'h3cd52148),
	.w4(32'hba85b35f),
	.w5(32'hbc2104f9),
	.w6(32'h3ae958fc),
	.w7(32'hbc60c278),
	.w8(32'h389933f6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29fe89),
	.w1(32'hba8d9b3a),
	.w2(32'hbb29fcb5),
	.w3(32'hb9a3515c),
	.w4(32'h3a8607b0),
	.w5(32'hbb680857),
	.w6(32'h3bfefaef),
	.w7(32'h3b05a75a),
	.w8(32'hbb9b6cb7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e119b),
	.w1(32'hbc1256aa),
	.w2(32'hbceea393),
	.w3(32'h3b685d7c),
	.w4(32'hbbfc8371),
	.w5(32'hbbc92443),
	.w6(32'hba9ff61a),
	.w7(32'h3a61fc12),
	.w8(32'hba55a817),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f3373),
	.w1(32'h3b18b17d),
	.w2(32'hbb977dfc),
	.w3(32'hbbc65b0c),
	.w4(32'h3a6f3244),
	.w5(32'h3ab6c077),
	.w6(32'h3b65a554),
	.w7(32'h399b7b32),
	.w8(32'h3b446f9d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69d872),
	.w1(32'hbb11d6e7),
	.w2(32'hbbb32d52),
	.w3(32'h3c781dea),
	.w4(32'h3c3a70f4),
	.w5(32'hb9c1431e),
	.w6(32'h3c387fbc),
	.w7(32'hbae6f729),
	.w8(32'hbc200cdb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42caef),
	.w1(32'h3a6f720f),
	.w2(32'h3b03b286),
	.w3(32'h3b233240),
	.w4(32'hbbd2436e),
	.w5(32'hbb406352),
	.w6(32'h3b2bdd1c),
	.w7(32'hb9f17a2a),
	.w8(32'hbb8cc498),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9800329),
	.w1(32'h39c52033),
	.w2(32'h3b812194),
	.w3(32'h3995c8d0),
	.w4(32'h3c72237b),
	.w5(32'h3cb65b43),
	.w6(32'h3b0bd75a),
	.w7(32'h3b3165c2),
	.w8(32'hb91782de),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaedd2b),
	.w1(32'h3c54709d),
	.w2(32'h3aec6142),
	.w3(32'hbb64177b),
	.w4(32'h3d5b42c5),
	.w5(32'hbc0777e7),
	.w6(32'hbbb08c83),
	.w7(32'h3c1da037),
	.w8(32'hbc5e2d44),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a243515),
	.w1(32'h3b5ef405),
	.w2(32'hbc1cb11c),
	.w3(32'h3d21ee8a),
	.w4(32'h3b2bdaed),
	.w5(32'hbbd9eb68),
	.w6(32'hbb852d30),
	.w7(32'hbc36ca4c),
	.w8(32'hbb651ca9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45f8e9),
	.w1(32'h3c328987),
	.w2(32'hbb8758ef),
	.w3(32'h3c032cb6),
	.w4(32'h3b94c972),
	.w5(32'hbc0d0c1c),
	.w6(32'hbb73eea1),
	.w7(32'h3b498cfa),
	.w8(32'hbba7eba2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17568c),
	.w1(32'h3ba85be5),
	.w2(32'h3be63118),
	.w3(32'hbb99eb91),
	.w4(32'h3bb7b066),
	.w5(32'h3b2cd07f),
	.w6(32'h3a9527d9),
	.w7(32'h3b47ceeb),
	.w8(32'h3b8dc01f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d755),
	.w1(32'h3a305ad4),
	.w2(32'h3b18f220),
	.w3(32'hbb5cfa3a),
	.w4(32'hbb2d56a7),
	.w5(32'h3c113eeb),
	.w6(32'h3b8650ab),
	.w7(32'hbaa80142),
	.w8(32'hbba629d8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67c6e6),
	.w1(32'hb99de814),
	.w2(32'hbc043a43),
	.w3(32'hba77fbe9),
	.w4(32'h3bd1e131),
	.w5(32'h3a84ad67),
	.w6(32'hb98ce73f),
	.w7(32'hbab7c140),
	.w8(32'hbaf3254c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58d7ee),
	.w1(32'h3b6b8806),
	.w2(32'h3a84f855),
	.w3(32'h3afbc793),
	.w4(32'hbac1ca73),
	.w5(32'h3b47234f),
	.w6(32'h3b6cbe5a),
	.w7(32'hbb4f29a4),
	.w8(32'hbac5967c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54932),
	.w1(32'hbca8d424),
	.w2(32'h3ababe42),
	.w3(32'h3c495f13),
	.w4(32'hbb3cca19),
	.w5(32'h3b7ca166),
	.w6(32'hbb2bdd55),
	.w7(32'h3cacad31),
	.w8(32'hbb316729),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae371da),
	.w1(32'h3bb12e65),
	.w2(32'h3af7edc6),
	.w3(32'hba02d90d),
	.w4(32'hbb1715c8),
	.w5(32'h3bcd5bad),
	.w6(32'h38406858),
	.w7(32'hba554ee1),
	.w8(32'hba5aedd4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f10a4),
	.w1(32'hbb487e1c),
	.w2(32'h3add4568),
	.w3(32'h3bccddd5),
	.w4(32'h3c16944d),
	.w5(32'hbbe8ae45),
	.w6(32'h3baed818),
	.w7(32'hbabf412b),
	.w8(32'h3c41c66a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd8b38),
	.w1(32'hb9e30a4c),
	.w2(32'hbb6f3a32),
	.w3(32'h3974ba6d),
	.w4(32'h3a3785f6),
	.w5(32'h3bac4536),
	.w6(32'h3c1f5bf1),
	.w7(32'hb9dafa10),
	.w8(32'hbbbc1f12),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7945),
	.w1(32'h39f64b15),
	.w2(32'hbb708f72),
	.w3(32'hbc3f3903),
	.w4(32'hbaab0c39),
	.w5(32'hbaf5043e),
	.w6(32'h3bae657a),
	.w7(32'hbc0ba636),
	.w8(32'h39ed3f8e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab1a00),
	.w1(32'hb903a3f8),
	.w2(32'h3cd406f6),
	.w3(32'hbb7741db),
	.w4(32'h3b8731ef),
	.w5(32'hbb3e8473),
	.w6(32'hba885c37),
	.w7(32'h3a78f499),
	.w8(32'h3b4fc97c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2e043),
	.w1(32'h3b339784),
	.w2(32'hbcaf51b4),
	.w3(32'h3bd16a92),
	.w4(32'h3c2468a0),
	.w5(32'hbb3ee143),
	.w6(32'hbbd9082d),
	.w7(32'h3aa66472),
	.w8(32'hbc31e802),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb534952),
	.w1(32'hbb2f450b),
	.w2(32'hbb8ef70c),
	.w3(32'hbac5e618),
	.w4(32'h3a9d4b06),
	.w5(32'hbb34c55a),
	.w6(32'hbad81fdf),
	.w7(32'hbc1f0f8d),
	.w8(32'hbb9cdab8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e3d3f),
	.w1(32'hb9e6076f),
	.w2(32'hba4a71e5),
	.w3(32'h3aed7f63),
	.w4(32'h3c1df1a8),
	.w5(32'h3c3cd97f),
	.w6(32'hbbad3c4f),
	.w7(32'hbb20ce40),
	.w8(32'h3c513c83),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50166e),
	.w1(32'hbc677bac),
	.w2(32'hbc30cc5c),
	.w3(32'h3bfdac20),
	.w4(32'hbb5d2ef0),
	.w5(32'hbb2efbff),
	.w6(32'hba99fa98),
	.w7(32'h3b5cbef1),
	.w8(32'hba9fc13b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ca64f),
	.w1(32'hbb17ff0a),
	.w2(32'hb9a581a4),
	.w3(32'h3a650d3c),
	.w4(32'h3c1b1151),
	.w5(32'h3c20605a),
	.w6(32'hbc0537a9),
	.w7(32'h3c8bc925),
	.w8(32'h3c1950f4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b4f06),
	.w1(32'hba0f5826),
	.w2(32'h3b261f9f),
	.w3(32'h3ba07d91),
	.w4(32'hbb9aa17a),
	.w5(32'hbb00b49b),
	.w6(32'h3c8f9ad2),
	.w7(32'hbace02ff),
	.w8(32'h3bccd58f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855ed4),
	.w1(32'hbab38159),
	.w2(32'hbb1827fb),
	.w3(32'h3a40a7d8),
	.w4(32'h38066e06),
	.w5(32'hbc47b1ee),
	.w6(32'h3c0fb511),
	.w7(32'hba4e1d19),
	.w8(32'hb73a2f98),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f2b57),
	.w1(32'hb886d604),
	.w2(32'h3bc29a8b),
	.w3(32'h3bbde6f7),
	.w4(32'h3bd268cf),
	.w5(32'h39cc422a),
	.w6(32'h3990d743),
	.w7(32'hbb97a204),
	.w8(32'hbad6172b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6a1be),
	.w1(32'h381cc363),
	.w2(32'h3b9afa4e),
	.w3(32'h3a33dd86),
	.w4(32'hbad2d8b2),
	.w5(32'h3ba4ab0d),
	.w6(32'h3b38c9c3),
	.w7(32'h3a6475da),
	.w8(32'h3b961cc1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08b59c),
	.w1(32'hbc282a1d),
	.w2(32'hbc59f3ed),
	.w3(32'h3bbe6ecf),
	.w4(32'hba9b9329),
	.w5(32'hbc12cf4b),
	.w6(32'h3b755ad7),
	.w7(32'h3c2f648b),
	.w8(32'hbb8f5cec),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb266b8f),
	.w1(32'hbc398f32),
	.w2(32'hbc032f5d),
	.w3(32'hbbaf488c),
	.w4(32'hba19d08b),
	.w5(32'h3a697f1b),
	.w6(32'h3a991900),
	.w7(32'h3c2efa8e),
	.w8(32'hbb898871),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfed45),
	.w1(32'hbbc99886),
	.w2(32'hbc0d4f86),
	.w3(32'h3b93cbcb),
	.w4(32'h3bf1054b),
	.w5(32'hbbf35fc1),
	.w6(32'h3b707d6e),
	.w7(32'h3ad2a882),
	.w8(32'hbb37f109),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a709f27),
	.w1(32'hbbc01405),
	.w2(32'hbb6f5282),
	.w3(32'hbb621e1d),
	.w4(32'hbb570b43),
	.w5(32'hbc03dec2),
	.w6(32'hba611ac0),
	.w7(32'h3bd2de89),
	.w8(32'hba2d67f1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43297e),
	.w1(32'hbba710ec),
	.w2(32'h3b8c8471),
	.w3(32'h3a77e4dd),
	.w4(32'h3b854aec),
	.w5(32'hba249e93),
	.w6(32'h3aea1769),
	.w7(32'h3c970c51),
	.w8(32'hba8f17ef),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37833dae),
	.w1(32'h3b08c2fc),
	.w2(32'h3a1782af),
	.w3(32'h3b9f4efd),
	.w4(32'h39f8f965),
	.w5(32'hbafc34ff),
	.w6(32'hbafc77be),
	.w7(32'hbb442a4b),
	.w8(32'h3b8b9fef),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50b1ab),
	.w1(32'h3a7ddef6),
	.w2(32'hbb21b459),
	.w3(32'hbb47038e),
	.w4(32'hba76cd10),
	.w5(32'h3b596c54),
	.w6(32'h3bd213f0),
	.w7(32'h3d22250b),
	.w8(32'h3bbed6aa),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00e307),
	.w1(32'hbbfbf729),
	.w2(32'hbc03a6ef),
	.w3(32'h3a978b65),
	.w4(32'h3b85a86d),
	.w5(32'h3a05b96b),
	.w6(32'hba24abba),
	.w7(32'h3b36ee8f),
	.w8(32'hbbfe3a90),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c8bbb),
	.w1(32'h3c109bce),
	.w2(32'hbb5320b7),
	.w3(32'hba3cf78c),
	.w4(32'hba7f206f),
	.w5(32'hb9f8ba0a),
	.w6(32'h3a2a7d31),
	.w7(32'h3b2c7048),
	.w8(32'h3c0a2401),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9f95c),
	.w1(32'h3beddddf),
	.w2(32'hbacdb54e),
	.w3(32'hbc05c836),
	.w4(32'hbad52d97),
	.w5(32'h3b61cefc),
	.w6(32'h3b294f18),
	.w7(32'hbbeabd79),
	.w8(32'hbafd556f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba855de6),
	.w1(32'hbadbb44c),
	.w2(32'h3c249aad),
	.w3(32'hba5556f6),
	.w4(32'h3b8fa2be),
	.w5(32'h3c72314c),
	.w6(32'hbb58bbdc),
	.w7(32'h3c0ee841),
	.w8(32'hb8c6b04d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa36992),
	.w1(32'h3c9d08d0),
	.w2(32'hbb887a1e),
	.w3(32'hbae8d4de),
	.w4(32'h3ba1c72f),
	.w5(32'hbb8eb3a7),
	.w6(32'hba5bf98d),
	.w7(32'h3bce5609),
	.w8(32'hba87f100),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea9454),
	.w1(32'hbb28e72f),
	.w2(32'hbb7aa547),
	.w3(32'h3c0a8375),
	.w4(32'h3c04e92a),
	.w5(32'h3c0bbd0a),
	.w6(32'h3c337d8a),
	.w7(32'h39a36fed),
	.w8(32'hbaf0e6c0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2f69e),
	.w1(32'hba1efd3d),
	.w2(32'hbb021474),
	.w3(32'hbb6394fe),
	.w4(32'hbb8390eb),
	.w5(32'h3a061985),
	.w6(32'h3c729a00),
	.w7(32'h3b181fb0),
	.w8(32'hbb7126af),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fcf31),
	.w1(32'hbc04b37e),
	.w2(32'hbc2804ce),
	.w3(32'h3ce86a0f),
	.w4(32'hbb20340f),
	.w5(32'h3b9e6de7),
	.w6(32'h36bd80a0),
	.w7(32'hbbc134cf),
	.w8(32'h387a0998),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42a89c),
	.w1(32'hb85d0efa),
	.w2(32'h3a50c054),
	.w3(32'hbb19aab1),
	.w4(32'h3be4773b),
	.w5(32'h3ad07418),
	.w6(32'h3ab24337),
	.w7(32'hbb82528f),
	.w8(32'h3a595282),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b543),
	.w1(32'h397687a4),
	.w2(32'h3b670ca5),
	.w3(32'h3c22c30a),
	.w4(32'h3ac6bb92),
	.w5(32'h3a9c5872),
	.w6(32'h3b35e665),
	.w7(32'h3b2fa835),
	.w8(32'hbb85699e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule