module layer_8_featuremap_204(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd345ccd),
	.w1(32'hbbd98035),
	.w2(32'hba8e50d2),
	.w3(32'hbd19c38a),
	.w4(32'hbaa45b24),
	.w5(32'hbabd730f),
	.w6(32'hbaa40fd0),
	.w7(32'hb90cc6e2),
	.w8(32'h3c21a749),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375d918d),
	.w1(32'h3b6e566c),
	.w2(32'h3b9c1e46),
	.w3(32'h3961fc71),
	.w4(32'h3bffa307),
	.w5(32'h3bf5fa62),
	.w6(32'h3c24c055),
	.w7(32'h3c526ae5),
	.w8(32'h3ba11b21),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80dd9a),
	.w1(32'h398c9ba0),
	.w2(32'h3ba0251e),
	.w3(32'hba78fa8a),
	.w4(32'hb9320932),
	.w5(32'h3b81cc1a),
	.w6(32'h3ba26505),
	.w7(32'h3b8e93cd),
	.w8(32'h3b01360c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f62a3),
	.w1(32'hbbf83060),
	.w2(32'hbb019138),
	.w3(32'h3a143df8),
	.w4(32'hba6525b6),
	.w5(32'hbc09a076),
	.w6(32'h3b9cf430),
	.w7(32'h3b486573),
	.w8(32'h3bfdba08),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d96dc8),
	.w1(32'hbcb9e905),
	.w2(32'hba0c1981),
	.w3(32'hbc0ec2ea),
	.w4(32'hbc95c466),
	.w5(32'hbaede7d5),
	.w6(32'hbc1b55a1),
	.w7(32'h3b8f2504),
	.w8(32'h3c7a55b5),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c818ad7),
	.w1(32'h39aa073a),
	.w2(32'h3beed3c3),
	.w3(32'h3c1e30fb),
	.w4(32'hbc0bb04b),
	.w5(32'h3a89c044),
	.w6(32'hbc1b70a0),
	.w7(32'h3c104548),
	.w8(32'h3c04501b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e5d46),
	.w1(32'hbb5ac1ec),
	.w2(32'hb9693184),
	.w3(32'h3c8cf02a),
	.w4(32'hbb8f5dcd),
	.w5(32'hb8ab562a),
	.w6(32'hbb854b87),
	.w7(32'hbb1429a3),
	.w8(32'h3a9886f0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ed68d),
	.w1(32'hbc2d8730),
	.w2(32'hbad31172),
	.w3(32'hb8dc6c1e),
	.w4(32'hbc323b50),
	.w5(32'hbb00a8cf),
	.w6(32'hbb607036),
	.w7(32'h3bf53cc4),
	.w8(32'h3c5ea850),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c6e34),
	.w1(32'hbd0f72b6),
	.w2(32'h3bfd8a68),
	.w3(32'hbb04898b),
	.w4(32'hbceb092d),
	.w5(32'h3bd15012),
	.w6(32'hbc68dcf1),
	.w7(32'h3c6e8464),
	.w8(32'h3d17aab4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebee45),
	.w1(32'h3bed8818),
	.w2(32'h3b169c79),
	.w3(32'h3cdc939a),
	.w4(32'h3b9794de),
	.w5(32'h3b03fb25),
	.w6(32'hbb6749a3),
	.w7(32'hbc1c5984),
	.w8(32'hb7277020),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ff349),
	.w1(32'hbc304f9c),
	.w2(32'hbbb851a0),
	.w3(32'hbc85d079),
	.w4(32'hbc697fe4),
	.w5(32'hbbf0a289),
	.w6(32'hbc3ca4a4),
	.w7(32'hbb970e73),
	.w8(32'h3c30837b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c946e1b),
	.w1(32'h3b56ee1b),
	.w2(32'hbb0fc640),
	.w3(32'h3c6bc42d),
	.w4(32'h3bec6b4e),
	.w5(32'hba4786b7),
	.w6(32'h3b069964),
	.w7(32'h3b14e2df),
	.w8(32'hbb22f229),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e1445),
	.w1(32'hbac439c0),
	.w2(32'h3b975d76),
	.w3(32'hbc599226),
	.w4(32'h3b57c957),
	.w5(32'h3c0cd80f),
	.w6(32'hbbd049d1),
	.w7(32'hbc2271ad),
	.w8(32'h3b7f0ab0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc9fc3),
	.w1(32'hb880ee04),
	.w2(32'hbb6870d9),
	.w3(32'hbbb29e10),
	.w4(32'h3c0a8224),
	.w5(32'hbb95fd00),
	.w6(32'h38ac96e1),
	.w7(32'hbbff5d0e),
	.w8(32'hbb9b96b0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38c2bc),
	.w1(32'hbca0133d),
	.w2(32'hbacfa813),
	.w3(32'hbc2c5471),
	.w4(32'hbcb05c54),
	.w5(32'hbbb8664b),
	.w6(32'hbc61313f),
	.w7(32'hba63230c),
	.w8(32'h3ca079bf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9eb7f8),
	.w1(32'h3b3040af),
	.w2(32'hbc2b6ffa),
	.w3(32'h3c5899a0),
	.w4(32'hb8504592),
	.w5(32'hbc315012),
	.w6(32'hbb16ec84),
	.w7(32'hbb0b8d21),
	.w8(32'hbbf68066),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5d2f1),
	.w1(32'h36b51fa3),
	.w2(32'hbbccf9e5),
	.w3(32'hbb9eb54c),
	.w4(32'hbb8e99c7),
	.w5(32'h3b2244e8),
	.w6(32'h3be0c0da),
	.w7(32'h398da6f7),
	.w8(32'h39879cfd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe962e7),
	.w1(32'hba8cbf96),
	.w2(32'hbb688d82),
	.w3(32'h3a28d090),
	.w4(32'h3a2f918f),
	.w5(32'hbb294ccf),
	.w6(32'hbb50e209),
	.w7(32'hbc3370d2),
	.w8(32'hbba129f5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d5528),
	.w1(32'hbba03eea),
	.w2(32'hbc8be482),
	.w3(32'hbc060820),
	.w4(32'hbb5cb7ad),
	.w5(32'hbc5553d4),
	.w6(32'hbc500564),
	.w7(32'hbcba0086),
	.w8(32'hbc6a91ed),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5eb2f0),
	.w1(32'hbbc46176),
	.w2(32'hbb2ffd5d),
	.w3(32'hbc8b4092),
	.w4(32'hbc4250e4),
	.w5(32'hbbc68c64),
	.w6(32'hbbddfd6b),
	.w7(32'hbb34d3ee),
	.w8(32'h3b9144e8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cd2f6),
	.w1(32'h3c37f8d5),
	.w2(32'h3c9a3486),
	.w3(32'h3c02a8d5),
	.w4(32'h3b505b91),
	.w5(32'h3c805182),
	.w6(32'h3b67f0b9),
	.w7(32'h3c45fe07),
	.w8(32'h3c362e4b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77db8d),
	.w1(32'h3bdb9a9b),
	.w2(32'h3c500870),
	.w3(32'h3c1da852),
	.w4(32'h3c2b09ec),
	.w5(32'h3c4694ed),
	.w6(32'h3b3a528a),
	.w7(32'h3b9e5231),
	.w8(32'h3c21cf91),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0da263),
	.w1(32'hbbe4125e),
	.w2(32'hbb8d328d),
	.w3(32'h3c2072f0),
	.w4(32'h3ad11f7d),
	.w5(32'h3c13f285),
	.w6(32'hbc13054d),
	.w7(32'hbc5b8816),
	.w8(32'h3b2359d0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15c225),
	.w1(32'h3ba92d00),
	.w2(32'h3bc9143f),
	.w3(32'h3c20f883),
	.w4(32'h3b95c551),
	.w5(32'h3b3103a5),
	.w6(32'h3b65bd62),
	.w7(32'hbabbb4af),
	.w8(32'h3be76e42),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6cd65),
	.w1(32'h3a851cfc),
	.w2(32'hbc2f4326),
	.w3(32'hbb2da543),
	.w4(32'h3bcc43a5),
	.w5(32'hbaa7ce0e),
	.w6(32'h3b58ada4),
	.w7(32'h3bd7e433),
	.w8(32'hba541e2b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bfd5),
	.w1(32'h3b157964),
	.w2(32'h3c67bb6c),
	.w3(32'hbbc1e21d),
	.w4(32'hb9e65c76),
	.w5(32'h3bee0d28),
	.w6(32'h3c5069ad),
	.w7(32'h3c1280a2),
	.w8(32'hbaf37bcf),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c919ed2),
	.w1(32'h3bdc94aa),
	.w2(32'h3c267446),
	.w3(32'h3c5ff2a9),
	.w4(32'h3bf012b5),
	.w5(32'h3aa694a5),
	.w6(32'h3c44c7f0),
	.w7(32'h3c23b6c9),
	.w8(32'h3ad9b4ee),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaedc90),
	.w1(32'hbc7688a8),
	.w2(32'hbc66c140),
	.w3(32'hbccce446),
	.w4(32'hbc7e1457),
	.w5(32'hbc588074),
	.w6(32'hbb893d8c),
	.w7(32'h39203156),
	.w8(32'h3bdb32bf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085013),
	.w1(32'hbd17bc14),
	.w2(32'hbd32c222),
	.w3(32'hbc892d58),
	.w4(32'hbd1ed010),
	.w5(32'hbd1aea4f),
	.w6(32'hbcbfc9f0),
	.w7(32'hbcc1b544),
	.w8(32'hbcedf6e5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3c5cee),
	.w1(32'hbad9fff6),
	.w2(32'h3a868f64),
	.w3(32'hbd2a337f),
	.w4(32'h3b9de897),
	.w5(32'h3b9f684d),
	.w6(32'h3a4748b0),
	.w7(32'hba1e8aaf),
	.w8(32'h3c9f1b8b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94d4d4),
	.w1(32'h3bc13bca),
	.w2(32'hb9745a71),
	.w3(32'h3ccfb5a6),
	.w4(32'hbbb48891),
	.w5(32'h3b71c753),
	.w6(32'h3c1df99d),
	.w7(32'h3ba643fd),
	.w8(32'hbc27b6e3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35c75f),
	.w1(32'hbbd160de),
	.w2(32'h3bbbaf44),
	.w3(32'h3b713c22),
	.w4(32'hbb62e72d),
	.w5(32'h3bb51534),
	.w6(32'hbbc1f3d5),
	.w7(32'h3b2b8bb5),
	.w8(32'h3c12e846),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5d5df),
	.w1(32'h3b92e8a7),
	.w2(32'hbae03fbc),
	.w3(32'h3bee8db1),
	.w4(32'h3b92784b),
	.w5(32'hbbb7e789),
	.w6(32'h3b8e2132),
	.w7(32'h3b01d13c),
	.w8(32'hbbd91a33),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d0063),
	.w1(32'h3a95cf87),
	.w2(32'h3a80a62a),
	.w3(32'hbc5a705c),
	.w4(32'h3ba2e5b9),
	.w5(32'h3b8ada7b),
	.w6(32'h3be4ee92),
	.w7(32'hb9f93291),
	.w8(32'hbbf44077),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82eb66),
	.w1(32'hbbdf9d4f),
	.w2(32'hbad11100),
	.w3(32'h3b1617e3),
	.w4(32'h3c2dde1d),
	.w5(32'hba94854f),
	.w6(32'h39814e4d),
	.w7(32'h38e3e8c9),
	.w8(32'hbb3e3448),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc42ea6),
	.w1(32'hbbecdfbb),
	.w2(32'h3b225c12),
	.w3(32'hbc4b035d),
	.w4(32'hbb82f603),
	.w5(32'h3b01c396),
	.w6(32'h3b332b0d),
	.w7(32'h3ac7a92c),
	.w8(32'hb831527f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018264),
	.w1(32'hbd16886f),
	.w2(32'hbd18136f),
	.w3(32'h3bfec5d2),
	.w4(32'hbd008a81),
	.w5(32'hbd082fd4),
	.w6(32'hbce3c955),
	.w7(32'hbcd95a5e),
	.w8(32'hbcd66770),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c4769),
	.w1(32'hbcba2156),
	.w2(32'hbc167271),
	.w3(32'hbd0f1d43),
	.w4(32'hbca7fb4a),
	.w5(32'hbc50388a),
	.w6(32'hbc398d1c),
	.w7(32'hbb2b505a),
	.w8(32'h3c512d2b),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04229a),
	.w1(32'h3b8bb1f8),
	.w2(32'hbad50152),
	.w3(32'h3b21cb96),
	.w4(32'h3b62a09c),
	.w5(32'hbb3847c5),
	.w6(32'hbadae21e),
	.w7(32'hbb8f2a50),
	.w8(32'h3ab1488c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e9f31),
	.w1(32'h3b3d5341),
	.w2(32'hbad8d6ef),
	.w3(32'h3a3842e0),
	.w4(32'hbb51bdc2),
	.w5(32'hbba03b5c),
	.w6(32'hba86a9ab),
	.w7(32'h38a775df),
	.w8(32'h3b70ee41),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35302e),
	.w1(32'h399ae285),
	.w2(32'hbbda20e9),
	.w3(32'hb8870421),
	.w4(32'h3bad24e0),
	.w5(32'hbb514461),
	.w6(32'h3b089566),
	.w7(32'hbb0061e6),
	.w8(32'hba17794e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dd7f5),
	.w1(32'h3d6d22ec),
	.w2(32'h3d4dff6f),
	.w3(32'hbb9e980c),
	.w4(32'h3d317d00),
	.w5(32'h3d254d77),
	.w6(32'h3d274e7e),
	.w7(32'h3ced64e0),
	.w8(32'h3c09c16e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd6d88e),
	.w1(32'hbcc010dd),
	.w2(32'hbd05aa84),
	.w3(32'h3cda5732),
	.w4(32'hbc3ac04a),
	.w5(32'hbc9d4092),
	.w6(32'hbc353fc1),
	.w7(32'hbc960fb3),
	.w8(32'hbcadbd2b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd056262),
	.w1(32'hba95e9b3),
	.w2(32'hbc1d451e),
	.w3(32'hbcd1ad35),
	.w4(32'h3a11917d),
	.w5(32'hbb34453b),
	.w6(32'hbb871d3a),
	.w7(32'hbbf6b6ba),
	.w8(32'hbb4ff0db),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba22fa2),
	.w1(32'hbb9ea512),
	.w2(32'h3b90d1b8),
	.w3(32'hbb9e009a),
	.w4(32'h3a6b5a4f),
	.w5(32'hba8b6384),
	.w6(32'h3c819cc3),
	.w7(32'h3c234360),
	.w8(32'h3c3232fe),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b980c),
	.w1(32'hbb9e1fd7),
	.w2(32'h3a286ee0),
	.w3(32'hbbfb846c),
	.w4(32'hbb253893),
	.w5(32'h3b06e349),
	.w6(32'hbaf905d3),
	.w7(32'h3a684362),
	.w8(32'h38b249d1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb201f),
	.w1(32'hbbf69543),
	.w2(32'hbbf4e496),
	.w3(32'h3a72e802),
	.w4(32'hbc28b88a),
	.w5(32'hbc30c449),
	.w6(32'hbb5aea30),
	.w7(32'hbb3c8fcb),
	.w8(32'hbba0af86),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8161f9),
	.w1(32'hbba0623d),
	.w2(32'hbc1ac371),
	.w3(32'hbc57d485),
	.w4(32'hbbec31f1),
	.w5(32'hbbb27349),
	.w6(32'hbbaf1681),
	.w7(32'hbb294c1f),
	.w8(32'hbc0bb1ab),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a225b),
	.w1(32'h3ab53ce0),
	.w2(32'h3a197c1d),
	.w3(32'h3a9efbe8),
	.w4(32'hbb0c6ab8),
	.w5(32'hb9fbd810),
	.w6(32'hbb263da4),
	.w7(32'hbbd1f3cc),
	.w8(32'hbb63f252),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6bcff),
	.w1(32'h3abbec8b),
	.w2(32'h3bc29b37),
	.w3(32'hbb265a75),
	.w4(32'hbc08a10b),
	.w5(32'h3c2740b4),
	.w6(32'hbc22472f),
	.w7(32'h3b55196a),
	.w8(32'h3c4f255a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80b2e9),
	.w1(32'hbc01781a),
	.w2(32'hbc3dca9d),
	.w3(32'h3c5b7ba0),
	.w4(32'h3b00ca8c),
	.w5(32'h3aaf642d),
	.w6(32'h3a4ed0cf),
	.w7(32'h3a0b4439),
	.w8(32'h3bb9f065),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe454c),
	.w1(32'h3cabfec8),
	.w2(32'h3cda62d6),
	.w3(32'hbbcf7a80),
	.w4(32'h3c0ca8db),
	.w5(32'h3c9430d7),
	.w6(32'h3c12e4e2),
	.w7(32'h3c18d6d7),
	.w8(32'h3c81f066),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0cbeae),
	.w1(32'hbc930792),
	.w2(32'hba54fa27),
	.w3(32'h3ce3890f),
	.w4(32'hbc41fcc8),
	.w5(32'h3b221228),
	.w6(32'hbb98a188),
	.w7(32'h3bec72bc),
	.w8(32'h3c7e0609),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c427b9f),
	.w1(32'hbb9249d1),
	.w2(32'hbc365b31),
	.w3(32'h3c4bd09b),
	.w4(32'hba7d2c70),
	.w5(32'hbb284280),
	.w6(32'h3b9017c0),
	.w7(32'hbba7a87d),
	.w8(32'hbb69f3de),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf50885),
	.w1(32'h3c02af58),
	.w2(32'hbc0994a0),
	.w3(32'hbbe243b1),
	.w4(32'h3bbb3a58),
	.w5(32'hbc20646a),
	.w6(32'h3c7516f7),
	.w7(32'hbb982258),
	.w8(32'hbc5937bd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2217bd),
	.w1(32'hbb75a858),
	.w2(32'h3a82a7e6),
	.w3(32'hbb8f9f28),
	.w4(32'h3a0b45c4),
	.w5(32'h3b92db0b),
	.w6(32'h3b825c5d),
	.w7(32'h3b8d394b),
	.w8(32'h3c2f53d7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf6a8),
	.w1(32'h3ba7c0cd),
	.w2(32'hbc312979),
	.w3(32'h3bfe7164),
	.w4(32'h3bb1e988),
	.w5(32'hbb1ec6f1),
	.w6(32'hba9d20b1),
	.w7(32'hbb9fe632),
	.w8(32'hbc8bfb20),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab7a89),
	.w1(32'hbd410e2f),
	.w2(32'hbd802091),
	.w3(32'hbc9bf558),
	.w4(32'hbd3318f8),
	.w5(32'hbd6c3003),
	.w6(32'hbd1d836d),
	.w7(32'hbd41790d),
	.w8(32'hbcfed02c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3798d6),
	.w1(32'h3b8afb90),
	.w2(32'hbb69668b),
	.w3(32'hbd31bdd7),
	.w4(32'h3b86d407),
	.w5(32'hbad15df3),
	.w6(32'h3bc75c21),
	.w7(32'h3ac02cc2),
	.w8(32'hbbb3c229),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ce18),
	.w1(32'h3b265f43),
	.w2(32'h3bda40c9),
	.w3(32'hbc0ae60c),
	.w4(32'h3b699df3),
	.w5(32'h3b4006c2),
	.w6(32'h3945ab46),
	.w7(32'h3b3badc8),
	.w8(32'hb95c1f2f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6a167),
	.w1(32'h3a44252e),
	.w2(32'h3a013407),
	.w3(32'h3aaa75ca),
	.w4(32'hbb55c90c),
	.w5(32'h3b0e54b1),
	.w6(32'hba91e681),
	.w7(32'h3b4f31de),
	.w8(32'hbbfcaa51),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce37fc),
	.w1(32'hbc9eb731),
	.w2(32'hbbf2212f),
	.w3(32'hbbfabb4c),
	.w4(32'hbbcfd19e),
	.w5(32'hbbb8d0cc),
	.w6(32'hbcc3e27b),
	.w7(32'hbb731eff),
	.w8(32'h3b8f3a92),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b757879),
	.w1(32'hbc3ae7d8),
	.w2(32'hbc218916),
	.w3(32'hbc245a76),
	.w4(32'hbc1bdbca),
	.w5(32'hbc3b48ec),
	.w6(32'hbc229441),
	.w7(32'hbc61549b),
	.w8(32'hbc371fcc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b8686),
	.w1(32'hbba8ac8a),
	.w2(32'hbc8b7fe8),
	.w3(32'hbc0ec7a0),
	.w4(32'hb93fadcd),
	.w5(32'hbc63492c),
	.w6(32'hb90d47ce),
	.w7(32'hbc4e7764),
	.w8(32'hbc60e5c2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb500be),
	.w1(32'h3c3b1aed),
	.w2(32'hba0c1096),
	.w3(32'hbc8b34d8),
	.w4(32'h3c1a5b87),
	.w5(32'h39a2a5df),
	.w6(32'h3c144c28),
	.w7(32'h3acb3c5b),
	.w8(32'hbc084818),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc433177),
	.w1(32'h3ab9e2e0),
	.w2(32'h3a4152eb),
	.w3(32'hbbc93b35),
	.w4(32'h3a870af6),
	.w5(32'h3b1761e3),
	.w6(32'h3bb1466c),
	.w7(32'hbb330442),
	.w8(32'hbaeb7fca),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53c848),
	.w1(32'h3bc58bfe),
	.w2(32'h3c1d1365),
	.w3(32'h3b533835),
	.w4(32'h3bb392bc),
	.w5(32'h3c0cc687),
	.w6(32'h3c1b669e),
	.w7(32'h3c80802a),
	.w8(32'h3c4601e0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4673aa),
	.w1(32'hbb0a498c),
	.w2(32'h3bacee2a),
	.w3(32'h3c7b7818),
	.w4(32'hbba179fc),
	.w5(32'h3b437295),
	.w6(32'h3c002257),
	.w7(32'h3a200ef7),
	.w8(32'hba94cc71),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8408a),
	.w1(32'h3ba7abfb),
	.w2(32'h3c3957d7),
	.w3(32'h3b859f3e),
	.w4(32'h3bdb9762),
	.w5(32'h3b572f15),
	.w6(32'hbac1266e),
	.w7(32'h3bde0831),
	.w8(32'h3a57845d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f4c6a),
	.w1(32'hbacfad4d),
	.w2(32'hbbc89dec),
	.w3(32'hbacfd6de),
	.w4(32'h3b010f0e),
	.w5(32'h3c021182),
	.w6(32'h3a8bd9f8),
	.w7(32'hbbaac3b5),
	.w8(32'hbc333dce),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72444b),
	.w1(32'h3d257cf3),
	.w2(32'h3d69685a),
	.w3(32'h3a304740),
	.w4(32'h3ce87620),
	.w5(32'h3d3ff519),
	.w6(32'h3cf8f83a),
	.w7(32'h3d1f6b61),
	.w8(32'h3d14b2d3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d42b410),
	.w1(32'hbb724c50),
	.w2(32'hbb297c1f),
	.w3(32'h3d46cc45),
	.w4(32'h3bc577da),
	.w5(32'h3b3e2898),
	.w6(32'h3b8534ba),
	.w7(32'hbaf540b6),
	.w8(32'hba3b1ee3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee5db),
	.w1(32'h3b5a2126),
	.w2(32'h3b7eddf7),
	.w3(32'h3b116d69),
	.w4(32'h3ba37f9e),
	.w5(32'h3a6e7b42),
	.w6(32'h3ae8134c),
	.w7(32'h3be584c2),
	.w8(32'hb9f95335),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb022c),
	.w1(32'h3a021631),
	.w2(32'hbcaec5af),
	.w3(32'h3b98cea5),
	.w4(32'h3b1b81a3),
	.w5(32'hbc8ef7f7),
	.w6(32'hba85bea2),
	.w7(32'hbbdaa1e8),
	.w8(32'h3b8b79b6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d75ea),
	.w1(32'h3d0de706),
	.w2(32'h3cf897d5),
	.w3(32'hbbeb2995),
	.w4(32'h3d012203),
	.w5(32'h3cf274b2),
	.w6(32'h3cb13eb6),
	.w7(32'h3c84b8a5),
	.w8(32'h3c553c6b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2a499),
	.w1(32'hbb723d04),
	.w2(32'h3bbf1f35),
	.w3(32'h3c9152bd),
	.w4(32'h39191b19),
	.w5(32'h3afd76dd),
	.w6(32'hbb083e77),
	.w7(32'h3b5b794d),
	.w8(32'hbbb6b944),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29137f),
	.w1(32'hbc25cdd4),
	.w2(32'hbcaa0fda),
	.w3(32'hb9e1a788),
	.w4(32'hbbee33a1),
	.w5(32'hbc68becc),
	.w6(32'hbc0a855d),
	.w7(32'hbc436696),
	.w8(32'hbc4d86fb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3ab4d),
	.w1(32'hbcf5ed60),
	.w2(32'hbd317fa4),
	.w3(32'hbc9f5491),
	.w4(32'hbcd69145),
	.w5(32'hbd107e4a),
	.w6(32'hbc9e9918),
	.w7(32'hbd038bab),
	.w8(32'hbcd8cb10),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd043e5f),
	.w1(32'h3cb71f12),
	.w2(32'h3c7fc4a1),
	.w3(32'hbd0a84c8),
	.w4(32'h3be1d3d5),
	.w5(32'h3c4d4e21),
	.w6(32'h3b8d236b),
	.w7(32'h3c477c42),
	.w8(32'h3bd18745),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c438d65),
	.w1(32'hba00f429),
	.w2(32'h3b8e59f5),
	.w3(32'h3c1b4263),
	.w4(32'hbbbe275f),
	.w5(32'h3b7f2950),
	.w6(32'hbb3693d5),
	.w7(32'hb9ab5afb),
	.w8(32'h3b8a30f8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72322e),
	.w1(32'hbb2e29f0),
	.w2(32'h3aed5e00),
	.w3(32'hbb411520),
	.w4(32'h3c01b3d1),
	.w5(32'h3b696453),
	.w6(32'hbba1616f),
	.w7(32'h3b61ac2c),
	.w8(32'h39309116),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a4534),
	.w1(32'hbb8784dc),
	.w2(32'h3b27a7cb),
	.w3(32'hbbe7f722),
	.w4(32'h3a059d68),
	.w5(32'h3bafe1f4),
	.w6(32'hb9fd8007),
	.w7(32'h3ae1d5de),
	.w8(32'h3b643a9d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc618f3),
	.w1(32'hbb760eb4),
	.w2(32'hbbd36d9f),
	.w3(32'hb84bb456),
	.w4(32'h3ae90006),
	.w5(32'hbc23c8ca),
	.w6(32'hbb985bee),
	.w7(32'hbc241d82),
	.w8(32'hbad173ad),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e014e),
	.w1(32'h3c6321d4),
	.w2(32'hbc282c96),
	.w3(32'h3926e96f),
	.w4(32'h3c59b9b0),
	.w5(32'hbc3f3744),
	.w6(32'h3b6864fe),
	.w7(32'hbb052c8c),
	.w8(32'hbab02a6d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb788530),
	.w1(32'hb8b9a22f),
	.w2(32'hbc0b3ffa),
	.w3(32'hbbfffe3c),
	.w4(32'hbb8a3d0f),
	.w5(32'hba685ef9),
	.w6(32'hbb3fc043),
	.w7(32'h3b043198),
	.w8(32'h3b41f7c6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefc11),
	.w1(32'h3a955b48),
	.w2(32'h3a9cc385),
	.w3(32'hbbb925c1),
	.w4(32'h3a8fe453),
	.w5(32'h3b5734f2),
	.w6(32'h3b585584),
	.w7(32'h3a605bbd),
	.w8(32'h3bc80fdf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ed997),
	.w1(32'h3c733a9e),
	.w2(32'h3c207aa1),
	.w3(32'h3c3a2c57),
	.w4(32'h3c094afa),
	.w5(32'h3c316ceb),
	.w6(32'h3c8c42f7),
	.w7(32'h3c28f359),
	.w8(32'h3c059032),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10e895),
	.w1(32'hbc10cf1b),
	.w2(32'hbc786abc),
	.w3(32'h3c6a836f),
	.w4(32'h3c0af446),
	.w5(32'hbbbf5371),
	.w6(32'hbc29bbcc),
	.w7(32'hbb7e029d),
	.w8(32'hbb3cd8fb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c655),
	.w1(32'hbc0a50ad),
	.w2(32'hbc1e9c9d),
	.w3(32'hbc7e23d5),
	.w4(32'h3b165ee0),
	.w5(32'h39d68f2d),
	.w6(32'h3b54b630),
	.w7(32'h3aa452b4),
	.w8(32'hbb12f37a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba496b3),
	.w1(32'h3b90f5ea),
	.w2(32'h3ad772d3),
	.w3(32'hbba71d93),
	.w4(32'h3b38bd80),
	.w5(32'hbb912438),
	.w6(32'hbb131aba),
	.w7(32'h38df6d0c),
	.w8(32'h3ae2eb78),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2191a9),
	.w1(32'h3ae23a01),
	.w2(32'hbb458c0d),
	.w3(32'hba701d43),
	.w4(32'h3b496788),
	.w5(32'h3bafb28e),
	.w6(32'h3bbc5131),
	.w7(32'h3bb3a3f9),
	.w8(32'h3b99c6f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12c398),
	.w1(32'hba31938a),
	.w2(32'hb9e41e4a),
	.w3(32'h3aa743f3),
	.w4(32'hbac5274e),
	.w5(32'h3a09ca79),
	.w6(32'hbb0c5b03),
	.w7(32'h3afec053),
	.w8(32'hbb2564e8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87cc2d),
	.w1(32'h3bc12297),
	.w2(32'h3b182700),
	.w3(32'h3b7f35f0),
	.w4(32'h3b8d1f66),
	.w5(32'h393f3db2),
	.w6(32'h3b921f91),
	.w7(32'hba2b240c),
	.w8(32'hbbb933c7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd99ce),
	.w1(32'h3c3622c0),
	.w2(32'h3b56b1a5),
	.w3(32'hbbfc53d9),
	.w4(32'h3c256243),
	.w5(32'h3bb0c688),
	.w6(32'h3c2a2a61),
	.w7(32'h3befec48),
	.w8(32'hbad8a4f6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e1f56),
	.w1(32'hbc4fa9dd),
	.w2(32'hbb4b2132),
	.w3(32'hbb415747),
	.w4(32'hbc46794a),
	.w5(32'h3aa3a44f),
	.w6(32'hbbeeb8e3),
	.w7(32'h3c6643cc),
	.w8(32'h3c9d2979),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd23ef),
	.w1(32'hbd24095f),
	.w2(32'hbd1da058),
	.w3(32'h3b8c90ea),
	.w4(32'hbd134c26),
	.w5(32'hbd0d6bee),
	.w6(32'hbcdb1d6d),
	.w7(32'hbcc8baa3),
	.w8(32'hbcf25012),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2a70b4),
	.w1(32'h39bbca43),
	.w2(32'hbc11e598),
	.w3(32'hbd286c0a),
	.w4(32'hbba638a4),
	.w5(32'hbba1ee0a),
	.w6(32'h3b1236b9),
	.w7(32'hbb9bcd85),
	.w8(32'hbc8016de),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae7c20),
	.w1(32'h3b1b452e),
	.w2(32'hbab3885a),
	.w3(32'hbc08ea09),
	.w4(32'h3bb22923),
	.w5(32'hbb1eb4c3),
	.w6(32'hbbfed0c2),
	.w7(32'hba5dd191),
	.w8(32'hbb69c7fa),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49f58d),
	.w1(32'hbc138731),
	.w2(32'hbbcf31ca),
	.w3(32'hbbeec11a),
	.w4(32'hbb8a7e98),
	.w5(32'hba874ba4),
	.w6(32'hbbca98bd),
	.w7(32'hbbd88a36),
	.w8(32'h3adf7691),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1cfa8),
	.w1(32'hbb8d5578),
	.w2(32'hbb82ec37),
	.w3(32'h3b5b80fa),
	.w4(32'hbc84b9a8),
	.w5(32'hbb96955d),
	.w6(32'h3a95b2ab),
	.w7(32'hbb0d0929),
	.w8(32'hbc1130fc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ba74),
	.w1(32'hbb30a127),
	.w2(32'hbc0cc79b),
	.w3(32'h3ab0c310),
	.w4(32'h3b873c84),
	.w5(32'hbc2889a9),
	.w6(32'h3acc93b1),
	.w7(32'hbb189a14),
	.w8(32'h3b996d3e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dce7a),
	.w1(32'h3aef9402),
	.w2(32'h3bc10f6a),
	.w3(32'hbc0b8bc3),
	.w4(32'h3bcfcdff),
	.w5(32'h3bf1bbd5),
	.w6(32'h3bdae9ce),
	.w7(32'h3bb5d7d3),
	.w8(32'h3c4cd078),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33fb54),
	.w1(32'h3bb791fa),
	.w2(32'h3b03242b),
	.w3(32'h3be49297),
	.w4(32'hbad79d44),
	.w5(32'h3ae787f2),
	.w6(32'hbb1520eb),
	.w7(32'h3b1165ee),
	.w8(32'hb9473f16),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b5c66),
	.w1(32'h3c57b488),
	.w2(32'h3c700b27),
	.w3(32'hbaa52e4b),
	.w4(32'h3c84da9f),
	.w5(32'h3b961eae),
	.w6(32'h3c57e17e),
	.w7(32'h3bd5305d),
	.w8(32'hbb399955),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94ff2c),
	.w1(32'hbad84701),
	.w2(32'hbb56d2aa),
	.w3(32'h3bb7c7a8),
	.w4(32'hbaf95353),
	.w5(32'hbc06ec15),
	.w6(32'h3ab454eb),
	.w7(32'hba788937),
	.w8(32'h3ac69556),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093e74),
	.w1(32'hbb9d4c31),
	.w2(32'h3bada8c9),
	.w3(32'h3bcba993),
	.w4(32'hbbd1f56e),
	.w5(32'h3b6b66b3),
	.w6(32'hbaac9564),
	.w7(32'h3b968168),
	.w8(32'h3bf54f0b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51215f),
	.w1(32'hbc3a9b78),
	.w2(32'hbc64c2f5),
	.w3(32'h3c3a7ebd),
	.w4(32'hbc32c19b),
	.w5(32'hbbc2c1b3),
	.w6(32'h3b9ba7f9),
	.w7(32'hb9a4053d),
	.w8(32'hbc125375),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19d4cb),
	.w1(32'hbca5c12f),
	.w2(32'hbd0b5ae2),
	.w3(32'hbbaab8f2),
	.w4(32'hbc6744ef),
	.w5(32'hbcc3ed23),
	.w6(32'hbc4e9fd0),
	.w7(32'hbc960840),
	.w8(32'hbc61beb2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca16836),
	.w1(32'hbb856f47),
	.w2(32'hbb9d7d19),
	.w3(32'hbcabb0bd),
	.w4(32'hbaac1017),
	.w5(32'hbc22f2af),
	.w6(32'hbace7b2e),
	.w7(32'hbb7c5bc8),
	.w8(32'hbb2f24cd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fcc36),
	.w1(32'h3bef0d1d),
	.w2(32'h3b982939),
	.w3(32'hbb89998a),
	.w4(32'h3c10e83a),
	.w5(32'h3b961d2f),
	.w6(32'h3bf946ce),
	.w7(32'h3bd9a901),
	.w8(32'hbaaa0501),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa7018),
	.w1(32'hbb3e1c2d),
	.w2(32'hbba68d7e),
	.w3(32'hbbb8a823),
	.w4(32'h3b2a1fd8),
	.w5(32'hb94ed90e),
	.w6(32'h3b86692b),
	.w7(32'hb93941a4),
	.w8(32'h3b89acca),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae7cfa),
	.w1(32'h3ca14fde),
	.w2(32'h3bd4df3f),
	.w3(32'hba37b970),
	.w4(32'h3c9e295a),
	.w5(32'h3c2a0757),
	.w6(32'h3c6fbbd5),
	.w7(32'h3c008668),
	.w8(32'hbbd7d99a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f91de),
	.w1(32'hba8caa9f),
	.w2(32'h3b795f99),
	.w3(32'hbb8287bd),
	.w4(32'hbb94165a),
	.w5(32'h3bee2939),
	.w6(32'hbaa49085),
	.w7(32'h3ae8f7f3),
	.w8(32'h3b1630ab),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9e6fb),
	.w1(32'h3b8ee0fe),
	.w2(32'h3ab20758),
	.w3(32'hbbe1ed49),
	.w4(32'h3b106e12),
	.w5(32'h3c04c3fc),
	.w6(32'hbaa53372),
	.w7(32'hb7caa736),
	.w8(32'h3a3e6e5a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f2f4),
	.w1(32'h3cb0a024),
	.w2(32'h3ccfda06),
	.w3(32'h3c44677c),
	.w4(32'h3c98cc79),
	.w5(32'h3cbb6b82),
	.w6(32'h3c51db08),
	.w7(32'h3c808c11),
	.w8(32'h3c765c9f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc09643),
	.w1(32'h3bae1c91),
	.w2(32'hbaed9a28),
	.w3(32'h3cc1bf18),
	.w4(32'h3bc2c425),
	.w5(32'hb8967770),
	.w6(32'h3bb9b023),
	.w7(32'h3b2c78f0),
	.w8(32'hbbb9f73f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2475f3),
	.w1(32'h3b84cfc7),
	.w2(32'h3c10c438),
	.w3(32'hbbe3baf1),
	.w4(32'hbc547fff),
	.w5(32'h3c16d3a9),
	.w6(32'h3b6e3d92),
	.w7(32'h3bf0304a),
	.w8(32'h3bcc1465),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fb6dd),
	.w1(32'hbaa458c5),
	.w2(32'hb991ddb5),
	.w3(32'h3ca4ae5c),
	.w4(32'h3ab50eda),
	.w5(32'hbaed6801),
	.w6(32'hbb8e0bdc),
	.w7(32'hbb2dbd84),
	.w8(32'hb86b9423),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd8c43),
	.w1(32'h3b822b41),
	.w2(32'hbbfc2027),
	.w3(32'h3b0cc647),
	.w4(32'h3b92c219),
	.w5(32'hbab2c9b5),
	.w6(32'hbc29236a),
	.w7(32'hbb6fd9c0),
	.w8(32'h3b1fa625),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b565929),
	.w1(32'h3ca8ce5d),
	.w2(32'h3c8fc1cf),
	.w3(32'hbbf1ad4e),
	.w4(32'h3c5af31a),
	.w5(32'h3c310e3d),
	.w6(32'h3c4ee89d),
	.w7(32'h3bfc6245),
	.w8(32'h3ba2c5fe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c749bf8),
	.w1(32'h3c235e4d),
	.w2(32'h3c203f2b),
	.w3(32'h3c5ac445),
	.w4(32'h3b995b81),
	.w5(32'h3c86d147),
	.w6(32'h3bb759a4),
	.w7(32'h3ba28e91),
	.w8(32'h3b93df00),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09de18),
	.w1(32'hbb58ef09),
	.w2(32'hba72692e),
	.w3(32'h3b165364),
	.w4(32'h3a4635b9),
	.w5(32'hbba0a9eb),
	.w6(32'hbb377c38),
	.w7(32'h3987a5d3),
	.w8(32'h3aa2ffc0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f067a),
	.w1(32'hbbad0793),
	.w2(32'hbb8f2861),
	.w3(32'hbba82629),
	.w4(32'hbb0d09ef),
	.w5(32'hbb74ab7d),
	.w6(32'hb8cd4c16),
	.w7(32'hbafc57bf),
	.w8(32'hbbf48ea9),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38a32f),
	.w1(32'h3b2f15a1),
	.w2(32'h3b925320),
	.w3(32'hbc10928d),
	.w4(32'h3b89aa8b),
	.w5(32'hba95d643),
	.w6(32'hba1c7f17),
	.w7(32'h3a76d720),
	.w8(32'h3a92d176),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd24904),
	.w1(32'h3a39d945),
	.w2(32'hbb2b4760),
	.w3(32'h3be2b16a),
	.w4(32'h3b3bc9a0),
	.w5(32'h3b3df073),
	.w6(32'hbadd288d),
	.w7(32'hbb406a0c),
	.w8(32'hbb9c1b10),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7606),
	.w1(32'hbb2ffd9e),
	.w2(32'hbb6a1457),
	.w3(32'h3b3b6536),
	.w4(32'hbbb0c6c0),
	.w5(32'h3ab44f9a),
	.w6(32'hbb47c5e1),
	.w7(32'hbb39c1c1),
	.w8(32'hbbbc9787),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895123a),
	.w1(32'h3a154dec),
	.w2(32'h3b204ac1),
	.w3(32'h3b841330),
	.w4(32'h3ab65c04),
	.w5(32'h3bb17861),
	.w6(32'h3b0d2fa4),
	.w7(32'h3b7dae06),
	.w8(32'h3aaac59e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133b24),
	.w1(32'h3c114360),
	.w2(32'h3bee8823),
	.w3(32'hba454c74),
	.w4(32'h3c2680c1),
	.w5(32'h3ac6dc83),
	.w6(32'h3bb9e03c),
	.w7(32'h3b640dc4),
	.w8(32'hbba1df4d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule