module layer_10_featuremap_444(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac07fc),
	.w1(32'hbb3e7df2),
	.w2(32'hbbd54816),
	.w3(32'hbad1fc07),
	.w4(32'h3af9e8eb),
	.w5(32'h3b5c8739),
	.w6(32'h39adb08f),
	.w7(32'h39fa6c9d),
	.w8(32'h3c04c841),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1e577),
	.w1(32'h3a4a99ce),
	.w2(32'h3b45ce66),
	.w3(32'h3b77840e),
	.w4(32'h3b423cad),
	.w5(32'h3b8803b1),
	.w6(32'h3bacb0e7),
	.w7(32'h3ae612e1),
	.w8(32'h3bc7e293),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf180db),
	.w1(32'h393d0ad2),
	.w2(32'hbb7a6a2f),
	.w3(32'hbb36da57),
	.w4(32'h3b6f7f71),
	.w5(32'h3b093b4a),
	.w6(32'hbb88401c),
	.w7(32'h3a3f1cb3),
	.w8(32'h39c2fce5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba497961),
	.w1(32'hbbc01dff),
	.w2(32'hbbe81de3),
	.w3(32'h3beb8437),
	.w4(32'hbbaf4f92),
	.w5(32'hbc126add),
	.w6(32'h3b3335f2),
	.w7(32'h3b4a6865),
	.w8(32'h3b38a745),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dd2cd),
	.w1(32'hbaf36cce),
	.w2(32'hbb22676e),
	.w3(32'h3b4fac84),
	.w4(32'hbbda331d),
	.w5(32'h3b012e4f),
	.w6(32'hba539171),
	.w7(32'hbb1e8973),
	.w8(32'hba9134e7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fb98ef),
	.w1(32'h3b150a51),
	.w2(32'h3a381147),
	.w3(32'h3b0cd674),
	.w4(32'h3b9b882c),
	.w5(32'hbbd51b1b),
	.w6(32'h3a2661a9),
	.w7(32'hbba5255e),
	.w8(32'hba152eb5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17ee47),
	.w1(32'hbbb0d9da),
	.w2(32'hbc823486),
	.w3(32'hbae91749),
	.w4(32'hbc1da071),
	.w5(32'hbc850734),
	.w6(32'hbbf6b580),
	.w7(32'hbc55c4cc),
	.w8(32'hbc7bcea6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83f18b),
	.w1(32'hbaff9457),
	.w2(32'h3a2bdcfb),
	.w3(32'hba45e051),
	.w4(32'hbc16c950),
	.w5(32'h3bbb6e7c),
	.w6(32'hba06f1d1),
	.w7(32'h3a5053a2),
	.w8(32'h3c084a58),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae00eef),
	.w1(32'h3a877ca0),
	.w2(32'h3b2d9c69),
	.w3(32'h3b0d56b4),
	.w4(32'hbacfa384),
	.w5(32'hbb0538d5),
	.w6(32'hb882b4b5),
	.w7(32'h3acb7898),
	.w8(32'h3bc8da5e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d6291),
	.w1(32'hbb9adf16),
	.w2(32'hbbe38612),
	.w3(32'h3c6f333b),
	.w4(32'hbacba61b),
	.w5(32'hbbe43eb2),
	.w6(32'h3b7e3359),
	.w7(32'hbba04f38),
	.w8(32'hbafa10d8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c08b25),
	.w1(32'hbb36d9a7),
	.w2(32'hbb113ffc),
	.w3(32'h3a3cc5ea),
	.w4(32'hbb226902),
	.w5(32'h3a5d0629),
	.w6(32'hbb827697),
	.w7(32'hb9bf44fb),
	.w8(32'hba025045),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947c35),
	.w1(32'hbb4f0117),
	.w2(32'hbba3439d),
	.w3(32'h3bd6d38d),
	.w4(32'hbb98d939),
	.w5(32'hbc099e5f),
	.w6(32'hbb05e544),
	.w7(32'hbc4b03be),
	.w8(32'hbc88ac07),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4237ea),
	.w1(32'hbc0fc5d9),
	.w2(32'hbb636d7e),
	.w3(32'h3adb73b7),
	.w4(32'hbc7a519c),
	.w5(32'hbc04631c),
	.w6(32'hbafcfe2b),
	.w7(32'hbc8b3e5f),
	.w8(32'hbc114396),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe75a4b),
	.w1(32'hbb9a3742),
	.w2(32'h3a1ff886),
	.w3(32'hbbc10ddb),
	.w4(32'hbbfaaed4),
	.w5(32'hbbbd708d),
	.w6(32'hbc381f35),
	.w7(32'hbb9b3353),
	.w8(32'hbb4c263a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6a938),
	.w1(32'hbbd81744),
	.w2(32'h39ce18e7),
	.w3(32'h3b164a8a),
	.w4(32'hbaedd332),
	.w5(32'h3b35b73b),
	.w6(32'h3ac7fc2e),
	.w7(32'h3ad6f934),
	.w8(32'hbacdb3a3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dc788),
	.w1(32'hba9e509b),
	.w2(32'h3c38e3dd),
	.w3(32'h3aa48f9d),
	.w4(32'hbb893e79),
	.w5(32'h3c7058ee),
	.w6(32'h3b8038fe),
	.w7(32'h3be550a6),
	.w8(32'h3c08e5f8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d31a6),
	.w1(32'hbb062bcd),
	.w2(32'hba61617e),
	.w3(32'hbaa87727),
	.w4(32'hbadd7711),
	.w5(32'hbb1b3e05),
	.w6(32'hbaf32645),
	.w7(32'hba80ca44),
	.w8(32'hbac72d8c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd5390),
	.w1(32'hbbf69ab1),
	.w2(32'hbc0fca85),
	.w3(32'hbb6a0f72),
	.w4(32'hbc4050f1),
	.w5(32'hbc002388),
	.w6(32'hbb5f370d),
	.w7(32'hbbb62d12),
	.w8(32'h3b2af7a2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7dd8c),
	.w1(32'hbbdde497),
	.w2(32'hbbbc2caa),
	.w3(32'hba500597),
	.w4(32'hbc6a7187),
	.w5(32'hbc1b1471),
	.w6(32'h3b56832a),
	.w7(32'hbc42612f),
	.w8(32'hbb939716),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb978533),
	.w1(32'hbba5d6ed),
	.w2(32'hba436d91),
	.w3(32'hba6a6b10),
	.w4(32'hbb959a68),
	.w5(32'hb9a7fc32),
	.w6(32'hbaf5678f),
	.w7(32'hba0c5625),
	.w8(32'h3b77b3d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf8a9),
	.w1(32'h3aeb9401),
	.w2(32'hba01fc5d),
	.w3(32'hbb6da98b),
	.w4(32'h3b388d7b),
	.w5(32'hbbc028c6),
	.w6(32'hbb0be5dd),
	.w7(32'hba31b536),
	.w8(32'hb9cc474f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ba8bd),
	.w1(32'hba6d827c),
	.w2(32'h3bbcbee8),
	.w3(32'hb95036bb),
	.w4(32'h3b68345f),
	.w5(32'h3b9620b5),
	.w6(32'hbabf8b2f),
	.w7(32'h3ba21b7e),
	.w8(32'hbada8a45),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d437),
	.w1(32'h3be31218),
	.w2(32'hbb8d8ea9),
	.w3(32'h3a04c09d),
	.w4(32'h3b9798b8),
	.w5(32'hbc1793f2),
	.w6(32'hbb7c43ea),
	.w7(32'hbc8187d5),
	.w8(32'hbc84f6dc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dc7e7),
	.w1(32'hb98fde00),
	.w2(32'hb8f2d790),
	.w3(32'hbae74b87),
	.w4(32'h39f8171b),
	.w5(32'hbb24a1d5),
	.w6(32'hb979f6e9),
	.w7(32'hbbbae1e5),
	.w8(32'hbade73d6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917586),
	.w1(32'h3ac9dd1a),
	.w2(32'hbb2a89c7),
	.w3(32'h3b855f55),
	.w4(32'h3b928522),
	.w5(32'h3b8540b0),
	.w6(32'h3b9a38a2),
	.w7(32'hbaecac7e),
	.w8(32'h3b439c41),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2930bf),
	.w1(32'h3aff90e4),
	.w2(32'hbb1832bc),
	.w3(32'h3a829abd),
	.w4(32'h3b0d0b64),
	.w5(32'hbad9792a),
	.w6(32'hbb1567a4),
	.w7(32'h3ab059f0),
	.w8(32'hbb96655e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44b5ef),
	.w1(32'h3b49d075),
	.w2(32'h3b16321e),
	.w3(32'hbac991e1),
	.w4(32'h3a8f0b27),
	.w5(32'hba6ca75c),
	.w6(32'hbba15ef7),
	.w7(32'h3928e7be),
	.w8(32'h3a14e4ed),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c31f9),
	.w1(32'hbaf8ae3c),
	.w2(32'hbbfab777),
	.w3(32'h3bc6c592),
	.w4(32'hbbfe799a),
	.w5(32'hbb901fcd),
	.w6(32'h3bbec653),
	.w7(32'h3b9bd78d),
	.w8(32'hbc05af5e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39888787),
	.w1(32'h3b9a25bc),
	.w2(32'h3bb4900c),
	.w3(32'hba883b8a),
	.w4(32'h3bbab584),
	.w5(32'h3adb7568),
	.w6(32'hbac37e84),
	.w7(32'hba82f2ec),
	.w8(32'h3b9f3c14),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d9e1),
	.w1(32'h3b172b53),
	.w2(32'h3acd153c),
	.w3(32'hbadbba21),
	.w4(32'hbb41bb23),
	.w5(32'h3b3c50a0),
	.w6(32'hbbd6e374),
	.w7(32'hbbaa1a27),
	.w8(32'h3b50bcc7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944648),
	.w1(32'hba8f2ed6),
	.w2(32'hbad7d451),
	.w3(32'hba31b8ef),
	.w4(32'hba7d6ac2),
	.w5(32'hbb2798f8),
	.w6(32'h3b4450c3),
	.w7(32'hbb27e2e9),
	.w8(32'h3a851302),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb293a6d),
	.w1(32'h3b06722f),
	.w2(32'hbae1e1f8),
	.w3(32'hbb8530cf),
	.w4(32'h3b92ed07),
	.w5(32'hba750e00),
	.w6(32'hbb705899),
	.w7(32'h3b6fd5b2),
	.w8(32'h3af3dc74),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e3cc7e),
	.w1(32'hba4f043f),
	.w2(32'hbb0f075b),
	.w3(32'h3accfe38),
	.w4(32'hbb12c21e),
	.w5(32'hbb66404e),
	.w6(32'h3b079489),
	.w7(32'hba6b15a7),
	.w8(32'hbb89fd27),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e035),
	.w1(32'h3c041819),
	.w2(32'h3b898ff0),
	.w3(32'h3bbb492e),
	.w4(32'h3b0fafff),
	.w5(32'h39e3fe86),
	.w6(32'hbae974d4),
	.w7(32'h3bc76cc6),
	.w8(32'h3a7978ea),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95cb47a),
	.w1(32'h3b02bca1),
	.w2(32'hba425fba),
	.w3(32'h3b986bb9),
	.w4(32'hbb3a171a),
	.w5(32'hbb067586),
	.w6(32'h3a37d32e),
	.w7(32'hba8b28d2),
	.w8(32'h3b2d4c39),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa5681),
	.w1(32'hbbb14624),
	.w2(32'hbba26ed9),
	.w3(32'h3a09c1cf),
	.w4(32'hbb12c76b),
	.w5(32'hbbf89892),
	.w6(32'h3a62d6d6),
	.w7(32'hbb74d753),
	.w8(32'hbb9e8e91),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4af3b6),
	.w1(32'h3c1b7b5c),
	.w2(32'hba404424),
	.w3(32'h3b9b2666),
	.w4(32'h3ca52b4c),
	.w5(32'h37b72d44),
	.w6(32'h3c21cf2b),
	.w7(32'h3c2a7d7f),
	.w8(32'hbc9be28d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00205),
	.w1(32'h3a9c184b),
	.w2(32'hbbbbad65),
	.w3(32'hbc25344f),
	.w4(32'h3c270e2e),
	.w5(32'h3c201d78),
	.w6(32'hbc2e8af6),
	.w7(32'h3b9518a1),
	.w8(32'h3bf49046),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc3bcf),
	.w1(32'hbc48f7ca),
	.w2(32'hbc5d57db),
	.w3(32'hbcb1a28c),
	.w4(32'hbb8223bd),
	.w5(32'h3b841743),
	.w6(32'hbc8db1e9),
	.w7(32'hb9a323cb),
	.w8(32'h3b445870),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1023f1),
	.w1(32'h3b3a2610),
	.w2(32'hbb66ab07),
	.w3(32'h3b3abd78),
	.w4(32'h3be6d963),
	.w5(32'h39ad79eb),
	.w6(32'h3bb2b115),
	.w7(32'h3bca647e),
	.w8(32'h3b25933c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932711),
	.w1(32'hbb4b5b78),
	.w2(32'h3b836017),
	.w3(32'hbb211512),
	.w4(32'hbb83536c),
	.w5(32'h3b553373),
	.w6(32'hbb9faeac),
	.w7(32'hbb68e5fb),
	.w8(32'hbb73f293),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22b55c),
	.w1(32'h3a29c93d),
	.w2(32'h38c735f2),
	.w3(32'hbb6587b0),
	.w4(32'h3969d6c1),
	.w5(32'hbb4b8dda),
	.w6(32'hbb6f5f52),
	.w7(32'hba8a89b4),
	.w8(32'hbb92cea3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27caba),
	.w1(32'hba9a4f80),
	.w2(32'h3ab01210),
	.w3(32'hbb206a62),
	.w4(32'hbb679bf9),
	.w5(32'h3b122a13),
	.w6(32'h3a274505),
	.w7(32'h3a298de3),
	.w8(32'h3b526e88),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad24f),
	.w1(32'hbbd5a177),
	.w2(32'hbc1d828e),
	.w3(32'hbb1ad922),
	.w4(32'hbc4f6213),
	.w5(32'hbc55329e),
	.w6(32'h393416d9),
	.w7(32'hbc267c39),
	.w8(32'h3bdfebfd),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baaf9b1),
	.w1(32'hbb67fc3c),
	.w2(32'hbb3a3d65),
	.w3(32'h3bf9e0a9),
	.w4(32'hbb7cb657),
	.w5(32'hb9e54e47),
	.w6(32'h3c2e505d),
	.w7(32'hbab4c7ce),
	.w8(32'hbb0ca822),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb8d05),
	.w1(32'hbb45ca09),
	.w2(32'hbbb0c909),
	.w3(32'h3b6562be),
	.w4(32'hbb3c2af1),
	.w5(32'h3ade685a),
	.w6(32'h3911157c),
	.w7(32'h3ad742b4),
	.w8(32'h3ac8e243),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc06e3),
	.w1(32'h3aee68b7),
	.w2(32'hbab4331e),
	.w3(32'h3b1b4ec9),
	.w4(32'h3b8f622d),
	.w5(32'hbb4dd1c7),
	.w6(32'h3b016f07),
	.w7(32'hbb020c9f),
	.w8(32'hbbbeefa2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef9ad5),
	.w1(32'hbc351f84),
	.w2(32'hbc4b4021),
	.w3(32'h3b54fc58),
	.w4(32'hbc5f1310),
	.w5(32'hbc84a833),
	.w6(32'hbc102d65),
	.w7(32'hbc5b8972),
	.w8(32'hbc51f285),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43f645),
	.w1(32'hbaa701b6),
	.w2(32'hbacc60d7),
	.w3(32'h3b1996ce),
	.w4(32'hba88518f),
	.w5(32'hbbb943f5),
	.w6(32'h3b54c97b),
	.w7(32'hb9bb922d),
	.w8(32'h3a149e46),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5913db),
	.w1(32'h3b51db83),
	.w2(32'hbb1c2fdc),
	.w3(32'h3a768235),
	.w4(32'hba40a314),
	.w5(32'hbb10d0bc),
	.w6(32'h3b0182cd),
	.w7(32'h3ae51dfd),
	.w8(32'hbad91b06),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe3777),
	.w1(32'h3a35538f),
	.w2(32'h3b621cb3),
	.w3(32'hba2d2fee),
	.w4(32'hbb620197),
	.w5(32'h3a5eafd0),
	.w6(32'hbb280dbc),
	.w7(32'hbbcc0816),
	.w8(32'h3be6e145),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5611f7),
	.w1(32'hbadb945a),
	.w2(32'hba496b32),
	.w3(32'h3c5ca96b),
	.w4(32'hbb13f946),
	.w5(32'hbae01836),
	.w6(32'h3aba60b4),
	.w7(32'hbb29735b),
	.w8(32'hbb37fb97),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc0ea8),
	.w1(32'h3bd3f244),
	.w2(32'h3bb5c9e3),
	.w3(32'hbb1ea29f),
	.w4(32'h3b8fe135),
	.w5(32'h3acf2745),
	.w6(32'hba84278b),
	.w7(32'h3b84da24),
	.w8(32'h3a1d3e8d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e029),
	.w1(32'hbbf28fbe),
	.w2(32'hbba693ea),
	.w3(32'h39fd68a4),
	.w4(32'hbc0d7f2f),
	.w5(32'hbc55c443),
	.w6(32'hbb1d4cdc),
	.w7(32'hbc34e63d),
	.w8(32'hbb951f2c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c0bc4),
	.w1(32'hbbb0cc36),
	.w2(32'hbc0751cb),
	.w3(32'h3acb8dc4),
	.w4(32'hbb91f88a),
	.w5(32'hbb9bac8f),
	.w6(32'h3b4bd3b8),
	.w7(32'hbacd85da),
	.w8(32'h3b0194ac),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb822f4c),
	.w1(32'hbb139a58),
	.w2(32'h3b213b2d),
	.w3(32'h3a0e9caa),
	.w4(32'h3adc6a85),
	.w5(32'hba02ec7f),
	.w6(32'h3aad7c07),
	.w7(32'hbb3429dc),
	.w8(32'h3aa45f2e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b240673),
	.w1(32'h3b16b454),
	.w2(32'hbaa1702b),
	.w3(32'h3b94f0a9),
	.w4(32'hbac767da),
	.w5(32'h3bc54027),
	.w6(32'h389326e2),
	.w7(32'hb896ff61),
	.w8(32'h3c0678de),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26a44),
	.w1(32'hbb5076e8),
	.w2(32'hbafe3c0b),
	.w3(32'h3b8569ed),
	.w4(32'hbb35dd1b),
	.w5(32'hbbb2d7a7),
	.w6(32'h3b1ecab3),
	.w7(32'hba0761ea),
	.w8(32'hbba552c7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a927420),
	.w1(32'hbaac6903),
	.w2(32'h3a25628a),
	.w3(32'hbabf0f05),
	.w4(32'hbb296890),
	.w5(32'h3b963839),
	.w6(32'hbb79972b),
	.w7(32'hbb0a97b2),
	.w8(32'h38b8b5b5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2fa60),
	.w1(32'hbbde9430),
	.w2(32'hbbe29572),
	.w3(32'h3a1412fe),
	.w4(32'hbb516ef4),
	.w5(32'hbb527381),
	.w6(32'h3b9bfc70),
	.w7(32'hbbd316c5),
	.w8(32'hbbc367dd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37845695),
	.w1(32'h3b3a2547),
	.w2(32'h3b13a212),
	.w3(32'hbabca9b2),
	.w4(32'hba032e9d),
	.w5(32'hbbad9b88),
	.w6(32'hbc198663),
	.w7(32'hbb55fb9f),
	.w8(32'h3ac57d64),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba899dd9),
	.w1(32'h3aff92fd),
	.w2(32'h3987d57a),
	.w3(32'hbb6f2727),
	.w4(32'hbb92aac8),
	.w5(32'h3baa7178),
	.w6(32'hbaaf1121),
	.w7(32'h3b86712d),
	.w8(32'h3c3c3af5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba084fc2),
	.w1(32'hb955e93c),
	.w2(32'hbbbbab2e),
	.w3(32'h3b5aa536),
	.w4(32'hbb757ce0),
	.w5(32'hbb8be9cf),
	.w6(32'h3b778aaa),
	.w7(32'hbb6b7d99),
	.w8(32'hbaebbf90),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530d67),
	.w1(32'hbb39f601),
	.w2(32'h3a99d767),
	.w3(32'hb99ed197),
	.w4(32'hbaf55467),
	.w5(32'h3c385e10),
	.w6(32'h3aa26b30),
	.w7(32'h3a802358),
	.w8(32'h3bdabb76),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f3799),
	.w1(32'h3bae8632),
	.w2(32'h3ade6f25),
	.w3(32'h3b7efc23),
	.w4(32'h3b5069a5),
	.w5(32'h3b67ef11),
	.w6(32'hbb97a106),
	.w7(32'h3b9a2c0b),
	.w8(32'h3be0cd95),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f338c2),
	.w1(32'hbb1f4e1f),
	.w2(32'hbad7f472),
	.w3(32'h3b651039),
	.w4(32'hbafcd1e0),
	.w5(32'hbb6237d5),
	.w6(32'h3b999145),
	.w7(32'h3b4283a5),
	.w8(32'hba632615),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219d38),
	.w1(32'hbb84c2ac),
	.w2(32'hba49ae92),
	.w3(32'h3c0b480b),
	.w4(32'hbb630522),
	.w5(32'hbab29454),
	.w6(32'h3c0957b8),
	.w7(32'hbab992c5),
	.w8(32'h3b058c63),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39745c14),
	.w1(32'h3b10f847),
	.w2(32'hbb2de594),
	.w3(32'h3bbfc2fa),
	.w4(32'hbbbfaef5),
	.w5(32'hbc0dd2e2),
	.w6(32'h3b982085),
	.w7(32'hba0ca181),
	.w8(32'h3c5ac70e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9415a),
	.w1(32'hbb909327),
	.w2(32'hbb08302f),
	.w3(32'h3c2a8e97),
	.w4(32'hbc089c2d),
	.w5(32'hbb6f5417),
	.w6(32'h3c301400),
	.w7(32'hbbccb12c),
	.w8(32'h3bb4943e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13107d),
	.w1(32'hbbdab397),
	.w2(32'hbc795253),
	.w3(32'h3be6429e),
	.w4(32'hb9b930d2),
	.w5(32'h3be6b325),
	.w6(32'h3ba46bc7),
	.w7(32'hbc12c493),
	.w8(32'h38e898cf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba615f3),
	.w1(32'h3a77b0be),
	.w2(32'h3c88a8b3),
	.w3(32'h3a6aad74),
	.w4(32'h3c4ee524),
	.w5(32'h3c295f0d),
	.w6(32'h3b3ad1bb),
	.w7(32'h3c200c0c),
	.w8(32'hbc15948c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3cf94),
	.w1(32'h3c446764),
	.w2(32'h3b777bb3),
	.w3(32'hbc114592),
	.w4(32'h3c3ac2a9),
	.w5(32'hb9c241dd),
	.w6(32'hbbe2b6a8),
	.w7(32'h3baed002),
	.w8(32'hbb2f11f5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76a3e4),
	.w1(32'hbb8482cb),
	.w2(32'h3c408270),
	.w3(32'h3b40acb6),
	.w4(32'hbb271344),
	.w5(32'h3c8c39f0),
	.w6(32'h3bad4191),
	.w7(32'h3bf2c683),
	.w8(32'h3ca2ffb9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf94c90),
	.w1(32'hbb547f39),
	.w2(32'hbb920f11),
	.w3(32'h3ab7b765),
	.w4(32'hbb1cdd82),
	.w5(32'hbbf74822),
	.w6(32'h3c1fc43a),
	.w7(32'h3a3aa78c),
	.w8(32'h39f4bfb6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d84f),
	.w1(32'hbbd205d1),
	.w2(32'hbc32bb5e),
	.w3(32'h3b9094ef),
	.w4(32'hbc07660d),
	.w5(32'h3b89bf01),
	.w6(32'h3b69b471),
	.w7(32'hbc51a9f8),
	.w8(32'hbb239b5f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dbbab),
	.w1(32'hbba25669),
	.w2(32'hbb8d5e27),
	.w3(32'hbb76fa91),
	.w4(32'hbbdf54ca),
	.w5(32'h3a1174f4),
	.w6(32'hbad351fa),
	.w7(32'hbc1d27ee),
	.w8(32'hbc49d5e4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a11ea),
	.w1(32'h3c7892ef),
	.w2(32'h3c68b0df),
	.w3(32'hbb3abf6a),
	.w4(32'h3d09f4ad),
	.w5(32'hba94108f),
	.w6(32'h3bdda209),
	.w7(32'h3d147712),
	.w8(32'h3d055b2a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceab873),
	.w1(32'h3b892e0c),
	.w2(32'h3928d42d),
	.w3(32'h3cb8d288),
	.w4(32'h3afc03b7),
	.w5(32'h3c92f247),
	.w6(32'h3ce60604),
	.w7(32'hbbed427b),
	.w8(32'h3c044026),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaeeb80),
	.w1(32'h3aa73c6f),
	.w2(32'h3a273008),
	.w3(32'hb9eb58d3),
	.w4(32'hb9ccfd95),
	.w5(32'h3bb59920),
	.w6(32'h3c10d271),
	.w7(32'hbb42f1cf),
	.w8(32'hbaea0d3d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f5826),
	.w1(32'hbc5fe9cd),
	.w2(32'hbb4bad3f),
	.w3(32'h3c022f4f),
	.w4(32'hbb5aba00),
	.w5(32'hbcb6103d),
	.w6(32'h3bba653f),
	.w7(32'hbbdf1533),
	.w8(32'hbaabcd0a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0983be),
	.w1(32'hbacf34da),
	.w2(32'hbc0a8d25),
	.w3(32'h3b00d0b4),
	.w4(32'hbb96b90a),
	.w5(32'hbc83852d),
	.w6(32'h3b88fbde),
	.w7(32'h3b62f9bc),
	.w8(32'hba0a00a5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3eb5e),
	.w1(32'hbbc8ad3b),
	.w2(32'h3b1dfe9e),
	.w3(32'hbb7696d8),
	.w4(32'hbc0262de),
	.w5(32'hbb812138),
	.w6(32'hbb4dee63),
	.w7(32'hbc25ad20),
	.w8(32'hbb8f76ee),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa82b6c),
	.w1(32'hbb2d851a),
	.w2(32'h3ab4a3fb),
	.w3(32'h3b51983f),
	.w4(32'hbc05bf9a),
	.w5(32'h3ae54099),
	.w6(32'h3bf174e4),
	.w7(32'hbba0d9da),
	.w8(32'h3af640e7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2db746),
	.w1(32'hbb6150a0),
	.w2(32'h3b945710),
	.w3(32'hba7a0792),
	.w4(32'h3b50bd2a),
	.w5(32'h3cb3ff11),
	.w6(32'hba9f0882),
	.w7(32'hb97852ee),
	.w8(32'h3c7bc819),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37e40),
	.w1(32'h3be71387),
	.w2(32'h3bb5e2cf),
	.w3(32'h3c94b0b7),
	.w4(32'hbac97b8d),
	.w5(32'h3c3325cb),
	.w6(32'h3c13b0f6),
	.w7(32'hbb80957b),
	.w8(32'h3ba472f8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b86413),
	.w1(32'h3c262ace),
	.w2(32'h3bb6c602),
	.w3(32'hbac27eba),
	.w4(32'hbc516217),
	.w5(32'hbc22913a),
	.w6(32'h3c2938f3),
	.w7(32'hbbad81ba),
	.w8(32'hbc13a9f5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdfb79),
	.w1(32'h3b0e1338),
	.w2(32'hbb0a161c),
	.w3(32'hbc209eae),
	.w4(32'hb9ecfba6),
	.w5(32'hbc8bdea0),
	.w6(32'h3b04024c),
	.w7(32'h3b9ccabc),
	.w8(32'hbc381875),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8f7d1),
	.w1(32'hbb8e9220),
	.w2(32'hbc085410),
	.w3(32'h3b448b20),
	.w4(32'hbc380ceb),
	.w5(32'hbc4ac626),
	.w6(32'hbb90712c),
	.w7(32'hbae6478c),
	.w8(32'hbbad8986),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2014),
	.w1(32'h39cd1abc),
	.w2(32'h3bdccea0),
	.w3(32'hbb98118a),
	.w4(32'h3c22a392),
	.w5(32'h3b11a085),
	.w6(32'hbc3ec194),
	.w7(32'h3b6c5335),
	.w8(32'h3b575336),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b8336),
	.w1(32'hbc59233b),
	.w2(32'hbbe88e06),
	.w3(32'h3c885809),
	.w4(32'hbc38adcc),
	.w5(32'hbb338eb9),
	.w6(32'hbae7b5cd),
	.w7(32'hbc604922),
	.w8(32'hbc109609),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde70f5),
	.w1(32'h396faa5f),
	.w2(32'h3c3c4310),
	.w3(32'hbbe5d4ef),
	.w4(32'hbc0c387f),
	.w5(32'h39bd37e2),
	.w6(32'hbb4644b4),
	.w7(32'hbbd999cf),
	.w8(32'hb9f5b406),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cab7e),
	.w1(32'h3be90af1),
	.w2(32'h3a0d2a34),
	.w3(32'h3cfba2f9),
	.w4(32'hbc2e978e),
	.w5(32'hbc93ceb3),
	.w6(32'h3c3705c3),
	.w7(32'hbbeac0c5),
	.w8(32'hbcbd1f4d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb479311),
	.w1(32'hbb7a21d4),
	.w2(32'hbb125bef),
	.w3(32'hbc2973d5),
	.w4(32'hbaf45374),
	.w5(32'h3c24c1b0),
	.w6(32'hbc40d94e),
	.w7(32'hbc01dc68),
	.w8(32'hbae6b44e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0edd0a),
	.w1(32'hbaa263d8),
	.w2(32'h3c043147),
	.w3(32'h3c2ea43d),
	.w4(32'h3ba1ebad),
	.w5(32'h3bcef2b6),
	.w6(32'h3984c3d9),
	.w7(32'h3c2e334f),
	.w8(32'h3cb64abc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61cc3e),
	.w1(32'h3b5d6589),
	.w2(32'h3bfd5046),
	.w3(32'h3ab62175),
	.w4(32'hbc0fae50),
	.w5(32'hbc5b986f),
	.w6(32'h399a3f71),
	.w7(32'h3b42a0f2),
	.w8(32'hbbcf2cfe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08a332),
	.w1(32'hbc218eea),
	.w2(32'hbbc81a85),
	.w3(32'h3b85dcec),
	.w4(32'hbab4c25e),
	.w5(32'hbbf9416d),
	.w6(32'hbaa77b53),
	.w7(32'hbb04df6d),
	.w8(32'hbbc82f2f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f4ae2),
	.w1(32'h3b350068),
	.w2(32'h3b77de1e),
	.w3(32'h3b20607f),
	.w4(32'hb96d767d),
	.w5(32'hbbed27a7),
	.w6(32'hbb3034eb),
	.w7(32'h3b5436b3),
	.w8(32'h3b2503a7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba68692),
	.w1(32'h3b1ba2d8),
	.w2(32'h387d1626),
	.w3(32'hbbbd6079),
	.w4(32'h3b4d3ae2),
	.w5(32'hbc2aa48d),
	.w6(32'hb842ddea),
	.w7(32'hbb73bde6),
	.w8(32'h3ba59dc9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca4a9),
	.w1(32'h3a80059a),
	.w2(32'hb966d4e0),
	.w3(32'hbb3d6c29),
	.w4(32'hbba09308),
	.w5(32'hbc311e55),
	.w6(32'h3af5d08c),
	.w7(32'h3be3f387),
	.w8(32'hb8cf3690),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadadb12),
	.w1(32'hbb2b2dbe),
	.w2(32'hbc549b15),
	.w3(32'h3ba765c3),
	.w4(32'h3cb14989),
	.w5(32'h3c04ae44),
	.w6(32'h3c40a09b),
	.w7(32'h3b7dad50),
	.w8(32'hbb1ef0a2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31b32a),
	.w1(32'hba9df18c),
	.w2(32'hbbbc54df),
	.w3(32'hbc311c7c),
	.w4(32'h3b827554),
	.w5(32'hbb72d016),
	.w6(32'h3b7b2b5d),
	.w7(32'h3c6b1053),
	.w8(32'h3c0ff1f8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e3539),
	.w1(32'hbbcb144e),
	.w2(32'hbb7f1e5c),
	.w3(32'h3ab22304),
	.w4(32'hbb2ea0c8),
	.w5(32'h3c825aa1),
	.w6(32'h3ae9c37e),
	.w7(32'hbc045e58),
	.w8(32'h3a0f8199),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb1077),
	.w1(32'h3bbbcecb),
	.w2(32'hba68f5c0),
	.w3(32'hbbe1df30),
	.w4(32'h3c0d4712),
	.w5(32'hbb15859b),
	.w6(32'h3bb7f370),
	.w7(32'hbb2159d3),
	.w8(32'hbc678a83),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93aaa5),
	.w1(32'h3b838395),
	.w2(32'h3b9d1ce0),
	.w3(32'h3b955287),
	.w4(32'h3b9af179),
	.w5(32'h3c98443d),
	.w6(32'h3bcb4c6d),
	.w7(32'h3c087d75),
	.w8(32'h3c16961f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f510),
	.w1(32'hbc2fb498),
	.w2(32'h3b0ee40b),
	.w3(32'hbbab5f2c),
	.w4(32'h3a367b78),
	.w5(32'hbc03924b),
	.w6(32'h3bdf60be),
	.w7(32'h3b973ee7),
	.w8(32'h3be56acd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c754c9a),
	.w1(32'hbbe2e4c3),
	.w2(32'hbac445f0),
	.w3(32'h3bf3e5cd),
	.w4(32'hbc837b9b),
	.w5(32'hbc932aad),
	.w6(32'hba21e9da),
	.w7(32'hbc32944a),
	.w8(32'hbc05c851),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beef8ea),
	.w1(32'hbb418ecf),
	.w2(32'hba39015e),
	.w3(32'h3bdd6e3c),
	.w4(32'hb9d19a12),
	.w5(32'h3ba2dd75),
	.w6(32'h3bc97985),
	.w7(32'hbb9d5694),
	.w8(32'hbb546699),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc170511),
	.w1(32'hbbd60652),
	.w2(32'hbc2203a5),
	.w3(32'hbc20a243),
	.w4(32'h3b13ca34),
	.w5(32'hbbefd8f6),
	.w6(32'hbb4c5e3a),
	.w7(32'hbbf611d6),
	.w8(32'hbc5cf9ef),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7ec05),
	.w1(32'hba0ce4c7),
	.w2(32'hbaca8f4f),
	.w3(32'h3b0bf193),
	.w4(32'hbbe10a66),
	.w5(32'hbb782a48),
	.w6(32'hbbdd8efb),
	.w7(32'hbc08b18c),
	.w8(32'hbc259073),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6637be),
	.w1(32'hbbc95874),
	.w2(32'h3b8c8ba2),
	.w3(32'h3bb3ec1e),
	.w4(32'hbaac11f6),
	.w5(32'hbc840862),
	.w6(32'h3afc0603),
	.w7(32'hbc2257bd),
	.w8(32'hbaeae4a0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6b48),
	.w1(32'hbc1db77b),
	.w2(32'hbbcf6cd6),
	.w3(32'hba2de340),
	.w4(32'hbc41199f),
	.w5(32'hbc6f27de),
	.w6(32'hbc61163d),
	.w7(32'hbae9b646),
	.w8(32'hbb3e3e31),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b221eaa),
	.w1(32'h3bdacbfc),
	.w2(32'h3c20b6ee),
	.w3(32'h39d44d17),
	.w4(32'hbbf07db5),
	.w5(32'h3c7a3a63),
	.w6(32'hbb4fe2fb),
	.w7(32'hb9adf512),
	.w8(32'hbb1897dc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a9912),
	.w1(32'h3ba69d5b),
	.w2(32'hbbbdb3e3),
	.w3(32'h3a4d3b53),
	.w4(32'h3b5370ef),
	.w5(32'hbc677875),
	.w6(32'h3c062468),
	.w7(32'h3b8c337a),
	.w8(32'hba823816),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4005a2),
	.w1(32'h3bdd7760),
	.w2(32'h3aece8d8),
	.w3(32'h3b89952d),
	.w4(32'h3c26097a),
	.w5(32'h3b748e01),
	.w6(32'hba78c5d4),
	.w7(32'h3b5cb5c0),
	.w8(32'h3c41bb2f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00d1b3),
	.w1(32'hbb3c28b6),
	.w2(32'hbb2ea01a),
	.w3(32'h3c2279cf),
	.w4(32'hbc243dee),
	.w5(32'hbc024102),
	.w6(32'h3ac72ed8),
	.w7(32'hbbc45283),
	.w8(32'hbc3a8226),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e689f),
	.w1(32'h3c35f557),
	.w2(32'h3c19d63b),
	.w3(32'h3b2479ab),
	.w4(32'h3b9fabf8),
	.w5(32'h3c8a454d),
	.w6(32'hbb0df706),
	.w7(32'h3bc1d671),
	.w8(32'h3c60251a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9e05),
	.w1(32'h3b888b29),
	.w2(32'h3c655621),
	.w3(32'h3b1653fd),
	.w4(32'h3b7c2ca9),
	.w5(32'h3bb2bb00),
	.w6(32'h3c103a0d),
	.w7(32'h3b2a653e),
	.w8(32'hbb2265e1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ddd8),
	.w1(32'h3b2f7620),
	.w2(32'h3b283a83),
	.w3(32'h3c511441),
	.w4(32'h3b8bfbda),
	.w5(32'hba25141e),
	.w6(32'h3ae97487),
	.w7(32'hbaf95a99),
	.w8(32'h3a9d35a0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06bd09),
	.w1(32'h3a475308),
	.w2(32'hbc58ec31),
	.w3(32'h3bd7008b),
	.w4(32'hb9bf15ad),
	.w5(32'h3bf42d26),
	.w6(32'hbb952b31),
	.w7(32'hbb9ba2a9),
	.w8(32'hba8beb95),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c411),
	.w1(32'h3bef20b7),
	.w2(32'h3a6e81c4),
	.w3(32'h3a31ec32),
	.w4(32'h3bb839a1),
	.w5(32'hbc401f17),
	.w6(32'h3b26fd4f),
	.w7(32'h3b476887),
	.w8(32'h3ba2cf4b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a8a7),
	.w1(32'h3c35d1d0),
	.w2(32'h39d8d1dc),
	.w3(32'h37431f75),
	.w4(32'h3c1dde0e),
	.w5(32'hbbaed8d9),
	.w6(32'hbb3bd2ba),
	.w7(32'h3c29ef5b),
	.w8(32'h3c8e959d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c2ee8),
	.w1(32'hbc0afe5f),
	.w2(32'hbc6fabe3),
	.w3(32'h3c85bd2a),
	.w4(32'hbc55c73b),
	.w5(32'hbc569afe),
	.w6(32'h3c8a383b),
	.w7(32'hbc9a8dc4),
	.w8(32'hbca910ad),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3377),
	.w1(32'h3b44a93c),
	.w2(32'h3b9b61a0),
	.w3(32'hbbf0e93c),
	.w4(32'h3c372093),
	.w5(32'h3c0f2894),
	.w6(32'hbc00eda8),
	.w7(32'h3bff34c2),
	.w8(32'h3c4bd962),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67b635),
	.w1(32'hbb08bb84),
	.w2(32'hbbb42324),
	.w3(32'hbc6044db),
	.w4(32'hbc8c708a),
	.w5(32'h3ba2c94d),
	.w6(32'hbc161a18),
	.w7(32'hbc625e0b),
	.w8(32'hbc1dae59),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554043),
	.w1(32'h3c05c460),
	.w2(32'h3b02b111),
	.w3(32'hbbe15964),
	.w4(32'h3a6afb7d),
	.w5(32'h3c8c516f),
	.w6(32'hbc15ade6),
	.w7(32'hbbe2bf75),
	.w8(32'hba02fabd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc806371),
	.w1(32'h3b8bceb0),
	.w2(32'h3a0f4b14),
	.w3(32'hbb3135ec),
	.w4(32'h3ad07d5c),
	.w5(32'h3b17cba5),
	.w6(32'hb9a2ca47),
	.w7(32'h3b089f43),
	.w8(32'hbb509184),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36060e),
	.w1(32'hbc106d60),
	.w2(32'hba0def91),
	.w3(32'h3b73510b),
	.w4(32'hbc369103),
	.w5(32'hbb2329be),
	.w6(32'hbc0f34b3),
	.w7(32'hbb975fe3),
	.w8(32'hbab0c6b4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90e51f),
	.w1(32'hbb175362),
	.w2(32'hb9e7723b),
	.w3(32'hbab83796),
	.w4(32'hbbad3917),
	.w5(32'hbc856ead),
	.w6(32'h3a9f59d9),
	.w7(32'hba61983d),
	.w8(32'h3b78b123),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5f3dc),
	.w1(32'h3b70eb9d),
	.w2(32'h389d5b5c),
	.w3(32'hbc01d9fd),
	.w4(32'h3b8357e8),
	.w5(32'hbcaa9571),
	.w6(32'hbbae250b),
	.w7(32'h3c336033),
	.w8(32'h3be0643c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d3e11),
	.w1(32'h3b59ab27),
	.w2(32'hbb7cafe4),
	.w3(32'h3b4581a6),
	.w4(32'h3b0c1faa),
	.w5(32'hba8c49c4),
	.w6(32'h3bc6db40),
	.w7(32'hbaffb7cf),
	.w8(32'hbc2734f9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03fa45),
	.w1(32'h3b603747),
	.w2(32'hbb888dda),
	.w3(32'hbbd59318),
	.w4(32'hba2e8021),
	.w5(32'hbaced2b1),
	.w6(32'hbbf54177),
	.w7(32'h39f40674),
	.w8(32'h3be978fd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dbc80),
	.w1(32'h3b454f1a),
	.w2(32'hbbb6de9b),
	.w3(32'hb9b54a20),
	.w4(32'hbb8d2505),
	.w5(32'hbb9cbe79),
	.w6(32'h3b32e424),
	.w7(32'h3a4dd00b),
	.w8(32'h3a22a220),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0c05),
	.w1(32'h3982a9ae),
	.w2(32'hbb5232b7),
	.w3(32'h3bb9729c),
	.w4(32'hbba82c81),
	.w5(32'hbbc308f9),
	.w6(32'hbaaf37c9),
	.w7(32'hbb0685a0),
	.w8(32'hbb007061),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03d6f),
	.w1(32'hbaf72752),
	.w2(32'hbb975c1c),
	.w3(32'hbc12e18c),
	.w4(32'hbc176fd8),
	.w5(32'h3c477e68),
	.w6(32'h3b0905d9),
	.w7(32'hbc0c8ee2),
	.w8(32'hbc2b891b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb480e69),
	.w1(32'h3a261e49),
	.w2(32'hbbc37afa),
	.w3(32'h3ad19273),
	.w4(32'hbbcf1a3b),
	.w5(32'hbc2e169d),
	.w6(32'hbbb8b75a),
	.w7(32'hbc5f6f4b),
	.w8(32'hbc74916c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3148eb),
	.w1(32'h3bea920c),
	.w2(32'hb9dde574),
	.w3(32'h3c4b2f2f),
	.w4(32'h3bd1c488),
	.w5(32'h3bf2c9fa),
	.w6(32'h3c1266a4),
	.w7(32'h3abfb3d2),
	.w8(32'h3c20d814),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb301b4),
	.w1(32'h39fd4f0f),
	.w2(32'h3bc9ca3e),
	.w3(32'h3bb35013),
	.w4(32'hbb25e7fe),
	.w5(32'hbbb62439),
	.w6(32'h3bc634ae),
	.w7(32'h3beff9a1),
	.w8(32'hbb058cd9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09b092),
	.w1(32'hbc5b8874),
	.w2(32'hbc87175c),
	.w3(32'h3aa15007),
	.w4(32'hbc49ca5d),
	.w5(32'hbc803890),
	.w6(32'hb959dc95),
	.w7(32'hbc06a05a),
	.w8(32'hbbe3cfa8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ba1b9),
	.w1(32'h3b975bca),
	.w2(32'hbb8fde70),
	.w3(32'h3c37ee3a),
	.w4(32'h3a82e31c),
	.w5(32'hb98f7044),
	.w6(32'h3a01450e),
	.w7(32'hbb5b0010),
	.w8(32'hbc58ea47),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba06107),
	.w1(32'h3bf9a50c),
	.w2(32'h3b960fc0),
	.w3(32'h3ae19648),
	.w4(32'h3c650f01),
	.w5(32'h3b315544),
	.w6(32'hbbdb9bc8),
	.w7(32'h3bb89cf6),
	.w8(32'h3c6eac76),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47af24),
	.w1(32'hbbf0fb58),
	.w2(32'h3b589581),
	.w3(32'h3bd57cbb),
	.w4(32'hbc083b93),
	.w5(32'h3b638e35),
	.w6(32'h3cab3f81),
	.w7(32'hbb529d32),
	.w8(32'h3bdb2dee),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dca8a),
	.w1(32'hbbddec8a),
	.w2(32'hbb9ace10),
	.w3(32'hbc731dba),
	.w4(32'hbc3ff818),
	.w5(32'h3ac45b7d),
	.w6(32'hbba921f0),
	.w7(32'hbc057db8),
	.w8(32'hbbd24660),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba4052),
	.w1(32'h3b8e3554),
	.w2(32'h3c1578ee),
	.w3(32'hbb7c8c34),
	.w4(32'h3b9b83b7),
	.w5(32'h3c853b31),
	.w6(32'hbb3d7486),
	.w7(32'h3c2cd713),
	.w8(32'h3b38e09f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46d6f1),
	.w1(32'h3b146b40),
	.w2(32'hbb493e02),
	.w3(32'hbbb8fc0b),
	.w4(32'h3c10f9be),
	.w5(32'h3c07341d),
	.w6(32'h3bb23684),
	.w7(32'h3c21aabe),
	.w8(32'h3c94569d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807ab8),
	.w1(32'h3caf886f),
	.w2(32'h3cb31b30),
	.w3(32'hbc0a1cf8),
	.w4(32'h3c9b2720),
	.w5(32'h3ce23b2f),
	.w6(32'h3c4b1b5b),
	.w7(32'hbbb1be64),
	.w8(32'h3c54f0f9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ee471),
	.w1(32'h3c08c8a6),
	.w2(32'hbb364315),
	.w3(32'h3ca6ae36),
	.w4(32'h3c27a56a),
	.w5(32'hbb6a7f9d),
	.w6(32'h3c978ded),
	.w7(32'h3b2a6d1a),
	.w8(32'hbc34f227),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2145e0),
	.w1(32'h389266de),
	.w2(32'hbaec2db7),
	.w3(32'h3acecf66),
	.w4(32'h39beaf7a),
	.w5(32'h3c2d28bf),
	.w6(32'hbb3e3128),
	.w7(32'h3b92be88),
	.w8(32'h3bbb286f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada0165),
	.w1(32'h3bb9439f),
	.w2(32'h3cbdc527),
	.w3(32'h3b8011df),
	.w4(32'h3a90d555),
	.w5(32'h3c952ae7),
	.w6(32'h3c04ac6a),
	.w7(32'hbb3032f8),
	.w8(32'h3c2003ac),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf23df),
	.w1(32'hbc3c377e),
	.w2(32'hbbf63335),
	.w3(32'h3c680dab),
	.w4(32'hbbbb3528),
	.w5(32'hbb507342),
	.w6(32'h3cb272b6),
	.w7(32'hbc36fdea),
	.w8(32'hbc1dc1df),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada8fa4),
	.w1(32'hbb3b830a),
	.w2(32'h3c82e196),
	.w3(32'hbb5da23f),
	.w4(32'h3b0979b5),
	.w5(32'h3c2746cc),
	.w6(32'hbc1ff33b),
	.w7(32'h3b0108a1),
	.w8(32'hbb179467),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98f800),
	.w1(32'hbb2e7caa),
	.w2(32'hbc3b71f1),
	.w3(32'hbc5d6000),
	.w4(32'h3adc81f8),
	.w5(32'h3ac041f8),
	.w6(32'hbba69d7d),
	.w7(32'hbb1f357a),
	.w8(32'hbb7e0607),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37cff0),
	.w1(32'hbc403f18),
	.w2(32'hbbada1de),
	.w3(32'h3c52ab7f),
	.w4(32'hbc191c1a),
	.w5(32'hbc61be44),
	.w6(32'hbc42b7e2),
	.w7(32'hbc321347),
	.w8(32'hbc818840),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a189),
	.w1(32'hbcc2af7b),
	.w2(32'hbaddb45b),
	.w3(32'hbc16baa2),
	.w4(32'hbcf6aab4),
	.w5(32'hbc20c94e),
	.w6(32'hbc13b4cf),
	.w7(32'hbcaacfde),
	.w8(32'hbc63d863),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e65f1),
	.w1(32'hb99accc7),
	.w2(32'h39737fea),
	.w3(32'h394d7973),
	.w4(32'h3bcb3425),
	.w5(32'h3c7e1f39),
	.w6(32'hbc13f09d),
	.w7(32'hbbcf19b0),
	.w8(32'h3b34cee6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6bc22),
	.w1(32'hbb8c63a9),
	.w2(32'h3b6ea060),
	.w3(32'hbc1f54ec),
	.w4(32'h3bd651d9),
	.w5(32'h3aba89d3),
	.w6(32'hbbf26e42),
	.w7(32'h3c216bdb),
	.w8(32'h3b05cf72),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becec4f),
	.w1(32'hbb79ca96),
	.w2(32'hbc20578a),
	.w3(32'hbbee5d60),
	.w4(32'hbbd49705),
	.w5(32'hbc6dd1a2),
	.w6(32'hbbefa361),
	.w7(32'h391ea28a),
	.w8(32'hbc704f22),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba68d06),
	.w1(32'hbba83f91),
	.w2(32'h3bbd0bbd),
	.w3(32'hbc2d551b),
	.w4(32'h3c05ee7f),
	.w5(32'h3c29c009),
	.w6(32'hbc13cca3),
	.w7(32'h3c408806),
	.w8(32'h3bef93c0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c914f86),
	.w1(32'hbbb59b81),
	.w2(32'hb9c6cfbf),
	.w3(32'h3bb09785),
	.w4(32'hba755d87),
	.w5(32'h3be5be92),
	.w6(32'hbbdd267a),
	.w7(32'hbc23f34e),
	.w8(32'hbb6dd3eb),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97a358),
	.w1(32'h3c55bb4b),
	.w2(32'h3b997193),
	.w3(32'hbb9865b6),
	.w4(32'h3ca9caba),
	.w5(32'h3c32f21f),
	.w6(32'hbad8e12c),
	.w7(32'hbb4ed2d4),
	.w8(32'hbbee7155),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6d70),
	.w1(32'h3bcc37ff),
	.w2(32'h3c09214b),
	.w3(32'h3c9cd2f0),
	.w4(32'h3b592e07),
	.w5(32'h3bfa56cc),
	.w6(32'h3b55651c),
	.w7(32'hb99d09f4),
	.w8(32'h3b21be3b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835b74),
	.w1(32'h3b241611),
	.w2(32'hbb37e38b),
	.w3(32'h3c222528),
	.w4(32'hbb5cdb1d),
	.w5(32'hbc5d4455),
	.w6(32'h3ba4ad16),
	.w7(32'h3b698e97),
	.w8(32'hbc139b5c),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb825ff4),
	.w1(32'h3b81d316),
	.w2(32'hbbb833e5),
	.w3(32'h3bc02c2d),
	.w4(32'h39bcee8b),
	.w5(32'hbba94a1c),
	.w6(32'h3b8829e6),
	.w7(32'h3aacf8fe),
	.w8(32'hb8591703),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eaf62),
	.w1(32'h3bca258d),
	.w2(32'h3b9f668f),
	.w3(32'h3c015a93),
	.w4(32'hbae35f61),
	.w5(32'h3b92017a),
	.w6(32'h387fcde1),
	.w7(32'h3b84aeca),
	.w8(32'h3c235414),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e36a2),
	.w1(32'h3b5b2b6c),
	.w2(32'h3b46d206),
	.w3(32'hbae45617),
	.w4(32'h3c0ec0c9),
	.w5(32'hbb9cfcb1),
	.w6(32'hbba6813e),
	.w7(32'h3a2569c5),
	.w8(32'hbae95931),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28c033),
	.w1(32'hbbde153b),
	.w2(32'hbc2450e6),
	.w3(32'h3c0bf077),
	.w4(32'hbc7c0e6c),
	.w5(32'hbc20c86d),
	.w6(32'hbb562814),
	.w7(32'hbc202624),
	.w8(32'hbbff158b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078ad3),
	.w1(32'h3b292772),
	.w2(32'h3b90cd0c),
	.w3(32'hbaf35fbe),
	.w4(32'hbc3e1fe2),
	.w5(32'hbae04b75),
	.w6(32'hbbc659ec),
	.w7(32'hbc2a0a98),
	.w8(32'hbbb81b64),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4afdcd),
	.w1(32'hbbbf3c8b),
	.w2(32'hbbcf874b),
	.w3(32'h3b99702e),
	.w4(32'h3a9c5d8e),
	.w5(32'hbca6a5eb),
	.w6(32'h3b3b5d50),
	.w7(32'h3c0c797e),
	.w8(32'h3b6a0dc6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43dfa3),
	.w1(32'hba518a4c),
	.w2(32'hb9fed7d0),
	.w3(32'hbb0ebb2c),
	.w4(32'hbb8b5648),
	.w5(32'hbb416cb4),
	.w6(32'hbb86c30e),
	.w7(32'hbade26ae),
	.w8(32'hbbe62ce9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c002e),
	.w1(32'hbb5181d3),
	.w2(32'hbbcec991),
	.w3(32'h3bded405),
	.w4(32'h3be2c54d),
	.w5(32'hbbc156dd),
	.w6(32'h3b80d143),
	.w7(32'h3bbf95c1),
	.w8(32'h3bc34aae),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f88b83),
	.w1(32'hba858d1b),
	.w2(32'hbb3afd50),
	.w3(32'hbb94ca4e),
	.w4(32'hbb8cf411),
	.w5(32'hba91aeea),
	.w6(32'h3c27efcd),
	.w7(32'hbbf29d7f),
	.w8(32'hbbbe1938),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b1751),
	.w1(32'hbb08e54f),
	.w2(32'h3b488cc0),
	.w3(32'hbbb4aa17),
	.w4(32'hbb26b9b8),
	.w5(32'h3b3b9ecd),
	.w6(32'hba82501d),
	.w7(32'h39e773bf),
	.w8(32'h3b3043f0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde7063),
	.w1(32'h3b643135),
	.w2(32'hbc007a37),
	.w3(32'h3ac153a6),
	.w4(32'h3bd52950),
	.w5(32'hbc5686d5),
	.w6(32'h39eabde4),
	.w7(32'h3c24a1b3),
	.w8(32'h396cb049),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba05d3c),
	.w1(32'hbb0b24a0),
	.w2(32'hbb970fb2),
	.w3(32'h3b1e4447),
	.w4(32'hbbf1c75a),
	.w5(32'h3b294a6a),
	.w6(32'h3bda891f),
	.w7(32'hbb0b90af),
	.w8(32'h3bd8b9cf),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7e31a),
	.w1(32'h3be82abe),
	.w2(32'h3bb88cb4),
	.w3(32'hba3538b0),
	.w4(32'h3cab20a6),
	.w5(32'h3cd84d16),
	.w6(32'hbbcff767),
	.w7(32'h3c2fc5c2),
	.w8(32'h3ca9b398),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2052c1),
	.w1(32'hbbe61a7d),
	.w2(32'hbbb1c7e6),
	.w3(32'hb9c90c2b),
	.w4(32'hbc1226ba),
	.w5(32'hbcca322a),
	.w6(32'h3ca773b8),
	.w7(32'hbc550617),
	.w8(32'hbc4da640),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24d964),
	.w1(32'h3b5b5ff4),
	.w2(32'hbba4e508),
	.w3(32'hbc4e8191),
	.w4(32'hbb6221c1),
	.w5(32'hbc2a9b5a),
	.w6(32'hbc53ee6e),
	.w7(32'hbb799835),
	.w8(32'h3af0a97f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb27e33),
	.w1(32'hb9326d94),
	.w2(32'h3c3bdcb0),
	.w3(32'hbbdc0a1b),
	.w4(32'hbbbb69d7),
	.w5(32'h3af8e87a),
	.w6(32'hba6da913),
	.w7(32'h3a1f9524),
	.w8(32'hbc652a87),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25d5ea),
	.w1(32'h3c0d7a78),
	.w2(32'h3c148ad1),
	.w3(32'h3be5888d),
	.w4(32'h3be3786e),
	.w5(32'h3b38ae21),
	.w6(32'h39a04f25),
	.w7(32'h3b107d88),
	.w8(32'hbb808d04),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cf404),
	.w1(32'hbbaba425),
	.w2(32'hbbf28d65),
	.w3(32'h3beef6da),
	.w4(32'hbb2d728c),
	.w5(32'hbba24d66),
	.w6(32'hba0b189a),
	.w7(32'hbafb5c88),
	.w8(32'hbbad7299),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a9f14),
	.w1(32'h3c1f9ed4),
	.w2(32'h3bec7541),
	.w3(32'hbc8ddca5),
	.w4(32'h3c5ab650),
	.w5(32'h3b29e900),
	.w6(32'hbc23e253),
	.w7(32'hbb3c77c6),
	.w8(32'h3b879db2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b8a83),
	.w1(32'h3b175a94),
	.w2(32'h3b04ef2b),
	.w3(32'h3c06a177),
	.w4(32'hbad366a3),
	.w5(32'h3c581854),
	.w6(32'h3c5cdd6f),
	.w7(32'hbb8f9e27),
	.w8(32'hbb55fba0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ba57),
	.w1(32'h3b9cd6c7),
	.w2(32'h3ba59f73),
	.w3(32'h3bae773e),
	.w4(32'h3b397eb0),
	.w5(32'h39534dd6),
	.w6(32'h3883e13f),
	.w7(32'h3a4b75a8),
	.w8(32'h3b63a89d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c618d91),
	.w1(32'hbb698b6e),
	.w2(32'h39ae4240),
	.w3(32'h3b5b0c86),
	.w4(32'hbc5aede4),
	.w5(32'hbb69a0e9),
	.w6(32'hbb3a9895),
	.w7(32'hbbac3614),
	.w8(32'hbb786d13),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24d0ce),
	.w1(32'h3b738112),
	.w2(32'hbb5208ee),
	.w3(32'hb9472cac),
	.w4(32'h3a82cea3),
	.w5(32'h3c13e196),
	.w6(32'hba598e6f),
	.w7(32'h3b47dda9),
	.w8(32'h3b01fc2e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39796),
	.w1(32'h3a8aac31),
	.w2(32'hbc14e886),
	.w3(32'hbb83d9cd),
	.w4(32'h3b9d993b),
	.w5(32'hbb999f57),
	.w6(32'hbb478cac),
	.w7(32'hbb66c62a),
	.w8(32'hbbcb8922),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c32e5),
	.w1(32'hbc0cb7df),
	.w2(32'hbc5f7763),
	.w3(32'hbc9ab8a1),
	.w4(32'h39829b8c),
	.w5(32'h3b0a195e),
	.w6(32'hbc669b61),
	.w7(32'hba7350ca),
	.w8(32'hbc452dad),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8412d),
	.w1(32'hbb731e5c),
	.w2(32'h3a99853a),
	.w3(32'hbb9b35e9),
	.w4(32'h3980fd52),
	.w5(32'h3bc6cc06),
	.w6(32'h3bb74767),
	.w7(32'h3adaa043),
	.w8(32'h3c023645),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc80d75),
	.w1(32'hbc466896),
	.w2(32'hbb88063b),
	.w3(32'h3ba3d61f),
	.w4(32'hbcfeb747),
	.w5(32'hbcf0d47a),
	.w6(32'h3c28737c),
	.w7(32'hbcba7ba0),
	.w8(32'hbcb9b655),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00deac),
	.w1(32'h3ad814ba),
	.w2(32'hbb8b38b3),
	.w3(32'hbb99785f),
	.w4(32'h39fc62ac),
	.w5(32'hbb82cfc2),
	.w6(32'hbc5da1eb),
	.w7(32'h3c0cf3e3),
	.w8(32'hbb83a52b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacff7e),
	.w1(32'hbb2f7072),
	.w2(32'hbac52cd0),
	.w3(32'hbb9dd0d5),
	.w4(32'hbc122cbd),
	.w5(32'hbc8f703e),
	.w6(32'hbc50099e),
	.w7(32'hbba17d81),
	.w8(32'hbc204609),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73741),
	.w1(32'hbc74b6bc),
	.w2(32'hbc9fe993),
	.w3(32'h3c4f4ba6),
	.w4(32'hbbd3e8d1),
	.w5(32'hbc5d6cf9),
	.w6(32'hbad1aad0),
	.w7(32'hbb998caf),
	.w8(32'hbb89ea73),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b680e),
	.w1(32'h3c16ff64),
	.w2(32'hbb3f003e),
	.w3(32'hbb82fcbc),
	.w4(32'h3b9be113),
	.w5(32'hbbc05e32),
	.w6(32'hbbf91fb5),
	.w7(32'h3c759f47),
	.w8(32'h3c80bba0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2df71),
	.w1(32'hba1c5407),
	.w2(32'hbb9a37c6),
	.w3(32'h3b21c548),
	.w4(32'hb9086e74),
	.w5(32'hbb60e91c),
	.w6(32'h3c0f4a41),
	.w7(32'h3ae9a494),
	.w8(32'h3a8fb434),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1c103),
	.w1(32'hbbc6a8c9),
	.w2(32'hbbf81070),
	.w3(32'hba209e1c),
	.w4(32'h3b494428),
	.w5(32'hbbd59cfa),
	.w6(32'hbb8f3d02),
	.w7(32'hbb28937e),
	.w8(32'hbbd224c5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af23a50),
	.w1(32'hbabeb462),
	.w2(32'h3c116d22),
	.w3(32'h3b900866),
	.w4(32'hbab7a3fe),
	.w5(32'hbc619b4b),
	.w6(32'hbc008578),
	.w7(32'hbbfb4236),
	.w8(32'hbbd0f1c5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42b056),
	.w1(32'h3acde525),
	.w2(32'h3caff6ef),
	.w3(32'h3b44f7ce),
	.w4(32'hbbb209aa),
	.w5(32'hb9f82734),
	.w6(32'hbb94ae88),
	.w7(32'hbb9d2ff5),
	.w8(32'h3bad7660),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14a681),
	.w1(32'h3b838769),
	.w2(32'hb95da718),
	.w3(32'h3cb0db51),
	.w4(32'hbc202ac5),
	.w5(32'hbc60768b),
	.w6(32'h3c281fb7),
	.w7(32'h3c03822a),
	.w8(32'h3bbcffee),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad87f3),
	.w1(32'h3c315870),
	.w2(32'h38dfb57c),
	.w3(32'h3bab0151),
	.w4(32'hbb36ab13),
	.w5(32'hbc3f76c5),
	.w6(32'h3bf4d7c0),
	.w7(32'hbba4265b),
	.w8(32'hbc1f39cb),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c606a10),
	.w1(32'h3ad2e90e),
	.w2(32'hbc52748e),
	.w3(32'h3c522d11),
	.w4(32'h3abde890),
	.w5(32'hbbd78120),
	.w6(32'h3c432215),
	.w7(32'hba600c83),
	.w8(32'hbc58823c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc160a21),
	.w1(32'hba1dccc9),
	.w2(32'hbb990acd),
	.w3(32'hbb8ace05),
	.w4(32'h3bcaea1b),
	.w5(32'h3d4897af),
	.w6(32'hbb8b9cc8),
	.w7(32'hbc16cd13),
	.w8(32'hbc9f9b95),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c37d6),
	.w1(32'h3b816fae),
	.w2(32'h3c23f600),
	.w3(32'h3be01e64),
	.w4(32'hbb9924ab),
	.w5(32'h3ba480c7),
	.w6(32'hbb1d51a1),
	.w7(32'h3ad6cf95),
	.w8(32'hb9e855b3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d1f2f),
	.w1(32'hbb6aa193),
	.w2(32'hbb569dc2),
	.w3(32'hbb5ff14a),
	.w4(32'h3a72d888),
	.w5(32'hbb6f7420),
	.w6(32'hb9b613b3),
	.w7(32'hbbed4712),
	.w8(32'hba34ab61),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c150ab5),
	.w1(32'h3c024b41),
	.w2(32'hbb828b10),
	.w3(32'h3c38d831),
	.w4(32'hbb1fb419),
	.w5(32'hbb1f437a),
	.w6(32'h3bf6fae4),
	.w7(32'hbb416189),
	.w8(32'h3b197ef5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c447676),
	.w1(32'hbb74c8ef),
	.w2(32'hbc4f206d),
	.w3(32'h3b3247b3),
	.w4(32'h3c52d53b),
	.w5(32'h3cd6ed61),
	.w6(32'h3a98bb2b),
	.w7(32'hbba948b5),
	.w8(32'hbc5e0da9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7be9f),
	.w1(32'h3b93c2b8),
	.w2(32'h3aa47a03),
	.w3(32'h3ae820ae),
	.w4(32'h3c11b32f),
	.w5(32'hbc105db4),
	.w6(32'hbbe5ac92),
	.w7(32'h3c0568ef),
	.w8(32'h3be1a120),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3ba03),
	.w1(32'hbbde323b),
	.w2(32'h3c1b5796),
	.w3(32'hba0cf5cc),
	.w4(32'hbaf82c0c),
	.w5(32'hbcd1bf6e),
	.w6(32'h3b80643b),
	.w7(32'h3bfd4cd3),
	.w8(32'h3c9ca0a0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b973864),
	.w1(32'hbb77d1ba),
	.w2(32'hbacbbfd4),
	.w3(32'hbbe291a2),
	.w4(32'hbb04ab25),
	.w5(32'hbc0761fb),
	.w6(32'h3bc0ea50),
	.w7(32'hbb9ad018),
	.w8(32'h39ddd334),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1be996),
	.w1(32'hba5ce549),
	.w2(32'h3bb4c1de),
	.w3(32'h3acc2424),
	.w4(32'h3a5a88dc),
	.w5(32'hbb17b8ea),
	.w6(32'h3bbc2786),
	.w7(32'hbb5c7f79),
	.w8(32'hbaf55e71),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c978af3),
	.w1(32'h3c4a4f2c),
	.w2(32'h3bc6586c),
	.w3(32'h3c4564d4),
	.w4(32'h3b392063),
	.w5(32'hbb036977),
	.w6(32'h3be04613),
	.w7(32'h386ccae0),
	.w8(32'hbb09a7b1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4447d1),
	.w1(32'h39e27b73),
	.w2(32'h3b7b350c),
	.w3(32'h3b793f54),
	.w4(32'h3b6a513c),
	.w5(32'h3b2c0cb1),
	.w6(32'h3ae587e5),
	.w7(32'hb9392ffa),
	.w8(32'h3ac7783d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad8ff2),
	.w1(32'hb99b4ae7),
	.w2(32'hbc04f18a),
	.w3(32'hba2ecd37),
	.w4(32'hbb8197ca),
	.w5(32'h3b8ef980),
	.w6(32'h3a8a396f),
	.w7(32'hbb5faa4f),
	.w8(32'hbc1059ac),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28068e),
	.w1(32'hbb222265),
	.w2(32'hbba8c9e8),
	.w3(32'h3bc2b5b9),
	.w4(32'hbb260095),
	.w5(32'h3a538edb),
	.w6(32'hbae20ddb),
	.w7(32'hbb833ce6),
	.w8(32'hbc1fd65f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57116a),
	.w1(32'hbb82cf84),
	.w2(32'hb88a62f8),
	.w3(32'h3c124b5f),
	.w4(32'hbb3fa8c0),
	.w5(32'h3c113018),
	.w6(32'h3b900a48),
	.w7(32'hbb4ef5ba),
	.w8(32'hbbbdc037),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff2de9),
	.w1(32'hbad0535e),
	.w2(32'hbc07f8be),
	.w3(32'h3c2c435f),
	.w4(32'h3b7e8d74),
	.w5(32'h3b5afc6f),
	.w6(32'h3b28eabc),
	.w7(32'hbb946717),
	.w8(32'hbc5c9728),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bde236),
	.w1(32'hbbc81f29),
	.w2(32'h3ba6601a),
	.w3(32'h3bdd1841),
	.w4(32'h3b45cd0b),
	.w5(32'hbc5fcffb),
	.w6(32'h3bc34bc4),
	.w7(32'h39bdeb71),
	.w8(32'h3bbb1d51),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a818dbc),
	.w1(32'hbbdf3ca6),
	.w2(32'h3c0adf99),
	.w3(32'hbbae2ed0),
	.w4(32'hbbb20077),
	.w5(32'hbb9ffede),
	.w6(32'h3b1ae556),
	.w7(32'h3c222db1),
	.w8(32'h3ce3f192),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6e346),
	.w1(32'h3987942c),
	.w2(32'hbaa29966),
	.w3(32'hbc3d7f2c),
	.w4(32'hbad24e0a),
	.w5(32'hbb56f115),
	.w6(32'h3c627642),
	.w7(32'h3b2a2878),
	.w8(32'h3a0df3c4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80f62),
	.w1(32'hbc63fa62),
	.w2(32'hbc29f82d),
	.w3(32'hbb9fb386),
	.w4(32'hbbb78044),
	.w5(32'hbcb9fe87),
	.w6(32'hbb9e3fce),
	.w7(32'hbc12570f),
	.w8(32'hbc60407c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30afb7),
	.w1(32'hbbb60211),
	.w2(32'hbc8e8178),
	.w3(32'h3bef1844),
	.w4(32'hbc55f085),
	.w5(32'hbc934c55),
	.w6(32'h3b7c5c27),
	.w7(32'hbc3d02e8),
	.w8(32'hbc806ba9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20f2fd),
	.w1(32'hbc0e7de3),
	.w2(32'hbc1d5f34),
	.w3(32'h3b9cc86c),
	.w4(32'hbb51ce9a),
	.w5(32'hbbcfdd6a),
	.w6(32'hba2002d1),
	.w7(32'hbc607637),
	.w8(32'hbc98556b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba571776),
	.w1(32'h3ba80ced),
	.w2(32'hbbb88bfb),
	.w3(32'hb9fb6076),
	.w4(32'h3c0da183),
	.w5(32'h3d60e392),
	.w6(32'hbbf008d1),
	.w7(32'hbc5aa042),
	.w8(32'hbcb8d0b4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460622),
	.w1(32'h3c294539),
	.w2(32'h3c351360),
	.w3(32'h3b99f772),
	.w4(32'h3ba29e33),
	.w5(32'h3c9d6957),
	.w6(32'hbcac4cce),
	.w7(32'hbc0c1489),
	.w8(32'hbc243bd3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ffc8),
	.w1(32'hbb21a9e8),
	.w2(32'h39a001e6),
	.w3(32'h3bb3402d),
	.w4(32'hbb85d33b),
	.w5(32'hbaa50c55),
	.w6(32'hbbe73900),
	.w7(32'hbb86b2f7),
	.w8(32'hbbe7d15b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcaa87),
	.w1(32'hba91a8af),
	.w2(32'hba5d02ef),
	.w3(32'h3bf8eed2),
	.w4(32'hbba49f32),
	.w5(32'hbc9ec95c),
	.w6(32'h3b65f1d6),
	.w7(32'hbb366683),
	.w8(32'hbb1056da),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022fcd),
	.w1(32'h39efee2f),
	.w2(32'h3b4364db),
	.w3(32'h3ad07de3),
	.w4(32'h3b56c7ce),
	.w5(32'hbc4a6526),
	.w6(32'h3b8abbc3),
	.w7(32'hba5d37d0),
	.w8(32'h39826575),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a708b),
	.w1(32'h3b43fabc),
	.w2(32'hbbec2062),
	.w3(32'h3870d4f0),
	.w4(32'h3c121a96),
	.w5(32'hbb37f848),
	.w6(32'h3b52795d),
	.w7(32'hbb97b5cf),
	.w8(32'hbb583fce),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5434b7),
	.w1(32'hbb789806),
	.w2(32'hbacd155c),
	.w3(32'hbc1c98bb),
	.w4(32'hbbf4d311),
	.w5(32'hbbd1a25b),
	.w6(32'hbb4311f6),
	.w7(32'hbaab80cd),
	.w8(32'hbbf29ce5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d25de),
	.w1(32'hbc5da498),
	.w2(32'hbc06ae76),
	.w3(32'h3c141656),
	.w4(32'hbc0795a8),
	.w5(32'hbc8e7bc5),
	.w6(32'h3bf43215),
	.w7(32'hbc0657cd),
	.w8(32'hba91abf4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a53d9),
	.w1(32'hbb8bb22b),
	.w2(32'hbb1b1463),
	.w3(32'hbbd83a2c),
	.w4(32'h3aab2c95),
	.w5(32'h3bc5c3ab),
	.w6(32'h3bbeaa9a),
	.w7(32'h3b2f844d),
	.w8(32'h3b4c811b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8684a9),
	.w1(32'h3bf57fd0),
	.w2(32'h3ba3e098),
	.w3(32'h3ac3d580),
	.w4(32'hbbf8429c),
	.w5(32'h3c0a36b7),
	.w6(32'hba612bfc),
	.w7(32'hbb9e8ac6),
	.w8(32'hbb115dda),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835b52),
	.w1(32'hbbdbf698),
	.w2(32'h3b0c3153),
	.w3(32'h3bc2ec8d),
	.w4(32'hbc9706cb),
	.w5(32'hbcc845da),
	.w6(32'hb96fe0f0),
	.w7(32'hbaaa1db2),
	.w8(32'h3bef4771),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12a72a),
	.w1(32'hbc88b7e6),
	.w2(32'hba0c6857),
	.w3(32'hbb503b31),
	.w4(32'hbc0001b2),
	.w5(32'hbc95d66d),
	.w6(32'h3c21006c),
	.w7(32'hbbabcac6),
	.w8(32'hbb04b3ed),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f52c5),
	.w1(32'hbb940cde),
	.w2(32'hbc71b2c1),
	.w3(32'hbbd1ebab),
	.w4(32'hba715476),
	.w5(32'h3d48b222),
	.w6(32'hbb26fc5a),
	.w7(32'hbaacbc55),
	.w8(32'hbc7677d5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3e0d7),
	.w1(32'hbbc5c128),
	.w2(32'hbba74e59),
	.w3(32'h3c10e005),
	.w4(32'hbb527955),
	.w5(32'h3b82f4b9),
	.w6(32'hbb7390a4),
	.w7(32'hbb349b17),
	.w8(32'h3ae578f8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2af94c),
	.w1(32'hbae2d3c0),
	.w2(32'hb9daa4c6),
	.w3(32'h3bbc92bd),
	.w4(32'hb99952ae),
	.w5(32'h39ddd890),
	.w6(32'h3b86ec81),
	.w7(32'hbacce1b5),
	.w8(32'hbb4ac49e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7e2d4),
	.w1(32'hbae2821e),
	.w2(32'hbbeb7a93),
	.w3(32'hbb3e0637),
	.w4(32'h3a8aeb8b),
	.w5(32'h3b859f24),
	.w6(32'h3a3ce2b5),
	.w7(32'hbb2ecef3),
	.w8(32'hbc17b697),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd3013),
	.w1(32'h3aac6447),
	.w2(32'hbbfc84e3),
	.w3(32'hbae1b39a),
	.w4(32'h3ba0dacb),
	.w5(32'h3d77f2d2),
	.w6(32'hbbe363fa),
	.w7(32'hbbb83a15),
	.w8(32'hbc9ca1aa),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2c991),
	.w1(32'hbbacbef0),
	.w2(32'hbcaf08c7),
	.w3(32'h3c31694a),
	.w4(32'hbbc3407d),
	.w5(32'h3d303f4a),
	.w6(32'hbaa2b37f),
	.w7(32'hba4a4ab0),
	.w8(32'hbc09c961),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74553),
	.w1(32'hbbeb5922),
	.w2(32'hbbc081e6),
	.w3(32'hbaba08ee),
	.w4(32'hbafd3e68),
	.w5(32'h3bd72e82),
	.w6(32'hbbd3235d),
	.w7(32'hba3c149f),
	.w8(32'h3ad96ff5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390e21),
	.w1(32'hbbab4921),
	.w2(32'hb95bbc01),
	.w3(32'h3b06a65d),
	.w4(32'hbbd867b8),
	.w5(32'hbbbcacc6),
	.w6(32'hbb34cffa),
	.w7(32'hbb67a54f),
	.w8(32'hbbc72b0e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392323e8),
	.w1(32'h3a4f9f34),
	.w2(32'h3b132b52),
	.w3(32'h3b9933fc),
	.w4(32'hbc7e6f2b),
	.w5(32'hbd037b30),
	.w6(32'h3ab52fb0),
	.w7(32'h3b8e518a),
	.w8(32'h3cbd2526),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf769),
	.w1(32'hbc85e9d0),
	.w2(32'hbce2cbd4),
	.w3(32'hba89c83f),
	.w4(32'hbb018ed7),
	.w5(32'h3c770111),
	.w6(32'h3c32e6d8),
	.w7(32'hbc9e161b),
	.w8(32'hbc68b132),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18aee0),
	.w1(32'hbaa5e905),
	.w2(32'hbb50940c),
	.w3(32'hb8c135e8),
	.w4(32'hba5916c1),
	.w5(32'h3b838f74),
	.w6(32'h3bdd6c2c),
	.w7(32'hbbd8e680),
	.w8(32'hbbd7b664),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046a6c),
	.w1(32'h3b626ebd),
	.w2(32'hbace66b3),
	.w3(32'h3bad4bf5),
	.w4(32'h3bdce0b0),
	.w5(32'hbb846156),
	.w6(32'hb9ee40a6),
	.w7(32'h3c20b066),
	.w8(32'h3ba37df2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab67d73),
	.w1(32'h3a1bab91),
	.w2(32'hbc45e8ed),
	.w3(32'hbb6f74fc),
	.w4(32'h3b3ad8a7),
	.w5(32'h3c5b18f5),
	.w6(32'h3b584434),
	.w7(32'h3b09f822),
	.w8(32'hbc085d5c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656780),
	.w1(32'h3c85098c),
	.w2(32'h3c23ba29),
	.w3(32'h3bf8d102),
	.w4(32'hbb01e11f),
	.w5(32'h3cc0d4dc),
	.w6(32'hbc2bfdb4),
	.w7(32'hbc6a8011),
	.w8(32'hbccd2dfd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33f8a7),
	.w1(32'hbc82f753),
	.w2(32'hbb9b733f),
	.w3(32'h3b4a5c3f),
	.w4(32'hbc47f26d),
	.w5(32'hbbc96a49),
	.w6(32'hbc42d8cc),
	.w7(32'hbc55cd7c),
	.w8(32'h3c37541d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61c955),
	.w1(32'hbb583e58),
	.w2(32'hbb954c98),
	.w3(32'hbc2d2195),
	.w4(32'hbc223866),
	.w5(32'hbbcdeb90),
	.w6(32'hbb90ba00),
	.w7(32'hbba65dfb),
	.w8(32'hbba18e5d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc174c41),
	.w1(32'h3a8a9d96),
	.w2(32'hbb6860c2),
	.w3(32'h3abf3a06),
	.w4(32'h3bab431d),
	.w5(32'hbb9c8071),
	.w6(32'hbb8a5538),
	.w7(32'h387cc237),
	.w8(32'hbb0d1f08),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab56867),
	.w1(32'hbba26dc2),
	.w2(32'hbbf435d2),
	.w3(32'hbae613c0),
	.w4(32'hbbf8c701),
	.w5(32'h3b79c079),
	.w6(32'hba1c16d1),
	.w7(32'hbadf4fb9),
	.w8(32'hbae08634),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc031512),
	.w1(32'h3b032c4f),
	.w2(32'h3b8dc21f),
	.w3(32'hbb3b6795),
	.w4(32'hbbfe3ea8),
	.w5(32'hbcd509d9),
	.w6(32'hbb7ed96d),
	.w7(32'h3b9143cd),
	.w8(32'h3c0a4287),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3d33),
	.w1(32'h3ac385e6),
	.w2(32'h3b910bf3),
	.w3(32'hbb27a960),
	.w4(32'h3b4defb4),
	.w5(32'h3be974bd),
	.w6(32'h3b257c27),
	.w7(32'hba2099cd),
	.w8(32'hbc1de9c3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26f535),
	.w1(32'hba8752b8),
	.w2(32'hbb97ea0e),
	.w3(32'h3bdbc7a5),
	.w4(32'h3b00ce4d),
	.w5(32'h3d907baf),
	.w6(32'hbc17083e),
	.w7(32'hbbf5d4b5),
	.w8(32'hbc9140d6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ae1c2),
	.w1(32'hbb9cde97),
	.w2(32'hbc468969),
	.w3(32'h3ba34efc),
	.w4(32'hbc00c650),
	.w5(32'h3d1eaa2a),
	.w6(32'hbb388b63),
	.w7(32'hbc66798a),
	.w8(32'hbba79b5a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc240284),
	.w1(32'hbc1224c5),
	.w2(32'hbbbe695b),
	.w3(32'h3b7b6405),
	.w4(32'hbb31772b),
	.w5(32'hbb6a2f13),
	.w6(32'h3b58c9eb),
	.w7(32'hbc1b3e20),
	.w8(32'hbc13ff73),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac93da3),
	.w1(32'h3b8b155d),
	.w2(32'h3b05ed4a),
	.w3(32'hba714b73),
	.w4(32'hbab54dbe),
	.w5(32'hba46ac6b),
	.w6(32'hbc2eab03),
	.w7(32'h3b2c8df6),
	.w8(32'h39244187),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule