module Layer_1(data_in, valid_in, data_out, valid_out, Clk, Rst, En);
    parameter DATA_WIDTH = 8;

    input Clk, Rst, En, valid_in;
    input [DATA_WIDTH - 1:0] data_in;
    output valid_out;
    output [DATA_WIDTH - 1:0] data_out;

    wire    Conv_valid_out0, Conv_valid_out1, Conv_valid_out2, Conv_valid_out3, Conv_valid_out4, Conv_valid_out5, Conv_valid_out6, 
            Conv_valid_out7, Conv_valid_out8, Conv_valid_out9, Conv_valid_out10, Conv_valid_out11, Conv_valid_out12, Conv_valid_out13, 
            Conv_valid_out14, Conv_valid_out15, Conv_valid_out16, Conv_valid_out17, Conv_valid_out18, Conv_valid_out19, Conv_valid_out20, 
            Conv_valid_out21, Conv_valid_out22, Conv_valid_out23, Conv_valid_out24, Conv_valid_out25, Conv_valid_out26, Conv_valid_out27, 
            Conv_valid_out28, Conv_valid_out29, Conv_valid_out30, Conv_valid_out31, Conv_valid_out32, Conv_valid_out33, Conv_valid_out34, 
            Conv_valid_out35, Conv_valid_out36, Conv_valid_out37, Conv_valid_out38, Conv_valid_out39, Conv_valid_out40, Conv_valid_out41, 
            Conv_valid_out42, Conv_valid_out43, Conv_valid_out44, Conv_valid_out45, Conv_valid_out46, Conv_valid_out47, Conv_valid_out48, 
            Conv_valid_out49, Conv_valid_out50, Conv_valid_out51, Conv_valid_out52, Conv_valid_out53, Conv_valid_out54, Conv_valid_out55, 
            Conv_valid_out56, Conv_valid_out57, Conv_valid_out58, Conv_valid_out59, Conv_valid_out60, Conv_valid_out61, Conv_valid_out62, 
            Conv_valid_out63, Conv_valid_out64, Conv_valid_out65, Conv_valid_out66, Conv_valid_out67, Conv_valid_out68, Conv_valid_out69, 
            Conv_valid_out70, Conv_valid_out71, Conv_valid_out72, Conv_valid_out73, Conv_valid_out74, Conv_valid_out75, Conv_valid_out76, 
            Conv_valid_out77, Conv_valid_out78, Conv_valid_out79, Conv_valid_out80, Conv_valid_out81, Conv_valid_out82, Conv_valid_out83, 
            Conv_valid_out84, Conv_valid_out85, Conv_valid_out86, Conv_valid_out87, Conv_valid_out88, Conv_valid_out89, Conv_valid_out90, 
            Conv_valid_out91, Conv_valid_out92, Conv_valid_out93, Conv_valid_out94, Conv_valid_out95, Conv_valid_out96, Conv_valid_out97, 
            Conv_valid_out98, Conv_valid_out99, Conv_valid_out100, Conv_valid_out101, Conv_valid_out102, Conv_valid_out103, Conv_valid_out104, 
            Conv_valid_out105, Conv_valid_out106, Conv_valid_out107, Conv_valid_out108, Conv_valid_out109, Conv_valid_out110, Conv_valid_out111, 
            Conv_valid_out112, Conv_valid_out113, Conv_valid_out114, Conv_valid_out115, Conv_valid_out116, Conv_valid_out117, Conv_valid_out118, 
            Conv_valid_out119, Conv_valid_out120, Conv_valid_out121, Conv_valid_out122, Conv_valid_out123, Conv_valid_out124, Conv_valid_out125, 
            Conv_valid_out126, Conv_valid_out127, Conv_valid_out128, Conv_valid_out129, Conv_valid_out130, Conv_valid_out131, Conv_valid_out132, 
            Conv_valid_out133, Conv_valid_out134, Conv_valid_out135, Conv_valid_out136, Conv_valid_out137, Conv_valid_out138, Conv_valid_out139, 
            Conv_valid_out140, Conv_valid_out141, Conv_valid_out142, Conv_valid_out143, Conv_valid_out144, Conv_valid_out145, Conv_valid_out146, 
            Conv_valid_out147, Conv_valid_out148, Conv_valid_out149, Conv_valid_out150, Conv_valid_out151, Conv_valid_out152, Conv_valid_out153, 
            Conv_valid_out154, Conv_valid_out155, Conv_valid_out156, Conv_valid_out157, Conv_valid_out158, Conv_valid_out159, Conv_valid_out160, 
            Conv_valid_out161, Conv_valid_out162, Conv_valid_out163, Conv_valid_out164, Conv_valid_out165, Conv_valid_out166, Conv_valid_out167, 
            Conv_valid_out168, Conv_valid_out169, Conv_valid_out170, Conv_valid_out171, Conv_valid_out172, Conv_valid_out173, Conv_valid_out174, 
            Conv_valid_out175, Conv_valid_out176, Conv_valid_out177, Conv_valid_out178, Conv_valid_out179, Conv_valid_out180, Conv_valid_out181, 
            Conv_valid_out182, Conv_valid_out183, Conv_valid_out184, Conv_valid_out185, Conv_valid_out186, Conv_valid_out187, Conv_valid_out188, 
            Conv_valid_out189, Conv_valid_out190, Conv_valid_out191;

    wire [DATA_WIDTH - 1:0]
        ConvUnit_Out0, ConvUnit_Out1, ConvUnit_Out2, ConvUnit_Out3, ConvUnit_Out4, ConvUnit_Out5, ConvUnit_Out6, 
        ConvUnit_Out7, ConvUnit_Out8, ConvUnit_Out9, ConvUnit_Out10, ConvUnit_Out11, ConvUnit_Out12, ConvUnit_Out13, 
        ConvUnit_Out14, ConvUnit_Out15, ConvUnit_Out16, ConvUnit_Out17, ConvUnit_Out18, ConvUnit_Out19, ConvUnit_Out20, 
        ConvUnit_Out21, ConvUnit_Out22, ConvUnit_Out23, ConvUnit_Out24, ConvUnit_Out25, ConvUnit_Out26, ConvUnit_Out27, 
        ConvUnit_Out28, ConvUnit_Out29, ConvUnit_Out30, ConvUnit_Out31, ConvUnit_Out32, ConvUnit_Out33, ConvUnit_Out34, 
        ConvUnit_Out35, ConvUnit_Out36, ConvUnit_Out37, ConvUnit_Out38, ConvUnit_Out39, ConvUnit_Out40, ConvUnit_Out41, 
        ConvUnit_Out42, ConvUnit_Out43, ConvUnit_Out44, ConvUnit_Out45, ConvUnit_Out46, ConvUnit_Out47, ConvUnit_Out48, 
        ConvUnit_Out49, ConvUnit_Out50, ConvUnit_Out51, ConvUnit_Out52, ConvUnit_Out53, ConvUnit_Out54, ConvUnit_Out55, 
        ConvUnit_Out56, ConvUnit_Out57, ConvUnit_Out58, ConvUnit_Out59, ConvUnit_Out60, ConvUnit_Out61, ConvUnit_Out62, 
        ConvUnit_Out63, ConvUnit_Out64, ConvUnit_Out65, ConvUnit_Out66, ConvUnit_Out67, ConvUnit_Out68, ConvUnit_Out69, 
        ConvUnit_Out70, ConvUnit_Out71, ConvUnit_Out72, ConvUnit_Out73, ConvUnit_Out74, ConvUnit_Out75, ConvUnit_Out76, 
        ConvUnit_Out77, ConvUnit_Out78, ConvUnit_Out79, ConvUnit_Out80, ConvUnit_Out81, ConvUnit_Out82, ConvUnit_Out83, 
        ConvUnit_Out84, ConvUnit_Out85, ConvUnit_Out86, ConvUnit_Out87, ConvUnit_Out88, ConvUnit_Out89, ConvUnit_Out90, 
        ConvUnit_Out91, ConvUnit_Out92, ConvUnit_Out93, ConvUnit_Out94, ConvUnit_Out95, ConvUnit_Out96, ConvUnit_Out97, 
        ConvUnit_Out98, ConvUnit_Out99, ConvUnit_Out100, ConvUnit_Out101, ConvUnit_Out102, ConvUnit_Out103, ConvUnit_Out104, 
        ConvUnit_Out105, ConvUnit_Out106, ConvUnit_Out107, ConvUnit_Out108, ConvUnit_Out109, ConvUnit_Out110, ConvUnit_Out111, 
        ConvUnit_Out112, ConvUnit_Out113, ConvUnit_Out114, ConvUnit_Out115, ConvUnit_Out116, ConvUnit_Out117, ConvUnit_Out118, 
        ConvUnit_Out119, ConvUnit_Out120, ConvUnit_Out121, ConvUnit_Out122, ConvUnit_Out123, ConvUnit_Out124, ConvUnit_Out125, 
        ConvUnit_Out126, ConvUnit_Out127, ConvUnit_Out128, ConvUnit_Out129, ConvUnit_Out130, ConvUnit_Out131, ConvUnit_Out132, 
        ConvUnit_Out133, ConvUnit_Out134, ConvUnit_Out135, ConvUnit_Out136, ConvUnit_Out137, ConvUnit_Out138, ConvUnit_Out139, 
        ConvUnit_Out140, ConvUnit_Out141, ConvUnit_Out142, ConvUnit_Out143, ConvUnit_Out144, ConvUnit_Out145, ConvUnit_Out146, 
        ConvUnit_Out147, ConvUnit_Out148, ConvUnit_Out149, ConvUnit_Out150, ConvUnit_Out151, ConvUnit_Out152, ConvUnit_Out153, 
        ConvUnit_Out154, ConvUnit_Out155, ConvUnit_Out156, ConvUnit_Out157, ConvUnit_Out158, ConvUnit_Out159, ConvUnit_Out160, 
        ConvUnit_Out161, ConvUnit_Out162, ConvUnit_Out163, ConvUnit_Out164, ConvUnit_Out165, ConvUnit_Out166, ConvUnit_Out167, 
        ConvUnit_Out168, ConvUnit_Out169, ConvUnit_Out170, ConvUnit_Out171, ConvUnit_Out172, ConvUnit_Out173, ConvUnit_Out174, 
        ConvUnit_Out175, ConvUnit_Out176, ConvUnit_Out177, ConvUnit_Out178, ConvUnit_Out179, ConvUnit_Out180, ConvUnit_Out181, 
        ConvUnit_Out182, ConvUnit_Out183, ConvUnit_Out184, ConvUnit_Out185, ConvUnit_Out186, ConvUnit_Out187, ConvUnit_Out188, 
        ConvUnit_Out189, ConvUnit_Out190, ConvUnit_Out191;

    Maxpool Maxpool_Inst0(
        .data_in(Adder_Out),
        .data_out(),
        .Clk(Clk),
        .valid_in(),
        .valid_out(),
        .Rst(Rst)
    );

    ConvUnit Conv_Unit_Inst0 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out0), .data_out(ConvUnit_Out0)
    );
    ConvUnit Conv_Unit_Inst1 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out1), .data_out(ConvUnit_Out1)
    );
    ConvUnit Conv_Unit_Inst2 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out2), .data_out(ConvUnit_Out2)
    );
    ConvUnit Conv_Unit_Inst3 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out3), .data_out(ConvUnit_Out3)
    );
    ConvUnit Conv_Unit_Inst4 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out4), .data_out(ConvUnit_Out4)
    );
    ConvUnit Conv_Unit_Inst5 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out5), .data_out(ConvUnit_Out5)
    );
    ConvUnit Conv_Unit_Inst6 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out6), .data_out(ConvUnit_Out6)
    );
    ConvUnit Conv_Unit_Inst7 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out7), .data_out(ConvUnit_Out7)
    );
    ConvUnit Conv_Unit_Inst8 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out8), .data_out(ConvUnit_Out8)
    );
    ConvUnit Conv_Unit_Inst9 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out9), .data_out(ConvUnit_Out9)
    );
    ConvUnit Conv_Unit_Inst10 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out10), .data_out(ConvUnit_Out10)
    );
    ConvUnit Conv_Unit_Inst11 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out11), .data_out(ConvUnit_Out11)
    );
    ConvUnit Conv_Unit_Inst12 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out12), .data_out(ConvUnit_Out12)
    );
    ConvUnit Conv_Unit_Inst13 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out13), .data_out(ConvUnit_Out13)
    );
    ConvUnit Conv_Unit_Inst14 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out14), .data_out(ConvUnit_Out14)
    );
    ConvUnit Conv_Unit_Inst15 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out15), .data_out(ConvUnit_Out15)
    );
    ConvUnit Conv_Unit_Inst16 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out16), .data_out(ConvUnit_Out16)
    );
    ConvUnit Conv_Unit_Inst17 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out17), .data_out(ConvUnit_Out17)
    );
    ConvUnit Conv_Unit_Inst18 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out18), .data_out(ConvUnit_Out18)
    );
    ConvUnit Conv_Unit_Inst19 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out19), .data_out(ConvUnit_Out19)
    );
    ConvUnit Conv_Unit_Inst20 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out20), .data_out(ConvUnit_Out20)
    );
    ConvUnit Conv_Unit_Inst21 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out21), .data_out(ConvUnit_Out21)
    );
    ConvUnit Conv_Unit_Inst22 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out22), .data_out(ConvUnit_Out22)
    );
    ConvUnit Conv_Unit_Inst23 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out23), .data_out(ConvUnit_Out23)
    );
    ConvUnit Conv_Unit_Inst24 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out24), .data_out(ConvUnit_Out24)
    );
    ConvUnit Conv_Unit_Inst25 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out25), .data_out(ConvUnit_Out25)
    );
    ConvUnit Conv_Unit_Inst26 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out26), .data_out(ConvUnit_Out26)
    );
    ConvUnit Conv_Unit_Inst27 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out27), .data_out(ConvUnit_Out27)
    );
    ConvUnit Conv_Unit_Inst28 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out28), .data_out(ConvUnit_Out28)
    );
    ConvUnit Conv_Unit_Inst29 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out29), .data_out(ConvUnit_Out29)
    );
    ConvUnit Conv_Unit_Inst30 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out30), .data_out(ConvUnit_Out30)
    );
    ConvUnit Conv_Unit_Inst31 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out31), .data_out(ConvUnit_Out31)
    );
    ConvUnit Conv_Unit_Inst32 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out32), .data_out(ConvUnit_Out32)
    );
    ConvUnit Conv_Unit_Inst33 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out33), .data_out(ConvUnit_Out33)
    );
    ConvUnit Conv_Unit_Inst34 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out34), .data_out(ConvUnit_Out34)
    );
    ConvUnit Conv_Unit_Inst35 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out35), .data_out(ConvUnit_Out35)
    );
    ConvUnit Conv_Unit_Inst36 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out36), .data_out(ConvUnit_Out36)
    );
    ConvUnit Conv_Unit_Inst37 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out37), .data_out(ConvUnit_Out37)
    );
    ConvUnit Conv_Unit_Inst38 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out38), .data_out(ConvUnit_Out38)
    );
    ConvUnit Conv_Unit_Inst39 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out39), .data_out(ConvUnit_Out39)
    );
    ConvUnit Conv_Unit_Inst40 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out40), .data_out(ConvUnit_Out40)
    );
    ConvUnit Conv_Unit_Inst41 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out41), .data_out(ConvUnit_Out41)
    );
    ConvUnit Conv_Unit_Inst42 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out42), .data_out(ConvUnit_Out42)
    );
    ConvUnit Conv_Unit_Inst43 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out43), .data_out(ConvUnit_Out43)
    );
    ConvUnit Conv_Unit_Inst44 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out44), .data_out(ConvUnit_Out44)
    );
    ConvUnit Conv_Unit_Inst45 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out45), .data_out(ConvUnit_Out45)
    );
    ConvUnit Conv_Unit_Inst46 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out46), .data_out(ConvUnit_Out46)
    );
    ConvUnit Conv_Unit_Inst47 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out47), .data_out(ConvUnit_Out47)
    );
    ConvUnit Conv_Unit_Inst48 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out48), .data_out(ConvUnit_Out48)
    );
    ConvUnit Conv_Unit_Inst49 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out49), .data_out(ConvUnit_Out49)
    );
    ConvUnit Conv_Unit_Inst50 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out50), .data_out(ConvUnit_Out50)
    );
    ConvUnit Conv_Unit_Inst51 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out51), .data_out(ConvUnit_Out51)
    );
    ConvUnit Conv_Unit_Inst52 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out52), .data_out(ConvUnit_Out52)
    );
    ConvUnit Conv_Unit_Inst53 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out53), .data_out(ConvUnit_Out53)
    );
    ConvUnit Conv_Unit_Inst54 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out54), .data_out(ConvUnit_Out54)
    );
    ConvUnit Conv_Unit_Inst55 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out55), .data_out(ConvUnit_Out55)
    );
    ConvUnit Conv_Unit_Inst56 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out56), .data_out(ConvUnit_Out56)
    );
    ConvUnit Conv_Unit_Inst57 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out57), .data_out(ConvUnit_Out57)
    );
    ConvUnit Conv_Unit_Inst58 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out58), .data_out(ConvUnit_Out58)
    );
    ConvUnit Conv_Unit_Inst59 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out59), .data_out(ConvUnit_Out59)
    );
    ConvUnit Conv_Unit_Inst60 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out60), .data_out(ConvUnit_Out60)
    );
    ConvUnit Conv_Unit_Inst61 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out61), .data_out(ConvUnit_Out61)
    );
    ConvUnit Conv_Unit_Inst62 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out62), .data_out(ConvUnit_Out62)
    );
    ConvUnit Conv_Unit_Inst63 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out63), .data_out(ConvUnit_Out63)
    );
    ConvUnit Conv_Unit_Inst64 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out64), .data_out(ConvUnit_Out64)
    );
    ConvUnit Conv_Unit_Inst65 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out65), .data_out(ConvUnit_Out65)
    );
    ConvUnit Conv_Unit_Inst66 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out66), .data_out(ConvUnit_Out66)
    );
    ConvUnit Conv_Unit_Inst67 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out67), .data_out(ConvUnit_Out67)
    );
    ConvUnit Conv_Unit_Inst68 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out68), .data_out(ConvUnit_Out68)
    );
    ConvUnit Conv_Unit_Inst69 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out69), .data_out(ConvUnit_Out69)
    );
    ConvUnit Conv_Unit_Inst70 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out70), .data_out(ConvUnit_Out70)
    );
    ConvUnit Conv_Unit_Inst71 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out71), .data_out(ConvUnit_Out71)
    );
    ConvUnit Conv_Unit_Inst72 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out72), .data_out(ConvUnit_Out72)
    );
    ConvUnit Conv_Unit_Inst73 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out73), .data_out(ConvUnit_Out73)
    );
    ConvUnit Conv_Unit_Inst74 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out74), .data_out(ConvUnit_Out74)
    );
    ConvUnit Conv_Unit_Inst75 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out75), .data_out(ConvUnit_Out75)
    );
    ConvUnit Conv_Unit_Inst76 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out76), .data_out(ConvUnit_Out76)
    );
    ConvUnit Conv_Unit_Inst77 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out77), .data_out(ConvUnit_Out77)
    );
    ConvUnit Conv_Unit_Inst78 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out78), .data_out(ConvUnit_Out78)
    );
    ConvUnit Conv_Unit_Inst79 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out79), .data_out(ConvUnit_Out79)
    );
    ConvUnit Conv_Unit_Inst80 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out80), .data_out(ConvUnit_Out80)
    );
    ConvUnit Conv_Unit_Inst81 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out81), .data_out(ConvUnit_Out81)
    );
    ConvUnit Conv_Unit_Inst82 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out82), .data_out(ConvUnit_Out82)
    );
    ConvUnit Conv_Unit_Inst83 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out83), .data_out(ConvUnit_Out83)
    );
    ConvUnit Conv_Unit_Inst84 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out84), .data_out(ConvUnit_Out84)
    );
    ConvUnit Conv_Unit_Inst85 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out85), .data_out(ConvUnit_Out85)
    );
    ConvUnit Conv_Unit_Inst86 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out86), .data_out(ConvUnit_Out86)
    );
    ConvUnit Conv_Unit_Inst87 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out87), .data_out(ConvUnit_Out87)
    );
    ConvUnit Conv_Unit_Inst88 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out88), .data_out(ConvUnit_Out88)
    );
    ConvUnit Conv_Unit_Inst89 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out89), .data_out(ConvUnit_Out89)
    );
    ConvUnit Conv_Unit_Inst90 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out90), .data_out(ConvUnit_Out90)
    );
    ConvUnit Conv_Unit_Inst91 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out91), .data_out(ConvUnit_Out91)
    );
    ConvUnit Conv_Unit_Inst92 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out92), .data_out(ConvUnit_Out92)
    );
    ConvUnit Conv_Unit_Inst93 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out93), .data_out(ConvUnit_Out93)
    );
    ConvUnit Conv_Unit_Inst94 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out94), .data_out(ConvUnit_Out94)
    );
    ConvUnit Conv_Unit_Inst95 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out95), .data_out(ConvUnit_Out95)
    );
    ConvUnit Conv_Unit_Inst96 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out96), .data_out(ConvUnit_Out96)
    );
    ConvUnit Conv_Unit_Inst97 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out97), .data_out(ConvUnit_Out97)
    );
    ConvUnit Conv_Unit_Inst98 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out98), .data_out(ConvUnit_Out98)
    );
    ConvUnit Conv_Unit_Inst99 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out99), .data_out(ConvUnit_Out99)
    );
    ConvUnit Conv_Unit_Inst100 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out100), .data_out(ConvUnit_Out100)
    );
    ConvUnit Conv_Unit_Inst101 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out101), .data_out(ConvUnit_Out101)
    );
    ConvUnit Conv_Unit_Inst102 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out102), .data_out(ConvUnit_Out102)
    );
    ConvUnit Conv_Unit_Inst103 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out103), .data_out(ConvUnit_Out103)
    );
    ConvUnit Conv_Unit_Inst104 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out104), .data_out(ConvUnit_Out104)
    );
    ConvUnit Conv_Unit_Inst105 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out105), .data_out(ConvUnit_Out105)
    );
    ConvUnit Conv_Unit_Inst106 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out106), .data_out(ConvUnit_Out106)
    );
    ConvUnit Conv_Unit_Inst107 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out107), .data_out(ConvUnit_Out107)
    );
    ConvUnit Conv_Unit_Inst108 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out108), .data_out(ConvUnit_Out108)
    );
    ConvUnit Conv_Unit_Inst109 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out109), .data_out(ConvUnit_Out109)
    );
    ConvUnit Conv_Unit_Inst110 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out110), .data_out(ConvUnit_Out110)
    );
    ConvUnit Conv_Unit_Inst111 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out111), .data_out(ConvUnit_Out111)
    );
    ConvUnit Conv_Unit_Inst112 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out112), .data_out(ConvUnit_Out112)
    );
    ConvUnit Conv_Unit_Inst113 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out113), .data_out(ConvUnit_Out113)
    );
    ConvUnit Conv_Unit_Inst114 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out114), .data_out(ConvUnit_Out114)
    );
    ConvUnit Conv_Unit_Inst115 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out115), .data_out(ConvUnit_Out115)
    );
    ConvUnit Conv_Unit_Inst116 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out116), .data_out(ConvUnit_Out116)
    );
    ConvUnit Conv_Unit_Inst117 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out117), .data_out(ConvUnit_Out117)
    );
    ConvUnit Conv_Unit_Inst118 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out118), .data_out(ConvUnit_Out118)
    );
    ConvUnit Conv_Unit_Inst119 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out119), .data_out(ConvUnit_Out119)
    );
    ConvUnit Conv_Unit_Inst120 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out120), .data_out(ConvUnit_Out120)
    );
    ConvUnit Conv_Unit_Inst121 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out121), .data_out(ConvUnit_Out121)
    );
    ConvUnit Conv_Unit_Inst122 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out122), .data_out(ConvUnit_Out122)
    );
    ConvUnit Conv_Unit_Inst123 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out123), .data_out(ConvUnit_Out123)
    );
    ConvUnit Conv_Unit_Inst124 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out124), .data_out(ConvUnit_Out124)
    );
    ConvUnit Conv_Unit_Inst125 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out125), .data_out(ConvUnit_Out125)
    );
    ConvUnit Conv_Unit_Inst126 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out126), .data_out(ConvUnit_Out126)
    );
    ConvUnit Conv_Unit_Inst127 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out127), .data_out(ConvUnit_Out127)
    );
    ConvUnit Conv_Unit_Inst128 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out128), .data_out(ConvUnit_Out128)
    );
    ConvUnit Conv_Unit_Inst129 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out129), .data_out(ConvUnit_Out129)
    );
    ConvUnit Conv_Unit_Inst130 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out130), .data_out(ConvUnit_Out130)
    );
    ConvUnit Conv_Unit_Inst131 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out131), .data_out(ConvUnit_Out131)
    );
    ConvUnit Conv_Unit_Inst132 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out132), .data_out(ConvUnit_Out132)
    );
    ConvUnit Conv_Unit_Inst133 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out133), .data_out(ConvUnit_Out133)
    );
    ConvUnit Conv_Unit_Inst134 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out134), .data_out(ConvUnit_Out134)
    );
    ConvUnit Conv_Unit_Inst135 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out135), .data_out(ConvUnit_Out135)
    );
    ConvUnit Conv_Unit_Inst136 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out136), .data_out(ConvUnit_Out136)
    );
    ConvUnit Conv_Unit_Inst137 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out137), .data_out(ConvUnit_Out137)
    );
    ConvUnit Conv_Unit_Inst138 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out138), .data_out(ConvUnit_Out138)
    );
    ConvUnit Conv_Unit_Inst139 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out139), .data_out(ConvUnit_Out139)
    );
    ConvUnit Conv_Unit_Inst140 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out140), .data_out(ConvUnit_Out140)
    );
    ConvUnit Conv_Unit_Inst141 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out141), .data_out(ConvUnit_Out141)
    );
    ConvUnit Conv_Unit_Inst142 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out142), .data_out(ConvUnit_Out142)
    );
    ConvUnit Conv_Unit_Inst143 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out143), .data_out(ConvUnit_Out143)
    );
    ConvUnit Conv_Unit_Inst144 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out144), .data_out(ConvUnit_Out144)
    );
    ConvUnit Conv_Unit_Inst145 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out145), .data_out(ConvUnit_Out145)
    );
    ConvUnit Conv_Unit_Inst146 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out146), .data_out(ConvUnit_Out146)
    );
    ConvUnit Conv_Unit_Inst147 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out147), .data_out(ConvUnit_Out147)
    );
    ConvUnit Conv_Unit_Inst148 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out148), .data_out(ConvUnit_Out148)
    );
    ConvUnit Conv_Unit_Inst149 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out149), .data_out(ConvUnit_Out149)
    );
    ConvUnit Conv_Unit_Inst150 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out150), .data_out(ConvUnit_Out150)
    );
    ConvUnit Conv_Unit_Inst151 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out151), .data_out(ConvUnit_Out151)
    );
    ConvUnit Conv_Unit_Inst152 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out152), .data_out(ConvUnit_Out152)
    );
    ConvUnit Conv_Unit_Inst153 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out153), .data_out(ConvUnit_Out153)
    );
    ConvUnit Conv_Unit_Inst154 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out154), .data_out(ConvUnit_Out154)
    );
    ConvUnit Conv_Unit_Inst155 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out155), .data_out(ConvUnit_Out155)
    );
    ConvUnit Conv_Unit_Inst156 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out156), .data_out(ConvUnit_Out156)
    );
    ConvUnit Conv_Unit_Inst157 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out157), .data_out(ConvUnit_Out157)
    );
    ConvUnit Conv_Unit_Inst158 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out158), .data_out(ConvUnit_Out158)
    );
    ConvUnit Conv_Unit_Inst159 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out159), .data_out(ConvUnit_Out159)
    );
    ConvUnit Conv_Unit_Inst160 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out160), .data_out(ConvUnit_Out160)
    );
    ConvUnit Conv_Unit_Inst161 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out161), .data_out(ConvUnit_Out161)
    );
    ConvUnit Conv_Unit_Inst162 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out162), .data_out(ConvUnit_Out162)
    );
    ConvUnit Conv_Unit_Inst163 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out163), .data_out(ConvUnit_Out163)
    );
    ConvUnit Conv_Unit_Inst164 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out164), .data_out(ConvUnit_Out164)
    );
    ConvUnit Conv_Unit_Inst165 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out165), .data_out(ConvUnit_Out165)
    );
    ConvUnit Conv_Unit_Inst166 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out166), .data_out(ConvUnit_Out166)
    );
    ConvUnit Conv_Unit_Inst167 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out167), .data_out(ConvUnit_Out167)
    );
    ConvUnit Conv_Unit_Inst168 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out168), .data_out(ConvUnit_Out168)
    );
    ConvUnit Conv_Unit_Inst169 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out169), .data_out(ConvUnit_Out169)
    );
    ConvUnit Conv_Unit_Inst170 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out170), .data_out(ConvUnit_Out170)
    );
    ConvUnit Conv_Unit_Inst171 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out171), .data_out(ConvUnit_Out171)
    );
    ConvUnit Conv_Unit_Inst172 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out172), .data_out(ConvUnit_Out172)
    );
    ConvUnit Conv_Unit_Inst173 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out173), .data_out(ConvUnit_Out173)
    );
    ConvUnit Conv_Unit_Inst174 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out174), .data_out(ConvUnit_Out174)
    );
    ConvUnit Conv_Unit_Inst175 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out175), .data_out(ConvUnit_Out175)
    );
    ConvUnit Conv_Unit_Inst176 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out176), .data_out(ConvUnit_Out176)
    );
    ConvUnit Conv_Unit_Inst177 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out177), .data_out(ConvUnit_Out177)
    );
    ConvUnit Conv_Unit_Inst178 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out178), .data_out(ConvUnit_Out178)
    );
    ConvUnit Conv_Unit_Inst179 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out179), .data_out(ConvUnit_Out179)
    );
    ConvUnit Conv_Unit_Inst180 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out180), .data_out(ConvUnit_Out180)
    );
    ConvUnit Conv_Unit_Inst181 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out181), .data_out(ConvUnit_Out181)
    );
    ConvUnit Conv_Unit_Inst182 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out182), .data_out(ConvUnit_Out182)
    );
    ConvUnit Conv_Unit_Inst183 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out183), .data_out(ConvUnit_Out183)
    );
    ConvUnit Conv_Unit_Inst184 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out184), .data_out(ConvUnit_Out184)
    );
    ConvUnit Conv_Unit_Inst185 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out185), .data_out(ConvUnit_Out185)
    );
    ConvUnit Conv_Unit_Inst186 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out186), .data_out(ConvUnit_Out186)
    );
    ConvUnit Conv_Unit_Inst187 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out187), .data_out(ConvUnit_Out187)
    );
    ConvUnit Conv_Unit_Inst188 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out188), .data_out(ConvUnit_Out188)
    );
    ConvUnit Conv_Unit_Inst189 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out189), .data_out(ConvUnit_Out189)
    );
    ConvUnit Conv_Unit_Inst190 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out190), .data_out(ConvUnit_Out190)
    );
    ConvUnit Conv_Unit_Inst191 (
        .data_in(fifo_in_out), .Clk(Clk), .Rst(Rst), .valid_in(valid_in_signal), .valid_out(Conv_valid_out191), .data_out(ConvUnit_Out191)
    );
endmodule