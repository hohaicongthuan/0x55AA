module layer_10_featuremap_418(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4943b6),
	.w1(32'hbb840ef9),
	.w2(32'hbae2ce6d),
	.w3(32'hbbac0d13),
	.w4(32'hbb8fb7ea),
	.w5(32'h3ad4503e),
	.w6(32'hbb2799b7),
	.w7(32'hbab74e06),
	.w8(32'h3a280807),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c414e),
	.w1(32'hbc2d151c),
	.w2(32'h3b38563a),
	.w3(32'hbc00af60),
	.w4(32'h3c6e6f69),
	.w5(32'h3cba63ac),
	.w6(32'hbc13c8db),
	.w7(32'h3c28010a),
	.w8(32'h3c943d18),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6006b9),
	.w1(32'hbc07dd26),
	.w2(32'h3a9bf74d),
	.w3(32'hbb44aa1a),
	.w4(32'hbbcd4477),
	.w5(32'h3b3f52a8),
	.w6(32'hbc238d81),
	.w7(32'hbaa47c0c),
	.w8(32'h3bee2224),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc61b9b),
	.w1(32'hbad6dc42),
	.w2(32'hba2ac985),
	.w3(32'h3c0d44e0),
	.w4(32'h39842493),
	.w5(32'h3bd19482),
	.w6(32'h3bd74db3),
	.w7(32'hbb036513),
	.w8(32'h3b8b13ec),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870e5f),
	.w1(32'hbb17491a),
	.w2(32'h3afe096d),
	.w3(32'hba006dcb),
	.w4(32'h3b318cee),
	.w5(32'h3c1669f0),
	.w6(32'hbb1a4842),
	.w7(32'h3b57d8f0),
	.w8(32'h3ba48c15),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83e46e),
	.w1(32'hbaebc7a2),
	.w2(32'h3b6ef258),
	.w3(32'h3c3d42cb),
	.w4(32'hba8e2fca),
	.w5(32'hbb38dcd4),
	.w6(32'h3b0a9cee),
	.w7(32'hbb23bd63),
	.w8(32'h3b13e511),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899bdde),
	.w1(32'hbb0e4097),
	.w2(32'hbc396f2d),
	.w3(32'h3b4fc99d),
	.w4(32'hbb939c82),
	.w5(32'hbc862271),
	.w6(32'h3c24e661),
	.w7(32'hbb10bc1f),
	.w8(32'hbb5d9906),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc793eb1),
	.w1(32'hbc123302),
	.w2(32'hbc397ee5),
	.w3(32'hbc768cfb),
	.w4(32'hbc1e3586),
	.w5(32'hbc42fb2c),
	.w6(32'hbafd99f0),
	.w7(32'hbbeab30d),
	.w8(32'h3bb58a5e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bddc4),
	.w1(32'h3aac3c79),
	.w2(32'hbb62c4e0),
	.w3(32'hbb14acf1),
	.w4(32'hbb55b6e2),
	.w5(32'hbc1f98eb),
	.w6(32'h3b11ff6e),
	.w7(32'hbad97357),
	.w8(32'hbc0c9b3c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3552b0),
	.w1(32'h3b680316),
	.w2(32'hbc548d2c),
	.w3(32'hbc07d6dc),
	.w4(32'h3c16a214),
	.w5(32'hbc00c246),
	.w6(32'hbc008cc7),
	.w7(32'h3c686a02),
	.w8(32'hbb5f6f6d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1825fd),
	.w1(32'h3b1ca4ed),
	.w2(32'h3c3dfe71),
	.w3(32'hbc15cd9a),
	.w4(32'hbb8a850d),
	.w5(32'h3a89c132),
	.w6(32'hbbb71a01),
	.w7(32'hbbf3e982),
	.w8(32'hbbaf88d3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4bd057),
	.w1(32'h3ba6b2a9),
	.w2(32'h3bd34b42),
	.w3(32'hbc293d4e),
	.w4(32'h3a7eb30b),
	.w5(32'h3bbfd40f),
	.w6(32'hbac4eec4),
	.w7(32'h3bce2ad8),
	.w8(32'h3a3ec04a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4271e4),
	.w1(32'h3bac1033),
	.w2(32'hbc83866f),
	.w3(32'h3bdf1606),
	.w4(32'h3c8c2d28),
	.w5(32'h3c129edc),
	.w6(32'h3b99b73f),
	.w7(32'h3c766f32),
	.w8(32'h3a137cdc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1715a6),
	.w1(32'hba1a5e49),
	.w2(32'hbb8acf8c),
	.w3(32'hb97da14a),
	.w4(32'hbb9fc8f1),
	.w5(32'hbc0189ac),
	.w6(32'hbb7524b2),
	.w7(32'hba749346),
	.w8(32'hbbc16e26),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99901),
	.w1(32'hbc0dcedf),
	.w2(32'hbbb3bc35),
	.w3(32'hba85b478),
	.w4(32'hb81ecfe6),
	.w5(32'hbb24e657),
	.w6(32'hbc47805e),
	.w7(32'hbb5095a7),
	.w8(32'hbb973e6d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c1d51),
	.w1(32'hbbc2c972),
	.w2(32'hbc77bb96),
	.w3(32'hbbb821a9),
	.w4(32'hba17b2c2),
	.w5(32'hbc55d587),
	.w6(32'hbc726787),
	.w7(32'hbb900162),
	.w8(32'hbc2e3df5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af38743),
	.w1(32'hbafc7fa7),
	.w2(32'h3a50c91e),
	.w3(32'hbbb02682),
	.w4(32'hbbb599ad),
	.w5(32'hba511cd6),
	.w6(32'hbb920ff0),
	.w7(32'hbb282527),
	.w8(32'hbad17319),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1d319),
	.w1(32'hbb8452c3),
	.w2(32'hbce42ddc),
	.w3(32'hbbae5cce),
	.w4(32'h3acd998d),
	.w5(32'hbc95040b),
	.w6(32'hbaf64ac7),
	.w7(32'h39e08369),
	.w8(32'hbc8ce32a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6cc14),
	.w1(32'h3b89a261),
	.w2(32'hbc628d1b),
	.w3(32'hbb2d05bb),
	.w4(32'h3b5ccc1f),
	.w5(32'hbbb84193),
	.w6(32'h3a4d5bd1),
	.w7(32'h3bd022ee),
	.w8(32'hbbdcc006),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb138aba),
	.w1(32'hbaa153c6),
	.w2(32'h3ba2ae7f),
	.w3(32'h3b847703),
	.w4(32'hba38b58c),
	.w5(32'h3c332322),
	.w6(32'h3a08d163),
	.w7(32'h3b3157d2),
	.w8(32'h3bd69215),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff607),
	.w1(32'h3ab632e6),
	.w2(32'h3b1e0d73),
	.w3(32'hb93bccba),
	.w4(32'hb9b28fb0),
	.w5(32'hba8b9d30),
	.w6(32'hbb07c38f),
	.w7(32'h37d19dfc),
	.w8(32'hbb4cac63),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04f495),
	.w1(32'h39c80371),
	.w2(32'h3a584df1),
	.w3(32'hbba112cd),
	.w4(32'h3b16cfd4),
	.w5(32'h3ba00fc3),
	.w6(32'hbc313c0e),
	.w7(32'h3b04daa3),
	.w8(32'h3b634175),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1173e1),
	.w1(32'hbc7d5da9),
	.w2(32'hbc737d57),
	.w3(32'hbcca8afb),
	.w4(32'hbb17a442),
	.w5(32'hba7ce7f2),
	.w6(32'hbcae7d81),
	.w7(32'hbb4bcb58),
	.w8(32'hbc1574c6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e81a7),
	.w1(32'hbbec066d),
	.w2(32'hbbb4b52b),
	.w3(32'hbb53f23b),
	.w4(32'h3c7d37aa),
	.w5(32'h3c66c45c),
	.w6(32'hbc39005d),
	.w7(32'h3c0b8ad5),
	.w8(32'h3c385db4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd094bae),
	.w1(32'hbc0ee5be),
	.w2(32'hbae0ef11),
	.w3(32'hbc20ee8b),
	.w4(32'h3ba42753),
	.w5(32'h3c01f708),
	.w6(32'hbcbd6fe2),
	.w7(32'h3bcff045),
	.w8(32'h3c261a2e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ba528),
	.w1(32'h3b03ae98),
	.w2(32'h3b3ae0c9),
	.w3(32'hbba18170),
	.w4(32'h3b97962e),
	.w5(32'h3bc17ecd),
	.w6(32'hbb418f04),
	.w7(32'h3b2f4558),
	.w8(32'h3b3153b7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70f115),
	.w1(32'h3bf665df),
	.w2(32'h3bf880aa),
	.w3(32'h3b832ed2),
	.w4(32'h3b61f672),
	.w5(32'hbb11a096),
	.w6(32'h3b56fc37),
	.w7(32'h3b8a45fc),
	.w8(32'hba35b8bc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0547c0),
	.w1(32'hbc0bb98e),
	.w2(32'hbc25c6b9),
	.w3(32'hb93b3dca),
	.w4(32'hba791731),
	.w5(32'hbb3da677),
	.w6(32'hbbe6ad60),
	.w7(32'hbc1ed0b4),
	.w8(32'hbb9ab091),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b2b2),
	.w1(32'h3b751ffb),
	.w2(32'h3bef4252),
	.w3(32'hbc20241d),
	.w4(32'h3afe9b0d),
	.w5(32'h3ba65190),
	.w6(32'hbc365b78),
	.w7(32'hba37a2c1),
	.w8(32'h3aebf90b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b575f30),
	.w1(32'hbb603147),
	.w2(32'hb9517e4c),
	.w3(32'h3b70f4b7),
	.w4(32'h3b747d17),
	.w5(32'h3b8b75b3),
	.w6(32'h3b2ebad7),
	.w7(32'h3b11a5a3),
	.w8(32'h3b1677a7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e1df7),
	.w1(32'hb9643fce),
	.w2(32'hbaed76d3),
	.w3(32'hb921e294),
	.w4(32'hbba14852),
	.w5(32'hbb3fbaef),
	.w6(32'h39e86d04),
	.w7(32'hba174d91),
	.w8(32'h3afc5e01),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeee8fa),
	.w1(32'h3a28bc85),
	.w2(32'h3a2e5bad),
	.w3(32'hbb27d0f2),
	.w4(32'h3bd1ae01),
	.w5(32'hbaeaed54),
	.w6(32'hb9954ede),
	.w7(32'h3bde2389),
	.w8(32'h3a13b82e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c080a),
	.w1(32'hbb7a8140),
	.w2(32'hbbcea30a),
	.w3(32'hbb77b6ab),
	.w4(32'hb938aee4),
	.w5(32'hbb190a5c),
	.w6(32'hbabdd639),
	.w7(32'h3c0929fb),
	.w8(32'h3c291fdc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c65f9),
	.w1(32'hbbded568),
	.w2(32'hba083ea6),
	.w3(32'hbc29dec6),
	.w4(32'hbb71b9e2),
	.w5(32'h3a96bd22),
	.w6(32'hbbb5fa35),
	.w7(32'hbbe3b0a2),
	.w8(32'hbb94280a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac101de),
	.w1(32'h3af902cb),
	.w2(32'h3bd0362f),
	.w3(32'h3a90db87),
	.w4(32'hbab86735),
	.w5(32'hb9dd34ed),
	.w6(32'hbb8e179f),
	.w7(32'hba9c8664),
	.w8(32'hbb5840d7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e50a9),
	.w1(32'h3a50c8f9),
	.w2(32'h3b1edf92),
	.w3(32'hb950d402),
	.w4(32'hbba734bc),
	.w5(32'hbb6959b4),
	.w6(32'hbb33e273),
	.w7(32'hbbd3c470),
	.w8(32'hbc0e57a8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b55db),
	.w1(32'h3c145f41),
	.w2(32'h3c0ba19b),
	.w3(32'hbd120bb7),
	.w4(32'h3be0bbed),
	.w5(32'h3c30c1a5),
	.w6(32'hbca4c43e),
	.w7(32'h3a9326c9),
	.w8(32'h3b395718),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd23055c),
	.w1(32'hbc57bfec),
	.w2(32'h3ca9958f),
	.w3(32'hbca2efd6),
	.w4(32'h3c4105c9),
	.w5(32'h3d0bb11a),
	.w6(32'hbce66c90),
	.w7(32'h3c5d3609),
	.w8(32'h3cf3c204),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd004122),
	.w1(32'hbc9ae6cc),
	.w2(32'h3bc1b6ac),
	.w3(32'hbcbe70c1),
	.w4(32'hbbf8ba52),
	.w5(32'h3c06c043),
	.w6(32'hbd252f6e),
	.w7(32'hbc909aa5),
	.w8(32'hbc110098),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fe656),
	.w1(32'hb9bd24ee),
	.w2(32'h3bf0408c),
	.w3(32'hbb309a17),
	.w4(32'h3af343b1),
	.w5(32'h3c5c4394),
	.w6(32'hbc580e4d),
	.w7(32'h3aefda49),
	.w8(32'h3c3548c5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c39079),
	.w1(32'hbc18d224),
	.w2(32'h3af4b87b),
	.w3(32'hbadbcb42),
	.w4(32'h3c278e58),
	.w5(32'h3cab4375),
	.w6(32'h3a3dd572),
	.w7(32'hbb0b21e2),
	.w8(32'h3c423d94),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932a2c),
	.w1(32'hbbaa1206),
	.w2(32'hbaf0e9fb),
	.w3(32'h3c587f38),
	.w4(32'h39d2c332),
	.w5(32'hbbb2eecc),
	.w6(32'h3bb8ab87),
	.w7(32'hbb668891),
	.w8(32'hbb5297c2),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e45b),
	.w1(32'hbb72ce15),
	.w2(32'h3b0a2c92),
	.w3(32'hbc168e8a),
	.w4(32'hba8200f0),
	.w5(32'h3c9c571b),
	.w6(32'hbc32c46f),
	.w7(32'hbb8f0aa5),
	.w8(32'h3c5b80b2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5ebc),
	.w1(32'h38801eda),
	.w2(32'hbcc0d567),
	.w3(32'h3b991c3a),
	.w4(32'h3b3e12a8),
	.w5(32'hbc9453ee),
	.w6(32'hbba96d17),
	.w7(32'h3aa26d63),
	.w8(32'hbc5f1b66),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ce9b5),
	.w1(32'hbb4b6e8a),
	.w2(32'hbba8031a),
	.w3(32'hbc20a0d0),
	.w4(32'h3bf7733d),
	.w5(32'h3c3d8b7c),
	.w6(32'hbc3ace70),
	.w7(32'h3c3c4926),
	.w8(32'h3c82877f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8110dc),
	.w1(32'hbc205c09),
	.w2(32'hbc9b3650),
	.w3(32'h3b4f5a3d),
	.w4(32'h3b6ac649),
	.w5(32'hbc038307),
	.w6(32'h3af819e5),
	.w7(32'h3bfca58e),
	.w8(32'h3b230152),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca86196),
	.w1(32'hbb9dacf9),
	.w2(32'hb8ab2e9a),
	.w3(32'hbc938a1d),
	.w4(32'h3b95f234),
	.w5(32'h3b68d3e6),
	.w6(32'hbc9957bc),
	.w7(32'hbbde5134),
	.w8(32'hbb62d26a),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc068f8),
	.w1(32'h3b889392),
	.w2(32'hbc98207d),
	.w3(32'hbbf2e892),
	.w4(32'hbb83bf04),
	.w5(32'hbc9145f7),
	.w6(32'hbae1bf43),
	.w7(32'h3bf6e1f4),
	.w8(32'hbc29dfbd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2986d2),
	.w1(32'h39b67778),
	.w2(32'h39b3f338),
	.w3(32'hbbc3eace),
	.w4(32'hbb831ed8),
	.w5(32'hbb1eac19),
	.w6(32'hbb133fa1),
	.w7(32'hb9b390e0),
	.w8(32'hbb034564),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb674262),
	.w1(32'hbbd6e709),
	.w2(32'h3b8c4676),
	.w3(32'hbb800989),
	.w4(32'hbb99ee4d),
	.w5(32'hbb66d10a),
	.w6(32'hbc2de1f7),
	.w7(32'hbb76b17b),
	.w8(32'hbb6808a4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b371ccb),
	.w1(32'h3b03d79c),
	.w2(32'h3b3e0a9a),
	.w3(32'hba844cc4),
	.w4(32'hbafe09c2),
	.w5(32'hbb3b976a),
	.w6(32'hbbe86cc2),
	.w7(32'hbaa684ec),
	.w8(32'hbb54c8f0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1453aa),
	.w1(32'hbb844bbc),
	.w2(32'hbc58c4f4),
	.w3(32'h3b329a37),
	.w4(32'hb9c91cf9),
	.w5(32'hbc256c21),
	.w6(32'hbb8db5d0),
	.w7(32'h3ac6ec19),
	.w8(32'hbb1ba6b4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaaba2),
	.w1(32'h3aadc28d),
	.w2(32'h3a7fdf1d),
	.w3(32'hbb9ace72),
	.w4(32'hbb88faec),
	.w5(32'hbb2c27fb),
	.w6(32'hb90499c8),
	.w7(32'hbb1c6fc4),
	.w8(32'h3a9ca0d6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d15c1),
	.w1(32'hbaf5e7ab),
	.w2(32'hbcb420ec),
	.w3(32'hbc2cbb3e),
	.w4(32'hbbc1e19d),
	.w5(32'hbc86f5eb),
	.w6(32'hba51cfc0),
	.w7(32'h3a13162c),
	.w8(32'hbc88a50b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ba477),
	.w1(32'hbb621c77),
	.w2(32'hbc0fee92),
	.w3(32'hbbc7dff9),
	.w4(32'h3a2c7b13),
	.w5(32'h39ca4ca0),
	.w6(32'hbc45b842),
	.w7(32'h3bda1252),
	.w8(32'h3b0b37b1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b386d),
	.w1(32'hbc13913d),
	.w2(32'hbbafa002),
	.w3(32'hbb1fe3aa),
	.w4(32'hbb95271f),
	.w5(32'h3c01795e),
	.w6(32'hb9f470e2),
	.w7(32'h3b25d3ab),
	.w8(32'h3c094be4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1abcc),
	.w1(32'h379a4954),
	.w2(32'h3add69b9),
	.w3(32'h38cdc4e0),
	.w4(32'hba366b52),
	.w5(32'hba04ceba),
	.w6(32'hbb908661),
	.w7(32'hbb230594),
	.w8(32'hbb567f58),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388fb4f6),
	.w1(32'hbb79e8fe),
	.w2(32'hbb186494),
	.w3(32'h3b4cabc5),
	.w4(32'h393f9ae2),
	.w5(32'hbabba710),
	.w6(32'hbadd4e53),
	.w7(32'hbbc9cdfa),
	.w8(32'h3b6560e2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4af92),
	.w1(32'hbbebfedf),
	.w2(32'hbbb9735e),
	.w3(32'hbba7d31f),
	.w4(32'h3baf43d6),
	.w5(32'h3c6348cf),
	.w6(32'hbbc0f69b),
	.w7(32'hbb27c0b6),
	.w8(32'h3b375954),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc691fd1),
	.w1(32'h3b4c2a04),
	.w2(32'hbb7f64d6),
	.w3(32'hba167f29),
	.w4(32'h3bb40e83),
	.w5(32'h3b9ac68e),
	.w6(32'hbb744bbd),
	.w7(32'hbbbfeec8),
	.w8(32'hbb4dafff),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f4f3a),
	.w1(32'h3a0435ab),
	.w2(32'hbb92de90),
	.w3(32'hbc1ebe60),
	.w4(32'h3b3b591b),
	.w5(32'h3aab9838),
	.w6(32'hbb407480),
	.w7(32'h3ade7cf2),
	.w8(32'hbb2110c9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d8e5),
	.w1(32'hbc0774fd),
	.w2(32'hbc488450),
	.w3(32'hbbda4139),
	.w4(32'hbba07b6e),
	.w5(32'hbbab4b8e),
	.w6(32'hbc21fe89),
	.w7(32'hbbceea30),
	.w8(32'hbbaba041),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb449650),
	.w1(32'hbbb365d5),
	.w2(32'hba0c650f),
	.w3(32'h3c03c538),
	.w4(32'h3b49eb5e),
	.w5(32'h3c75490d),
	.w6(32'h396ad225),
	.w7(32'hbbae7924),
	.w8(32'h3b7ca58f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14eee5),
	.w1(32'hbae3cc9c),
	.w2(32'h3a5dfb1a),
	.w3(32'h3c169acf),
	.w4(32'hbb6b57c7),
	.w5(32'h3b4e975d),
	.w6(32'h3b5ae475),
	.w7(32'hbae1057a),
	.w8(32'h3b5c411b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e6989),
	.w1(32'h3c124ff1),
	.w2(32'h3c13fe94),
	.w3(32'h3c229978),
	.w4(32'h3b778054),
	.w5(32'hbab20017),
	.w6(32'h3bd32bfe),
	.w7(32'h3b62039b),
	.w8(32'hbb2d8164),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1717bb),
	.w1(32'hbbb605f8),
	.w2(32'hbb151457),
	.w3(32'hbc2668a7),
	.w4(32'hba96d753),
	.w5(32'h3a752d11),
	.w6(32'hbc1bb2f4),
	.w7(32'hbb987c2d),
	.w8(32'h3b104899),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3c72c),
	.w1(32'hbba6fbbb),
	.w2(32'hbcb7848f),
	.w3(32'h3abbd325),
	.w4(32'hbbf7c136),
	.w5(32'hbca74c4e),
	.w6(32'hbc0dc281),
	.w7(32'hbc91a6d3),
	.w8(32'hbc75b25d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce40df5),
	.w1(32'hbc570834),
	.w2(32'hbc91ab05),
	.w3(32'hbc1ab0b8),
	.w4(32'hb9ee828d),
	.w5(32'hbab1d4c6),
	.w6(32'hbc5e3297),
	.w7(32'h3b3a6a44),
	.w8(32'h3bf6f06f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0d43b),
	.w1(32'hbba59954),
	.w2(32'hbc91f44b),
	.w3(32'hbbfe827c),
	.w4(32'h3bf20020),
	.w5(32'hbbdb5e4f),
	.w6(32'hbc6d74bc),
	.w7(32'hba0aeed5),
	.w8(32'hbad78b51),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcb138),
	.w1(32'hbb6d2b43),
	.w2(32'h3bd06a10),
	.w3(32'hbc2878be),
	.w4(32'h3c803ed6),
	.w5(32'h3cd705e3),
	.w6(32'hbca58f72),
	.w7(32'h3c9877b5),
	.w8(32'h3cd09f5b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b880f3),
	.w1(32'h38527662),
	.w2(32'h3882414a),
	.w3(32'h39b94b21),
	.w4(32'h3737b8e0),
	.w5(32'h373caa03),
	.w6(32'h39c969f3),
	.w7(32'h37dc8bee),
	.w8(32'h382edf47),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cd965),
	.w1(32'h38aa0be1),
	.w2(32'h391266de),
	.w3(32'h3a041f3e),
	.w4(32'hb7ca0af2),
	.w5(32'h37f43ec5),
	.w6(32'h39fafcfb),
	.w7(32'h3820f19c),
	.w8(32'h38fe5931),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e49c1),
	.w1(32'h37644833),
	.w2(32'h3807c0a8),
	.w3(32'h3a1d42e8),
	.w4(32'hb8767579),
	.w5(32'hb8e25630),
	.w6(32'h39f8b24a),
	.w7(32'hb847e052),
	.w8(32'hb896cb5a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d63ab),
	.w1(32'h3a45e348),
	.w2(32'hbb5d3e2f),
	.w3(32'hba88a4e0),
	.w4(32'h3a684d46),
	.w5(32'hbb1ff9f8),
	.w6(32'h39cbad17),
	.w7(32'h3ae304ac),
	.w8(32'hbaead2e6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3512f),
	.w1(32'h3883789c),
	.w2(32'hb7886ceb),
	.w3(32'h39ae9eda),
	.w4(32'hb79c3c92),
	.w5(32'hb8230ea6),
	.w6(32'h39bf4523),
	.w7(32'h388cbcec),
	.w8(32'h3854cfdb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ab77),
	.w1(32'h3aca6e7e),
	.w2(32'hbb8db7bf),
	.w3(32'hbadbcc4f),
	.w4(32'h391f9fa2),
	.w5(32'hbaa879fa),
	.w6(32'h3c01f3df),
	.w7(32'h3b92a410),
	.w8(32'h3b3f505c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dae7b),
	.w1(32'hbae29368),
	.w2(32'hbba16ba9),
	.w3(32'hbbf8bd46),
	.w4(32'hba92eb56),
	.w5(32'h3b4be045),
	.w6(32'h3aae6e7a),
	.w7(32'h3b02c656),
	.w8(32'h3ba907af),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41ffc7),
	.w1(32'hbbd4a6fb),
	.w2(32'hbbeba2e9),
	.w3(32'hbba33704),
	.w4(32'h3b988004),
	.w5(32'h3b3a7195),
	.w6(32'hbbdf2123),
	.w7(32'h3bc7c433),
	.w8(32'h3c0ae344),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbaef2),
	.w1(32'hb902b4be),
	.w2(32'hbc0858d9),
	.w3(32'hbb918b05),
	.w4(32'h3b0d04b5),
	.w5(32'hbb9c13c2),
	.w6(32'hbbb3994b),
	.w7(32'h3a99e353),
	.w8(32'hbae24d8b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c7c2b),
	.w1(32'h3b39b25d),
	.w2(32'hbbd2d091),
	.w3(32'hb9f85fc3),
	.w4(32'h3b4412c2),
	.w5(32'hbb75005d),
	.w6(32'hb7a2a6c8),
	.w7(32'h3a913270),
	.w8(32'hb98ccf34),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae003c5),
	.w1(32'hbae88029),
	.w2(32'hbbaeca33),
	.w3(32'hba02d999),
	.w4(32'h3ad4d44d),
	.w5(32'hbac6e883),
	.w6(32'hbacba25c),
	.w7(32'h3b62f2c8),
	.w8(32'h3b1efd3d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18d5ec),
	.w1(32'h3b42967e),
	.w2(32'hbc18f4b3),
	.w3(32'h3a17b2dc),
	.w4(32'h3b3be47a),
	.w5(32'hbbdd5415),
	.w6(32'h3b8759f5),
	.w7(32'h3bc27696),
	.w8(32'hbaf6eedf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857713e),
	.w1(32'h377a6229),
	.w2(32'h380a2fa9),
	.w3(32'h37cc6b48),
	.w4(32'hb74dcf38),
	.w5(32'h3697d6dd),
	.w6(32'h373aa47e),
	.w7(32'hb741673f),
	.w8(32'h37280c47),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37899a2e),
	.w1(32'h36ac083b),
	.w2(32'hb7bf6115),
	.w3(32'hb68c0cf8),
	.w4(32'hb6adda10),
	.w5(32'hb68d11c8),
	.w6(32'hb6e0b1a6),
	.w7(32'hb811da63),
	.w8(32'hb7e13cd2),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e25df6),
	.w1(32'h38e9bee1),
	.w2(32'h388ba752),
	.w3(32'hb87a779e),
	.w4(32'hb83c104c),
	.w5(32'hb79c00a3),
	.w6(32'h3870a9cd),
	.w7(32'h38755858),
	.w8(32'hb87c8a21),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382196b0),
	.w1(32'hba8f2212),
	.w2(32'h38d6a9db),
	.w3(32'h3ab23b6a),
	.w4(32'hb873640f),
	.w5(32'h3a08b9f4),
	.w6(32'hb862fa9a),
	.w7(32'hba8c87b5),
	.w8(32'hb96ad52f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac01f9),
	.w1(32'hbc35ccf7),
	.w2(32'h3b9c59db),
	.w3(32'hbc45e5de),
	.w4(32'hbbae159a),
	.w5(32'h3c20e840),
	.w6(32'hbc73117d),
	.w7(32'hbb0eeb9c),
	.w8(32'h3c3492d3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b1e1b8),
	.w1(32'h39884318),
	.w2(32'h3ac3c8da),
	.w3(32'h3a48820f),
	.w4(32'h3a830f84),
	.w5(32'h3af6f428),
	.w6(32'hba428f4d),
	.w7(32'hba361bfe),
	.w8(32'h3a29289a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc248079),
	.w1(32'hbb6c4656),
	.w2(32'hbc0e7509),
	.w3(32'hbb8011ec),
	.w4(32'hba40df1e),
	.w5(32'hbb0d7c78),
	.w6(32'hbae0c92c),
	.w7(32'h3b8b9e2e),
	.w8(32'h3b297b4d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6badc9),
	.w1(32'hbbb1b4f9),
	.w2(32'hbc900c8c),
	.w3(32'hbc6c19ae),
	.w4(32'hbbea34b8),
	.w5(32'hbc54ea26),
	.w6(32'hbc08bc51),
	.w7(32'hbbedbd10),
	.w8(32'hbc22bc15),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201694),
	.w1(32'hbbccc343),
	.w2(32'h3b4f61eb),
	.w3(32'hbb9150c1),
	.w4(32'hbaa1404f),
	.w5(32'h3b4a545a),
	.w6(32'hbc3823e5),
	.w7(32'hbbcf5096),
	.w8(32'h3935d3ff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc406ef6),
	.w1(32'hbb508871),
	.w2(32'hbb050f7e),
	.w3(32'hbacec82f),
	.w4(32'h3ab58e59),
	.w5(32'h3bb9ef17),
	.w6(32'h39b0274a),
	.w7(32'h3a9b8bb7),
	.w8(32'h3a84256a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77ba0b),
	.w1(32'hbad5de75),
	.w2(32'h3b99053d),
	.w3(32'h3af203ec),
	.w4(32'h3bb4bfe9),
	.w5(32'h3c3ec239),
	.w6(32'hba950c7f),
	.w7(32'h3bd908c1),
	.w8(32'h3c294fb2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca46de9),
	.w1(32'hbb7ab9fa),
	.w2(32'hbc235354),
	.w3(32'hbc9c9224),
	.w4(32'hbb18308c),
	.w5(32'hbb8b9968),
	.w6(32'hbca55b6c),
	.w7(32'hbbaa046d),
	.w8(32'hbb5677ba),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47281a),
	.w1(32'hbbd70953),
	.w2(32'hbaf0c2fb),
	.w3(32'hbbad987e),
	.w4(32'h3b18395d),
	.w5(32'h3b9b9645),
	.w6(32'hbc2af5e2),
	.w7(32'hba806225),
	.w8(32'h3ba342bf),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53d9c1),
	.w1(32'hbbe3cf31),
	.w2(32'h3b27692e),
	.w3(32'hbbb3e905),
	.w4(32'h3b6377d8),
	.w5(32'h3c355993),
	.w6(32'hbc698ed7),
	.w7(32'hb9d3e887),
	.w8(32'h3c5d97f4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cfcf4),
	.w1(32'h3a1002c5),
	.w2(32'h36261141),
	.w3(32'h3a84d0bf),
	.w4(32'h3a4cd3ad),
	.w5(32'h3916da13),
	.w6(32'h3a98e274),
	.w7(32'h3a5e1932),
	.w8(32'h3a540ed1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33b829),
	.w1(32'h3ac47bed),
	.w2(32'hbc8f71f8),
	.w3(32'hbc136c32),
	.w4(32'h3bd4ce88),
	.w5(32'hbbb8645c),
	.w6(32'hbbc07af8),
	.w7(32'h3ba8b4d3),
	.w8(32'hbb898d01),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74cc63),
	.w1(32'hb97c9641),
	.w2(32'hbc0df5a4),
	.w3(32'hbb4f7006),
	.w4(32'h3bf5fe71),
	.w5(32'hb9b33f52),
	.w6(32'h3b84bcd7),
	.w7(32'h3bd7d32a),
	.w8(32'hb9dbc029),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1b6e8),
	.w1(32'hba51cbbf),
	.w2(32'hba414be2),
	.w3(32'hbc284a3d),
	.w4(32'h3b623106),
	.w5(32'h3c1e07e0),
	.w6(32'h3c5433cc),
	.w7(32'h3cc25754),
	.w8(32'h3c5b1498),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3b9c49),
	.w1(32'hbc542314),
	.w2(32'h3d125124),
	.w3(32'hbd025a15),
	.w4(32'hbc2ae87d),
	.w5(32'h3cfea888),
	.w6(32'hbd0e3f6b),
	.w7(32'hbc787883),
	.w8(32'h3cca3a1d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc336cfb),
	.w1(32'hbb99190c),
	.w2(32'hbbeb7444),
	.w3(32'hbb097f02),
	.w4(32'h3bb87007),
	.w5(32'h3b7b8e07),
	.w6(32'hbb0385d5),
	.w7(32'h3c3939b5),
	.w8(32'h3c0c3d35),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb94934),
	.w1(32'h3a0d210f),
	.w2(32'h3a462c5e),
	.w3(32'hbc7ec1e7),
	.w4(32'hba4c5afe),
	.w5(32'h3bc2de74),
	.w6(32'h3b31ee5b),
	.w7(32'h3c62b542),
	.w8(32'h3b5b6e07),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39911a82),
	.w1(32'h3a7dc8ef),
	.w2(32'h3a30c777),
	.w3(32'h3a1fa97c),
	.w4(32'hb7cbd392),
	.w5(32'h39bffb38),
	.w6(32'h39d03b90),
	.w7(32'h3a862f2d),
	.w8(32'h3a892dbb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcefc263),
	.w1(32'hbc285ec6),
	.w2(32'hbbaeb2fb),
	.w3(32'hbc5a9b64),
	.w4(32'hbb52e293),
	.w5(32'h3c8699f9),
	.w6(32'h3bd30dce),
	.w7(32'h3c067bbf),
	.w8(32'h3c1eb349),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc309b83),
	.w1(32'h3a8efa3a),
	.w2(32'h3c078a9f),
	.w3(32'hbada3049),
	.w4(32'hb90f674c),
	.w5(32'h3c2c6ea9),
	.w6(32'h3bb46cbf),
	.w7(32'h3b604fc9),
	.w8(32'h3c2a06ac),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7a7a0),
	.w1(32'h394b0ef9),
	.w2(32'h390dfa60),
	.w3(32'hb8f47e56),
	.w4(32'h3a08765d),
	.w5(32'h396754a9),
	.w6(32'hb9e7f7c6),
	.w7(32'h39058218),
	.w8(32'hb8ab8507),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69d8fa),
	.w1(32'hbb556eb8),
	.w2(32'hbb4eca7f),
	.w3(32'hb94f6d2b),
	.w4(32'h3a1e54a8),
	.w5(32'hbafa2274),
	.w6(32'hbb684ac6),
	.w7(32'hb963924c),
	.w8(32'hb9f2564a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0aa9c),
	.w1(32'hba5f4b14),
	.w2(32'hbc3b02f7),
	.w3(32'hbb9d81e0),
	.w4(32'hba895e19),
	.w5(32'hbc155677),
	.w6(32'hbb956ffe),
	.w7(32'h392bf2fd),
	.w8(32'hbbbfe348),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912e13),
	.w1(32'hba98759a),
	.w2(32'hbb5ba599),
	.w3(32'h3adf8705),
	.w4(32'h3bb91e2b),
	.w5(32'h3b8e2631),
	.w6(32'h389b0bab),
	.w7(32'h3c0a7736),
	.w8(32'h3bf57ef0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26452e),
	.w1(32'hbc4b001d),
	.w2(32'hbba4ae79),
	.w3(32'hbb8c0ce1),
	.w4(32'hbb81b530),
	.w5(32'h390ed364),
	.w6(32'hbc1d821d),
	.w7(32'hbbae6766),
	.w8(32'h39ffdda2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e2a7),
	.w1(32'hbb58ad43),
	.w2(32'hbb82dc8c),
	.w3(32'hbbc04868),
	.w4(32'h3a1f6b42),
	.w5(32'h3af5c896),
	.w6(32'hbb90b5d3),
	.w7(32'h3b1b6a64),
	.w8(32'h3b8f7690),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8131d6),
	.w1(32'h3abb22be),
	.w2(32'h3b475187),
	.w3(32'hbc06805f),
	.w4(32'h3b8f5c9d),
	.w5(32'h3b95c99a),
	.w6(32'hbb13c475),
	.w7(32'h3bfd7520),
	.w8(32'h3babaa84),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1a8c7),
	.w1(32'hbac3f202),
	.w2(32'hbc2ae1ed),
	.w3(32'hbbb61341),
	.w4(32'h3a02beab),
	.w5(32'hbbb86a01),
	.w6(32'hbbe44569),
	.w7(32'hbacd113a),
	.w8(32'hbbb4acff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82ac0e),
	.w1(32'hba3f9aa2),
	.w2(32'hbb312d9b),
	.w3(32'hbab4df73),
	.w4(32'h3b4da7b3),
	.w5(32'h3a090bc4),
	.w6(32'hbab371fa),
	.w7(32'h3ba3db19),
	.w8(32'h3b02b880),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907519e),
	.w1(32'hb90bd6a2),
	.w2(32'hb7d5eeee),
	.w3(32'hb904ed14),
	.w4(32'hb8299312),
	.w5(32'h37c8fe43),
	.w6(32'hb88805a2),
	.w7(32'hb7136fc2),
	.w8(32'h38e2157e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9a27d),
	.w1(32'hbaca7574),
	.w2(32'hba57ea78),
	.w3(32'hba9662ae),
	.w4(32'hba848ac1),
	.w5(32'hb898ad59),
	.w6(32'hbaf44802),
	.w7(32'hba893351),
	.w8(32'hba5b70e9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8304516),
	.w1(32'h38c0bf3b),
	.w2(32'h38d81794),
	.w3(32'hb9111578),
	.w4(32'h38d9132f),
	.w5(32'h38d3c0b5),
	.w6(32'hb8c0214e),
	.w7(32'h388e3b04),
	.w8(32'h3738881f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d81f8),
	.w1(32'h3a9e6661),
	.w2(32'h3a9099b3),
	.w3(32'h39b6d1d9),
	.w4(32'h3ab017dc),
	.w5(32'h3a48157b),
	.w6(32'h38b5966a),
	.w7(32'h3a74805f),
	.w8(32'h3a5d1698),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb31b8),
	.w1(32'h397c8078),
	.w2(32'hbb3645b1),
	.w3(32'hbabe9313),
	.w4(32'h3bc3c6a0),
	.w5(32'h3b3f3466),
	.w6(32'hbb261c3a),
	.w7(32'h3c0a7bf3),
	.w8(32'h3bbec87a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f374),
	.w1(32'hb83303b2),
	.w2(32'h38f383e7),
	.w3(32'hba0869c1),
	.w4(32'h3a766bc6),
	.w5(32'h39e8f619),
	.w6(32'hb9ce7593),
	.w7(32'h3a8acc8a),
	.w8(32'h3a54cf76),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd33754),
	.w1(32'h3a89359b),
	.w2(32'hbb31b1fd),
	.w3(32'hbaf71434),
	.w4(32'h3972e37a),
	.w5(32'hb8004370),
	.w6(32'h3ba861bd),
	.w7(32'h3b69d21a),
	.w8(32'hbac5366f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc982a43),
	.w1(32'hbc3ba021),
	.w2(32'h3ada5c1f),
	.w3(32'hbc2fe7d4),
	.w4(32'hb926ba4f),
	.w5(32'h3c1a9e03),
	.w6(32'hbc7a3fe3),
	.w7(32'hbb8fabdd),
	.w8(32'h3be63829),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab0ac1),
	.w1(32'hb6abfac3),
	.w2(32'hb93bf16f),
	.w3(32'h39e25179),
	.w4(32'h3988370d),
	.w5(32'h38baeb08),
	.w6(32'h39c18be9),
	.w7(32'h39d7632e),
	.w8(32'h396f668a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db5251),
	.w1(32'h39dcee08),
	.w2(32'hb8be87cc),
	.w3(32'hb9a263c8),
	.w4(32'h3a2e8e9c),
	.w5(32'hb72b84bf),
	.w6(32'hb9fe5332),
	.w7(32'hb8569304),
	.w8(32'hba04862f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390079c2),
	.w1(32'h38484111),
	.w2(32'h38aa25fb),
	.w3(32'h38b15d86),
	.w4(32'hb79f0d56),
	.w5(32'h381fe094),
	.w6(32'h387f20ed),
	.w7(32'hb8395ec4),
	.w8(32'h3655fef4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ddd33),
	.w1(32'hbaebc4f7),
	.w2(32'hba50301c),
	.w3(32'hbb82e387),
	.w4(32'hbb117354),
	.w5(32'hbaa831f5),
	.w6(32'hbb6fab95),
	.w7(32'hbb033705),
	.w8(32'hbaa55212),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ba8e7),
	.w1(32'hbab1a572),
	.w2(32'hbc2a3d1e),
	.w3(32'h3b9a3af9),
	.w4(32'h3a4c3d9b),
	.w5(32'hbc0699cf),
	.w6(32'h3c3979b3),
	.w7(32'h3c16ee7a),
	.w8(32'hbb57851d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8878ee),
	.w1(32'h3b48cf7a),
	.w2(32'hbc8569bd),
	.w3(32'hbbbbb8a8),
	.w4(32'h3b81c0d3),
	.w5(32'hbc371c5d),
	.w6(32'hba63f15e),
	.w7(32'h3b9e3691),
	.w8(32'hbbe11f88),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0961ad),
	.w1(32'hba1f92fd),
	.w2(32'hba67f57b),
	.w3(32'hba529c3f),
	.w4(32'hba8311ec),
	.w5(32'h399fffd1),
	.w6(32'h3ae92423),
	.w7(32'h39d3acb7),
	.w8(32'hb95553a1),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb202b),
	.w1(32'hbb1d37ce),
	.w2(32'hbb365f41),
	.w3(32'hbb98da0d),
	.w4(32'hba84c817),
	.w5(32'hba36d04d),
	.w6(32'hbb568230),
	.w7(32'h3907167c),
	.w8(32'h393140d1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbab6a8),
	.w1(32'hbac6ab01),
	.w2(32'hba0a7b76),
	.w3(32'hbb5e56cf),
	.w4(32'h3ae758a6),
	.w5(32'h3afabab4),
	.w6(32'hbb927847),
	.w7(32'h3ab885a4),
	.w8(32'h3b34d99b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6da62d),
	.w1(32'hb9a95c52),
	.w2(32'hbb9c6d1c),
	.w3(32'hbb8d74e2),
	.w4(32'hb9c8b0ae),
	.w5(32'hbb1ad84c),
	.w6(32'hbb773af8),
	.w7(32'hbab3b7df),
	.w8(32'h3892a935),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01f4f8),
	.w1(32'hbba57aad),
	.w2(32'hbbaed156),
	.w3(32'hbb1f7a30),
	.w4(32'h3a7caf57),
	.w5(32'hbb34a853),
	.w6(32'hbbe9f8ee),
	.w7(32'hbad661ad),
	.w8(32'hb9ac3c1c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb971d35),
	.w1(32'h3a3da9ed),
	.w2(32'hbca42351),
	.w3(32'hbba078ef),
	.w4(32'h3b987d24),
	.w5(32'hbc451e91),
	.w6(32'h3ba38c9d),
	.w7(32'h3af5278c),
	.w8(32'hbc1cb22c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d173a),
	.w1(32'hbb818288),
	.w2(32'h39d5e60a),
	.w3(32'hbbf1f9fc),
	.w4(32'hba32e812),
	.w5(32'h3bae6eee),
	.w6(32'hbc3ad3db),
	.w7(32'hba8cacdd),
	.w8(32'h3b934e68),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ffa1b),
	.w1(32'hbbad5717),
	.w2(32'hbbeabf9a),
	.w3(32'hbb90d76c),
	.w4(32'h3af14b79),
	.w5(32'h3a68db76),
	.w6(32'hbb556edb),
	.w7(32'h3aa71eca),
	.w8(32'h389a13de),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4711d8),
	.w1(32'h3aa5d705),
	.w2(32'hbc8522f8),
	.w3(32'hbc78a617),
	.w4(32'hba375669),
	.w5(32'hbc37665b),
	.w6(32'h3b2bb15f),
	.w7(32'h3c01de6d),
	.w8(32'hbc172576),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e8341),
	.w1(32'hbb9b2657),
	.w2(32'h3ae5d512),
	.w3(32'hbbc304e3),
	.w4(32'h3a2146ed),
	.w5(32'h3bd1bed8),
	.w6(32'hbbe18e67),
	.w7(32'h3b06696c),
	.w8(32'h3bccba19),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba661cf),
	.w1(32'hb8fec166),
	.w2(32'hbbc81c5c),
	.w3(32'hbbb715bc),
	.w4(32'hb9a0dec4),
	.w5(32'hbb4e3da9),
	.w6(32'hbb2b56f2),
	.w7(32'hbb164fbd),
	.w8(32'hbb524d74),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad78417),
	.w1(32'hb6ecc0c4),
	.w2(32'hbafb27d0),
	.w3(32'h380c1a0e),
	.w4(32'h3b08ace7),
	.w5(32'h39c2079b),
	.w6(32'hb9a83137),
	.w7(32'h3b2df360),
	.w8(32'h3acb97f5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc680021),
	.w1(32'hbc043611),
	.w2(32'h3af74319),
	.w3(32'hbbcb795f),
	.w4(32'hbab40b96),
	.w5(32'h3bb267c2),
	.w6(32'hbc716532),
	.w7(32'hbb3be7f0),
	.w8(32'h3bfa69ef),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc189ffd),
	.w1(32'hbbb6c896),
	.w2(32'hba7d1680),
	.w3(32'hbbb9400b),
	.w4(32'hbac10bd3),
	.w5(32'h3b512acb),
	.w6(32'hbb8df6db),
	.w7(32'h39c3731b),
	.w8(32'h3b90382c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999d3eb),
	.w1(32'hb92a7447),
	.w2(32'hb9b5d513),
	.w3(32'h39a06be4),
	.w4(32'h37eeeb99),
	.w5(32'hb98de216),
	.w6(32'h394e7094),
	.w7(32'h3890c9a7),
	.w8(32'hb959dc8c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e9e615),
	.w1(32'h38097c9d),
	.w2(32'h3811fd43),
	.w3(32'hb89f27d2),
	.w4(32'hb8cda3ac),
	.w5(32'hb8e100dd),
	.w6(32'h391910e5),
	.w7(32'h38462d6b),
	.w8(32'h38f5ee2b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96c854),
	.w1(32'hbaab0176),
	.w2(32'h3b031247),
	.w3(32'hbb4f3e37),
	.w4(32'h39b9ba15),
	.w5(32'h3baff015),
	.w6(32'hb960c443),
	.w7(32'h39b7618c),
	.w8(32'h3b9f6cc1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe1173),
	.w1(32'hbc1a4c5b),
	.w2(32'hbaa34324),
	.w3(32'hbc57ae74),
	.w4(32'hbad8c29b),
	.w5(32'h3c076e0c),
	.w6(32'hbc4edcf6),
	.w7(32'hbb27e7d0),
	.w8(32'h3c0cfef5),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7709a),
	.w1(32'h3ae67439),
	.w2(32'hbc567795),
	.w3(32'hba95a8ff),
	.w4(32'h3c22bd2f),
	.w5(32'hbb360e38),
	.w6(32'h3aa1a328),
	.w7(32'h3c504a1e),
	.w8(32'h3ab85e8a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38931016),
	.w1(32'h37a963ba),
	.w2(32'hb8e3e43e),
	.w3(32'hb88a339d),
	.w4(32'hb8b02831),
	.w5(32'hb91a8e22),
	.w6(32'hb96e2c6f),
	.w7(32'hb9616b15),
	.w8(32'hb8ed44f5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c864),
	.w1(32'hba1ab793),
	.w2(32'hbc5a28d4),
	.w3(32'hbb89130c),
	.w4(32'h3b80b8c6),
	.w5(32'hbc026902),
	.w6(32'hbb06d586),
	.w7(32'h3bc30c03),
	.w8(32'hba7d7c4c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c001),
	.w1(32'hbb14544f),
	.w2(32'hbbcaa5fc),
	.w3(32'hbb90f062),
	.w4(32'h3ac62d69),
	.w5(32'hbafe6a54),
	.w6(32'hbb8c20e4),
	.w7(32'h3b53ee7a),
	.w8(32'h3a602784),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24f2b4),
	.w1(32'h3ad78f0a),
	.w2(32'hbc240e01),
	.w3(32'hbbc4a834),
	.w4(32'h3ba77326),
	.w5(32'hbb56b5fa),
	.w6(32'h389f04f3),
	.w7(32'h3bf64a9e),
	.w8(32'hbbbcbcfd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40c0f6),
	.w1(32'hbb4feb42),
	.w2(32'hbbda33b3),
	.w3(32'h3c0d95b4),
	.w4(32'h3c848ee6),
	.w5(32'h3bc31831),
	.w6(32'hbaa5749b),
	.w7(32'h3c786a70),
	.w8(32'h3c37b918),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a9422),
	.w1(32'hbc02be78),
	.w2(32'hbb010134),
	.w3(32'hbc0ee242),
	.w4(32'hbbe2295d),
	.w5(32'hbacdd1d2),
	.w6(32'hbc0fbcf3),
	.w7(32'hbbb46b79),
	.w8(32'hbadf4bee),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a685634),
	.w1(32'h3a4ce67b),
	.w2(32'h3ae2bfe1),
	.w3(32'h3993702a),
	.w4(32'hb87fece8),
	.w5(32'h3a751ce9),
	.w6(32'h38d9c3af),
	.w7(32'h3942bb2d),
	.w8(32'h3a9ab9f6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e119f),
	.w1(32'hbb0a65f0),
	.w2(32'h3abb19c7),
	.w3(32'hbbf6e58e),
	.w4(32'h3aead68a),
	.w5(32'h3ba0a7c8),
	.w6(32'hbc1490a5),
	.w7(32'h3b16aaa0),
	.w8(32'h3b9437d7),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0a24b),
	.w1(32'hbc0887c0),
	.w2(32'h3ab573ae),
	.w3(32'hbc2e9cf4),
	.w4(32'hbb825421),
	.w5(32'h3b0df94b),
	.w6(32'hbc740b90),
	.w7(32'hbb95a914),
	.w8(32'hb9abd806),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbd061),
	.w1(32'h3a77515d),
	.w2(32'h3ba1a31c),
	.w3(32'hbb88d411),
	.w4(32'h3b72690e),
	.w5(32'h3bce70f8),
	.w6(32'hbbfc04a9),
	.w7(32'h3b0fe6c5),
	.w8(32'h3ba2452a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba976cc8),
	.w1(32'h39ec4d69),
	.w2(32'hbb29b018),
	.w3(32'hba8924d0),
	.w4(32'hba37fcd2),
	.w5(32'hbb105be1),
	.w6(32'h3b0491b0),
	.w7(32'h3a3625e4),
	.w8(32'hbb080fc3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f6fbc),
	.w1(32'hba8de644),
	.w2(32'hbabf0d8f),
	.w3(32'hbab5843e),
	.w4(32'hba8b31ec),
	.w5(32'hba97ac53),
	.w6(32'hba74f0aa),
	.w7(32'hbaaa6dfb),
	.w8(32'hba914b36),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37f0f8),
	.w1(32'hbae72f31),
	.w2(32'hbc077ec0),
	.w3(32'hbbfba631),
	.w4(32'h39c5ef24),
	.w5(32'hbab71601),
	.w6(32'hbb9d1eb3),
	.w7(32'h3ac617d0),
	.w8(32'hbab41f33),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecd2fc),
	.w1(32'h3ab23e5f),
	.w2(32'hb9da2692),
	.w3(32'h3ae4bfcb),
	.w4(32'h3aad39fc),
	.w5(32'hb9ae1845),
	.w6(32'h3b049551),
	.w7(32'h3ae69be0),
	.w8(32'h39ce97b2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ec1c0),
	.w1(32'hbac6318c),
	.w2(32'hbabdb095),
	.w3(32'hb931cf0d),
	.w4(32'h3b48d894),
	.w5(32'h3ad4af45),
	.w6(32'hbabefd13),
	.w7(32'h3b9d9b59),
	.w8(32'h3baa0deb),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e73bd6),
	.w1(32'h38940f05),
	.w2(32'hb832a92b),
	.w3(32'hb8f3e9b1),
	.w4(32'h39b10960),
	.w5(32'h39717b7a),
	.w6(32'hb7b927d9),
	.w7(32'hb78d39cf),
	.w8(32'h3956e7a6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b056868),
	.w1(32'h3bf4e183),
	.w2(32'hba31d832),
	.w3(32'h3b559f5f),
	.w4(32'h3c288e9b),
	.w5(32'h3b3ca339),
	.w6(32'h3b5bb142),
	.w7(32'h3c20ebc1),
	.w8(32'h3adf144d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ca07f),
	.w1(32'hb8037a2f),
	.w2(32'hb8294223),
	.w3(32'h3813575d),
	.w4(32'hb8ab3757),
	.w5(32'hb8ed683e),
	.w6(32'hb7b4121a),
	.w7(32'hb94ed080),
	.w8(32'hb91fe85d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7399ff),
	.w1(32'hb96567f9),
	.w2(32'hb9e8f326),
	.w3(32'hba6825ff),
	.w4(32'hb9c28b11),
	.w5(32'hba0ba2d1),
	.w6(32'hba387314),
	.w7(32'hb9b79648),
	.w8(32'hba75cd12),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2431b9),
	.w1(32'hbbaa0ca2),
	.w2(32'hba8f9b5e),
	.w3(32'hbc095d55),
	.w4(32'hbae58699),
	.w5(32'h3a9e3412),
	.w6(32'hbc2f45ce),
	.w7(32'hbaf040e6),
	.w8(32'h3b581b5a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9800b3),
	.w1(32'hbb5302ed),
	.w2(32'hbc2d8230),
	.w3(32'hbbaa5844),
	.w4(32'h3b04bf28),
	.w5(32'hbbb57878),
	.w6(32'hba7feaad),
	.w7(32'h3c38691d),
	.w8(32'h3b4ddb2c),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb972235),
	.w1(32'h3af6e3c3),
	.w2(32'h3b187c23),
	.w3(32'hbb9eee69),
	.w4(32'h3afd310e),
	.w5(32'h3b0179ac),
	.w6(32'hbbd4027a),
	.w7(32'h38be7468),
	.w8(32'hba1b75e2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ea54),
	.w1(32'hba159944),
	.w2(32'hbb5adce9),
	.w3(32'hbb69c77c),
	.w4(32'h3b53f585),
	.w5(32'h3adadd2b),
	.w6(32'hbbaec648),
	.w7(32'h3b62a057),
	.w8(32'h3b5e0b25),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba041cd3),
	.w1(32'h38c77ade),
	.w2(32'hbaa77efb),
	.w3(32'h3a374c4c),
	.w4(32'h3b36cba2),
	.w5(32'h3a7366c9),
	.w6(32'hbb4d1290),
	.w7(32'h3a776490),
	.w8(32'h3aa6d26f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc692807),
	.w1(32'h3ada790c),
	.w2(32'hbc8e194f),
	.w3(32'hbc20d5c0),
	.w4(32'h3bf3c732),
	.w5(32'hbbc8de84),
	.w6(32'hbc7593ee),
	.w7(32'h3bb04029),
	.w8(32'hbb9d17ef),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45f2f4),
	.w1(32'hbb197b77),
	.w2(32'hbbf32816),
	.w3(32'hbbc874d3),
	.w4(32'h3b4beb88),
	.w5(32'h3a844788),
	.w6(32'hbba82a7a),
	.w7(32'h3b5865e1),
	.w8(32'h3adb5752),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9a22),
	.w1(32'h3b555857),
	.w2(32'hbc94fdc8),
	.w3(32'hbb1d1394),
	.w4(32'h3b86e6d3),
	.w5(32'hbc4a3363),
	.w6(32'h3a815b2c),
	.w7(32'h3c08c0fa),
	.w8(32'hbbc9d3ee),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2cbe2),
	.w1(32'h39814d7d),
	.w2(32'h39cd3038),
	.w3(32'h3927329d),
	.w4(32'h39bc39bd),
	.w5(32'h3a1499d0),
	.w6(32'h3a02e13a),
	.w7(32'h39af1432),
	.w8(32'h3a62327b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbc0d9),
	.w1(32'hba37e581),
	.w2(32'hbc0d834e),
	.w3(32'hbbe96a55),
	.w4(32'hbaa45b60),
	.w5(32'hbba34d5b),
	.w6(32'hbba7748b),
	.w7(32'h3ac619fc),
	.w8(32'hbb06e544),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a5b5a),
	.w1(32'h38ddd308),
	.w2(32'h37ca4548),
	.w3(32'h3976c560),
	.w4(32'h37f36780),
	.w5(32'hb818045c),
	.w6(32'h3964724c),
	.w7(32'h384c21ba),
	.w8(32'hb830adc5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad40f7),
	.w1(32'h3a6c2c4c),
	.w2(32'hbb8d4687),
	.w3(32'h3b216e1f),
	.w4(32'h3aec2de5),
	.w5(32'hbacbc379),
	.w6(32'h3afcd252),
	.w7(32'h3ada5acc),
	.w8(32'hbaa94fc1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6804b6),
	.w1(32'hb97528a6),
	.w2(32'h3a0887ff),
	.w3(32'hbb35fbea),
	.w4(32'h3a166966),
	.w5(32'h3ad66cc1),
	.w6(32'hbb0bbefe),
	.w7(32'h39d6ee39),
	.w8(32'h3a9f6258),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb3bce),
	.w1(32'h3a07696d),
	.w2(32'hbb609dde),
	.w3(32'hbb6c4f4e),
	.w4(32'h3b31a18e),
	.w5(32'hbab65d91),
	.w6(32'hbc00640e),
	.w7(32'h3a882d0b),
	.w8(32'hba98b694),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6f322),
	.w1(32'h378d5543),
	.w2(32'h3607d9ef),
	.w3(32'h38c374a1),
	.w4(32'h360e5144),
	.w5(32'hb70c5200),
	.w6(32'h38b0dc5d),
	.w7(32'h38050a88),
	.w8(32'h3826a2cf),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38716c72),
	.w1(32'h3935a1b5),
	.w2(32'h36825a3d),
	.w3(32'hb8de4e8e),
	.w4(32'hb857170d),
	.w5(32'hb71e4ef4),
	.w6(32'hb81beac7),
	.w7(32'h37bf1418),
	.w8(32'h387562c4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91887),
	.w1(32'hbb1332b6),
	.w2(32'hb9c615eb),
	.w3(32'hbadac821),
	.w4(32'h3acb0bd6),
	.w5(32'h3b3eadd1),
	.w6(32'hbb34bc59),
	.w7(32'h3acced4c),
	.w8(32'h3af084f5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9644b6),
	.w1(32'hbbdbbd8f),
	.w2(32'hb9ad3835),
	.w3(32'hbc3aa3f4),
	.w4(32'hbaa70283),
	.w5(32'h3b85be85),
	.w6(32'hbc84c02f),
	.w7(32'hbb9cc8b8),
	.w8(32'hbaed9a2c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc512dd7),
	.w1(32'h3b9d9857),
	.w2(32'h3c12b013),
	.w3(32'hbc2e4a98),
	.w4(32'h3a3f139d),
	.w5(32'h3c435182),
	.w6(32'h3aebccc1),
	.w7(32'h3b0bf386),
	.w8(32'h3bbc6ec9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba868c3c),
	.w1(32'h3a0acdd7),
	.w2(32'hba1f8888),
	.w3(32'hba4194ce),
	.w4(32'h39c8d829),
	.w5(32'hba48f31d),
	.w6(32'hbab6a6c1),
	.w7(32'h3a144b04),
	.w8(32'hba1fdd65),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48ffb8),
	.w1(32'h3b7b911e),
	.w2(32'hbcfd7543),
	.w3(32'hbbcc2186),
	.w4(32'h3c6d8fe6),
	.w5(32'hbc63d5fd),
	.w6(32'h3b0d75d2),
	.w7(32'h3ccc13fa),
	.w8(32'hbbf4e84a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc27d5e),
	.w1(32'hbc65196b),
	.w2(32'hbba8fe70),
	.w3(32'hbc0e1622),
	.w4(32'h3b1baa3d),
	.w5(32'h3b051696),
	.w6(32'hbcb3b459),
	.w7(32'h3a921963),
	.w8(32'h3c173252),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69b473),
	.w1(32'h3ae569ee),
	.w2(32'h3a1fc082),
	.w3(32'h3ae477b8),
	.w4(32'h3a1494ea),
	.w5(32'h39f9cdfa),
	.w6(32'h3baf5132),
	.w7(32'h3ab37596),
	.w8(32'h39657657),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923f1f3),
	.w1(32'hb77d583f),
	.w2(32'hb8e9d2ed),
	.w3(32'h388a9c35),
	.w4(32'hb8f7072f),
	.w5(32'hb9836585),
	.w6(32'h37c5006e),
	.w7(32'hb9712cc8),
	.w8(32'hb8d5ca92),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb700bb05),
	.w1(32'hb90c8467),
	.w2(32'h388dcfdc),
	.w3(32'hb92c1488),
	.w4(32'hb9d2cce7),
	.w5(32'hb987b2d2),
	.w6(32'hb9096a02),
	.w7(32'hb9ad6aa2),
	.w8(32'hb840fee2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ff0bc),
	.w1(32'h38125494),
	.w2(32'h3788b40f),
	.w3(32'h39026e14),
	.w4(32'hb7859f1e),
	.w5(32'hb82e9336),
	.w6(32'h3930e936),
	.w7(32'hb693625b),
	.w8(32'hb76672ba),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafe61f),
	.w1(32'hbaae8ddb),
	.w2(32'hba8e12b5),
	.w3(32'hbb3ae088),
	.w4(32'hb4e5bf80),
	.w5(32'h3a12623b),
	.w6(32'h3b107e6c),
	.w7(32'hbb16692b),
	.w8(32'hbb2c7de3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47e84c),
	.w1(32'hbbc6d63d),
	.w2(32'hbc02c84a),
	.w3(32'hbbb8bc49),
	.w4(32'h39bdbe0b),
	.w5(32'hbab84e68),
	.w6(32'hbb094664),
	.w7(32'h3ad850ec),
	.w8(32'hba110eea),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bfdc9),
	.w1(32'hbb893a5b),
	.w2(32'hbbd85252),
	.w3(32'hbbd2af8f),
	.w4(32'h3be13006),
	.w5(32'h3bb60f5d),
	.w6(32'hbc18682f),
	.w7(32'h3bddf4e9),
	.w8(32'h3c038d0a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8489ad),
	.w1(32'hba1f9697),
	.w2(32'hba0e5d0f),
	.w3(32'hbaef717c),
	.w4(32'h3ab6f9ab),
	.w5(32'h3b01e0c0),
	.w6(32'hbadb6cdd),
	.w7(32'h3adca5a0),
	.w8(32'h3a99afa3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd22bb),
	.w1(32'hbac1d1ac),
	.w2(32'hbc74a25a),
	.w3(32'hbb403eb4),
	.w4(32'h3933236d),
	.w5(32'hbc04a9b5),
	.w6(32'hba9b7055),
	.w7(32'h3ab34144),
	.w8(32'hbb209d24),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd595e),
	.w1(32'hbb9a8b06),
	.w2(32'hbb34471d),
	.w3(32'hbbec0a00),
	.w4(32'h3b48aaab),
	.w5(32'h3c8d797c),
	.w6(32'h3b936ccd),
	.w7(32'h3bcab60c),
	.w8(32'hbbdcba4d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf9644),
	.w1(32'hbb179e74),
	.w2(32'h3a6bc99b),
	.w3(32'h3b4d7e5c),
	.w4(32'hbbab3c3f),
	.w5(32'hbb10fb66),
	.w6(32'hbbc05dda),
	.w7(32'hbc0ce24d),
	.w8(32'hbb31d688),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16c83b),
	.w1(32'hbacabe91),
	.w2(32'hbaa6c3e5),
	.w3(32'hbbb8da3e),
	.w4(32'hbc04c227),
	.w5(32'h3a40c94f),
	.w6(32'h3c2a03e1),
	.w7(32'hbbc42e65),
	.w8(32'h3b7ecaeb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e7a2),
	.w1(32'hbb422144),
	.w2(32'hbb922ea3),
	.w3(32'hbbc49547),
	.w4(32'hbadd01b9),
	.w5(32'h3c61c8da),
	.w6(32'hba7fb06a),
	.w7(32'hb9147f59),
	.w8(32'hb9077b70),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ecd01),
	.w1(32'hbbb8bed2),
	.w2(32'hbb86efcc),
	.w3(32'h3a865948),
	.w4(32'hba4f0bb5),
	.w5(32'h3c097e90),
	.w6(32'hbc005937),
	.w7(32'h3c10d89a),
	.w8(32'h3c1e7414),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bb496),
	.w1(32'hbbe3b66e),
	.w2(32'h3a67e4cc),
	.w3(32'hbbccb27b),
	.w4(32'hbb970bc8),
	.w5(32'h3c28a80c),
	.w6(32'hbca2ce34),
	.w7(32'hbbbd6934),
	.w8(32'h3a0cbf30),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bf679),
	.w1(32'hbbb5f051),
	.w2(32'h3a6e754d),
	.w3(32'hbc0baa7d),
	.w4(32'h3a0a7a57),
	.w5(32'h3c0509e0),
	.w6(32'hbc7a5fda),
	.w7(32'h3b9a5ee5),
	.w8(32'h3c28d8dd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30d9b3),
	.w1(32'hbbbbfd18),
	.w2(32'hba863a74),
	.w3(32'hbaca54f3),
	.w4(32'hbbf70461),
	.w5(32'hbc0e1543),
	.w6(32'h3a33fbdf),
	.w7(32'h3aeeb814),
	.w8(32'h3afc01cd),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb16b77),
	.w1(32'hbc5af838),
	.w2(32'hba4fb203),
	.w3(32'hbca31f61),
	.w4(32'hbb07a405),
	.w5(32'hbaa6960a),
	.w6(32'hbca7f422),
	.w7(32'hbba672b6),
	.w8(32'h3c0608fa),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ff526),
	.w1(32'h3b077a6a),
	.w2(32'hb905d086),
	.w3(32'h3ac90c5c),
	.w4(32'h3bad8c80),
	.w5(32'h3ad3c0f3),
	.w6(32'h3aa28610),
	.w7(32'hbb155267),
	.w8(32'h3bb49f93),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2964d),
	.w1(32'h3c497359),
	.w2(32'hbac35e69),
	.w3(32'h3a594f24),
	.w4(32'h3c8915ca),
	.w5(32'hba2db893),
	.w6(32'h3bda32c5),
	.w7(32'h3c60be72),
	.w8(32'h3bb03f0f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3587f),
	.w1(32'hbb147e14),
	.w2(32'h3b4ced98),
	.w3(32'h3c0354f9),
	.w4(32'h3a0ddd2d),
	.w5(32'h3b741395),
	.w6(32'h3c0d01f2),
	.w7(32'h3b40578a),
	.w8(32'h3b985f3e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5213f4),
	.w1(32'hbb812d79),
	.w2(32'h3ac436d5),
	.w3(32'h3b6f2631),
	.w4(32'h3b5d68dc),
	.w5(32'h3a361910),
	.w6(32'h3b29339d),
	.w7(32'hbb13c8f5),
	.w8(32'h3b490766),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bdc98),
	.w1(32'hbaac18c8),
	.w2(32'h3b819186),
	.w3(32'hbba12944),
	.w4(32'h3c185ff4),
	.w5(32'h3c20522c),
	.w6(32'hbb37f3a2),
	.w7(32'h3cc56cb3),
	.w8(32'h3c635f0b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab42933),
	.w1(32'h3a3f0495),
	.w2(32'hbc5c8031),
	.w3(32'h3c0d8bf3),
	.w4(32'h3b7c2df1),
	.w5(32'hbb962c46),
	.w6(32'hbb3ea66d),
	.w7(32'h3c4c078d),
	.w8(32'h3bf69c8b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc894ceb),
	.w1(32'hbc2c64ef),
	.w2(32'hbc513d1e),
	.w3(32'hbbe26cb4),
	.w4(32'h3b82bc79),
	.w5(32'h3c428331),
	.w6(32'hbbed931c),
	.w7(32'h3b97a542),
	.w8(32'h3a86c2c0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab38907),
	.w1(32'h38a865ce),
	.w2(32'hbc16cf91),
	.w3(32'hbbd2a508),
	.w4(32'hbb6cc783),
	.w5(32'hbc4d3463),
	.w6(32'hbc1018f5),
	.w7(32'hbb2f881a),
	.w8(32'hbc488c08),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11844e),
	.w1(32'hbb3b1987),
	.w2(32'hbc2b6a32),
	.w3(32'h39c41cac),
	.w4(32'h39edd75f),
	.w5(32'h3c56beb9),
	.w6(32'h3b139f7c),
	.w7(32'h3b922437),
	.w8(32'hbae7ae3e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f4b3a),
	.w1(32'hbb4d0304),
	.w2(32'hba9c7014),
	.w3(32'h3ba71577),
	.w4(32'hbbefcec8),
	.w5(32'hba9cee06),
	.w6(32'hbaebe898),
	.w7(32'h3bd19af0),
	.w8(32'h3c2a70cd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a90f),
	.w1(32'h3bc59ceb),
	.w2(32'h3bccc7dd),
	.w3(32'h3be8479a),
	.w4(32'h3aec1ecb),
	.w5(32'hba93ac2c),
	.w6(32'h3c5550eb),
	.w7(32'h3c59ca41),
	.w8(32'h3c214358),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ff907),
	.w1(32'hbb481816),
	.w2(32'hbcd345d3),
	.w3(32'hbc1cac4a),
	.w4(32'hb9da44cb),
	.w5(32'hbc11b512),
	.w6(32'hbabdda3d),
	.w7(32'h3bd9389f),
	.w8(32'hbbc0ed17),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c953a),
	.w1(32'hbc06bbfd),
	.w2(32'hbc2a10c1),
	.w3(32'hbbc7115f),
	.w4(32'h3b489066),
	.w5(32'h3c4c129e),
	.w6(32'h3c06d330),
	.w7(32'h3c75424d),
	.w8(32'h39e90c19),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74cea8),
	.w1(32'hbb38bab2),
	.w2(32'h3c59e55a),
	.w3(32'h3ba0a518),
	.w4(32'h3bc299e9),
	.w5(32'hb9bfa9cb),
	.w6(32'hbc471571),
	.w7(32'hbb39bae0),
	.w8(32'h3bee5800),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc570dc6),
	.w1(32'hbbe9fed6),
	.w2(32'hbbdd2864),
	.w3(32'hbc274b73),
	.w4(32'h3982da60),
	.w5(32'h38b98180),
	.w6(32'hbbbfd46a),
	.w7(32'hbaae5790),
	.w8(32'h3b86b9d8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc98670),
	.w1(32'hbb7729fd),
	.w2(32'hbb9c2ada),
	.w3(32'hbb2a8624),
	.w4(32'hbba56506),
	.w5(32'hbb004dff),
	.w6(32'hbb8757e7),
	.w7(32'h3bf32433),
	.w8(32'h3c0eb8ce),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7abd6e),
	.w1(32'h39e4d8b9),
	.w2(32'hbbee25d8),
	.w3(32'h3c1f3d75),
	.w4(32'h3b1cffd2),
	.w5(32'h3cd1c02e),
	.w6(32'h3b0592c3),
	.w7(32'h3b1c1be1),
	.w8(32'hbba253fe),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee255),
	.w1(32'hbacb9ed8),
	.w2(32'hbc10d6cf),
	.w3(32'h3b896e45),
	.w4(32'hbaeaf738),
	.w5(32'h3c9354c3),
	.w6(32'h3a6cf768),
	.w7(32'h3c7f8846),
	.w8(32'h3c291bed),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b995190),
	.w1(32'h39552ed6),
	.w2(32'h3bcdbcf9),
	.w3(32'h3c637bae),
	.w4(32'h3aef868b),
	.w5(32'h3b96cd33),
	.w6(32'hba9b6d37),
	.w7(32'hb9b75b45),
	.w8(32'h3b5c99ac),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf80c),
	.w1(32'hb9a451d2),
	.w2(32'h3a7892f5),
	.w3(32'hbb01fe30),
	.w4(32'hbbe81dd4),
	.w5(32'hbb000ad7),
	.w6(32'h3b1d513c),
	.w7(32'hbbb664d3),
	.w8(32'hba5c99c1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45d729),
	.w1(32'hbb4aded4),
	.w2(32'hbc06454e),
	.w3(32'hbbab7d3c),
	.w4(32'h3b83d3b2),
	.w5(32'hbba4fdfd),
	.w6(32'hbbef6a64),
	.w7(32'h3c1b4903),
	.w8(32'hbaf26e5d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ce7c1),
	.w1(32'hbbe125f5),
	.w2(32'hbba539b1),
	.w3(32'hbc4c6acc),
	.w4(32'hbc0d704e),
	.w5(32'h3be1ffa5),
	.w6(32'hbb75c38d),
	.w7(32'h3b0160ad),
	.w8(32'h3b92867d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03c05d),
	.w1(32'hbb36a37e),
	.w2(32'h39a3aa2a),
	.w3(32'h3c367f9a),
	.w4(32'hbb3a4484),
	.w5(32'h3b926d71),
	.w6(32'h3a830b4e),
	.w7(32'hb9d7f250),
	.w8(32'h3bc84d46),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63c6b0),
	.w1(32'h3b470023),
	.w2(32'hbb941a9b),
	.w3(32'hbc532c51),
	.w4(32'hbacbdc3d),
	.w5(32'h3c6ad87b),
	.w6(32'h3c06a737),
	.w7(32'h3c675ee4),
	.w8(32'hbc2c3413),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d1f3),
	.w1(32'h3b03b6e0),
	.w2(32'hbbc81f50),
	.w3(32'hba3fcd14),
	.w4(32'h3b8c89b7),
	.w5(32'h3a714bbd),
	.w6(32'h3af5429d),
	.w7(32'h3baf5b2c),
	.w8(32'hbb0ef32c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d1fe2),
	.w1(32'hbc615eab),
	.w2(32'h3a94ca1d),
	.w3(32'h3aade24b),
	.w4(32'hbb2b243d),
	.w5(32'h3b41eb8c),
	.w6(32'hbabc77ef),
	.w7(32'hba443b2f),
	.w8(32'h3ba83270),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb43cb),
	.w1(32'h3b40c3b1),
	.w2(32'hbbee6735),
	.w3(32'h3b6ba110),
	.w4(32'hbb085844),
	.w5(32'hbc042786),
	.w6(32'h39c89025),
	.w7(32'h3bd00492),
	.w8(32'h3bc5db99),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67189),
	.w1(32'h3ab11b8f),
	.w2(32'h3b1b9d5f),
	.w3(32'h3ba8db43),
	.w4(32'h3b7bdc28),
	.w5(32'hba875d52),
	.w6(32'h3be5b19a),
	.w7(32'h3a1d40ca),
	.w8(32'hbb6810e5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe68cf5),
	.w1(32'h3b8e8c30),
	.w2(32'h3949e990),
	.w3(32'hbb898a11),
	.w4(32'h3bd81b9a),
	.w5(32'h3be5469d),
	.w6(32'hbba185b7),
	.w7(32'hbabc582e),
	.w8(32'h3bd1eb79),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3efb2b),
	.w1(32'hba1c5c07),
	.w2(32'h3b82b961),
	.w3(32'hbb3c0009),
	.w4(32'h3b437eb7),
	.w5(32'h3a907f6c),
	.w6(32'hbb115b49),
	.w7(32'hbb95639b),
	.w8(32'hbb90a432),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57699b),
	.w1(32'hbbb4bd61),
	.w2(32'hbb5ef53c),
	.w3(32'hbb03946c),
	.w4(32'h3b9a0ce8),
	.w5(32'hbbed2771),
	.w6(32'h3b61b771),
	.w7(32'h3a8040ca),
	.w8(32'hbb3bc79c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38cc0e),
	.w1(32'h3b1d5a46),
	.w2(32'h3c16dbaf),
	.w3(32'hbc031b6f),
	.w4(32'h3c630cfd),
	.w5(32'h3c9575fd),
	.w6(32'hbbe1564b),
	.w7(32'h3bbfb84d),
	.w8(32'hbafd8f39),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72d13),
	.w1(32'h3b0c7d80),
	.w2(32'hbcb8f348),
	.w3(32'h3b4fb27d),
	.w4(32'hba6d5546),
	.w5(32'hbc9f8ee9),
	.w6(32'hbc26e890),
	.w7(32'h3ba72f6e),
	.w8(32'hbbbf3ca5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72ea91),
	.w1(32'h3b1b9e23),
	.w2(32'hbc502921),
	.w3(32'hbb81621b),
	.w4(32'h3b9031f5),
	.w5(32'h3bdac5c7),
	.w6(32'hbac98b3d),
	.w7(32'h3bbb03ab),
	.w8(32'hbbb30057),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3b7a8),
	.w1(32'hb9925fc8),
	.w2(32'hbc9dd063),
	.w3(32'hbad1761a),
	.w4(32'h3b54c31c),
	.w5(32'hbc80b152),
	.w6(32'hbb6167e2),
	.w7(32'hbad860c0),
	.w8(32'hbc5765bb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4889),
	.w1(32'hbb699841),
	.w2(32'h3a167c38),
	.w3(32'hbb26d9d5),
	.w4(32'hb92bb702),
	.w5(32'hb9afc815),
	.w6(32'hbb8ec140),
	.w7(32'hbb96c275),
	.w8(32'h3bb5687e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58afe9),
	.w1(32'hb8e85a55),
	.w2(32'h39a97759),
	.w3(32'h3bd0cbb4),
	.w4(32'h3b6e4034),
	.w5(32'h3c233e97),
	.w6(32'h3c14a769),
	.w7(32'h3b369ac6),
	.w8(32'h3bc304bd),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1cf0c),
	.w1(32'h3a9ac666),
	.w2(32'hbabb04b0),
	.w3(32'h399efa62),
	.w4(32'h3b038369),
	.w5(32'hbb82f4cf),
	.w6(32'h3a3c8b9c),
	.w7(32'hb9f42a4b),
	.w8(32'hbb5e7b7c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba107e2a),
	.w1(32'h3aba638f),
	.w2(32'h3a48f279),
	.w3(32'hbb813876),
	.w4(32'h3a6699e1),
	.w5(32'hbc22125a),
	.w6(32'hbb16f6c7),
	.w7(32'hbbbc5332),
	.w8(32'h3b93bde1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcca131c),
	.w1(32'hbbf9d255),
	.w2(32'hbc834ec5),
	.w3(32'hbcaa95c7),
	.w4(32'hbb432c20),
	.w5(32'h3c780ce7),
	.w6(32'hbc11ab9e),
	.w7(32'h3c168e7c),
	.w8(32'hbb1626fc),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07a9e),
	.w1(32'h3b2f1f23),
	.w2(32'hbb8d9063),
	.w3(32'h3b898b61),
	.w4(32'h3b475f9b),
	.w5(32'h38cbbe11),
	.w6(32'hba06d715),
	.w7(32'hbb82cdcd),
	.w8(32'hbb7c2523),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c1def),
	.w1(32'h3aa429aa),
	.w2(32'h3bc1b603),
	.w3(32'hbbf29b14),
	.w4(32'hbade904c),
	.w5(32'hbaf766f1),
	.w6(32'hbb1b8d8d),
	.w7(32'hba909dd4),
	.w8(32'h3a375da4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba685593),
	.w1(32'hbabc2180),
	.w2(32'hbb14cf89),
	.w3(32'hbb463bc1),
	.w4(32'hb8c7106f),
	.w5(32'h3be21a7c),
	.w6(32'hbbfd3ebf),
	.w7(32'hbb5bb887),
	.w8(32'hbb5aa003),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf61b90),
	.w1(32'hbbe0800b),
	.w2(32'hbbfbd099),
	.w3(32'hb9caae40),
	.w4(32'hbb8d3984),
	.w5(32'h3c753b6f),
	.w6(32'hbb714d9e),
	.w7(32'h3b7d7764),
	.w8(32'hbb685f72),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb5043),
	.w1(32'hbb8f5d46),
	.w2(32'hbc44db7b),
	.w3(32'h3ae4978c),
	.w4(32'hbbbd17e7),
	.w5(32'hb9111d3a),
	.w6(32'hbbb7b72b),
	.w7(32'hbbaf2f47),
	.w8(32'hbba93181),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4298ab),
	.w1(32'h3ae7bb54),
	.w2(32'h3b32708b),
	.w3(32'h3b7ff582),
	.w4(32'hbb4c5393),
	.w5(32'hbbfecdae),
	.w6(32'hbb9aae4f),
	.w7(32'hbbdd27d3),
	.w8(32'h3a203255),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65dab8),
	.w1(32'hbc560b8b),
	.w2(32'hbc89229d),
	.w3(32'hbc760af1),
	.w4(32'hba8769be),
	.w5(32'hbb8d8f7b),
	.w6(32'hbc25bf75),
	.w7(32'hbb8bcec7),
	.w8(32'hbb679c3d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670861),
	.w1(32'h3aa8878e),
	.w2(32'hbbb952aa),
	.w3(32'h3b8412e5),
	.w4(32'hbba79e7f),
	.w5(32'hbbab6d55),
	.w6(32'h39c5b29b),
	.w7(32'hb7244c9c),
	.w8(32'hb907ee73),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e6b8e),
	.w1(32'hbbea24e3),
	.w2(32'hbac7092e),
	.w3(32'hbc21be87),
	.w4(32'h3bb9c935),
	.w5(32'h3cf8037f),
	.w6(32'hbc7e6d23),
	.w7(32'h3c3c051a),
	.w8(32'h3c98d799),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule