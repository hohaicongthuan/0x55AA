module layer_8_featuremap_205(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb907ebb),
	.w1(32'hbc8469f3),
	.w2(32'hbc94a299),
	.w3(32'h3ba5077f),
	.w4(32'h3aa3d215),
	.w5(32'hbb2b4bf0),
	.w6(32'hbac76cb6),
	.w7(32'hbc224c91),
	.w8(32'hbc6e8d6e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90b267),
	.w1(32'hbb341503),
	.w2(32'h3bb3ad19),
	.w3(32'hbc44d38a),
	.w4(32'hbbd00303),
	.w5(32'h3a4821ad),
	.w6(32'h3b0ad48d),
	.w7(32'h3c234b45),
	.w8(32'h3be3f4dc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec18c5),
	.w1(32'hbaebc899),
	.w2(32'h3b8e222e),
	.w3(32'h3bb55757),
	.w4(32'hb91a572b),
	.w5(32'h3baa5467),
	.w6(32'h3b02402a),
	.w7(32'h3b85d242),
	.w8(32'h3b1b8ad9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c218684),
	.w1(32'hbae8d655),
	.w2(32'h3b504fa6),
	.w3(32'hba5c47cd),
	.w4(32'hba5fb034),
	.w5(32'h3ae5c931),
	.w6(32'h3baf33a0),
	.w7(32'hbbcd5dcf),
	.w8(32'hbc4cc16e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3be5c),
	.w1(32'hbabd06a8),
	.w2(32'hbb5544a5),
	.w3(32'h3b33bc4e),
	.w4(32'hb9eb610f),
	.w5(32'h3bb7e607),
	.w6(32'hbb14e767),
	.w7(32'hbb87d31a),
	.w8(32'hbc36dbe3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc290410),
	.w1(32'hba4cf3a6),
	.w2(32'h3b84f60a),
	.w3(32'hba401396),
	.w4(32'h3ba12e42),
	.w5(32'h3c6d8a50),
	.w6(32'h3bd65548),
	.w7(32'hbae03cb2),
	.w8(32'h3b06460d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94406d),
	.w1(32'hbae5a398),
	.w2(32'hbbec13e2),
	.w3(32'h3b722db8),
	.w4(32'hbb817fbc),
	.w5(32'hbbd4f435),
	.w6(32'hbb8eb1ce),
	.w7(32'hbc222f2c),
	.w8(32'hbbe5f288),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0811f0),
	.w1(32'hbb694f0e),
	.w2(32'hbba2f4f4),
	.w3(32'hbbcbc605),
	.w4(32'hbc102fc9),
	.w5(32'hbc34ce67),
	.w6(32'hbb2c52df),
	.w7(32'h3a44e572),
	.w8(32'hbb80157e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e799),
	.w1(32'h3b61b577),
	.w2(32'hbbcee808),
	.w3(32'h3b501c13),
	.w4(32'h3c2448b8),
	.w5(32'h3c807861),
	.w6(32'hbbdaa381),
	.w7(32'hbc936fab),
	.w8(32'hbcffc14c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdfbc62),
	.w1(32'hbc0314f9),
	.w2(32'hbcb8b660),
	.w3(32'hbb185471),
	.w4(32'hbbf328e7),
	.w5(32'hbc3708ef),
	.w6(32'hbc38864d),
	.w7(32'hbc868022),
	.w8(32'hbb9e5bdb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc765194),
	.w1(32'hbc32cfd9),
	.w2(32'h3c1b5ba6),
	.w3(32'hbc29e884),
	.w4(32'hbc321ef4),
	.w5(32'h3adea871),
	.w6(32'hbb9c302f),
	.w7(32'h3c4065d3),
	.w8(32'h3b612416),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e5e54),
	.w1(32'hbb174500),
	.w2(32'hbbd732b7),
	.w3(32'h3c0de39d),
	.w4(32'hbab9a293),
	.w5(32'hbb98ad4e),
	.w6(32'hbae4eca0),
	.w7(32'h39f3f9c1),
	.w8(32'h3c410e12),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badadb2),
	.w1(32'hbc7e4ec8),
	.w2(32'hbca90f0a),
	.w3(32'hbb6d3c78),
	.w4(32'hbc1940dd),
	.w5(32'hbc12a5cc),
	.w6(32'hbbc58425),
	.w7(32'hbb897358),
	.w8(32'hbc1e2ac0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5ca34),
	.w1(32'hbb8d494d),
	.w2(32'hbc2ad18e),
	.w3(32'hbbf56a11),
	.w4(32'hbba4ca19),
	.w5(32'hbc19534d),
	.w6(32'hbbfab481),
	.w7(32'hbb9d1ecc),
	.w8(32'hbbe7cf4f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb58570),
	.w1(32'h398bf885),
	.w2(32'hbc2d5ec1),
	.w3(32'hbc20254e),
	.w4(32'h38ff32d9),
	.w5(32'hbb9b6bef),
	.w6(32'hbb6b23c8),
	.w7(32'hbc4cfdd7),
	.w8(32'hbc404d16),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ef1db),
	.w1(32'hbb6e6b51),
	.w2(32'h3a9ca8ca),
	.w3(32'hbc1ca908),
	.w4(32'hbb779e87),
	.w5(32'hbb803e5a),
	.w6(32'h3ac0e696),
	.w7(32'hbb99e76d),
	.w8(32'hbbf2f69d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b5430),
	.w1(32'hbc277b12),
	.w2(32'hbb3fa432),
	.w3(32'hbbb0b2e1),
	.w4(32'hbbae6b19),
	.w5(32'hbbbb7640),
	.w6(32'h39315ea2),
	.w7(32'h3b03a091),
	.w8(32'h3b3c2035),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18e7f7),
	.w1(32'hbbeb0e08),
	.w2(32'hbc338d81),
	.w3(32'h3b5c26dc),
	.w4(32'hbc29a897),
	.w5(32'hbc436331),
	.w6(32'hbb9cb7ad),
	.w7(32'hbbc7bdd9),
	.w8(32'hbc02785e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd85e16),
	.w1(32'hbc8ce394),
	.w2(32'hbcea0907),
	.w3(32'hbc1bcf2a),
	.w4(32'hbc4d42b2),
	.w5(32'hbcc1ac06),
	.w6(32'h3b0e8351),
	.w7(32'hbc0683d3),
	.w8(32'hbbc67ee6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96e344),
	.w1(32'h3bd667ea),
	.w2(32'h3b0c5e26),
	.w3(32'hbca3c7c5),
	.w4(32'h3c1ccdd8),
	.w5(32'h3c198b5f),
	.w6(32'h3baa47ed),
	.w7(32'hbaf8f924),
	.w8(32'hbb932f8b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb860fa7),
	.w1(32'h3c34a3ff),
	.w2(32'h3c80ee4c),
	.w3(32'h3b39c3f3),
	.w4(32'h39e56363),
	.w5(32'h3c00aa87),
	.w6(32'h3b4bed9a),
	.w7(32'h3b508ba7),
	.w8(32'h3bdb525e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb801),
	.w1(32'hba6c62ef),
	.w2(32'h39951e6e),
	.w3(32'hbb3ab9c7),
	.w4(32'hbb4ba068),
	.w5(32'hbb51c040),
	.w6(32'h3bc393fe),
	.w7(32'h3aa3663b),
	.w8(32'h3a5a9a81),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f2e95),
	.w1(32'hbb52d113),
	.w2(32'hbb56e4be),
	.w3(32'hbacb6bb4),
	.w4(32'hbbd26c6d),
	.w5(32'hbbf972e9),
	.w6(32'hbc27d116),
	.w7(32'hbc47215c),
	.w8(32'hbc151134),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5debfc),
	.w1(32'h3bdc4e29),
	.w2(32'h3b6330ce),
	.w3(32'hbb8f4086),
	.w4(32'hbb8654eb),
	.w5(32'hbabbebb8),
	.w6(32'h3b740231),
	.w7(32'h3b68352e),
	.w8(32'hb8190733),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62e304),
	.w1(32'hbae74b82),
	.w2(32'h3c1040e8),
	.w3(32'h3b77ea36),
	.w4(32'hba459ab3),
	.w5(32'h3c76e70e),
	.w6(32'h3b841d7d),
	.w7(32'h3bb91c86),
	.w8(32'h3b6a60c7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb52668),
	.w1(32'hbbc2cbd3),
	.w2(32'h3bb7505d),
	.w3(32'h3c166272),
	.w4(32'h3b3cbcd4),
	.w5(32'h3b3a8b00),
	.w6(32'hba9f49df),
	.w7(32'hbab63c06),
	.w8(32'h3a61cf42),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3533c),
	.w1(32'h3b14fdc2),
	.w2(32'h3c0979a2),
	.w3(32'hbbf91781),
	.w4(32'h3ba249f1),
	.w5(32'h3c662fe1),
	.w6(32'h3bdb9677),
	.w7(32'h3c109834),
	.w8(32'h3b4ca5ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03b3d5),
	.w1(32'hbb1b5fd4),
	.w2(32'hbc11dafe),
	.w3(32'h3c496a04),
	.w4(32'hbb9ff247),
	.w5(32'hb9b9e4a4),
	.w6(32'hbc1b3774),
	.w7(32'hbc88d1b7),
	.w8(32'hbbfceeaa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc939570),
	.w1(32'hbb21ad35),
	.w2(32'h3c93d8c9),
	.w3(32'hbc8c0c62),
	.w4(32'hbb97f716),
	.w5(32'h3b774480),
	.w6(32'hbbe5ee05),
	.w7(32'h3c539c72),
	.w8(32'h3b61ab12),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a32f7),
	.w1(32'h3b18b067),
	.w2(32'h3ba6add0),
	.w3(32'h3bdade28),
	.w4(32'h3c77b62b),
	.w5(32'h3cb0d061),
	.w6(32'hbaf8562b),
	.w7(32'h3b240f0d),
	.w8(32'h3c4bc372),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c225f21),
	.w1(32'hbc5529dd),
	.w2(32'hbc9428ad),
	.w3(32'h3cbe5f33),
	.w4(32'hbc2cf622),
	.w5(32'hbc6a6c41),
	.w6(32'hbc2acc3b),
	.w7(32'hbbae9cf8),
	.w8(32'h3a25ceb1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1fa66),
	.w1(32'hbbae2962),
	.w2(32'h3c0528b3),
	.w3(32'hbc3b5803),
	.w4(32'hbb50d3a6),
	.w5(32'hbbb754fb),
	.w6(32'h3b426eb1),
	.w7(32'h3c708096),
	.w8(32'h3bfe612c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e9fce),
	.w1(32'hbb6be720),
	.w2(32'hb9e09572),
	.w3(32'h3a9ed471),
	.w4(32'hbb0edcab),
	.w5(32'hba661b2c),
	.w6(32'hbbbd676e),
	.w7(32'hbbe25331),
	.w8(32'hbc3c56db),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8711b),
	.w1(32'h3a089b41),
	.w2(32'hbbc2c603),
	.w3(32'h3a431c7d),
	.w4(32'h3b6588f1),
	.w5(32'hb9f23c92),
	.w6(32'h3b926ee9),
	.w7(32'h3b156222),
	.w8(32'h3b8f8e3f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4460b5),
	.w1(32'h3a951ce1),
	.w2(32'hbc29e432),
	.w3(32'hb90386d5),
	.w4(32'h3ab0366d),
	.w5(32'h3a3531ea),
	.w6(32'h3b913eab),
	.w7(32'h3ab4e443),
	.w8(32'h3a41c552),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcacbce0),
	.w1(32'h3b9aa412),
	.w2(32'h3bd3fbe5),
	.w3(32'hbacce9e3),
	.w4(32'h3ba497e5),
	.w5(32'h3ae5d8ec),
	.w6(32'h3c0402cc),
	.w7(32'h3b850797),
	.w8(32'h3acaae2b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1baa5),
	.w1(32'h3c98a975),
	.w2(32'h3cc66850),
	.w3(32'hb982122b),
	.w4(32'h3c5c6847),
	.w5(32'h3cc17a92),
	.w6(32'h3c7a9ee0),
	.w7(32'h3c90296a),
	.w8(32'h3c0c1a99),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f43ac),
	.w1(32'h3ae03060),
	.w2(32'hbbf00e5e),
	.w3(32'h3cb55658),
	.w4(32'h3ac0306e),
	.w5(32'h3aa35b0a),
	.w6(32'hbb470e4d),
	.w7(32'hbc37debb),
	.w8(32'hbc865e71),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc893bf9),
	.w1(32'h3c0369c8),
	.w2(32'h3c8dc108),
	.w3(32'hbbfe05df),
	.w4(32'hba8eb2a5),
	.w5(32'h3bcaa147),
	.w6(32'h3c122969),
	.w7(32'h3c25246d),
	.w8(32'h3c75fd6c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b30b0),
	.w1(32'hbbd07163),
	.w2(32'hbb9ee0f1),
	.w3(32'h3b6d5cb2),
	.w4(32'hbb88f448),
	.w5(32'hbc063bed),
	.w6(32'hbb860c89),
	.w7(32'hbbd57c11),
	.w8(32'hbb8ac2c2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2baecb),
	.w1(32'hbb86985d),
	.w2(32'hbc23cb27),
	.w3(32'hbb5439ea),
	.w4(32'hbb9cbc2a),
	.w5(32'hbc477c7f),
	.w6(32'hbb4d74f8),
	.w7(32'hbbe668d8),
	.w8(32'hbbbad4d3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2fbfc),
	.w1(32'hbc7a7009),
	.w2(32'hbd0ab1c8),
	.w3(32'hbb7ec51d),
	.w4(32'hbc3f89f7),
	.w5(32'hbcee9774),
	.w6(32'hbb97c222),
	.w7(32'hbc98414d),
	.w8(32'h3bec51c8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4729d6),
	.w1(32'h3c449c4a),
	.w2(32'h3ce7eabd),
	.w3(32'hbc139e1b),
	.w4(32'h3bd17b83),
	.w5(32'h3c2841e9),
	.w6(32'h3b8c6723),
	.w7(32'h3c8c7b69),
	.w8(32'h3c1f6635),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0aa7d),
	.w1(32'hbc302a9d),
	.w2(32'hbb0274b0),
	.w3(32'h3c4e60fd),
	.w4(32'hbbbb2bfe),
	.w5(32'hbb8c3c1a),
	.w6(32'hbbb3c8aa),
	.w7(32'hba78dd25),
	.w8(32'h3b64c87c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba980bce),
	.w1(32'h3b3b86c4),
	.w2(32'hbbe18e0c),
	.w3(32'hbb84c0fd),
	.w4(32'hbb10f47a),
	.w5(32'hbb4274c9),
	.w6(32'h3be011c2),
	.w7(32'h3ba5c590),
	.w8(32'h39c2f415),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc39b2f),
	.w1(32'h398d0c34),
	.w2(32'hbb448a8a),
	.w3(32'hbc32c48e),
	.w4(32'h3aad0b0c),
	.w5(32'h373af8ba),
	.w6(32'h3bba9ede),
	.w7(32'h3b410425),
	.w8(32'h3aea5a69),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5e2c),
	.w1(32'hbc7dd6cc),
	.w2(32'hbbeb5c96),
	.w3(32'h39e612f5),
	.w4(32'hbcc0461d),
	.w5(32'hbc9d927f),
	.w6(32'hbc101070),
	.w7(32'h3b0f803a),
	.w8(32'h3c7c44e2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae10341),
	.w1(32'hb8cd5829),
	.w2(32'h3b221e0a),
	.w3(32'hbc070807),
	.w4(32'h3b74e943),
	.w5(32'h3c039edb),
	.w6(32'hbb7e59fe),
	.w7(32'h3b1c74b0),
	.w8(32'h3bdefb55),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9f395),
	.w1(32'h3b250adb),
	.w2(32'h3bcaca35),
	.w3(32'h3bf420b8),
	.w4(32'h3c140146),
	.w5(32'h3b569eda),
	.w6(32'h3ac33251),
	.w7(32'h3b52147d),
	.w8(32'h3c005f08),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36646),
	.w1(32'hbbd8ae35),
	.w2(32'hbc1f0a03),
	.w3(32'h3aedc393),
	.w4(32'hbbb6ba95),
	.w5(32'hbc4ca1a4),
	.w6(32'hbb9373ae),
	.w7(32'hbae1cbe0),
	.w8(32'hbbc342d8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc185c54),
	.w1(32'hba95fae9),
	.w2(32'hbc17d584),
	.w3(32'hbc3d2def),
	.w4(32'hba4a3781),
	.w5(32'hbc81b1e0),
	.w6(32'hbaab12ca),
	.w7(32'hbc0a64fe),
	.w8(32'hb9a26547),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96c128),
	.w1(32'hbcc7b706),
	.w2(32'hbceb6d9d),
	.w3(32'hbaf8adfe),
	.w4(32'hbc90ad72),
	.w5(32'hbcc6f136),
	.w6(32'hbc2e0dfc),
	.w7(32'hbc8b51cf),
	.w8(32'hbc0cac7c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8754d),
	.w1(32'h3b0ae056),
	.w2(32'h3a5d068c),
	.w3(32'hbc2a3e19),
	.w4(32'hbb4e8d75),
	.w5(32'hb7a3697a),
	.w6(32'h3b3e9b4c),
	.w7(32'h3b88b22a),
	.w8(32'hbb373809),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadd41f),
	.w1(32'h3c32a515),
	.w2(32'h3b8396ec),
	.w3(32'hbb310df7),
	.w4(32'h3c098daa),
	.w5(32'hbb853bdc),
	.w6(32'h3a58705d),
	.w7(32'hbb143583),
	.w8(32'h398ff24f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dbb53),
	.w1(32'h3a5fdc10),
	.w2(32'hb9b7c068),
	.w3(32'h3bce6973),
	.w4(32'h3beb0108),
	.w5(32'h3bb1b3cc),
	.w6(32'hbb89e81d),
	.w7(32'hbbab779d),
	.w8(32'hbaa7b1de),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919191),
	.w1(32'h3a9b4c2f),
	.w2(32'hbbff481c),
	.w3(32'hbbe3ee36),
	.w4(32'hbb8f3d26),
	.w5(32'hbc1e45e7),
	.w6(32'hbc0ded5a),
	.w7(32'hbc067560),
	.w8(32'hbb3d95bc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46fa5b),
	.w1(32'h3bf51f34),
	.w2(32'h3be785b0),
	.w3(32'h3b1b9974),
	.w4(32'hbb5ead9b),
	.w5(32'hbbb7b2dc),
	.w6(32'hbac29761),
	.w7(32'h3c6600f1),
	.w8(32'h3c42339f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e3acb),
	.w1(32'h3c7448c8),
	.w2(32'h3cdd0d09),
	.w3(32'h3bc70f90),
	.w4(32'h3c4035ab),
	.w5(32'h3cd3caac),
	.w6(32'h3be6abc6),
	.w7(32'h3c6dd55c),
	.w8(32'h3c56a8c1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d5f66),
	.w1(32'hbb2f8dfa),
	.w2(32'hbb3428db),
	.w3(32'h3c1bce28),
	.w4(32'hbbd2a703),
	.w5(32'hbc062650),
	.w6(32'hbb4a4b75),
	.w7(32'hb9c15da2),
	.w8(32'h3b1b423e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3f1f7),
	.w1(32'h3b41b697),
	.w2(32'h3a8bcda5),
	.w3(32'hbba237e5),
	.w4(32'hbac40a2a),
	.w5(32'hbb3775ef),
	.w6(32'h3a4ebb4d),
	.w7(32'h3a9e1872),
	.w8(32'hba9a06d0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b089be1),
	.w1(32'hbb22562e),
	.w2(32'h3c6f042f),
	.w3(32'h39b6f99b),
	.w4(32'h3b405947),
	.w5(32'h3ca3fff4),
	.w6(32'hbb14779d),
	.w7(32'h3ba5c2a3),
	.w8(32'h3c56a700),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cdf57),
	.w1(32'h3c3a9826),
	.w2(32'h3ccab40e),
	.w3(32'h3c81d573),
	.w4(32'h3c72fa4c),
	.w5(32'h3d19f672),
	.w6(32'h3c0dd5dd),
	.w7(32'h3c0bbf15),
	.w8(32'hbb2f4b94),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd99f52),
	.w1(32'h3bbdb791),
	.w2(32'h3c612dfd),
	.w3(32'h3cdfc843),
	.w4(32'h3c82d4e2),
	.w5(32'h3ca720ef),
	.w6(32'hbae751b5),
	.w7(32'h3b8ec7e6),
	.w8(32'hba828c0d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7127e),
	.w1(32'hbb94baad),
	.w2(32'hbc038f9d),
	.w3(32'h3c6e266d),
	.w4(32'hbc02f51e),
	.w5(32'hbc30bf93),
	.w6(32'hbb5dbe92),
	.w7(32'hbb81f9f1),
	.w8(32'hbb41930f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd05fc),
	.w1(32'hbb93f31c),
	.w2(32'h3b45aed8),
	.w3(32'hbc19d763),
	.w4(32'hbc65cdc8),
	.w5(32'hbc27b8b5),
	.w6(32'hbb05ee63),
	.w7(32'h3c0e13b1),
	.w8(32'h3c661b81),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47286a),
	.w1(32'hbb90a25f),
	.w2(32'hbc0e4139),
	.w3(32'hbb8a061f),
	.w4(32'hbb1b11eb),
	.w5(32'hbc2158b9),
	.w6(32'h3a91339d),
	.w7(32'hbbc8f93a),
	.w8(32'h3a71c90d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc843e),
	.w1(32'h3abb8a42),
	.w2(32'h3b05d3a2),
	.w3(32'h3a7df250),
	.w4(32'hbaaa62b2),
	.w5(32'h3c4a1ea2),
	.w6(32'h3bbf1177),
	.w7(32'hbb5bcbcf),
	.w8(32'hbb9092b8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bcbdb),
	.w1(32'hbb023e3d),
	.w2(32'h3c1e1661),
	.w3(32'h3c2b29c8),
	.w4(32'hbb83976b),
	.w5(32'hbb474337),
	.w6(32'h3a3beffa),
	.w7(32'h389b0129),
	.w8(32'h3c0c48ac),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8c24b),
	.w1(32'h3aa9500b),
	.w2(32'hbc20663b),
	.w3(32'h3afc5aa3),
	.w4(32'h3b796fa6),
	.w5(32'hb9526576),
	.w6(32'h3abdf87f),
	.w7(32'h3b26f0a8),
	.w8(32'h3b99622a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27e744),
	.w1(32'h3a52cc87),
	.w2(32'h3bbbb212),
	.w3(32'hbb2c022c),
	.w4(32'h3b34b2a2),
	.w5(32'h3c34af8f),
	.w6(32'hbb65b522),
	.w7(32'hbab39399),
	.w8(32'h3b22aa92),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be71f34),
	.w1(32'hbd05db0d),
	.w2(32'hbd39a96d),
	.w3(32'h3c1d9da1),
	.w4(32'hbce3e599),
	.w5(32'hbd0b6a13),
	.w6(32'hbcc15ff5),
	.w7(32'hbd1099c0),
	.w8(32'hbc93f20e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd19973d),
	.w1(32'h3a0c3d24),
	.w2(32'h3aec78cb),
	.w3(32'hbd070bd3),
	.w4(32'hba43a126),
	.w5(32'hbb47cd87),
	.w6(32'h3c1292d7),
	.w7(32'h3c108259),
	.w8(32'h3c341397),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c867),
	.w1(32'h3b15df51),
	.w2(32'h3c62eda1),
	.w3(32'hbb383071),
	.w4(32'h3bbb13c1),
	.w5(32'h3c387732),
	.w6(32'h3c0afa31),
	.w7(32'h3c7e9c66),
	.w8(32'h3c5c4fe2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2df33b),
	.w1(32'hbb16ff99),
	.w2(32'h3c10d4e7),
	.w3(32'h3aa96119),
	.w4(32'hbaa5d572),
	.w5(32'h3c0aef7b),
	.w6(32'h3afb8e70),
	.w7(32'h3baf8a9b),
	.w8(32'hbb2fe65d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e8dfe),
	.w1(32'hbc12411f),
	.w2(32'hbc372de0),
	.w3(32'hbb400dc7),
	.w4(32'hbba56a64),
	.w5(32'hbb3c36e5),
	.w6(32'h3ba4e201),
	.w7(32'hbb0d4836),
	.w8(32'h3c3b934c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b5261),
	.w1(32'h3b64a442),
	.w2(32'h3bd3f660),
	.w3(32'h3c151a9f),
	.w4(32'h3a8d3eec),
	.w5(32'h3bcee1c1),
	.w6(32'h39f28c10),
	.w7(32'h39f6b25d),
	.w8(32'hbb8f5056),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb673654),
	.w1(32'h3b3d7b27),
	.w2(32'h3c085ee1),
	.w3(32'h3b149a69),
	.w4(32'h3a71f454),
	.w5(32'hba66c63c),
	.w6(32'h3b77e5c9),
	.w7(32'h3c2e9d42),
	.w8(32'h3bb24c8f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392219c8),
	.w1(32'h3c7a5059),
	.w2(32'h3c93472e),
	.w3(32'h3b1c18f4),
	.w4(32'h3c22a43e),
	.w5(32'h3b6bb01c),
	.w6(32'h3c16bdfb),
	.w7(32'h3c6b8259),
	.w8(32'h3c1440ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4aafe3),
	.w1(32'hbcef0dfd),
	.w2(32'hbd2ff72c),
	.w3(32'h3c486194),
	.w4(32'hbcb274c8),
	.w5(32'hbce17bb2),
	.w6(32'hbc7baa08),
	.w7(32'hbcd147df),
	.w8(32'hbcb11478),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced0c45),
	.w1(32'hbc7f001a),
	.w2(32'hbc43f488),
	.w3(32'hbc8862db),
	.w4(32'hbbe5276d),
	.w5(32'hbbd226de),
	.w6(32'hbc4dde51),
	.w7(32'hbc120d96),
	.w8(32'hbb1889c5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1053),
	.w1(32'h3b1acf84),
	.w2(32'h3c1ae30c),
	.w3(32'hbb8dd6b1),
	.w4(32'h3ba37c99),
	.w5(32'h3bc877de),
	.w6(32'hba173394),
	.w7(32'h382b2fea),
	.w8(32'h3b59b434),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78f22f),
	.w1(32'h3bcf1d60),
	.w2(32'h3aa0e643),
	.w3(32'hbae663a7),
	.w4(32'h3bfdcd7d),
	.w5(32'h3bc390ea),
	.w6(32'h3c0edf47),
	.w7(32'h3bb23f67),
	.w8(32'h3b2d76b4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803295),
	.w1(32'hbab7a2dc),
	.w2(32'hbb333e63),
	.w3(32'hbaa55bba),
	.w4(32'hbb8c2c1c),
	.w5(32'h3b65a4b0),
	.w6(32'h3a15a50c),
	.w7(32'h3a9c8e83),
	.w8(32'hbb101a49),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc77ac),
	.w1(32'h3c0b932b),
	.w2(32'hb9afadad),
	.w3(32'hbc2a78e2),
	.w4(32'h3b4a09a3),
	.w5(32'h3af56fa1),
	.w6(32'h3c1e72a0),
	.w7(32'h3b8de369),
	.w8(32'h3c051485),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b925289),
	.w1(32'hbb1a5454),
	.w2(32'hbc55636a),
	.w3(32'hbb22c001),
	.w4(32'hbc933464),
	.w5(32'hbbbb2ec8),
	.w6(32'hbc6ea455),
	.w7(32'hbc53a231),
	.w8(32'hbbb3d3fe),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd6959),
	.w1(32'h3ab47e25),
	.w2(32'h3c5d1464),
	.w3(32'hbcbe1bad),
	.w4(32'h3bfb8bf5),
	.w5(32'h3c251cba),
	.w6(32'h3ba3cd10),
	.w7(32'h3b8f17c3),
	.w8(32'hbbc88acc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c85a0),
	.w1(32'hbcd0ce5a),
	.w2(32'hbd0b6e49),
	.w3(32'hbb426509),
	.w4(32'hbca1bc27),
	.w5(32'hbcdd57c0),
	.w6(32'hbca8d728),
	.w7(32'hbcc8b4d5),
	.w8(32'hbc9fe137),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0ea63),
	.w1(32'hbb4cf361),
	.w2(32'h3cdc8938),
	.w3(32'hbcd0e569),
	.w4(32'hbc23cb36),
	.w5(32'h3c729cd0),
	.w6(32'h3bd80d08),
	.w7(32'h3ca81e48),
	.w8(32'h3c064362),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0625e),
	.w1(32'hbcc72948),
	.w2(32'hbd0d954f),
	.w3(32'h3c90ef7f),
	.w4(32'hbc8a2f3e),
	.w5(32'hbcbd9864),
	.w6(32'hbc6a132f),
	.w7(32'hbc9a4f0c),
	.w8(32'hbc80990a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd001319),
	.w1(32'hbc099a3c),
	.w2(32'h3b394149),
	.w3(32'hbcb9a229),
	.w4(32'h3aa5596d),
	.w5(32'h3c135687),
	.w6(32'hbb90f52f),
	.w7(32'h3a0cef87),
	.w8(32'h3c0c96cd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0966c3),
	.w1(32'h3c05d40f),
	.w2(32'h3c5e9784),
	.w3(32'h3c1e32ea),
	.w4(32'h3c45ad80),
	.w5(32'h3bc55d6c),
	.w6(32'h399265fa),
	.w7(32'h3c3aa983),
	.w8(32'h3c0c11f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf31c23),
	.w1(32'h3b8650f1),
	.w2(32'hbadf2247),
	.w3(32'hbb85ab70),
	.w4(32'h3b48580c),
	.w5(32'hbc0d741a),
	.w6(32'h3af09765),
	.w7(32'h3b5eb08e),
	.w8(32'h3b525f0f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af61eb3),
	.w1(32'h3a773318),
	.w2(32'h3a6d6138),
	.w3(32'hbbb661c8),
	.w4(32'h3aae28d6),
	.w5(32'h3b5ba6d5),
	.w6(32'h3b93d158),
	.w7(32'h3be2d7a1),
	.w8(32'h3ba410f9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac1d05),
	.w1(32'hbc2de57b),
	.w2(32'hb9ed559b),
	.w3(32'h3b9e2381),
	.w4(32'hbc659ece),
	.w5(32'hbbe77536),
	.w6(32'hbbb020d5),
	.w7(32'h3b89dce4),
	.w8(32'h3beb34bb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc368d3),
	.w1(32'h3b565ebd),
	.w2(32'h3c42137b),
	.w3(32'h38f5cc3a),
	.w4(32'h3c076cc6),
	.w5(32'h3c3f8b0f),
	.w6(32'h3bcaec5a),
	.w7(32'h3c4a9000),
	.w8(32'h3bd46d30),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4e16f),
	.w1(32'h3bed1490),
	.w2(32'h3b0e31d2),
	.w3(32'h3bb90678),
	.w4(32'h3c05db64),
	.w5(32'hbb31ed4d),
	.w6(32'h3be0eb43),
	.w7(32'h3b39ef66),
	.w8(32'h3a9c7daf),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ccc21),
	.w1(32'hba55a22c),
	.w2(32'h3b53b8dd),
	.w3(32'hb9d1215e),
	.w4(32'hbc1da74c),
	.w5(32'hbba16c42),
	.w6(32'h3a9397e1),
	.w7(32'hbabbcf33),
	.w8(32'hba7027a1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba947b6),
	.w1(32'h3bf76865),
	.w2(32'h3c38a41b),
	.w3(32'hba6396fe),
	.w4(32'h3b7608e8),
	.w5(32'h3b4e16cb),
	.w6(32'h3b846e97),
	.w7(32'h3a3d9641),
	.w8(32'h3bae16df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bbe7a),
	.w1(32'h3c1d1e5d),
	.w2(32'h3c33d820),
	.w3(32'h3b8c3600),
	.w4(32'h3bb7558d),
	.w5(32'hb9954e54),
	.w6(32'h3aa34b68),
	.w7(32'h3c323e03),
	.w8(32'h3c73a122),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08fad9),
	.w1(32'hbc20de25),
	.w2(32'h3b9405d4),
	.w3(32'h3b67a35a),
	.w4(32'hbad01cd1),
	.w5(32'hbc3a36a2),
	.w6(32'hbc4da709),
	.w7(32'h37266030),
	.w8(32'hb9bcd4bd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62fb891),
	.w1(32'hbc4679b2),
	.w2(32'hbba1b3b2),
	.w3(32'hbbb875d4),
	.w4(32'hba491dd4),
	.w5(32'hbbb17ce8),
	.w6(32'hbc25349d),
	.w7(32'hbb2d24d6),
	.w8(32'h3b3dcfda),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedd7c9),
	.w1(32'h3ba44adb),
	.w2(32'hbc883a08),
	.w3(32'hbb902661),
	.w4(32'h3c300490),
	.w5(32'hbaa4a620),
	.w6(32'h3bdbf2a4),
	.w7(32'hb9a2efa1),
	.w8(32'h3ab2ed09),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25cc14),
	.w1(32'hbad6e4bd),
	.w2(32'hbb934fcd),
	.w3(32'hbc1e843b),
	.w4(32'hbbd0f86f),
	.w5(32'hb78a5fe6),
	.w6(32'h3a9e89a8),
	.w7(32'h3aceab01),
	.w8(32'h3bd0a113),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe89ea3),
	.w1(32'h3a819486),
	.w2(32'h3b077b01),
	.w3(32'hbc12c4b7),
	.w4(32'h3b7b61de),
	.w5(32'h3c0a4175),
	.w6(32'hbaa925dc),
	.w7(32'h3c54d862),
	.w8(32'h3c5bf081),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c157409),
	.w1(32'h3c013fc2),
	.w2(32'h3c3847ac),
	.w3(32'h3c3096f7),
	.w4(32'h3bff6d61),
	.w5(32'h3c78af18),
	.w6(32'h3c13f481),
	.w7(32'h3c2e5a1e),
	.w8(32'h3c82a3d7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c171e8c),
	.w1(32'h3aa967cf),
	.w2(32'h3ab8a0f1),
	.w3(32'h3c02ed92),
	.w4(32'hbaab32f0),
	.w5(32'hbb0501dd),
	.w6(32'h3bccd867),
	.w7(32'h3c01b6b8),
	.w8(32'h3c0d1177),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b603b64),
	.w1(32'hbc85b6a6),
	.w2(32'hbcc627a9),
	.w3(32'h3a117490),
	.w4(32'hbc06c427),
	.w5(32'hbc53ea22),
	.w6(32'hbb2a0a90),
	.w7(32'hbc4515bf),
	.w8(32'hbbf425d4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc796548),
	.w1(32'h3c45b554),
	.w2(32'h3c92914f),
	.w3(32'hbb968b5f),
	.w4(32'h3bdbec91),
	.w5(32'h3ca469e3),
	.w6(32'h3b8133b9),
	.w7(32'h3c0d7310),
	.w8(32'h3b04cab9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73071d),
	.w1(32'hbb9c0c35),
	.w2(32'hbc0baeaf),
	.w3(32'h3c4da16a),
	.w4(32'hbbcecdb7),
	.w5(32'hbc2129bb),
	.w6(32'hbb9c88db),
	.w7(32'hbc1a3c88),
	.w8(32'hbc1b48c2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc673185),
	.w1(32'hbbbd7c33),
	.w2(32'h3a8c6410),
	.w3(32'hbc3b42ce),
	.w4(32'hbc0a89f7),
	.w5(32'hbb8b8941),
	.w6(32'hbb539fca),
	.w7(32'h3b84106d),
	.w8(32'h3b9c1041),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5376c),
	.w1(32'hbb947414),
	.w2(32'hb8f496a1),
	.w3(32'h3adc5de2),
	.w4(32'h38e833f4),
	.w5(32'hbbd4b14f),
	.w6(32'h3c1ee15b),
	.w7(32'h3b7a0fa9),
	.w8(32'hbada90e3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac64faf),
	.w1(32'hbb9b5084),
	.w2(32'h3ac4084b),
	.w3(32'hbc052271),
	.w4(32'hbc3f60fa),
	.w5(32'hbc06532d),
	.w6(32'hbab6783b),
	.w7(32'h3bf0d2d6),
	.w8(32'h3be6677b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d461),
	.w1(32'h3c211312),
	.w2(32'h3c851320),
	.w3(32'hbad1aec6),
	.w4(32'h3c04740f),
	.w5(32'h3c39d1ec),
	.w6(32'hbaada377),
	.w7(32'h3c77d6d4),
	.w8(32'hbbd5bef8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a846058),
	.w1(32'h3b3e01a4),
	.w2(32'h3c5c8b5a),
	.w3(32'h3b7d5fee),
	.w4(32'h3a8e1f4c),
	.w5(32'h3bbc3634),
	.w6(32'hbbddfc30),
	.w7(32'h3b808200),
	.w8(32'h3ba0185d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a0867),
	.w1(32'hbcc7f5d1),
	.w2(32'hbd3c154a),
	.w3(32'h3bf64237),
	.w4(32'hbc833af2),
	.w5(32'hbcead962),
	.w6(32'hbc8b2c59),
	.w7(32'hbcf48eaf),
	.w8(32'hbc950202),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03a8c7),
	.w1(32'hb9af8664),
	.w2(32'h3bf3c385),
	.w3(32'hbcb60e29),
	.w4(32'hbba0acf3),
	.w5(32'hbab6b7b7),
	.w6(32'h3a6979f4),
	.w7(32'h3c2cea23),
	.w8(32'h3c2e56ba),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4632fd),
	.w1(32'hbb2d41d8),
	.w2(32'h3a8f260e),
	.w3(32'h3b9d7340),
	.w4(32'h3bc06974),
	.w5(32'h3c018287),
	.w6(32'h3a8fcf17),
	.w7(32'h3b8753ec),
	.w8(32'hbbda3924),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05a79c),
	.w1(32'h3babd2f3),
	.w2(32'h3c15e4a8),
	.w3(32'h3c849c24),
	.w4(32'h3b352368),
	.w5(32'h3c0f1353),
	.w6(32'h3b6cf904),
	.w7(32'h3bf28d5d),
	.w8(32'h3b2b5a6f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24b9fc),
	.w1(32'hbce409ff),
	.w2(32'hbd28f45c),
	.w3(32'h3bccccb4),
	.w4(32'hbcb37509),
	.w5(32'hbcaae2d5),
	.w6(32'hbc7c3cd7),
	.w7(32'hbca5494a),
	.w8(32'hbc97a1c1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdde3b1),
	.w1(32'hbc1e3d7d),
	.w2(32'hbc74e676),
	.w3(32'hbc9a85f6),
	.w4(32'h39b4b082),
	.w5(32'hbb8aead6),
	.w6(32'h3a00e515),
	.w7(32'hbb99de60),
	.w8(32'h3c1e1c0d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b686f),
	.w1(32'h3b1a3839),
	.w2(32'hb9f48558),
	.w3(32'hba7f8594),
	.w4(32'h3bcf4ec4),
	.w5(32'hbb22293a),
	.w6(32'hbb418480),
	.w7(32'hb9dbf364),
	.w8(32'h3c1cf488),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0fa72),
	.w1(32'hbc0d1274),
	.w2(32'hbc7b22eb),
	.w3(32'hbb9b1926),
	.w4(32'hbbb075c3),
	.w5(32'hbc7d0150),
	.w6(32'hbbd64d83),
	.w7(32'hbb0c94d5),
	.w8(32'h3a36fe47),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae52983),
	.w1(32'hbb5119b0),
	.w2(32'h3a226bb7),
	.w3(32'h3a2095f7),
	.w4(32'hbbc9e284),
	.w5(32'hbb3ce73a),
	.w6(32'hba93cd93),
	.w7(32'h3b8090cf),
	.w8(32'h3b4584de),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dab50c),
	.w1(32'h3b769f6f),
	.w2(32'h3c3e7573),
	.w3(32'h39fb9e57),
	.w4(32'h3af988d5),
	.w5(32'h3c637c10),
	.w6(32'h39dbb067),
	.w7(32'h3c0e7a15),
	.w8(32'hbbc0af83),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbda7),
	.w1(32'h3a37c37f),
	.w2(32'hbbe00a2e),
	.w3(32'h3aee9cd3),
	.w4(32'hbb36a595),
	.w5(32'h3b8515d0),
	.w6(32'hbb94e819),
	.w7(32'hbc30d6ac),
	.w8(32'hb92a5521),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d3886),
	.w1(32'h3a29e88c),
	.w2(32'hbac90a9a),
	.w3(32'hbb96b342),
	.w4(32'hba85a09b),
	.w5(32'h3b8d39bc),
	.w6(32'hbb898697),
	.w7(32'hbac50409),
	.w8(32'h3b900f1e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a0452),
	.w1(32'hbad1288e),
	.w2(32'hba979744),
	.w3(32'h3bfecb48),
	.w4(32'hb9b00d6d),
	.w5(32'hb9a6524c),
	.w6(32'h3a3e814b),
	.w7(32'hb60e7b58),
	.w8(32'h395a3b25),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39415725),
	.w1(32'h38f94819),
	.w2(32'h3c25bd37),
	.w3(32'h3a71f66d),
	.w4(32'h3bb87ee7),
	.w5(32'h3bc530c7),
	.w6(32'hbbc69547),
	.w7(32'hbabd3851),
	.w8(32'hba156dc2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule