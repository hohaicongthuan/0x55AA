module layer_10_featuremap_398(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ffeee),
	.w1(32'hbaf5ac17),
	.w2(32'hb9680ccb),
	.w3(32'h3bb21f22),
	.w4(32'hba315226),
	.w5(32'h3b11df4f),
	.w6(32'h3c418b09),
	.w7(32'h3a0e3329),
	.w8(32'h3bae6944),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88418),
	.w1(32'hbafeff37),
	.w2(32'hb8639041),
	.w3(32'hba9ed7b7),
	.w4(32'h3b734bbe),
	.w5(32'h38fb8f63),
	.w6(32'hbb2033f9),
	.w7(32'hba157f04),
	.w8(32'hbb965a5d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdd81),
	.w1(32'hbb9f6f57),
	.w2(32'hbb4d47be),
	.w3(32'hbb68a1be),
	.w4(32'h3aed9bdf),
	.w5(32'h3b88a41a),
	.w6(32'hbb12c7b7),
	.w7(32'hbb98fe01),
	.w8(32'hbbd38e31),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6f09),
	.w1(32'hbbed1aed),
	.w2(32'hbba7ce27),
	.w3(32'hbbef7645),
	.w4(32'hbbc75c5a),
	.w5(32'hba5d49c5),
	.w6(32'hbb7d0e52),
	.w7(32'h3b0c190d),
	.w8(32'hbadc9be7),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa28c4),
	.w1(32'hbb04a941),
	.w2(32'hbb527982),
	.w3(32'hbc062fd6),
	.w4(32'h3beb85af),
	.w5(32'h3b243fe8),
	.w6(32'hbb9542d5),
	.w7(32'h3bafc686),
	.w8(32'h3b66b434),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ab1f8),
	.w1(32'h3ad8ac09),
	.w2(32'h3c0f7539),
	.w3(32'h3ab3d943),
	.w4(32'hbbc93ce9),
	.w5(32'h3b8ee62f),
	.w6(32'hba465ec1),
	.w7(32'h38172f20),
	.w8(32'hba5d3fd4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb362e),
	.w1(32'hbb3d9af7),
	.w2(32'h3b4e6e2d),
	.w3(32'hbb73d3a5),
	.w4(32'hba975d76),
	.w5(32'h3be3b763),
	.w6(32'hbbcb20ca),
	.w7(32'hbb5739f9),
	.w8(32'hbb349a8d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964284),
	.w1(32'hbc447807),
	.w2(32'hbc2342df),
	.w3(32'hbacd7978),
	.w4(32'h3ba5baff),
	.w5(32'h3c2454ec),
	.w6(32'hb9a1604b),
	.w7(32'hbb920c38),
	.w8(32'hbb07b394),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc017faf),
	.w1(32'hbaeba46a),
	.w2(32'hbb60422c),
	.w3(32'hbbe21c0c),
	.w4(32'h3a854eb9),
	.w5(32'hbb3086fa),
	.w6(32'hbaf0f0b1),
	.w7(32'h3ad19223),
	.w8(32'hbb50977a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b83d1),
	.w1(32'hbb222f84),
	.w2(32'hbb92c096),
	.w3(32'hbba79dbb),
	.w4(32'hbbad5273),
	.w5(32'h3b704c3f),
	.w6(32'hbae8cfa5),
	.w7(32'h3b04abdf),
	.w8(32'h3c284a04),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1938db),
	.w1(32'h39d0a5f8),
	.w2(32'hbbb170a7),
	.w3(32'h3c3f93ea),
	.w4(32'h3b901e8f),
	.w5(32'hbbf31b70),
	.w6(32'h3bc9cdca),
	.w7(32'h3c5a3b01),
	.w8(32'h3bf36e90),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95455),
	.w1(32'h3a8c55fc),
	.w2(32'h3bc18ce6),
	.w3(32'hbb367a7f),
	.w4(32'h3b6a4c5c),
	.w5(32'h3b934b95),
	.w6(32'h3ba4b592),
	.w7(32'hbb3b603c),
	.w8(32'hbb0c37fc),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a45d7),
	.w1(32'hbb843ef7),
	.w2(32'hbbdeeefe),
	.w3(32'hbb930136),
	.w4(32'hbb30980c),
	.w5(32'h3b4d7e3d),
	.w6(32'h3b0e58a8),
	.w7(32'hbbf4298d),
	.w8(32'hbbffbb64),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe333e4),
	.w1(32'hbb227d73),
	.w2(32'hbadc30d5),
	.w3(32'hbb9b5f42),
	.w4(32'hbb87ebb0),
	.w5(32'hb8310aae),
	.w6(32'hba976cf0),
	.w7(32'hbbc6448e),
	.w8(32'hbae3cb0b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9e4b3),
	.w1(32'hbbb60c9c),
	.w2(32'h3b3a94cf),
	.w3(32'h3a134d01),
	.w4(32'hbb3fe216),
	.w5(32'h3c0c5f14),
	.w6(32'hbb9944eb),
	.w7(32'hbb5133e0),
	.w8(32'hbb9522c4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab4093),
	.w1(32'hb9c63c4f),
	.w2(32'h3893227e),
	.w3(32'h3a9ff434),
	.w4(32'hbac18da8),
	.w5(32'h3baa751b),
	.w6(32'hbb1ac50d),
	.w7(32'hbb3d6ffa),
	.w8(32'hbb58b434),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22f2fc),
	.w1(32'h3a994e6a),
	.w2(32'hba865d75),
	.w3(32'hba8067c3),
	.w4(32'h3b8b5566),
	.w5(32'hb925fedb),
	.w6(32'hba86fe24),
	.w7(32'h3bc050b6),
	.w8(32'hb9f32963),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24acb3),
	.w1(32'hbbbd25bf),
	.w2(32'hbb174233),
	.w3(32'h3ac7d9ed),
	.w4(32'h3ab562d0),
	.w5(32'h3b9aa7af),
	.w6(32'hb998a571),
	.w7(32'hb9bd736e),
	.w8(32'h3b82311b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3763c6),
	.w1(32'hbb428dcc),
	.w2(32'hbb43860e),
	.w3(32'hbba52373),
	.w4(32'h3920daba),
	.w5(32'h3b505a08),
	.w6(32'hbbc9918c),
	.w7(32'hbb74fa1a),
	.w8(32'hbbe18674),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cb13a),
	.w1(32'h3bd28494),
	.w2(32'h3c994642),
	.w3(32'hbaec5708),
	.w4(32'h3c05c52d),
	.w5(32'hbacaf751),
	.w6(32'h3b07a51b),
	.w7(32'h3bd9776d),
	.w8(32'hbbc525f0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5011f0),
	.w1(32'hba827025),
	.w2(32'h3bc9625a),
	.w3(32'h3c0ec6a8),
	.w4(32'h3bd0e1a9),
	.w5(32'h3c3bede8),
	.w6(32'hbbabf865),
	.w7(32'hbb24ba6f),
	.w8(32'h3a983eac),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3d370),
	.w1(32'hb8454cdb),
	.w2(32'hbb561f55),
	.w3(32'hbb362fd3),
	.w4(32'h3b53d15d),
	.w5(32'hbc30740f),
	.w6(32'h3b969b0f),
	.w7(32'h3ab4636e),
	.w8(32'hbb794acf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb968eec),
	.w1(32'hb9efe181),
	.w2(32'hbba8b43d),
	.w3(32'h3b4bfc0e),
	.w4(32'h39f80887),
	.w5(32'hbc0022e3),
	.w6(32'h3954ec91),
	.w7(32'h38e514ac),
	.w8(32'hbbc2891b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049752),
	.w1(32'h3c0710c8),
	.w2(32'h3bb67068),
	.w3(32'h3a2835af),
	.w4(32'h3bce6339),
	.w5(32'h3d44c0b4),
	.w6(32'h3b7994fb),
	.w7(32'h3bde584b),
	.w8(32'hbcbee5af),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64adbb),
	.w1(32'hbbb75593),
	.w2(32'hb9bde358),
	.w3(32'hbc4703b0),
	.w4(32'h3bdca90d),
	.w5(32'hbb492bfc),
	.w6(32'h3c213ced),
	.w7(32'hba92bf96),
	.w8(32'hbb9b684d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a439a62),
	.w1(32'h3c699fc1),
	.w2(32'h3c1c483e),
	.w3(32'hbc132d6a),
	.w4(32'h3be371ab),
	.w5(32'hbbe4eddc),
	.w6(32'h3aee41ac),
	.w7(32'h3bd12168),
	.w8(32'h3c414849),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc2362),
	.w1(32'h3c2159c1),
	.w2(32'hb8e16178),
	.w3(32'h3ac51721),
	.w4(32'hbb9241bf),
	.w5(32'hbbaa7440),
	.w6(32'h3b66e235),
	.w7(32'hbc2e2069),
	.w8(32'h398a23e0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f24a0),
	.w1(32'h3b05fe9e),
	.w2(32'h3a300476),
	.w3(32'h3bca1c94),
	.w4(32'h3b029b06),
	.w5(32'h3b8d08ee),
	.w6(32'h3be7ee30),
	.w7(32'hbb84cd4b),
	.w8(32'hbbaa6e0d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8f97),
	.w1(32'h3be53af5),
	.w2(32'h3c08a838),
	.w3(32'h3b0f20fa),
	.w4(32'h3bee3d60),
	.w5(32'hb9ab4dc6),
	.w6(32'hba8f1d4d),
	.w7(32'hbb8abc5e),
	.w8(32'h3b35236a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13dd1f),
	.w1(32'hbbcfe6c7),
	.w2(32'hb968a4ee),
	.w3(32'h3ad5f893),
	.w4(32'hbae37c55),
	.w5(32'h3ae109f5),
	.w6(32'h3ada6718),
	.w7(32'hbb1b9fca),
	.w8(32'h3b33fda4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0628f),
	.w1(32'hba094723),
	.w2(32'h3b9fe2ff),
	.w3(32'hbc0db432),
	.w4(32'h3acdfbf4),
	.w5(32'h3b8ca88f),
	.w6(32'hbb2c71f4),
	.w7(32'h3b009012),
	.w8(32'h3bbfe4da),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88eee8e),
	.w1(32'hbba88458),
	.w2(32'hba6c4fc9),
	.w3(32'h3b86471f),
	.w4(32'h3981e494),
	.w5(32'hb9f41192),
	.w6(32'h3b361724),
	.w7(32'h3a7bb6ab),
	.w8(32'hba114e56),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a29e6),
	.w1(32'hba9ab321),
	.w2(32'hbc01ad09),
	.w3(32'hba352b7a),
	.w4(32'hbc10063e),
	.w5(32'hbb93dc79),
	.w6(32'h3ae04203),
	.w7(32'h3b1327a5),
	.w8(32'h3b41ec9f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acb8d),
	.w1(32'hbb0571dc),
	.w2(32'hbb8071b0),
	.w3(32'h3bb6d554),
	.w4(32'hb914dfe2),
	.w5(32'h3b957aae),
	.w6(32'h3aafa03d),
	.w7(32'h3b8d5b08),
	.w8(32'h3c0426db),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8215d9),
	.w1(32'hbb569644),
	.w2(32'h3b5a2900),
	.w3(32'h3b821602),
	.w4(32'hb9412997),
	.w5(32'h3be9ad83),
	.w6(32'hb9be4ed7),
	.w7(32'hbc40ac74),
	.w8(32'hbc078b51),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7965e),
	.w1(32'hbbc19ac0),
	.w2(32'h3b5403d9),
	.w3(32'h3b05f87c),
	.w4(32'hbadec0f9),
	.w5(32'h3bd44f96),
	.w6(32'hbbefac9d),
	.w7(32'hba894619),
	.w8(32'h3922f08c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ecb6),
	.w1(32'hbb7e48c6),
	.w2(32'hbb9e9a81),
	.w3(32'hbbb67187),
	.w4(32'h3b180d27),
	.w5(32'hbc14664a),
	.w6(32'hbc04a4e3),
	.w7(32'h3bc41294),
	.w8(32'hba800f11),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaabc85),
	.w1(32'hbb27fd9c),
	.w2(32'hba1c47de),
	.w3(32'hbaa08de0),
	.w4(32'hb9b3ec2f),
	.w5(32'hbb9cd993),
	.w6(32'hba6852de),
	.w7(32'h38fe3f40),
	.w8(32'hbb735efa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8796d5),
	.w1(32'hbc0c2ad5),
	.w2(32'hbae8b9df),
	.w3(32'h3b4f2790),
	.w4(32'hbc2a3be7),
	.w5(32'h3b90a638),
	.w6(32'hbb3f8477),
	.w7(32'hbbe7cc65),
	.w8(32'hbb9f3723),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc177eea),
	.w1(32'h39aa7f0d),
	.w2(32'h3b046b81),
	.w3(32'hbaab79d6),
	.w4(32'h3b38f85a),
	.w5(32'h3b748519),
	.w6(32'hbc05a36e),
	.w7(32'h3a90bc0e),
	.w8(32'h3ba08d2c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb6f28),
	.w1(32'hbb61dcb4),
	.w2(32'hbc4ed049),
	.w3(32'h3bce74cf),
	.w4(32'hbc2ad886),
	.w5(32'h3af1fda3),
	.w6(32'h3b40060e),
	.w7(32'hba8a8e82),
	.w8(32'hbc3894b0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb767cd8),
	.w1(32'hbb016375),
	.w2(32'hba9d814d),
	.w3(32'hbc374115),
	.w4(32'h3a6c9ea1),
	.w5(32'h3b860158),
	.w6(32'h38ce5d29),
	.w7(32'hbafade44),
	.w8(32'hbb84da90),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab35a93),
	.w1(32'hbafaa56f),
	.w2(32'hbb905422),
	.w3(32'hbb7adabc),
	.w4(32'h3b2c3f28),
	.w5(32'h3b8b1576),
	.w6(32'h3ba9e72c),
	.w7(32'hbaa7beb4),
	.w8(32'hbb9e5311),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1939fa),
	.w1(32'hbbba25fd),
	.w2(32'hbbf59d27),
	.w3(32'hbb467bf6),
	.w4(32'hbb0c2839),
	.w5(32'h3b8ca4dd),
	.w6(32'h3b0076e1),
	.w7(32'hbb82153a),
	.w8(32'hbb207cca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a66ad),
	.w1(32'hbbe884cf),
	.w2(32'hbbb29718),
	.w3(32'hb9d90fab),
	.w4(32'hbbd3f3ff),
	.w5(32'hba5bdaa2),
	.w6(32'hbacf9625),
	.w7(32'hbbacb5c9),
	.w8(32'hbbbc1b8a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b68d8),
	.w1(32'h3a16e62c),
	.w2(32'hba064fa9),
	.w3(32'h3adb530b),
	.w4(32'hb99f1971),
	.w5(32'h3c24ddd6),
	.w6(32'h3b01032c),
	.w7(32'hbb9fd6d4),
	.w8(32'hbb8fc284),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb25874),
	.w1(32'h3bd2275a),
	.w2(32'h3c940e7c),
	.w3(32'hbab71a30),
	.w4(32'hbaedc490),
	.w5(32'h3c0ffaa9),
	.w6(32'hbb2449b9),
	.w7(32'hbb1e62ed),
	.w8(32'hbc259cd7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bed96f),
	.w1(32'hbad98720),
	.w2(32'h3ae062f8),
	.w3(32'hbb9cdc00),
	.w4(32'hbc18b2bf),
	.w5(32'hba933c2d),
	.w6(32'h3b21e2fb),
	.w7(32'hbba7dff8),
	.w8(32'hbb81a198),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c3033),
	.w1(32'hbb19b232),
	.w2(32'h3bde991b),
	.w3(32'h3bc647e9),
	.w4(32'hbb9a8bdc),
	.w5(32'h3b69c929),
	.w6(32'hbb901b4e),
	.w7(32'hbbfa4536),
	.w8(32'hbb81835a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c7aa),
	.w1(32'hbad763de),
	.w2(32'h3c035a88),
	.w3(32'hbc8bce60),
	.w4(32'hbb19c128),
	.w5(32'h3b1d0fd4),
	.w6(32'hbb79c483),
	.w7(32'hbb4256c4),
	.w8(32'h3a01f10f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfebbe),
	.w1(32'hbae264f3),
	.w2(32'hbaa4f1ce),
	.w3(32'hbc9020f1),
	.w4(32'hbba43665),
	.w5(32'hbb242d86),
	.w6(32'hbb8dd705),
	.w7(32'hbb332856),
	.w8(32'hbbe8c968),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb595c00),
	.w1(32'hbad34b22),
	.w2(32'hbb1ea43c),
	.w3(32'hbb5a6760),
	.w4(32'hb9d21ee8),
	.w5(32'h3c138e14),
	.w6(32'h3a88d921),
	.w7(32'hbb880eed),
	.w8(32'hbc1a2ef4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391eca83),
	.w1(32'hbae1a808),
	.w2(32'hbb07407d),
	.w3(32'hbad6928e),
	.w4(32'hbbbcb40d),
	.w5(32'h3b0f4147),
	.w6(32'hbb998e9b),
	.w7(32'h3ab1a80b),
	.w8(32'hbb312169),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba019ea7),
	.w1(32'h3b44d310),
	.w2(32'hbb3d1edb),
	.w3(32'hbbb3d3ea),
	.w4(32'h3a85e617),
	.w5(32'hbaba9ebe),
	.w6(32'hba921148),
	.w7(32'hbbe603b1),
	.w8(32'hbbcbb967),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb949f1a),
	.w1(32'hbbf47b56),
	.w2(32'h38d8ca35),
	.w3(32'hbb435f9b),
	.w4(32'hbac77128),
	.w5(32'h3b9f76f2),
	.w6(32'h3b0989f8),
	.w7(32'hbb5182ef),
	.w8(32'hba935da9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745435),
	.w1(32'h3af81e2f),
	.w2(32'h3a3b3719),
	.w3(32'h3ba7e165),
	.w4(32'h3b43ee77),
	.w5(32'h3b971796),
	.w6(32'hbc106965),
	.w7(32'hbb0d8354),
	.w8(32'h3b1ffc3c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401754),
	.w1(32'hbad77877),
	.w2(32'hbbd7ee63),
	.w3(32'hba608802),
	.w4(32'hba5cb5dd),
	.w5(32'hbbe303fc),
	.w6(32'hbb825cb0),
	.w7(32'hbb0f2c53),
	.w8(32'hbb9571d3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf654b),
	.w1(32'hba89a49f),
	.w2(32'h3b71eea4),
	.w3(32'hbb5b28f9),
	.w4(32'hbaed4259),
	.w5(32'h3c3205f0),
	.w6(32'h3b0f7eff),
	.w7(32'h3b2a8fe4),
	.w8(32'h3b6ff806),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0679a0),
	.w1(32'h3bc4fbe1),
	.w2(32'h3b748afe),
	.w3(32'h3b424568),
	.w4(32'h3bf20885),
	.w5(32'h3c5e7286),
	.w6(32'h39ca3bd2),
	.w7(32'h3b34e63b),
	.w8(32'h3a8f3b83),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19a995),
	.w1(32'hbb70bf83),
	.w2(32'h3bebe5ee),
	.w3(32'hbbe85b5e),
	.w4(32'h3a226b45),
	.w5(32'hb9a736cf),
	.w6(32'hbc690e9a),
	.w7(32'h3c05b5b7),
	.w8(32'h3a5df524),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4cfa6),
	.w1(32'h3b953eab),
	.w2(32'h3cbccace),
	.w3(32'h39dc8b0c),
	.w4(32'h3bbe2a34),
	.w5(32'h3c5890c2),
	.w6(32'hbb8c2274),
	.w7(32'hba95f784),
	.w8(32'h3c0ad00e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaea3fd),
	.w1(32'h3b8db079),
	.w2(32'h3a7a2996),
	.w3(32'h3c2d9077),
	.w4(32'h3ba87274),
	.w5(32'h3b74348d),
	.w6(32'h3b1ca8dd),
	.w7(32'h3b01a0f7),
	.w8(32'h3b57b79a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9f90),
	.w1(32'hbbb302a0),
	.w2(32'h3a946ca6),
	.w3(32'h3b6822f6),
	.w4(32'h3b603e9c),
	.w5(32'h3c82210e),
	.w6(32'h3b061d71),
	.w7(32'hbbcfab53),
	.w8(32'hbb1041fd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70c2bf),
	.w1(32'hbb10c5f2),
	.w2(32'hba534dc0),
	.w3(32'hbbb8a16a),
	.w4(32'hb9834763),
	.w5(32'h3a2bdfd7),
	.w6(32'hb984bb98),
	.w7(32'hbb716c73),
	.w8(32'hbb7555c9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a093),
	.w1(32'hbc9029d2),
	.w2(32'hbbe0690a),
	.w3(32'h3ad32099),
	.w4(32'hbbdccbf7),
	.w5(32'hba94eb67),
	.w6(32'hba32b54a),
	.w7(32'hbca87fa6),
	.w8(32'hbc684093),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e9f27),
	.w1(32'hbb038a19),
	.w2(32'hbaf3356f),
	.w3(32'hbc828f96),
	.w4(32'hbb96dee8),
	.w5(32'hb9e3c733),
	.w6(32'hbc5be3cc),
	.w7(32'hbaba809f),
	.w8(32'hbb481c31),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72b1f5),
	.w1(32'hbb141892),
	.w2(32'hbbdee6cf),
	.w3(32'hbc3df4cd),
	.w4(32'hbb1df311),
	.w5(32'hbc85a399),
	.w6(32'hbb9c8864),
	.w7(32'h3bbb5fd7),
	.w8(32'h3b022a19),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b5a77d),
	.w1(32'h3b428b77),
	.w2(32'h3c85fa99),
	.w3(32'hba93d6dd),
	.w4(32'h3c161048),
	.w5(32'h3b4b75a0),
	.w6(32'h39c3f88a),
	.w7(32'h3b4be884),
	.w8(32'h3a3df6d6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f25c3),
	.w1(32'h3b1f4c33),
	.w2(32'hba8a2aa3),
	.w3(32'hbbcc4ca0),
	.w4(32'h3bb26197),
	.w5(32'h3ad87594),
	.w6(32'hbbf7faa2),
	.w7(32'hbbbeb997),
	.w8(32'hbbaf6902),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3ff1),
	.w1(32'hbb6bca64),
	.w2(32'h39ed7202),
	.w3(32'h3b34593f),
	.w4(32'hbbf07901),
	.w5(32'hbb938e04),
	.w6(32'hbaf60adb),
	.w7(32'hbb10434c),
	.w8(32'h3ad90142),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119f4e),
	.w1(32'hbb39216e),
	.w2(32'hbac3a3a0),
	.w3(32'hbc8b7ae1),
	.w4(32'hbb81381f),
	.w5(32'hbbc7ed48),
	.w6(32'hbc220d64),
	.w7(32'hbba64f31),
	.w8(32'hbbfa4e3e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f596),
	.w1(32'h3ba78f14),
	.w2(32'h3ad2f087),
	.w3(32'hbc123d01),
	.w4(32'h3ba4ba91),
	.w5(32'hbc01ac65),
	.w6(32'hbbbf1d89),
	.w7(32'h3c1efe27),
	.w8(32'h3bb5ee89),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba37ac0),
	.w1(32'hba5a184b),
	.w2(32'h3a83fc16),
	.w3(32'h39fcf1a3),
	.w4(32'hbb929faa),
	.w5(32'h3bb4ce2d),
	.w6(32'hbb41487c),
	.w7(32'h3a7b0ea2),
	.w8(32'h3b231be4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69dc0c),
	.w1(32'h3bae8dfa),
	.w2(32'hba022849),
	.w3(32'hbba8c3a8),
	.w4(32'h3bd47030),
	.w5(32'hbb9f159c),
	.w6(32'hbb4fe9e5),
	.w7(32'h3b8f9f11),
	.w8(32'h3b84d62d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617349),
	.w1(32'hbc1037fb),
	.w2(32'hbbf592ec),
	.w3(32'h3bb13135),
	.w4(32'hbbf4f05c),
	.w5(32'hbc0c1894),
	.w6(32'h3b87f3f8),
	.w7(32'hbc4f5dfc),
	.w8(32'hbc1a252a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7b84),
	.w1(32'hbafa1228),
	.w2(32'hbba4675f),
	.w3(32'h3aa40f39),
	.w4(32'h3b5d7677),
	.w5(32'hbb1b9418),
	.w6(32'hbc1f9da3),
	.w7(32'hb92e9b54),
	.w8(32'h3a8007cd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a68ef),
	.w1(32'h3b4fcb56),
	.w2(32'hb9ef4ef5),
	.w3(32'hbb555ac0),
	.w4(32'h3ae4be6d),
	.w5(32'h3cd2243b),
	.w6(32'h3ae10150),
	.w7(32'h39e13a65),
	.w8(32'h3c976808),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04c8a5),
	.w1(32'hb9986ca8),
	.w2(32'hbbe94d1c),
	.w3(32'hbc028545),
	.w4(32'h3c29039c),
	.w5(32'hbbef8e23),
	.w6(32'h3b583c19),
	.w7(32'h3bb50ce2),
	.w8(32'h3b1b6b87),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eadcf),
	.w1(32'h3b84d38f),
	.w2(32'hbaf80204),
	.w3(32'h3b344089),
	.w4(32'h3bfd5ae0),
	.w5(32'hbb09f677),
	.w6(32'hbbab318b),
	.w7(32'h38edf1ec),
	.w8(32'h3b84d057),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15af33),
	.w1(32'h3c20c49d),
	.w2(32'hbc267cc5),
	.w3(32'h3ac98f20),
	.w4(32'hba9326d5),
	.w5(32'h3d1e6dcf),
	.w6(32'h39bf2e4d),
	.w7(32'hbbecd500),
	.w8(32'hb8863dd7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfcda),
	.w1(32'h3adfc4a3),
	.w2(32'hbb5c7568),
	.w3(32'hbb7c1f2b),
	.w4(32'h3ae0e646),
	.w5(32'hbc23e562),
	.w6(32'h3ba1f983),
	.w7(32'h3b0796d0),
	.w8(32'h3b61fcff),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4adfef),
	.w1(32'h3a1de218),
	.w2(32'h3ac33265),
	.w3(32'h3a4bb28d),
	.w4(32'h3b82b8b8),
	.w5(32'hbb77f2d3),
	.w6(32'h3b90112b),
	.w7(32'h3c088614),
	.w8(32'h3b8212d2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20451a),
	.w1(32'h3b58beff),
	.w2(32'h3b4ad5d1),
	.w3(32'h3b46f135),
	.w4(32'hba9458a1),
	.w5(32'h3aa2ef5d),
	.w6(32'h39ec0bce),
	.w7(32'hba687654),
	.w8(32'h3b009f7e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b0b18),
	.w1(32'hbba2063f),
	.w2(32'hbc443c90),
	.w3(32'hb71474af),
	.w4(32'h3ab7f031),
	.w5(32'hbc6a2411),
	.w6(32'h3b6097a7),
	.w7(32'hbbaa37f5),
	.w8(32'hbc2ddf3f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124c49),
	.w1(32'h3afccec1),
	.w2(32'h3b185341),
	.w3(32'h3bb37db2),
	.w4(32'hbb9dfdfe),
	.w5(32'h3bdf07ac),
	.w6(32'h3ac979ac),
	.w7(32'h3bf01169),
	.w8(32'h38cc5798),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2aa59),
	.w1(32'h3a0610db),
	.w2(32'hbc3c03a1),
	.w3(32'hbae9dd4e),
	.w4(32'h3b4e3705),
	.w5(32'hbcaba3ed),
	.w6(32'h3a12500e),
	.w7(32'hbb0407d1),
	.w8(32'hbc39784b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba89f26),
	.w1(32'hbadcc009),
	.w2(32'h3ba83e61),
	.w3(32'hbc3ce7bd),
	.w4(32'hbb80f570),
	.w5(32'h3ccfba68),
	.w6(32'hbc086d6a),
	.w7(32'h3a8025de),
	.w8(32'hbb93ef35),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45f753),
	.w1(32'h3b78cd2a),
	.w2(32'h3c116389),
	.w3(32'h3c101766),
	.w4(32'hbb57614f),
	.w5(32'hbb1ba3a0),
	.w6(32'hbb0ffb16),
	.w7(32'h3b86535e),
	.w8(32'hbb58ee6b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137ecf),
	.w1(32'hbace2dec),
	.w2(32'hbbf31898),
	.w3(32'h3b3c5cd6),
	.w4(32'h3c6cd1c6),
	.w5(32'h3af99e04),
	.w6(32'hbbe0389c),
	.w7(32'hb9d61fec),
	.w8(32'hbae32712),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf00478),
	.w1(32'hbba7d22a),
	.w2(32'hbbc016f4),
	.w3(32'hbbb05255),
	.w4(32'hb9e65aab),
	.w5(32'hba3b1d5d),
	.w6(32'hbb655c5c),
	.w7(32'h3b4caeac),
	.w8(32'hbb1318f0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43f717),
	.w1(32'hbc14baa1),
	.w2(32'hbb8e6dfa),
	.w3(32'h3b85b0db),
	.w4(32'hbbd970c7),
	.w5(32'hbb9f664b),
	.w6(32'hbbd500e2),
	.w7(32'hbb8bd96b),
	.w8(32'hbbb21088),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03e3ff),
	.w1(32'h3ba3d5cf),
	.w2(32'hba8d4a16),
	.w3(32'hbb16bfc6),
	.w4(32'h3b4f30e1),
	.w5(32'h3b7f4a2b),
	.w6(32'h3b2ba743),
	.w7(32'h3a1dd34c),
	.w8(32'hbb465786),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2783b6),
	.w1(32'h3c3b952c),
	.w2(32'h3bd6c6f4),
	.w3(32'h3b983bdc),
	.w4(32'h3b0a3a2a),
	.w5(32'h3a5d47e8),
	.w6(32'h3bacaf96),
	.w7(32'h3b34fbe4),
	.w8(32'hbb82ef9c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f92bc),
	.w1(32'h37a9ec34),
	.w2(32'h3937ed74),
	.w3(32'h3a498bb8),
	.w4(32'hbbee3ae0),
	.w5(32'hbbfb99c8),
	.w6(32'hbb094748),
	.w7(32'hbaae0ae5),
	.w8(32'h3b0d6273),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98411b),
	.w1(32'h3b96d262),
	.w2(32'hbc2d6368),
	.w3(32'hbb8b73ab),
	.w4(32'h3c0df800),
	.w5(32'h3cde2e98),
	.w6(32'h3b41dbe1),
	.w7(32'hbc3e6093),
	.w8(32'hbc0c672b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da9bf),
	.w1(32'h3af00b63),
	.w2(32'h3a16bf83),
	.w3(32'h3b6b5860),
	.w4(32'hbb6d9fe8),
	.w5(32'h3c20f63c),
	.w6(32'hb92c9a6f),
	.w7(32'hbb4de6a2),
	.w8(32'h3b0eb7eb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37813),
	.w1(32'hb9c5077d),
	.w2(32'h39b34402),
	.w3(32'hbb861735),
	.w4(32'h39c66db2),
	.w5(32'hbc30b085),
	.w6(32'hba817cdc),
	.w7(32'h3a201c3e),
	.w8(32'hbad5af3e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ff361),
	.w1(32'h3bb00ce9),
	.w2(32'h3b871c10),
	.w3(32'hb95e7b89),
	.w4(32'hbb05c98f),
	.w5(32'h3c5af3ab),
	.w6(32'hbb5de6ba),
	.w7(32'hbbc010f3),
	.w8(32'h3ae50f3c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3451a),
	.w1(32'hbc0b3b9f),
	.w2(32'hbb934c32),
	.w3(32'hbbac0cc7),
	.w4(32'hbb4fff3d),
	.w5(32'hbbf351ab),
	.w6(32'hbbbb6e22),
	.w7(32'hbb9b61d6),
	.w8(32'hbbfe64ce),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4238eb),
	.w1(32'hbc454c2c),
	.w2(32'hbc2cecef),
	.w3(32'hbbfdf049),
	.w4(32'h3ad2b650),
	.w5(32'hbbe92d6d),
	.w6(32'hbc4489df),
	.w7(32'hbbe5c335),
	.w8(32'h3a29385a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aacbe),
	.w1(32'h3bae10bf),
	.w2(32'hba5a31cc),
	.w3(32'h3ac9ac12),
	.w4(32'h3c1fcfd6),
	.w5(32'h3baaa2c4),
	.w6(32'hbc213efc),
	.w7(32'hba7a5852),
	.w8(32'h3b39f089),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba982840),
	.w1(32'h3ad4941c),
	.w2(32'hbb957d43),
	.w3(32'hb9f3d003),
	.w4(32'h3b26fbfd),
	.w5(32'h3c14cbe3),
	.w6(32'h398eb8a9),
	.w7(32'h3b19e11b),
	.w8(32'h3b0e2e64),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b1500),
	.w1(32'h3b848c58),
	.w2(32'hbbb8ad57),
	.w3(32'hbbfb88dd),
	.w4(32'h3b4b7f8d),
	.w5(32'hbb9d798f),
	.w6(32'hbb5c9f95),
	.w7(32'hbaa32f6e),
	.w8(32'hbb8e47f2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21724a),
	.w1(32'h39d16b5b),
	.w2(32'hbaa031bd),
	.w3(32'h38fcbf8f),
	.w4(32'hba6387e0),
	.w5(32'h3c168eb4),
	.w6(32'h3a5e3803),
	.w7(32'h3b1489d3),
	.w8(32'hba8c37aa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56511),
	.w1(32'h3b1823a6),
	.w2(32'hbb2dff60),
	.w3(32'hbb9e50f6),
	.w4(32'hbaa8a2c0),
	.w5(32'h3c7cae5a),
	.w6(32'hbb1985a6),
	.w7(32'h395a326c),
	.w8(32'h3c114735),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca70c2),
	.w1(32'h3b152af3),
	.w2(32'hbb700376),
	.w3(32'h3b8e87cc),
	.w4(32'hb9915209),
	.w5(32'hbaec3c54),
	.w6(32'h3bda7ca7),
	.w7(32'hba27fa65),
	.w8(32'hb9b32a91),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b171e1b),
	.w1(32'hba8050f2),
	.w2(32'h3b527b90),
	.w3(32'hbb59a638),
	.w4(32'h3ad5025e),
	.w5(32'hbbe01ae9),
	.w6(32'h39498871),
	.w7(32'h3b2ff90b),
	.w8(32'h3b0dc37d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30ea1f),
	.w1(32'h3ad7133e),
	.w2(32'h3a54ef7d),
	.w3(32'h3b94d651),
	.w4(32'hbc20330d),
	.w5(32'hbba66af4),
	.w6(32'hbabd51e4),
	.w7(32'hbc22885b),
	.w8(32'hbb85fe65),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc307701),
	.w1(32'h3b668061),
	.w2(32'hbb652d07),
	.w3(32'hb9f4367d),
	.w4(32'hbae478f7),
	.w5(32'h3ad75495),
	.w6(32'h3ba858aa),
	.w7(32'h3b35d0e0),
	.w8(32'hba410209),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4231e4),
	.w1(32'h3b511d6a),
	.w2(32'h3b6e7eb2),
	.w3(32'hbbc5b77c),
	.w4(32'hbbe3b6f6),
	.w5(32'h3d0ee2e8),
	.w6(32'hbbd9f214),
	.w7(32'h39c5845c),
	.w8(32'h3b489278),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68faf),
	.w1(32'hbbd64cc9),
	.w2(32'hbc0536ec),
	.w3(32'h3b3ae2ff),
	.w4(32'hbb1a61dd),
	.w5(32'hbbe15c47),
	.w6(32'hb94d0b75),
	.w7(32'hbb4cbe6e),
	.w8(32'hbbaa6a79),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d39b4),
	.w1(32'hbb1921a0),
	.w2(32'hbc4056b1),
	.w3(32'hbb15678b),
	.w4(32'h3b98adb5),
	.w5(32'hbb790a1e),
	.w6(32'hbbc17223),
	.w7(32'hbb1758ad),
	.w8(32'hbac7ffdd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aa1d6),
	.w1(32'h3ba22396),
	.w2(32'hbb246c8e),
	.w3(32'hbc1931be),
	.w4(32'h3bd55021),
	.w5(32'hbbe4d373),
	.w6(32'hbbf86af0),
	.w7(32'h3b1938bf),
	.w8(32'h3aae93e3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf95684),
	.w1(32'hbb5901d1),
	.w2(32'hbab40302),
	.w3(32'hba015bc2),
	.w4(32'h3bf2f26d),
	.w5(32'hbc2517e1),
	.w6(32'h3b125e75),
	.w7(32'hbb8385d1),
	.w8(32'hba10f468),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a145672),
	.w1(32'h3b86c516),
	.w2(32'h3b93876b),
	.w3(32'h3b0fba57),
	.w4(32'hbaa1d2ec),
	.w5(32'h3c166bb0),
	.w6(32'hbb77c9fc),
	.w7(32'hbb04d8f4),
	.w8(32'h394e5e13),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc392c60),
	.w1(32'hbaad09db),
	.w2(32'hbb159879),
	.w3(32'hbbc2a185),
	.w4(32'hbc07c2b8),
	.w5(32'hb9305907),
	.w6(32'h3b6f380b),
	.w7(32'hbb0a391b),
	.w8(32'hbb72d04f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaebaa),
	.w1(32'h3a8d6083),
	.w2(32'h3b945d1c),
	.w3(32'hbc498176),
	.w4(32'hbb9255c6),
	.w5(32'h3c8e0961),
	.w6(32'hbc1f8fe4),
	.w7(32'h3a326d61),
	.w8(32'hbb637020),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fa1f8),
	.w1(32'hb95316e2),
	.w2(32'hbab0a9de),
	.w3(32'hbb417615),
	.w4(32'hbb3a9df6),
	.w5(32'hba644d9a),
	.w6(32'h3abbb210),
	.w7(32'hbb5925fd),
	.w8(32'h3c083f00),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ee7de),
	.w1(32'h3baae9e3),
	.w2(32'hbacaade3),
	.w3(32'hbba983eb),
	.w4(32'h3bb0ce85),
	.w5(32'hbc1d5c16),
	.w6(32'h3b887584),
	.w7(32'h3b70daec),
	.w8(32'h3b460932),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b5e0),
	.w1(32'h38f40c83),
	.w2(32'hba1fca11),
	.w3(32'h3c20a9d4),
	.w4(32'hbaee075b),
	.w5(32'h3bb97a4b),
	.w6(32'h397149e1),
	.w7(32'hbbbc7b6e),
	.w8(32'hbc1b9e96),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0ce18),
	.w1(32'hbb9228ea),
	.w2(32'hbc213c9d),
	.w3(32'hba946f60),
	.w4(32'h3b6f7095),
	.w5(32'hbb345105),
	.w6(32'hbb65cb38),
	.w7(32'hb8af6e06),
	.w8(32'h3b87a08f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68dd30),
	.w1(32'hbc3af95f),
	.w2(32'h38ff476e),
	.w3(32'hbbc6a089),
	.w4(32'hbc4aa45c),
	.w5(32'hbc885913),
	.w6(32'hbb932ff1),
	.w7(32'hba88642c),
	.w8(32'hbaba5016),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7717f7),
	.w1(32'hb8b66326),
	.w2(32'hbaec4202),
	.w3(32'hbae91d9c),
	.w4(32'hbabfb9dc),
	.w5(32'hbbaebdde),
	.w6(32'hbb07f770),
	.w7(32'h3a8625f9),
	.w8(32'hbbd8526a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1550ef),
	.w1(32'hbbe86d6d),
	.w2(32'hbc0c98d6),
	.w3(32'h3a032354),
	.w4(32'hb9004fc3),
	.w5(32'hbc08fb66),
	.w6(32'hbb7fe8ed),
	.w7(32'h3bd4da8d),
	.w8(32'h3a38bac5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5efc75),
	.w1(32'h3c1ed2f3),
	.w2(32'h3b08774d),
	.w3(32'h3bb3379d),
	.w4(32'h3c0ae921),
	.w5(32'h3b501a68),
	.w6(32'h3b3a2127),
	.w7(32'h3c832508),
	.w8(32'h3be64983),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d9253),
	.w1(32'hbb7852b5),
	.w2(32'hbb910f09),
	.w3(32'h3a80bc89),
	.w4(32'h3b0bb8aa),
	.w5(32'hbc382844),
	.w6(32'h3a11bce3),
	.w7(32'hbb9ceb1b),
	.w8(32'hbb0f4ce8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eeacf),
	.w1(32'h3b8d4664),
	.w2(32'hbb7ab1db),
	.w3(32'hbba2cbe7),
	.w4(32'h3b9ec42a),
	.w5(32'h3cadb34c),
	.w6(32'hbbaa7379),
	.w7(32'hbb3ed92b),
	.w8(32'h3b994263),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3622c5),
	.w1(32'hbb2c80d8),
	.w2(32'hbb67e0a7),
	.w3(32'hbb81bde0),
	.w4(32'h3aede9f4),
	.w5(32'hbb8cd3dd),
	.w6(32'h3c1f7711),
	.w7(32'hbb461fb8),
	.w8(32'hbb9e5897),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8603993),
	.w1(32'hbbf50439),
	.w2(32'hbc2b2f96),
	.w3(32'hbafe2101),
	.w4(32'hbb5e404b),
	.w5(32'h3bc1ca10),
	.w6(32'hbb207a65),
	.w7(32'hbc48d991),
	.w8(32'hbb078430),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58095),
	.w1(32'hbbb69c9a),
	.w2(32'hbbbe4f80),
	.w3(32'hbaeb68b2),
	.w4(32'hbbc32f8d),
	.w5(32'hbb84d934),
	.w6(32'hbbe57e36),
	.w7(32'hbb91bb53),
	.w8(32'hbba56e19),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2dd6),
	.w1(32'hbb892ec1),
	.w2(32'hb732683b),
	.w3(32'hbc13c956),
	.w4(32'hbbd9e66b),
	.w5(32'h3c51c1b5),
	.w6(32'hbc2d991d),
	.w7(32'hbb8b7b94),
	.w8(32'hba3741f1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38bb9a),
	.w1(32'h39cdfd5d),
	.w2(32'h3b04ec98),
	.w3(32'hbb665ab0),
	.w4(32'h3c13fc61),
	.w5(32'hbbd1f7c1),
	.w6(32'h3a8af052),
	.w7(32'h3b9cf369),
	.w8(32'h3aed23d1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b3b0a),
	.w1(32'hbb39b381),
	.w2(32'hbc3b6ce0),
	.w3(32'h3ab29dbe),
	.w4(32'hbb906718),
	.w5(32'h3baf5ec8),
	.w6(32'h3a9c255c),
	.w7(32'hbb8eedcb),
	.w8(32'hbabb65a9),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32cd9),
	.w1(32'hbb0f9753),
	.w2(32'hbbcc0db5),
	.w3(32'hbbb02e89),
	.w4(32'h3b38cd85),
	.w5(32'hbb57ccb1),
	.w6(32'hbad18633),
	.w7(32'hbb2c2687),
	.w8(32'h3b5c929b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2abef),
	.w1(32'hbb2ffc2d),
	.w2(32'hbb13cad0),
	.w3(32'hbb900228),
	.w4(32'h3b362add),
	.w5(32'hbc2faa0e),
	.w6(32'hba28be38),
	.w7(32'h3b082bfd),
	.w8(32'h3abfc471),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e731e),
	.w1(32'hbafc42c6),
	.w2(32'h3ab1d320),
	.w3(32'h3b84311c),
	.w4(32'h3a9d2792),
	.w5(32'hbc29baf1),
	.w6(32'h3ac6e975),
	.w7(32'h3be64b2f),
	.w8(32'h3bf42d99),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03fef0),
	.w1(32'hba085496),
	.w2(32'h39019b32),
	.w3(32'h3b0be77f),
	.w4(32'hb949e7f7),
	.w5(32'hbb2905ab),
	.w6(32'h3c09da5b),
	.w7(32'hbb25b298),
	.w8(32'hbb971d02),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab20555),
	.w1(32'h3a767723),
	.w2(32'hbc0fed36),
	.w3(32'h3a5d738e),
	.w4(32'h3a532e14),
	.w5(32'hbc265bed),
	.w6(32'hbb181480),
	.w7(32'hbb554866),
	.w8(32'hbc1ccc71),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb45810),
	.w1(32'hba221d68),
	.w2(32'h3b712d3a),
	.w3(32'hbb40fe30),
	.w4(32'hbba3a1c1),
	.w5(32'h3b12d217),
	.w6(32'hbbdc5487),
	.w7(32'h3b98da3a),
	.w8(32'hbbd0b26a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eeca7),
	.w1(32'hbb3e8a5a),
	.w2(32'hbc36a260),
	.w3(32'h3b51753b),
	.w4(32'h3b8ad319),
	.w5(32'hbaf8e1a9),
	.w6(32'hbb8d326c),
	.w7(32'h3b862ecc),
	.w8(32'hba45ce91),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9aee),
	.w1(32'hbbcca8b7),
	.w2(32'hbbbe2435),
	.w3(32'hbb0d61f7),
	.w4(32'h3b4a007c),
	.w5(32'hbc3fe6cc),
	.w6(32'hbb406b74),
	.w7(32'h3b4c2964),
	.w8(32'h3b08b8a7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54207a),
	.w1(32'h3b0492e9),
	.w2(32'hb995aaf7),
	.w3(32'hbc25c9b8),
	.w4(32'hbb876617),
	.w5(32'h3cb58436),
	.w6(32'hbc104cbf),
	.w7(32'hba9de3a8),
	.w8(32'hbb129637),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2998aa),
	.w1(32'hbb92b257),
	.w2(32'hbbb82010),
	.w3(32'hbb0ba3f5),
	.w4(32'hbb3acaf2),
	.w5(32'h3ae27b2e),
	.w6(32'h3b4626f2),
	.w7(32'hba813c97),
	.w8(32'hbb2a7f78),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdb06f),
	.w1(32'h39ec6518),
	.w2(32'hbb7218d9),
	.w3(32'hbb6cefba),
	.w4(32'h3b925d1b),
	.w5(32'hba56a8fe),
	.w6(32'hbb22e924),
	.w7(32'h3ba1d944),
	.w8(32'hb8a38b52),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b57f),
	.w1(32'h3bad5ddc),
	.w2(32'h39d02605),
	.w3(32'hbb89c0c0),
	.w4(32'h3b097e13),
	.w5(32'h39ea8918),
	.w6(32'h3b123d94),
	.w7(32'h3a134298),
	.w8(32'hbc04f0a5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfeae9),
	.w1(32'h3ae34153),
	.w2(32'hbb933cf6),
	.w3(32'h3a910c44),
	.w4(32'h3a1b6ee4),
	.w5(32'h3c57db1a),
	.w6(32'hbc086d87),
	.w7(32'hbc4b3a46),
	.w8(32'h3b9a7d53),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc208b7c),
	.w1(32'hb8ddce6a),
	.w2(32'h3b2d7464),
	.w3(32'hb9bf7e7e),
	.w4(32'h3b5dba4d),
	.w5(32'hbb0783f5),
	.w6(32'h3b9903a4),
	.w7(32'h3b0bb472),
	.w8(32'hbbf1f7e0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5062fb),
	.w1(32'hbbb92310),
	.w2(32'h3aa45675),
	.w3(32'h3be2346d),
	.w4(32'hbb6cfcc8),
	.w5(32'hbb8308c1),
	.w6(32'hb8973f1f),
	.w7(32'h3b0d396a),
	.w8(32'h3b457c3b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a24f),
	.w1(32'hbb96431c),
	.w2(32'hb8507a5a),
	.w3(32'h3b96638a),
	.w4(32'hbbf5d66d),
	.w5(32'hbc2112f1),
	.w6(32'hbb9e6bf4),
	.w7(32'hbbb1abfd),
	.w8(32'hbb8b6551),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82834c),
	.w1(32'hbbf74d8c),
	.w2(32'hbba6bccd),
	.w3(32'hbbae8c41),
	.w4(32'hbbff7461),
	.w5(32'hbbc276fe),
	.w6(32'hbbc04237),
	.w7(32'hba05f700),
	.w8(32'h3ad16088),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03d53),
	.w1(32'h3aa8a75f),
	.w2(32'hba0e2884),
	.w3(32'hbb84ad29),
	.w4(32'h3b4a73d6),
	.w5(32'hbc2d02c6),
	.w6(32'hbb8d267d),
	.w7(32'h3b3ad093),
	.w8(32'h3c1aabfc),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfa169),
	.w1(32'h3a5a5c2f),
	.w2(32'hbb4c94b9),
	.w3(32'hbb8d6f52),
	.w4(32'h3bdb08a8),
	.w5(32'hbb6c81d9),
	.w6(32'hba1e524c),
	.w7(32'hba0303e0),
	.w8(32'hbbbb9a3a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe444),
	.w1(32'hbbbf43b9),
	.w2(32'h3bb01536),
	.w3(32'hbb2a9d03),
	.w4(32'hbc188f78),
	.w5(32'h3c704deb),
	.w6(32'hbc023b52),
	.w7(32'hbb9a0a3d),
	.w8(32'h39eb7e06),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7779b6),
	.w1(32'h3adb9bf6),
	.w2(32'h3c0399be),
	.w3(32'h3b8d6edd),
	.w4(32'h3b7edfef),
	.w5(32'hbc3acc5a),
	.w6(32'h3c117442),
	.w7(32'h3c0e3410),
	.w8(32'h3a73641a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c3afd),
	.w1(32'hbc0e2acc),
	.w2(32'hbb3cb39d),
	.w3(32'h3c22b1a7),
	.w4(32'hbb67e1e0),
	.w5(32'hbc27675a),
	.w6(32'h3c13d60b),
	.w7(32'hbb27b537),
	.w8(32'h3ad0ee59),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4db683),
	.w1(32'hbad38ebf),
	.w2(32'hb98feade),
	.w3(32'hbc358136),
	.w4(32'hba794f90),
	.w5(32'hbc280a4c),
	.w6(32'hbc2021db),
	.w7(32'h3b0db885),
	.w8(32'hbba5d551),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb518184),
	.w1(32'hbc489a07),
	.w2(32'h3b73eee1),
	.w3(32'hba3b9fc6),
	.w4(32'hbc76d84c),
	.w5(32'hbbf0ef35),
	.w6(32'h3bb7c1e4),
	.w7(32'hbb818301),
	.w8(32'hbb628e82),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb15533),
	.w1(32'hbba7d5b6),
	.w2(32'hbba24b31),
	.w3(32'hbc0a629e),
	.w4(32'h39de02b4),
	.w5(32'hbc5ae725),
	.w6(32'hbc0a4892),
	.w7(32'h3b9e1ec6),
	.w8(32'hbabcce32),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f52ad),
	.w1(32'hbaa43b1a),
	.w2(32'hbb55b061),
	.w3(32'h3bd5ba6b),
	.w4(32'h3c24af91),
	.w5(32'hbb9ccd7d),
	.w6(32'hbb700b67),
	.w7(32'h3c285e40),
	.w8(32'h3bdb2a5a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d2dd0),
	.w1(32'hbbc3b262),
	.w2(32'hbb48a50e),
	.w3(32'hbb2ed110),
	.w4(32'h3b9d37f7),
	.w5(32'h3a3f8c2e),
	.w6(32'hbb119f5c),
	.w7(32'h3bf28d1f),
	.w8(32'hbb093d1c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4779be),
	.w1(32'h3b3f9017),
	.w2(32'h3b1b79d9),
	.w3(32'hbb4bc822),
	.w4(32'h3bb1fc16),
	.w5(32'hba4898b4),
	.w6(32'hbc025819),
	.w7(32'h3bbe0de0),
	.w8(32'hb9a0e4b6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef63ab),
	.w1(32'h3b6c0901),
	.w2(32'hbb29c859),
	.w3(32'hbb5add1c),
	.w4(32'h3bbb828e),
	.w5(32'hbbc591ed),
	.w6(32'hbbfd1ea8),
	.w7(32'hbadb4884),
	.w8(32'h3a07c416),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cc2f0),
	.w1(32'h3a9a1647),
	.w2(32'hbbb3a6a0),
	.w3(32'hba472faa),
	.w4(32'hba8c448e),
	.w5(32'hbbbd273d),
	.w6(32'hb9689962),
	.w7(32'h389778ec),
	.w8(32'hbaf472a8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3717),
	.w1(32'h3c2cf024),
	.w2(32'hba54902b),
	.w3(32'hbbd96d10),
	.w4(32'h3b17338a),
	.w5(32'h3c56c3d3),
	.w6(32'h3b91d698),
	.w7(32'hbb95533b),
	.w8(32'h3b1775c8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07aecf),
	.w1(32'hbb8a4560),
	.w2(32'h3b848997),
	.w3(32'h3b29e3bd),
	.w4(32'hbc173d38),
	.w5(32'h3b019b90),
	.w6(32'h3bad6117),
	.w7(32'h3aac9d41),
	.w8(32'hbbae9914),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25909e),
	.w1(32'h3ace746f),
	.w2(32'hbb481bc8),
	.w3(32'h3c12a083),
	.w4(32'h3bc4ac2f),
	.w5(32'hb89815fa),
	.w6(32'h3acb2c8c),
	.w7(32'h3c1c4dba),
	.w8(32'h3c21089a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5d2f),
	.w1(32'h3ad030eb),
	.w2(32'h3b46d7a5),
	.w3(32'hbaa7e357),
	.w4(32'hbb99017c),
	.w5(32'h3cb0fdab),
	.w6(32'hbb8500d5),
	.w7(32'hbba52b8b),
	.w8(32'h3b3a897a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b3607),
	.w1(32'hbbec8b34),
	.w2(32'hbc04b3ce),
	.w3(32'h3b20385a),
	.w4(32'h3a33f91e),
	.w5(32'hbc8a76f6),
	.w6(32'h3b3ccb58),
	.w7(32'h3b526e5a),
	.w8(32'hbc0f04d3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306a7f),
	.w1(32'h3afdf95f),
	.w2(32'hbbd6d9fe),
	.w3(32'h3aecc11b),
	.w4(32'h3b7e846e),
	.w5(32'hbaf37087),
	.w6(32'hbbe1c099),
	.w7(32'hbb93dd97),
	.w8(32'hbb5b87cd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b575d91),
	.w1(32'h3b19b09e),
	.w2(32'hbb04497e),
	.w3(32'hbb1c18aa),
	.w4(32'h3c168d93),
	.w5(32'hba692d9e),
	.w6(32'h382a8e96),
	.w7(32'h3bafe33a),
	.w8(32'h3aba850f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba25bc5),
	.w1(32'h3a47f974),
	.w2(32'h3a86ab37),
	.w3(32'h3b75c40d),
	.w4(32'h3bad4c73),
	.w5(32'hbb54b9ce),
	.w6(32'h3b4a1aa4),
	.w7(32'h3a8f166e),
	.w8(32'hbbc4e135),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e91b2a),
	.w1(32'hbb592c7e),
	.w2(32'hbc013478),
	.w3(32'hbb202ff5),
	.w4(32'h3b80c40d),
	.w5(32'hbc5deba8),
	.w6(32'hbbcdd9ce),
	.w7(32'hbabc23ee),
	.w8(32'hbc44f67c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f60ed),
	.w1(32'h39959b96),
	.w2(32'h3bae0f41),
	.w3(32'h3ba6f06b),
	.w4(32'hbb7784e0),
	.w5(32'hbb878b77),
	.w6(32'hbbb5b1c1),
	.w7(32'h3ae89219),
	.w8(32'hbb07aab4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcc202),
	.w1(32'h3b09d90d),
	.w2(32'hbb8b6403),
	.w3(32'hbb317125),
	.w4(32'h3b97aed8),
	.w5(32'h3bc207ab),
	.w6(32'hbaf5eda6),
	.w7(32'h3b3acb96),
	.w8(32'h3a8bb143),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc02c0a),
	.w1(32'hba9830d7),
	.w2(32'h3c54c998),
	.w3(32'hbb853e3a),
	.w4(32'hbc4edb17),
	.w5(32'h3bb33738),
	.w6(32'h3903419b),
	.w7(32'hbbcfbff0),
	.w8(32'hbb2e1dfd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01ca56),
	.w1(32'hbb463fce),
	.w2(32'h3add68ae),
	.w3(32'hba025c29),
	.w4(32'hbbe2ff79),
	.w5(32'h3b149235),
	.w6(32'h3b006777),
	.w7(32'hbc09bdee),
	.w8(32'hbafcb81c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b2d7f),
	.w1(32'h3aacbe7b),
	.w2(32'hbb47d14c),
	.w3(32'hbbeda7c3),
	.w4(32'hbac9dd5f),
	.w5(32'h3a80725b),
	.w6(32'hbaa1cca5),
	.w7(32'h3b5e7d97),
	.w8(32'h3b5c1be0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0db488),
	.w1(32'h3ac1e4f6),
	.w2(32'hbb892086),
	.w3(32'hbc139f8f),
	.w4(32'h3babcb1f),
	.w5(32'hbb995997),
	.w6(32'hbb45c577),
	.w7(32'h3b5d626d),
	.w8(32'h3b99f542),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675f07),
	.w1(32'h3b5c8c2d),
	.w2(32'hbb935f57),
	.w3(32'h380dd848),
	.w4(32'hbb17fc6d),
	.w5(32'h3bc38943),
	.w6(32'h3b8c3121),
	.w7(32'hbbc47007),
	.w8(32'h3b77364a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dd022),
	.w1(32'h3b1ea9dd),
	.w2(32'h3bdddb63),
	.w3(32'hbc0308eb),
	.w4(32'hbb831af8),
	.w5(32'h3c6b38b3),
	.w6(32'h3bca1246),
	.w7(32'hbb0375a8),
	.w8(32'h3b8d5861),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4b6c7),
	.w1(32'h3bc86f78),
	.w2(32'h3bf4cb60),
	.w3(32'hbc05b6c8),
	.w4(32'h3bf82cbe),
	.w5(32'hbc14ef43),
	.w6(32'hbc360966),
	.w7(32'h3ba20c42),
	.w8(32'hbaeef5a3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba104d5),
	.w1(32'h3b9c040c),
	.w2(32'h3c3000c5),
	.w3(32'h3c2a0606),
	.w4(32'hbab23e92),
	.w5(32'h3bf0a53f),
	.w6(32'h3b8506a7),
	.w7(32'hbb31ce01),
	.w8(32'hba0d47e5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ffab7),
	.w1(32'hbbc5d7c2),
	.w2(32'h3b3724e5),
	.w3(32'h39736e3f),
	.w4(32'hba82defe),
	.w5(32'hbbff7569),
	.w6(32'h3b2a44f9),
	.w7(32'h3b4a038a),
	.w8(32'hbc0e5f11),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf106a8),
	.w1(32'hbb00e143),
	.w2(32'hbaa1371c),
	.w3(32'hbaa504f0),
	.w4(32'hb9cbc76d),
	.w5(32'h3acfa67f),
	.w6(32'hbb9a4709),
	.w7(32'hbac032e5),
	.w8(32'hbb356304),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a15f),
	.w1(32'hbb95f4ff),
	.w2(32'hbb4f10c4),
	.w3(32'h3b352120),
	.w4(32'h3a616a97),
	.w5(32'h39ad62c9),
	.w6(32'hbbe4d6b4),
	.w7(32'h3a0cf0df),
	.w8(32'h3b4761c5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820b2a),
	.w1(32'hbafc9b8d),
	.w2(32'hbb7594d8),
	.w3(32'hbab94ebd),
	.w4(32'h3b332105),
	.w5(32'hbb79051a),
	.w6(32'h3ac0194a),
	.w7(32'hbc236dbc),
	.w8(32'hba37e75d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc44ab),
	.w1(32'hbc3d6dff),
	.w2(32'hbc488483),
	.w3(32'hbbe1f830),
	.w4(32'hbb822023),
	.w5(32'hbc7f2193),
	.w6(32'hbc5fd83b),
	.w7(32'hbb45cfb8),
	.w8(32'hbc10525e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14dd90),
	.w1(32'h3c065326),
	.w2(32'h3ba4e398),
	.w3(32'hbc604b91),
	.w4(32'hbb98132d),
	.w5(32'h3caedfe4),
	.w6(32'hbc201f6a),
	.w7(32'hbb4b5fd3),
	.w8(32'hbc01e9b9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1f90),
	.w1(32'hbb70ab54),
	.w2(32'hbc34d31f),
	.w3(32'h3c90acbe),
	.w4(32'hba5a235d),
	.w5(32'hbc4ad62f),
	.w6(32'h3c47393a),
	.w7(32'h396e0d5e),
	.w8(32'h3ac407ea),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6283ff),
	.w1(32'hbbe3914f),
	.w2(32'hbb6f2b4e),
	.w3(32'hbc39c042),
	.w4(32'hb9d33204),
	.w5(32'hbbaa4b6c),
	.w6(32'h3965b09a),
	.w7(32'h3bac7da2),
	.w8(32'hbbe4fc74),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7811a8),
	.w1(32'hbb329c98),
	.w2(32'h3bb3275c),
	.w3(32'h3b39e815),
	.w4(32'hbbce14cd),
	.w5(32'h3bc8049a),
	.w6(32'hbb2e21f7),
	.w7(32'hbbf3340a),
	.w8(32'hbad0754a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acce109),
	.w1(32'hbad3fe58),
	.w2(32'hb9b30cfb),
	.w3(32'h3b3988d3),
	.w4(32'h3bd31575),
	.w5(32'h3c260b7d),
	.w6(32'h3a61b3ed),
	.w7(32'hb95954e3),
	.w8(32'h3b96f198),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2217),
	.w1(32'hbb503aed),
	.w2(32'hbb81668a),
	.w3(32'h3848055f),
	.w4(32'h3b04b4f1),
	.w5(32'hbb9bc139),
	.w6(32'h3b5b270b),
	.w7(32'hbad67e3e),
	.w8(32'h397e9e2a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1027a6),
	.w1(32'h3b5331bf),
	.w2(32'h3a2258d4),
	.w3(32'h3c052c95),
	.w4(32'hbb1bf0b4),
	.w5(32'h3c061d78),
	.w6(32'h3bc11ef0),
	.w7(32'h3b4f3707),
	.w8(32'hbae0575a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93239f),
	.w1(32'h3abd47b2),
	.w2(32'hbb82a05f),
	.w3(32'hb91f23e9),
	.w4(32'hbabbf3d1),
	.w5(32'hbaa8f779),
	.w6(32'hba494390),
	.w7(32'hbbecf562),
	.w8(32'hbb2ad9ab),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994d40),
	.w1(32'h39e27186),
	.w2(32'hbb13415a),
	.w3(32'hbbb1b05a),
	.w4(32'hbb7da277),
	.w5(32'hbb8a8acb),
	.w6(32'h3a0aa26b),
	.w7(32'hba1c56d5),
	.w8(32'hbb02ea15),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928bf6),
	.w1(32'h3b85a1ab),
	.w2(32'h3b7ff259),
	.w3(32'hbbba0a6d),
	.w4(32'hbc06806f),
	.w5(32'h3bfadeaf),
	.w6(32'h38837ac4),
	.w7(32'hbc3cdb73),
	.w8(32'h3bead662),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95b620),
	.w1(32'h3c5dce76),
	.w2(32'h3bd6530b),
	.w3(32'hbb65e992),
	.w4(32'hbb06bece),
	.w5(32'h3ad96643),
	.w6(32'hba835a66),
	.w7(32'hbc80f489),
	.w8(32'h3c418195),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c053),
	.w1(32'hbc7f21e9),
	.w2(32'hbcb3498a),
	.w3(32'hba5eb2d5),
	.w4(32'hbbeef3b6),
	.w5(32'hbb2a43b9),
	.w6(32'h3b1f5858),
	.w7(32'hbb91b3b6),
	.w8(32'h3b616c3e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84521f),
	.w1(32'hba9da856),
	.w2(32'h3ba396af),
	.w3(32'hba0b255a),
	.w4(32'hbb9e01cb),
	.w5(32'hbbf63d6f),
	.w6(32'hbaedf13a),
	.w7(32'h3bffa169),
	.w8(32'h3cba0121),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa9fb6),
	.w1(32'h3b4201e4),
	.w2(32'hbc990ee1),
	.w3(32'h39c3efd5),
	.w4(32'hbbbf250b),
	.w5(32'hbc22c30f),
	.w6(32'h3bc49a45),
	.w7(32'hbca79923),
	.w8(32'h39187f70),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92894f),
	.w1(32'hba3ccdc8),
	.w2(32'h3b20b389),
	.w3(32'h3b42c5cd),
	.w4(32'h39cda275),
	.w5(32'hba69b03f),
	.w6(32'h3c948217),
	.w7(32'h3c0286a3),
	.w8(32'hbb354a6c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c53d0),
	.w1(32'hbbe574e2),
	.w2(32'hbbc91f8c),
	.w3(32'hbbfc4010),
	.w4(32'hbc8d24b2),
	.w5(32'hbc8f1167),
	.w6(32'hbb0b903d),
	.w7(32'hbb5a7ce0),
	.w8(32'hbc3c7f6b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a54c),
	.w1(32'hbc646531),
	.w2(32'hbc77894e),
	.w3(32'hbc1b3a6d),
	.w4(32'hba033006),
	.w5(32'h3b63da4c),
	.w6(32'hbbb6fff5),
	.w7(32'hbaf479b2),
	.w8(32'h3baaf30d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c71c7),
	.w1(32'hba30eb06),
	.w2(32'hba571938),
	.w3(32'hbb464582),
	.w4(32'hbb8cdb83),
	.w5(32'hbaad05ef),
	.w6(32'h3a21e081),
	.w7(32'hbafbd138),
	.w8(32'h38c60f7b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7adf40),
	.w1(32'h3bc8297b),
	.w2(32'h3b19c10b),
	.w3(32'hbb3aedca),
	.w4(32'h3b0392be),
	.w5(32'hbb8fbe99),
	.w6(32'h3b499084),
	.w7(32'h3c1e6081),
	.w8(32'h3c40e2e3),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eb0bc),
	.w1(32'hbb489c2c),
	.w2(32'hbb9ceb82),
	.w3(32'hba953f08),
	.w4(32'hbba16057),
	.w5(32'hbb93564a),
	.w6(32'h3adb3edc),
	.w7(32'hbbaefc9d),
	.w8(32'hbb75e2da),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cf43b),
	.w1(32'hbc107b8e),
	.w2(32'hbb239e8b),
	.w3(32'hbb0c3d66),
	.w4(32'h3a90f367),
	.w5(32'hbb24b103),
	.w6(32'h3afe35b9),
	.w7(32'hbb0516b3),
	.w8(32'hba454f90),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39d697),
	.w1(32'h3cd857ee),
	.w2(32'h3d00432e),
	.w3(32'hbbae54ce),
	.w4(32'h3bc8d83d),
	.w5(32'h3b547955),
	.w6(32'hbbc97c55),
	.w7(32'hbca7a553),
	.w8(32'hbcc1f9f7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951466),
	.w1(32'h3ad5f635),
	.w2(32'h3bb5e47c),
	.w3(32'hba81e7f9),
	.w4(32'h370751be),
	.w5(32'h3bd452ca),
	.w6(32'hbc7747c5),
	.w7(32'hbc009e93),
	.w8(32'h3af8426f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205497),
	.w1(32'hb9ce8f98),
	.w2(32'hbc14d1d7),
	.w3(32'hba705346),
	.w4(32'h3b1d44b1),
	.w5(32'hbb9a61f1),
	.w6(32'hba2657f6),
	.w7(32'h3a8c800d),
	.w8(32'hbae67515),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc215a4b),
	.w1(32'hba228561),
	.w2(32'hbb9e48a0),
	.w3(32'hbb109248),
	.w4(32'hbba20d86),
	.w5(32'hbb6caf4a),
	.w6(32'hbad07f3a),
	.w7(32'hbbc70058),
	.w8(32'hbaaef648),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9b8b6),
	.w1(32'h3ae80140),
	.w2(32'hbba32775),
	.w3(32'hbb2099a9),
	.w4(32'h39ed5cbe),
	.w5(32'hba6c55e7),
	.w6(32'hbbc4b834),
	.w7(32'hba08e761),
	.w8(32'h3c0f352c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87f846),
	.w1(32'h3bf16445),
	.w2(32'h3aa053ce),
	.w3(32'hbb182137),
	.w4(32'h3ab3248e),
	.w5(32'h3ab98e42),
	.w6(32'h3c276117),
	.w7(32'h3ba3118c),
	.w8(32'hbbbfc010),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25227),
	.w1(32'hbbb2d3d5),
	.w2(32'hbc0b6a27),
	.w3(32'h3c22d6bc),
	.w4(32'hbbb0ded6),
	.w5(32'h3b63afd2),
	.w6(32'hbb05b098),
	.w7(32'h3ba3d75d),
	.w8(32'h3abe570d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bac25),
	.w1(32'h3c56004e),
	.w2(32'h39f5ff80),
	.w3(32'hbb843448),
	.w4(32'hbb1a7726),
	.w5(32'h3a9be87d),
	.w6(32'hbab794a0),
	.w7(32'h3be7ae1b),
	.w8(32'hba03bcf4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76db99),
	.w1(32'hbb7db033),
	.w2(32'hbc4d0927),
	.w3(32'hbc2b9313),
	.w4(32'h39af6aee),
	.w5(32'hba3b73a7),
	.w6(32'hbbf6edf0),
	.w7(32'h3b859ed8),
	.w8(32'h3bd1edc4),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51ad80),
	.w1(32'hbbb79c71),
	.w2(32'h3a7f5f3a),
	.w3(32'hbb92a710),
	.w4(32'hbb7ad5e1),
	.w5(32'hbb342312),
	.w6(32'h3a09a2d0),
	.w7(32'hbb929709),
	.w8(32'hbc364835),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9cdb8),
	.w1(32'hbaf09103),
	.w2(32'hbc5b4732),
	.w3(32'hbc004880),
	.w4(32'hb90d2ae8),
	.w5(32'h3aae31d7),
	.w6(32'hbc52acd1),
	.w7(32'h3b2941f7),
	.w8(32'h3bf3dedd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c275c),
	.w1(32'hbc5e3272),
	.w2(32'hbb7f6e23),
	.w3(32'hbbd7e119),
	.w4(32'hbb82bf02),
	.w5(32'hbc18fde7),
	.w6(32'h3be597fd),
	.w7(32'h3b84105c),
	.w8(32'hbbd88ef8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d6fdc),
	.w1(32'h3c365517),
	.w2(32'h3c32bfa0),
	.w3(32'hbc04b1e7),
	.w4(32'h3be137d7),
	.w5(32'h3bd18480),
	.w6(32'h3a718c34),
	.w7(32'hbc4d6430),
	.w8(32'hbc6c5827),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0c948),
	.w1(32'h3b358f2e),
	.w2(32'h3bb18ffa),
	.w3(32'hbb469abb),
	.w4(32'h3a2c9b83),
	.w5(32'h3c83ee39),
	.w6(32'hbc0c2a3a),
	.w7(32'hbbfd60d5),
	.w8(32'hbc04a292),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d7b1d),
	.w1(32'hbc010de7),
	.w2(32'hbc0b4efa),
	.w3(32'h3b3ac1fe),
	.w4(32'hbbaf556a),
	.w5(32'hbbc0a489),
	.w6(32'hbba38ff7),
	.w7(32'hbb810d32),
	.w8(32'hbc0caf86),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe66e75),
	.w1(32'h3b97895e),
	.w2(32'hbb301525),
	.w3(32'hbbcbd75d),
	.w4(32'hbb9c5289),
	.w5(32'hbbe92c56),
	.w6(32'hbc0d9e04),
	.w7(32'h3b8b015b),
	.w8(32'h3b5d90ed),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67d9cb),
	.w1(32'hb888264b),
	.w2(32'hbac714a5),
	.w3(32'h3b28f9ce),
	.w4(32'hbaf085a5),
	.w5(32'h3b1d7576),
	.w6(32'h3a949f87),
	.w7(32'h3ba8873e),
	.w8(32'h3bd833f1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc92294),
	.w1(32'hbc6b879e),
	.w2(32'hbb29cc53),
	.w3(32'hbb724234),
	.w4(32'hbb63c8f9),
	.w5(32'h3a764ea3),
	.w6(32'h3b480ca5),
	.w7(32'hb84693d6),
	.w8(32'h382194fa),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c5cdc),
	.w1(32'hbbca73a5),
	.w2(32'hbad9d142),
	.w3(32'hbb7f379e),
	.w4(32'hbb80b498),
	.w5(32'h3b8a3093),
	.w6(32'hbc981409),
	.w7(32'hbc4c61c1),
	.w8(32'hbc82f99e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc810da2),
	.w1(32'hbc1585d0),
	.w2(32'h3ac56d29),
	.w3(32'hbba56cd0),
	.w4(32'hbc169cb6),
	.w5(32'hbc26eba9),
	.w6(32'hbbba7793),
	.w7(32'hbbfadce0),
	.w8(32'hbc4c0e87),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30348),
	.w1(32'hbc16d8f0),
	.w2(32'hbc51b297),
	.w3(32'hbc11a4bd),
	.w4(32'hbc18dd76),
	.w5(32'hbc111a21),
	.w6(32'hbc73c5a4),
	.w7(32'hbb186691),
	.w8(32'hbc40f541),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f4aa),
	.w1(32'hbb6a9f14),
	.w2(32'hbb6b5e03),
	.w3(32'hbc06982d),
	.w4(32'hbb857c07),
	.w5(32'h3a8a3fa2),
	.w6(32'hbbda8b56),
	.w7(32'hbba96851),
	.w8(32'hbafbfb31),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7336),
	.w1(32'h3bed3592),
	.w2(32'h3a08e267),
	.w3(32'h3b830e77),
	.w4(32'hbb3d339e),
	.w5(32'hbb98fa5a),
	.w6(32'h3afc78ee),
	.w7(32'hbb1f435f),
	.w8(32'h3793794f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0940),
	.w1(32'hbb5fe942),
	.w2(32'hbb6e49fc),
	.w3(32'hba16991c),
	.w4(32'h3a70ff66),
	.w5(32'hbb9d14ae),
	.w6(32'h3b44236c),
	.w7(32'h3b4133cd),
	.w8(32'h3a23b076),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eb9f1),
	.w1(32'hbb922a0c),
	.w2(32'hbc74125b),
	.w3(32'h3abb4ac6),
	.w4(32'hbb816a99),
	.w5(32'hbc30f440),
	.w6(32'h3b9c3535),
	.w7(32'hbb9ee5fc),
	.w8(32'hbbb00635),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc9d7b),
	.w1(32'h3a3e4c9d),
	.w2(32'hba927067),
	.w3(32'hbaf0991e),
	.w4(32'hba26ddf3),
	.w5(32'h3b812a0b),
	.w6(32'hbb61294e),
	.w7(32'hbb09e11b),
	.w8(32'hbaa1303e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9769e),
	.w1(32'hbacfe05d),
	.w2(32'hbb728097),
	.w3(32'hbadbfca3),
	.w4(32'h3bc18649),
	.w5(32'h3adeb0e1),
	.w6(32'h39d2cc2a),
	.w7(32'h3b60e464),
	.w8(32'hb9534d01),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8195cc),
	.w1(32'h3c90ad06),
	.w2(32'h3b23c164),
	.w3(32'hbac0a59c),
	.w4(32'h3ca068e9),
	.w5(32'h37f4ff6b),
	.w6(32'hbbc8c6b9),
	.w7(32'h3c81f220),
	.w8(32'hba0c9bae),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae847ef),
	.w1(32'hbc355c7b),
	.w2(32'hbc629d8f),
	.w3(32'hbbc97915),
	.w4(32'hbc239575),
	.w5(32'hbc7f6545),
	.w6(32'h3be654bf),
	.w7(32'hbc6c0651),
	.w8(32'hbc8a29c5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375430),
	.w1(32'h3bcd0813),
	.w2(32'hbbfaa9ad),
	.w3(32'hbc3e0bf0),
	.w4(32'h3a3c5411),
	.w5(32'hbbc2bb95),
	.w6(32'hbc33313f),
	.w7(32'h3b75900c),
	.w8(32'hba8021dc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e923b),
	.w1(32'hbc7eb1b8),
	.w2(32'hbafeecd1),
	.w3(32'hbb83e8a2),
	.w4(32'h3b384197),
	.w5(32'h38bf3cdd),
	.w6(32'hbb5546cb),
	.w7(32'h3b9ec54e),
	.w8(32'hbb9e7626),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fb0e3),
	.w1(32'hbbc45b16),
	.w2(32'hbbc380d0),
	.w3(32'hba089547),
	.w4(32'hba884a12),
	.w5(32'hbb31a1c8),
	.w6(32'h3b54096f),
	.w7(32'h3b19653c),
	.w8(32'h3be9ed28),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43e7ac),
	.w1(32'hbb8edc91),
	.w2(32'hbc28943a),
	.w3(32'hb95640fd),
	.w4(32'hba095c0e),
	.w5(32'hbc12f1dc),
	.w6(32'h3a885f20),
	.w7(32'h3a8597e9),
	.w8(32'hbbb14471),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28afd),
	.w1(32'h3b6c9467),
	.w2(32'h393214e4),
	.w3(32'hbbcf5b52),
	.w4(32'h39093bd3),
	.w5(32'hbbf6d6b7),
	.w6(32'hbada072a),
	.w7(32'h3aceb438),
	.w8(32'h3c37f958),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2357),
	.w1(32'h3b055a47),
	.w2(32'h3b699588),
	.w3(32'hbb20e051),
	.w4(32'h3a2b8e99),
	.w5(32'hba40f882),
	.w6(32'h3b5335d3),
	.w7(32'hbbe51add),
	.w8(32'hbc78b355),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8e5ca),
	.w1(32'hbb8c8bd3),
	.w2(32'h3b93097f),
	.w3(32'hbb95e939),
	.w4(32'hbb52819b),
	.w5(32'h3b2de1f4),
	.w6(32'hbc1b8c6f),
	.w7(32'h3abe9b2b),
	.w8(32'h3b32e078),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99e9a1),
	.w1(32'hba18318f),
	.w2(32'hbb857bd9),
	.w3(32'h3b3c9640),
	.w4(32'h3ad477de),
	.w5(32'h3ab022e5),
	.w6(32'h3c1304d0),
	.w7(32'hbb92b84a),
	.w8(32'h3ab08f2b),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ac995),
	.w1(32'hba8b74a8),
	.w2(32'h3bb0ab7e),
	.w3(32'hba9fc2d9),
	.w4(32'h3bfa660d),
	.w5(32'h3c85ef53),
	.w6(32'h3a765923),
	.w7(32'h3c092535),
	.w8(32'h3c053822),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61b5a2),
	.w1(32'hbb92fa65),
	.w2(32'h3b416de6),
	.w3(32'hbaf3ac54),
	.w4(32'hbc18203e),
	.w5(32'hbc82bb28),
	.w6(32'hbb21eb15),
	.w7(32'h3a0a012e),
	.w8(32'hbb648f70),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c2e61),
	.w1(32'hbac5f2ae),
	.w2(32'hbb8bd724),
	.w3(32'hbb97534d),
	.w4(32'h3b5f846a),
	.w5(32'hbb722628),
	.w6(32'h3b158af1),
	.w7(32'h3b89d5d9),
	.w8(32'h3afc5b17),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1afc16),
	.w1(32'h3a93b207),
	.w2(32'hbbd0fdb9),
	.w3(32'h39f37b26),
	.w4(32'h39de2da1),
	.w5(32'h3b8f0e59),
	.w6(32'h3c0cb317),
	.w7(32'hba8ff00e),
	.w8(32'hbb6a322a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf03858),
	.w1(32'hbb8586d7),
	.w2(32'h3bc37fa8),
	.w3(32'hbba1af64),
	.w4(32'h3a8a3ee2),
	.w5(32'hbb9febea),
	.w6(32'hbb992acd),
	.w7(32'hbc743744),
	.w8(32'hbb9b2532),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea69b8),
	.w1(32'hbb28fa3c),
	.w2(32'hbc18daca),
	.w3(32'hbbadc797),
	.w4(32'hbab98642),
	.w5(32'h3a058bae),
	.w6(32'hbb022ce8),
	.w7(32'h3ad9c9fa),
	.w8(32'h3b7b90a9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb08cc6),
	.w1(32'h3b780fe6),
	.w2(32'hbb662b0d),
	.w3(32'hbb59d48b),
	.w4(32'h3b0ce740),
	.w5(32'hb58c5ca7),
	.w6(32'hbb45d6b6),
	.w7(32'hbbc80fcf),
	.w8(32'hbba12975),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82aff7),
	.w1(32'h3bb7a991),
	.w2(32'h3a39594d),
	.w3(32'hbb654cb1),
	.w4(32'hb916bedf),
	.w5(32'hbc090b21),
	.w6(32'hbbc6725d),
	.w7(32'h3bed49ad),
	.w8(32'h3bf1a1a1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183bdd),
	.w1(32'h3b79ba20),
	.w2(32'h3b15ace1),
	.w3(32'hbbed696f),
	.w4(32'hb9f42e7f),
	.w5(32'hbaefb9df),
	.w6(32'hbb87e2c0),
	.w7(32'hb86af68c),
	.w8(32'hbb833117),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1665bf),
	.w1(32'hbb3cf80c),
	.w2(32'hbbba5954),
	.w3(32'hbb0b6441),
	.w4(32'hbbba33de),
	.w5(32'hbbd72469),
	.w6(32'hbb8f9aa1),
	.w7(32'h3b98ddcc),
	.w8(32'h3bdaec22),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2983c7),
	.w1(32'hbb4758e7),
	.w2(32'hbb9e6048),
	.w3(32'hbc263202),
	.w4(32'hbbe79a5a),
	.w5(32'hbb1b1790),
	.w6(32'h3accbf22),
	.w7(32'hbb9add3a),
	.w8(32'hbb98cae2),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule