module layer_10_featuremap_200(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99eee04),
	.w1(32'h3a2e2d02),
	.w2(32'h3ab538af),
	.w3(32'hb98269fd),
	.w4(32'hb903b608),
	.w5(32'hb89f1a5f),
	.w6(32'hbaeb76be),
	.w7(32'hbad27f63),
	.w8(32'hb9ecefa8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3900b),
	.w1(32'h3aa07f97),
	.w2(32'h3a771519),
	.w3(32'h3a9274c6),
	.w4(32'h3a8bb4cd),
	.w5(32'h397f733b),
	.w6(32'h3a498fb1),
	.w7(32'h39ee7b18),
	.w8(32'hb93b63f3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d29ae),
	.w1(32'hba23f259),
	.w2(32'hb9dbfdf0),
	.w3(32'hb93f1c97),
	.w4(32'hb992be91),
	.w5(32'hb9f2aba1),
	.w6(32'hba0f621a),
	.w7(32'hb9fe01af),
	.w8(32'hba3b43f0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f458a5),
	.w1(32'hba9c0fc4),
	.w2(32'hbaa0bd64),
	.w3(32'hb93a3363),
	.w4(32'hba2267b3),
	.w5(32'hba7daaab),
	.w6(32'h3a71bd92),
	.w7(32'h3a7f5519),
	.w8(32'h3a9644c0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8beb81e),
	.w1(32'h3a4a7a63),
	.w2(32'hb9a9b4fc),
	.w3(32'h39ebdb96),
	.w4(32'h3a8f7d65),
	.w5(32'h3a5f8b9e),
	.w6(32'h3acda1cb),
	.w7(32'h3ab9e450),
	.w8(32'h3a90ce49),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52d852),
	.w1(32'hb9c67746),
	.w2(32'hba0cbbea),
	.w3(32'h38d7fcf8),
	.w4(32'hb9fef018),
	.w5(32'hba6afe2a),
	.w6(32'hb7731fe2),
	.w7(32'hba0d767e),
	.w8(32'hba1abee3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a158ad4),
	.w1(32'h398cae99),
	.w2(32'h398a8d32),
	.w3(32'h39f406e7),
	.w4(32'h3acb8ac4),
	.w5(32'h39f4f3df),
	.w6(32'h3ae2d8e4),
	.w7(32'h3a26a2cd),
	.w8(32'hba50cf4f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2c281),
	.w1(32'hba09384d),
	.w2(32'hbada7a37),
	.w3(32'hb90a1e76),
	.w4(32'hbb68da88),
	.w5(32'hbb0d4735),
	.w6(32'h3a226f72),
	.w7(32'hbab26258),
	.w8(32'hbadfba0a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e03a16),
	.w1(32'hba2329b2),
	.w2(32'hba7e31c9),
	.w3(32'h39ccf79d),
	.w4(32'hb939ae65),
	.w5(32'hb9e662aa),
	.w6(32'h39b35303),
	.w7(32'h3935080a),
	.w8(32'h393c7ad3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefc69b),
	.w1(32'hbace07b6),
	.w2(32'hba9117ca),
	.w3(32'hbae4f14f),
	.w4(32'h3935f319),
	.w5(32'hba1bfad3),
	.w6(32'hba11dcb6),
	.w7(32'hb8e9c85b),
	.w8(32'hba8110f6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb8f24),
	.w1(32'hba621ca5),
	.w2(32'hba400d5c),
	.w3(32'hb83ba30f),
	.w4(32'hba7320fc),
	.w5(32'hba924844),
	.w6(32'h392bce02),
	.w7(32'hb9d14993),
	.w8(32'hb919d881),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef4b37),
	.w1(32'hbac86f9b),
	.w2(32'hb9a9c447),
	.w3(32'h3b1aa3e1),
	.w4(32'hb934b314),
	.w5(32'hb8f5fad9),
	.w6(32'h3ae1b0fc),
	.w7(32'h3a6c72ed),
	.w8(32'h3a2a33d1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76ab68),
	.w1(32'hbb50fb90),
	.w2(32'hbb5d9ea9),
	.w3(32'hbb7bec95),
	.w4(32'hbb3460f9),
	.w5(32'hbb39fb3d),
	.w6(32'hbab413f6),
	.w7(32'hbab0a0ae),
	.w8(32'hbb0aa657),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d3a29),
	.w1(32'h399c18aa),
	.w2(32'hb99179ea),
	.w3(32'hba664b81),
	.w4(32'hba50c519),
	.w5(32'hba84568c),
	.w6(32'hba3177b4),
	.w7(32'hbab1b834),
	.w8(32'hba81d096),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aadae),
	.w1(32'hbb2efaf0),
	.w2(32'hbaf56d1a),
	.w3(32'h3a19d428),
	.w4(32'h3a8f674d),
	.w5(32'h39e43ebe),
	.w6(32'h381af440),
	.w7(32'h3b379281),
	.w8(32'h3b5314f1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1feab4),
	.w1(32'hb9ab6626),
	.w2(32'hbaa08913),
	.w3(32'hbb383a5f),
	.w4(32'hb8e971e0),
	.w5(32'hbac06ede),
	.w6(32'hbaba58c8),
	.w7(32'hbaab0681),
	.w8(32'hbad8b08d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79c97c),
	.w1(32'h3a1e960e),
	.w2(32'hb958b8e6),
	.w3(32'h3a325d6f),
	.w4(32'h3887ab4f),
	.w5(32'hba2ae275),
	.w6(32'h39f5a700),
	.w7(32'hbabf431e),
	.w8(32'hbb04196f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae37ad7),
	.w1(32'hbae37d8b),
	.w2(32'hbb168727),
	.w3(32'hba4387c5),
	.w4(32'hbb0e93dd),
	.w5(32'hbaed0973),
	.w6(32'h3b13c84d),
	.w7(32'hb9abdb9f),
	.w8(32'hbb2ffdef),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f9033),
	.w1(32'hbacb2d91),
	.w2(32'hbad8c663),
	.w3(32'hb9e4a3f5),
	.w4(32'hbb02e850),
	.w5(32'hbaf9ada9),
	.w6(32'hb7cc98f4),
	.w7(32'hba861237),
	.w8(32'hbaf28d1a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987bd5b),
	.w1(32'hba830d87),
	.w2(32'hba6789eb),
	.w3(32'hb9a27eb4),
	.w4(32'hba78cd3e),
	.w5(32'hba5278d0),
	.w6(32'hba4d5b0e),
	.w7(32'hba2260cf),
	.w8(32'hb9bf19a8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20664b),
	.w1(32'hba9237c8),
	.w2(32'hba83a3f3),
	.w3(32'hba00058e),
	.w4(32'hba1723e4),
	.w5(32'hba4f0535),
	.w6(32'hb82fe63d),
	.w7(32'hb9004cd3),
	.w8(32'h3949f60b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74047d),
	.w1(32'h3965d620),
	.w2(32'h3ab58f38),
	.w3(32'h3a9685cc),
	.w4(32'h39ca49d9),
	.w5(32'h3a72f3ff),
	.w6(32'hbaeb80d0),
	.w7(32'hbab2fa9f),
	.w8(32'hbaffbba6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8235d1),
	.w1(32'hbb928be1),
	.w2(32'hbb70dbe6),
	.w3(32'hbaf5d054),
	.w4(32'h3916044c),
	.w5(32'hbb15aa97),
	.w6(32'hbb4468c5),
	.w7(32'h3852a059),
	.w8(32'hba3ee6aa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661a40),
	.w1(32'hbaf6ba0b),
	.w2(32'hba9f038f),
	.w3(32'hbae2c927),
	.w4(32'hb9caa397),
	.w5(32'hb9cd4a38),
	.w6(32'hbadc1c19),
	.w7(32'hba340415),
	.w8(32'hb908ae19),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc9515),
	.w1(32'hb9377c76),
	.w2(32'hb93d3730),
	.w3(32'h38af16a6),
	.w4(32'h3a82c0a6),
	.w5(32'h39d7bf12),
	.w6(32'hbaccb344),
	.w7(32'hba125f3e),
	.w8(32'h3a2c7dac),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f8c17),
	.w1(32'h3a5928d9),
	.w2(32'h3ab71411),
	.w3(32'hba2617e2),
	.w4(32'h3a912e86),
	.w5(32'h3a2d4bf9),
	.w6(32'h396dc21d),
	.w7(32'h39e53cde),
	.w8(32'hb8a8a1d7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4afc20),
	.w1(32'hba9a7ee9),
	.w2(32'hba8ca061),
	.w3(32'h39ef4f8b),
	.w4(32'hba828d18),
	.w5(32'hba3f7e68),
	.w6(32'hba432ef9),
	.w7(32'hba0537d8),
	.w8(32'hb9e2ac81),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abc73c),
	.w1(32'hb9f15029),
	.w2(32'hbaf70eaa),
	.w3(32'hba505895),
	.w4(32'hbaaa75e1),
	.w5(32'hb9e27190),
	.w6(32'hb9161fbd),
	.w7(32'hbb69e8c9),
	.w8(32'hba6c20cc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38944557),
	.w1(32'hba166211),
	.w2(32'hba98de7e),
	.w3(32'h39b2f8d4),
	.w4(32'hb91cbbb2),
	.w5(32'hb9f40aa2),
	.w6(32'hb9922420),
	.w7(32'hba71b8a3),
	.w8(32'h3a5a9bcc),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d756e),
	.w1(32'hb8787372),
	.w2(32'hba92339b),
	.w3(32'hbae1d01b),
	.w4(32'h3ac3e8e0),
	.w5(32'hb9f7ce57),
	.w6(32'hba81b9f5),
	.w7(32'hba67a4cd),
	.w8(32'h39c8bc1b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21fe5c),
	.w1(32'hba4e8aa6),
	.w2(32'hba4cb8a6),
	.w3(32'h3a3d717a),
	.w4(32'hba073812),
	.w5(32'hba136799),
	.w6(32'hb98087b2),
	.w7(32'hb9810191),
	.w8(32'hb8dbd01c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01a6a3),
	.w1(32'hba7b1b38),
	.w2(32'hba7f400e),
	.w3(32'hb98513ce),
	.w4(32'hba2597dd),
	.w5(32'hba2fc0e3),
	.w6(32'hb9ed9af5),
	.w7(32'hb9dfdcc4),
	.w8(32'hb9939d4f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba256bde),
	.w1(32'h38236bfc),
	.w2(32'hba8b5126),
	.w3(32'h36e45515),
	.w4(32'h38d2e038),
	.w5(32'hba24b7aa),
	.w6(32'hb98871a0),
	.w7(32'hb9878a80),
	.w8(32'hb9d1d9b2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe988),
	.w1(32'hba7e8228),
	.w2(32'hb9d5e0a6),
	.w3(32'hba7c168e),
	.w4(32'hba12280a),
	.w5(32'h39c49c03),
	.w6(32'hbaf4323e),
	.w7(32'hba02234d),
	.w8(32'hba3752a9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9289ffc),
	.w1(32'h395d82b6),
	.w2(32'h39c873af),
	.w3(32'hb9b9c872),
	.w4(32'h38300daf),
	.w5(32'hb8870267),
	.w6(32'h3a213d5e),
	.w7(32'h39910dee),
	.w8(32'hb9e0236b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10a6ec),
	.w1(32'hbabb7715),
	.w2(32'hba92c31a),
	.w3(32'h39326ac0),
	.w4(32'hba9b971b),
	.w5(32'hbab11d5f),
	.w6(32'hb6ac5d19),
	.w7(32'hb988a579),
	.w8(32'hba035792),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e099b),
	.w1(32'hb93bc13a),
	.w2(32'h3acf5633),
	.w3(32'h3a528649),
	.w4(32'h3a7789f6),
	.w5(32'h39e3acac),
	.w6(32'h3b131095),
	.w7(32'h3b590abe),
	.w8(32'h3b0ba108),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ba891),
	.w1(32'h39b7700f),
	.w2(32'h3a4b1fd1),
	.w3(32'h3aab8f0e),
	.w4(32'h3b79b99d),
	.w5(32'h3b773dcc),
	.w6(32'h36b9ef97),
	.w7(32'h3ab040e4),
	.w8(32'h3b4232f0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf3c06),
	.w1(32'h3b1c02c6),
	.w2(32'h3b724ce9),
	.w3(32'h3b4a0628),
	.w4(32'h3b46db67),
	.w5(32'h3b875450),
	.w6(32'h3b33f7a8),
	.w7(32'h399ddb40),
	.w8(32'h3b5f974e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380bd38a),
	.w1(32'h3920fc76),
	.w2(32'h3960d206),
	.w3(32'h39bf1bc8),
	.w4(32'h3995ba54),
	.w5(32'h391fc429),
	.w6(32'hb80e3629),
	.w7(32'h39551b81),
	.w8(32'hb6983ae9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bcebe),
	.w1(32'hb8b517a4),
	.w2(32'hb9b374c3),
	.w3(32'hb9b4af83),
	.w4(32'h39957743),
	.w5(32'h3960088f),
	.w6(32'h3947eed2),
	.w7(32'h3882db82),
	.w8(32'h3971b725),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ffb683),
	.w1(32'hbac6d768),
	.w2(32'hba3c742c),
	.w3(32'h39a887c4),
	.w4(32'hbaaac2c2),
	.w5(32'hba76b222),
	.w6(32'hba2d5c0c),
	.w7(32'hba10191c),
	.w8(32'hba4c3803),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba830793),
	.w1(32'hba8f6053),
	.w2(32'hba7143c9),
	.w3(32'hbaab2fbf),
	.w4(32'hb9e71a15),
	.w5(32'hba49785b),
	.w6(32'hba191155),
	.w7(32'hb96fe786),
	.w8(32'hba34ca32),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad8974),
	.w1(32'h39ce69e6),
	.w2(32'hba0dfa58),
	.w3(32'hbb58cb19),
	.w4(32'h3b1c5792),
	.w5(32'h3aab0bef),
	.w6(32'h3abfc557),
	.w7(32'h392a17c0),
	.w8(32'h39c42f25),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b7413),
	.w1(32'hbb07de55),
	.w2(32'hba4633cb),
	.w3(32'hba1f3395),
	.w4(32'hb95d513c),
	.w5(32'h39962eb0),
	.w6(32'hbb319f84),
	.w7(32'hba113f6a),
	.w8(32'hb9424475),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782795),
	.w1(32'hbb4cf579),
	.w2(32'hba5791f8),
	.w3(32'hb9f4de03),
	.w4(32'hba4db812),
	.w5(32'h371b67e7),
	.w6(32'hbb56d2a8),
	.w7(32'hb9fd8ec9),
	.w8(32'hb908d50d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53957e),
	.w1(32'hbb92f19e),
	.w2(32'hbb1f5a97),
	.w3(32'hbad18a2b),
	.w4(32'hbb0fb916),
	.w5(32'hbae740cd),
	.w6(32'hbac99743),
	.w7(32'h3a1d5841),
	.w8(32'h3a86ad0e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1e15b),
	.w1(32'hbb8216f7),
	.w2(32'hbb9c5324),
	.w3(32'hbb0ecd80),
	.w4(32'hbb883d3e),
	.w5(32'hbb953cb6),
	.w6(32'h3ab1abfb),
	.w7(32'hbab7ce94),
	.w8(32'hbb423aea),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9837278),
	.w1(32'hbac2c629),
	.w2(32'hba942c69),
	.w3(32'hb94de38f),
	.w4(32'hbab16790),
	.w5(32'hba535a3c),
	.w6(32'hbac7d9c3),
	.w7(32'hbaa1c276),
	.w8(32'hba4ee790),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c7ea2),
	.w1(32'hbab4c325),
	.w2(32'hb9c7a284),
	.w3(32'hbb22c0af),
	.w4(32'hba8275f1),
	.w5(32'hba11fd90),
	.w6(32'hbacf3b3c),
	.w7(32'hb9a188a4),
	.w8(32'hb989732f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d3cfb),
	.w1(32'h3a0bae54),
	.w2(32'h3a2d2b1c),
	.w3(32'h39c8caa7),
	.w4(32'h3aa20b40),
	.w5(32'h3a9f5748),
	.w6(32'h38bdc44b),
	.w7(32'h3a56bf1a),
	.w8(32'h3a716df2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38cf90),
	.w1(32'hbb03407c),
	.w2(32'hbb2733e7),
	.w3(32'h3a0de63c),
	.w4(32'hba5c02d8),
	.w5(32'hba8441e9),
	.w6(32'hb741b9bd),
	.w7(32'hb830c6a5),
	.w8(32'h3a152f3c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91215c),
	.w1(32'hba032491),
	.w2(32'hba73bf24),
	.w3(32'h39efe88f),
	.w4(32'hb91ccfbf),
	.w5(32'hba57df41),
	.w6(32'h39f8c4cd),
	.w7(32'h38639007),
	.w8(32'h38baee81),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb922),
	.w1(32'hbb825919),
	.w2(32'hbb5b1c70),
	.w3(32'hbb6aebdb),
	.w4(32'hbb630964),
	.w5(32'hbae392ee),
	.w6(32'hba1ac35f),
	.w7(32'hba868d99),
	.w8(32'hbb0de3d7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4adc92),
	.w1(32'hb911f576),
	.w2(32'hb9a0ba22),
	.w3(32'hba9e1922),
	.w4(32'hb92d5872),
	.w5(32'hb98254ae),
	.w6(32'hb757670f),
	.w7(32'hba04889a),
	.w8(32'hba48b060),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16672e),
	.w1(32'h398c0c90),
	.w2(32'hb8f5faea),
	.w3(32'hb9511cb5),
	.w4(32'h3a394f1f),
	.w5(32'h394982d6),
	.w6(32'h3a734c98),
	.w7(32'h3a34ecc2),
	.w8(32'h3a4b33b5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39717a80),
	.w1(32'h3950ab56),
	.w2(32'h3a399f82),
	.w3(32'h3a1648fd),
	.w4(32'h3a0903ea),
	.w5(32'h3a7152af),
	.w6(32'h394688e8),
	.w7(32'h3a22b639),
	.w8(32'hb8139d50),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d8e9d0),
	.w1(32'hba7e63bc),
	.w2(32'hbada1489),
	.w3(32'h3a6bfb40),
	.w4(32'hba04d6a6),
	.w5(32'hb9d37c69),
	.w6(32'hba8c64f8),
	.w7(32'hba85a79b),
	.w8(32'hba39e496),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98365df),
	.w1(32'h3a5b94cf),
	.w2(32'h3a06de14),
	.w3(32'hba0b37bb),
	.w4(32'h3a4a4641),
	.w5(32'h39847b41),
	.w6(32'h3a307429),
	.w7(32'h39573498),
	.w8(32'hb7c58f62),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3855cffd),
	.w1(32'hba33eb72),
	.w2(32'hba39aa40),
	.w3(32'h3a1e6cc2),
	.w4(32'hb99e25f6),
	.w5(32'hb9936585),
	.w6(32'h398728d5),
	.w7(32'hb9bba160),
	.w8(32'h3783cae4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed3f51),
	.w1(32'hba9cd9bc),
	.w2(32'hbabd1672),
	.w3(32'hba8f9321),
	.w4(32'hba68a95e),
	.w5(32'hba7c5ead),
	.w6(32'hba2ad376),
	.w7(32'hba2784d0),
	.w8(32'hbae3ced9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e6cfe),
	.w1(32'hba28d27f),
	.w2(32'hba472e71),
	.w3(32'hbaf23142),
	.w4(32'hb9e4c9b2),
	.w5(32'hb996008e),
	.w6(32'hbaad2444),
	.w7(32'hbab4e85a),
	.w8(32'hba27297b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911d11a),
	.w1(32'hb88a0dfd),
	.w2(32'hba9f5fa4),
	.w3(32'h39bc36c5),
	.w4(32'hba2906de),
	.w5(32'hba8551f3),
	.w6(32'hbac6440f),
	.w7(32'hbac92546),
	.w8(32'hba5cd886),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a165077),
	.w1(32'h3ac1db7d),
	.w2(32'h3a436313),
	.w3(32'hb9172f5c),
	.w4(32'h3ae216b2),
	.w5(32'h3a77f3d3),
	.w6(32'h3adb831b),
	.w7(32'h3a620244),
	.w8(32'h39e8c0de),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1386e1),
	.w1(32'hb9588d42),
	.w2(32'hb9272537),
	.w3(32'h3a4d787d),
	.w4(32'hb8c422a6),
	.w5(32'hb9d2eb6e),
	.w6(32'h38fbb547),
	.w7(32'hb6c09dd1),
	.w8(32'hb9555b30),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0bff2),
	.w1(32'hba716027),
	.w2(32'hbaef1445),
	.w3(32'hb8a0d5de),
	.w4(32'hb9e6c2f4),
	.w5(32'hb98d462d),
	.w6(32'hba79f3cd),
	.w7(32'hba879ced),
	.w8(32'hba878759),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00d279),
	.w1(32'h397245ad),
	.w2(32'hba75c6a1),
	.w3(32'hbab16cda),
	.w4(32'h39fb42bc),
	.w5(32'h3aacb10b),
	.w6(32'h38a7aa9b),
	.w7(32'hbb3c27c5),
	.w8(32'hbb23664f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8281f7),
	.w1(32'hbaebac8f),
	.w2(32'hba8b7ad6),
	.w3(32'h3aea6f3a),
	.w4(32'hb82ce556),
	.w5(32'hba95acc4),
	.w6(32'h390c5622),
	.w7(32'h3a6a9d31),
	.w8(32'h39ee3eb9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba574ac8),
	.w1(32'hba7be8fa),
	.w2(32'hb9e20b3e),
	.w3(32'h3ad5dd5b),
	.w4(32'h3a713881),
	.w5(32'h39407e31),
	.w6(32'h39dd83bc),
	.w7(32'hba09bdd9),
	.w8(32'hb9961d5c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e01f),
	.w1(32'hbab52c42),
	.w2(32'hb8eac312),
	.w3(32'hba8f49b7),
	.w4(32'h3a58ad10),
	.w5(32'h3ab78aa7),
	.w6(32'hbb81acd8),
	.w7(32'hbb08b58d),
	.w8(32'h3a47403c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba645273),
	.w1(32'h39058035),
	.w2(32'h3939f9fa),
	.w3(32'hb8ddd80f),
	.w4(32'h3855c0ae),
	.w5(32'hb9397961),
	.w6(32'h399f2fe6),
	.w7(32'hb841e826),
	.w8(32'hb9a51f17),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971c213),
	.w1(32'hba2cfc81),
	.w2(32'hba53f2f6),
	.w3(32'hb93dd611),
	.w4(32'hba25c2df),
	.w5(32'hba3bc9b5),
	.w6(32'hb9b56c3f),
	.w7(32'hb9f86b3b),
	.w8(32'hb9390a2d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0425d7),
	.w1(32'hba26fee5),
	.w2(32'hba5348eb),
	.w3(32'hb9a51318),
	.w4(32'hba06b7f3),
	.w5(32'hba3209c5),
	.w6(32'hb971e5f0),
	.w7(32'hb9ed9deb),
	.w8(32'hb815b998),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd209e),
	.w1(32'hbafbfd3e),
	.w2(32'hbb025f1b),
	.w3(32'hb96e84b8),
	.w4(32'hbacc91f1),
	.w5(32'hbabb88f0),
	.w6(32'hb9ebd002),
	.w7(32'hba9171ad),
	.w8(32'hbaa444cb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9e565),
	.w1(32'hb859d175),
	.w2(32'h38fa9844),
	.w3(32'hba80bfc6),
	.w4(32'hb8bc70b1),
	.w5(32'hb9afa306),
	.w6(32'h399d30d9),
	.w7(32'h397de80b),
	.w8(32'hb7f939b0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7799cb),
	.w1(32'hbb3fc1e2),
	.w2(32'hbb087bad),
	.w3(32'hb9227141),
	.w4(32'hbb16782d),
	.w5(32'hbaf5cadf),
	.w6(32'h3ab5018f),
	.w7(32'h3a123882),
	.w8(32'hba8c6b4b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b6072),
	.w1(32'hba906eeb),
	.w2(32'hbb3e0519),
	.w3(32'h3a09c84c),
	.w4(32'hba66ca56),
	.w5(32'hbaa568c3),
	.w6(32'h3a539e35),
	.w7(32'hbabbf012),
	.w8(32'hbaaac648),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21429),
	.w1(32'hb9c547ff),
	.w2(32'hba6f9b52),
	.w3(32'hba1bcfdb),
	.w4(32'hb88c6e12),
	.w5(32'hba4a5791),
	.w6(32'hbae2b4e1),
	.w7(32'hba81a04e),
	.w8(32'hba26434c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2cb4a),
	.w1(32'hbad3a291),
	.w2(32'hbae3eb57),
	.w3(32'hba8ef936),
	.w4(32'hba9f6117),
	.w5(32'hbad5e276),
	.w6(32'hbaac4673),
	.w7(32'hbb1843bd),
	.w8(32'hbb441a50),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb948d067),
	.w1(32'hbad865c1),
	.w2(32'hbadb04ba),
	.w3(32'hba66ed39),
	.w4(32'hba8e0b66),
	.w5(32'hba3871f6),
	.w6(32'h39314a04),
	.w7(32'hbaa1022e),
	.w8(32'hba5f4aa7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef3b07),
	.w1(32'hba732dd8),
	.w2(32'hba05616f),
	.w3(32'hba8496af),
	.w4(32'h398e818a),
	.w5(32'h3a4399f5),
	.w6(32'hba5e8cf8),
	.w7(32'h39838d5d),
	.w8(32'h3a219770),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16aa80),
	.w1(32'h3a01ca9e),
	.w2(32'h39e74f6f),
	.w3(32'h3ac146a8),
	.w4(32'h393eacf6),
	.w5(32'h399d73e7),
	.w6(32'h3adb0df7),
	.w7(32'h3a586b87),
	.w8(32'hba438e46),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca0ee3),
	.w1(32'hb9c2510a),
	.w2(32'hb9b79826),
	.w3(32'h3960b2c6),
	.w4(32'hb95c094c),
	.w5(32'hb9c308e1),
	.w6(32'h3902d705),
	.w7(32'hb8b1b7a3),
	.w8(32'h394bbf50),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9088c61),
	.w1(32'h398a0e8b),
	.w2(32'h38de75a2),
	.w3(32'hb8e78334),
	.w4(32'h39d70c4c),
	.w5(32'hb865d02d),
	.w6(32'hb98998b1),
	.w7(32'hb9a80068),
	.w8(32'hba0852eb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99097e9),
	.w1(32'hba96d448),
	.w2(32'hba52f63d),
	.w3(32'hb9a1efc1),
	.w4(32'hba682a54),
	.w5(32'hb9a6044a),
	.w6(32'hba4d32f6),
	.w7(32'hb9f84372),
	.w8(32'h392c86cb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00f00e),
	.w1(32'h3a27f5ad),
	.w2(32'h3a6825e5),
	.w3(32'hb7a2c5c7),
	.w4(32'h3a66c526),
	.w5(32'h3a8df300),
	.w6(32'h3a14b39b),
	.w7(32'h3a19c3f8),
	.w8(32'h39eb01cf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c11b1),
	.w1(32'h39f48a8d),
	.w2(32'h3a354a7a),
	.w3(32'h3aba5c64),
	.w4(32'h3a3d4cde),
	.w5(32'h3aad4cc8),
	.w6(32'hb89fa47e),
	.w7(32'h370e57d6),
	.w8(32'h3a181b83),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398edf41),
	.w1(32'hba3eb5e3),
	.w2(32'hb9c0eace),
	.w3(32'h3a008f7c),
	.w4(32'hb97b38bf),
	.w5(32'hb7e01a3d),
	.w6(32'hb9d99030),
	.w7(32'hb9721091),
	.w8(32'h395e4573),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb4a59),
	.w1(32'hbacbc868),
	.w2(32'hba493468),
	.w3(32'hb909271d),
	.w4(32'hba3b2c3b),
	.w5(32'hbaaeb617),
	.w6(32'hb90628ff),
	.w7(32'h3a0819a6),
	.w8(32'hb9ebf9b2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa68ec6),
	.w1(32'hbb176f20),
	.w2(32'hbb2eb58b),
	.w3(32'hbaa0a0ca),
	.w4(32'hbb03f157),
	.w5(32'hbaccf8f9),
	.w6(32'hba2b3678),
	.w7(32'hbad4bc75),
	.w8(32'hbaf1d089),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aacc15),
	.w1(32'h39d465df),
	.w2(32'h3a516052),
	.w3(32'hb9e88f53),
	.w4(32'h39927881),
	.w5(32'h3a6c244a),
	.w6(32'hba278f7b),
	.w7(32'hb958bb50),
	.w8(32'h3accab32),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81de58),
	.w1(32'hba6c2c37),
	.w2(32'hbb09581c),
	.w3(32'h39cb7269),
	.w4(32'h3aeaa73d),
	.w5(32'h39005cb4),
	.w6(32'h3b2ba899),
	.w7(32'h3a97173f),
	.w8(32'hb9b9ddec),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88acc6),
	.w1(32'h3a7c1e08),
	.w2(32'h3a9173a1),
	.w3(32'h3b07ae4c),
	.w4(32'h3aa2ce49),
	.w5(32'h3a6d1106),
	.w6(32'h3ac48335),
	.w7(32'h3a9ad237),
	.w8(32'h3a76f874),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba011c2),
	.w1(32'hbb8fced1),
	.w2(32'hbb3b851d),
	.w3(32'hbb81bc67),
	.w4(32'hbb29de1d),
	.w5(32'hbb00a61a),
	.w6(32'hbb26f4ac),
	.w7(32'hbb405439),
	.w8(32'hbb2d6c8d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba958dc8),
	.w1(32'h3a5a5b61),
	.w2(32'h3995d3eb),
	.w3(32'h3a9a3beb),
	.w4(32'h3afcebf7),
	.w5(32'h3a729811),
	.w6(32'hb9a2e358),
	.w7(32'h3a5f46bb),
	.w8(32'h390f7a67),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada82ac),
	.w1(32'hba97cc4b),
	.w2(32'hb9e463ad),
	.w3(32'hba9e5362),
	.w4(32'hba81bcff),
	.w5(32'hb9a957a5),
	.w6(32'hbb0dcefb),
	.w7(32'hbb041de9),
	.w8(32'hb9e8a328),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07db03),
	.w1(32'h3995d537),
	.w2(32'hba488f2d),
	.w3(32'hba0c7b5f),
	.w4(32'hba3e3129),
	.w5(32'hba936a8a),
	.w6(32'hb99ce485),
	.w7(32'hb940b401),
	.w8(32'hbac0ebcc),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b9a8),
	.w1(32'hbb2f4152),
	.w2(32'hbb58f721),
	.w3(32'hbb55e9d5),
	.w4(32'hbaf25bd1),
	.w5(32'hbafc373e),
	.w6(32'hbb36cb97),
	.w7(32'hbb0558d6),
	.w8(32'h3787a0ef),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38153387),
	.w1(32'hba1a547d),
	.w2(32'h3aed5bde),
	.w3(32'h3af0c18e),
	.w4(32'h3ab2dee7),
	.w5(32'h3b31b8c1),
	.w6(32'h3aeec5c7),
	.w7(32'h39a2fff4),
	.w8(32'h39568e48),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548f24),
	.w1(32'hba23aab5),
	.w2(32'h37c57b96),
	.w3(32'h3ad91193),
	.w4(32'hba4a9c87),
	.w5(32'hbb2047e9),
	.w6(32'h399abceb),
	.w7(32'hb953b049),
	.w8(32'h39f370c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6e4a),
	.w1(32'hba8baf51),
	.w2(32'hbaa8d11f),
	.w3(32'hbacce4c5),
	.w4(32'h3afb5cc9),
	.w5(32'h3ad75d62),
	.w6(32'hbacf2243),
	.w7(32'h3b1a3195),
	.w8(32'h3b5c17c6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7537c),
	.w1(32'hbac985a6),
	.w2(32'hba5c8e43),
	.w3(32'hbb6357a3),
	.w4(32'hb981e354),
	.w5(32'h3a0f061f),
	.w6(32'hbb99bad4),
	.w7(32'hba2fdf14),
	.w8(32'hbaf11d9b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef1e39),
	.w1(32'hbb334188),
	.w2(32'hbae72721),
	.w3(32'h3afded33),
	.w4(32'h3a0a4935),
	.w5(32'hbb1955f1),
	.w6(32'h3af5c0e5),
	.w7(32'hb931aeb8),
	.w8(32'h391f6e77),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5767b1),
	.w1(32'h3a64857d),
	.w2(32'h39c1a238),
	.w3(32'h3ab6978c),
	.w4(32'h3a647493),
	.w5(32'h3a3f5bc7),
	.w6(32'h39a9bc30),
	.w7(32'h3a2fe43f),
	.w8(32'h3a9c43d1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a407d75),
	.w1(32'hbac83830),
	.w2(32'hbb08a81d),
	.w3(32'hbb005b07),
	.w4(32'hbb2b2dc8),
	.w5(32'hbb079f19),
	.w6(32'hba1f698d),
	.w7(32'hba936e2e),
	.w8(32'hba3587fb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbd535),
	.w1(32'hb9fdb12b),
	.w2(32'hba720be7),
	.w3(32'h3b116fd6),
	.w4(32'h397abcf4),
	.w5(32'h39518259),
	.w6(32'h3a035e47),
	.w7(32'h3a2324a3),
	.w8(32'h3a220b50),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9251880),
	.w1(32'hb9c0448a),
	.w2(32'hb924f88f),
	.w3(32'hb8a0452d),
	.w4(32'h38efc5be),
	.w5(32'hb83af2ce),
	.w6(32'hb9bf28ae),
	.w7(32'hba30f5cb),
	.w8(32'hba7cb6c4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8942a2),
	.w1(32'hbab08edf),
	.w2(32'hba810b93),
	.w3(32'hba57b044),
	.w4(32'hb9a22348),
	.w5(32'hba444f91),
	.w6(32'hba831aaf),
	.w7(32'hba387328),
	.w8(32'hb9eaaaad),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040ca1),
	.w1(32'hbad0548b),
	.w2(32'hbab3c0f4),
	.w3(32'hba545c93),
	.w4(32'hb95df4bd),
	.w5(32'hba0cd8f7),
	.w6(32'hba158be7),
	.w7(32'h37e6d2ef),
	.w8(32'h39c40da6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870951),
	.w1(32'hbae92dfb),
	.w2(32'hba7d140c),
	.w3(32'hbb125d63),
	.w4(32'hb987afd3),
	.w5(32'hba0492e1),
	.w6(32'hbb6c027e),
	.w7(32'hba7756cf),
	.w8(32'hb9ab6371),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7963f0),
	.w1(32'hba388608),
	.w2(32'hb9273748),
	.w3(32'hb9c096b3),
	.w4(32'hba133239),
	.w5(32'h39ff595a),
	.w6(32'hba515918),
	.w7(32'hb90895bf),
	.w8(32'h3b0ead5f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d657f),
	.w1(32'hbb11f242),
	.w2(32'hbadaf972),
	.w3(32'hbab42c0e),
	.w4(32'hbaf884c0),
	.w5(32'hba88c629),
	.w6(32'hbb447b30),
	.w7(32'hbb3d570d),
	.w8(32'hba99be55),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b5ed2),
	.w1(32'hb9b4c101),
	.w2(32'h39f5902e),
	.w3(32'h3a21bf4a),
	.w4(32'h37a08a70),
	.w5(32'h395cfa6b),
	.w6(32'h3a3af3c4),
	.w7(32'h3aafb45b),
	.w8(32'h3ab16828),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba497835),
	.w1(32'hb9f6bf24),
	.w2(32'hb9b8d518),
	.w3(32'hbaa21d98),
	.w4(32'hba132256),
	.w5(32'hbaa9f02a),
	.w6(32'hbad92e7c),
	.w7(32'hbb166f21),
	.w8(32'hbafe23e7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa07cbb),
	.w1(32'hbadff86d),
	.w2(32'hba8eb7a0),
	.w3(32'hba36375d),
	.w4(32'hba3d940a),
	.w5(32'hba11b7df),
	.w6(32'hba99d14a),
	.w7(32'hba1f2191),
	.w8(32'hb9664627),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c868b),
	.w1(32'hb982c1bc),
	.w2(32'hba39a1d4),
	.w3(32'hb9bdb074),
	.w4(32'h3892d6bf),
	.w5(32'hb95203b1),
	.w6(32'hb81c78f3),
	.w7(32'hb9dcc4a4),
	.w8(32'h39f78fc6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372ed91e),
	.w1(32'hb98b4537),
	.w2(32'hba23ff2a),
	.w3(32'h3a0791e5),
	.w4(32'hb9d35d5e),
	.w5(32'hba06310f),
	.w6(32'hb93a554c),
	.w7(32'hb9cc86a4),
	.w8(32'hb921899e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b36b),
	.w1(32'hb99eb058),
	.w2(32'hba0b296c),
	.w3(32'hb9002b25),
	.w4(32'hb973ac15),
	.w5(32'hb9fcd1ec),
	.w6(32'h38b6841c),
	.w7(32'hb91ed01a),
	.w8(32'h38eefcd2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec617f),
	.w1(32'hba18ce00),
	.w2(32'hb7c7e6da),
	.w3(32'h3a5f2360),
	.w4(32'hb9a3da0c),
	.w5(32'hb8374cbe),
	.w6(32'hbaef9568),
	.w7(32'hbabbebe1),
	.w8(32'hbb07fd5b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50ccf3),
	.w1(32'h332a2dc0),
	.w2(32'h385aeb80),
	.w3(32'hbae7cc90),
	.w4(32'h3a0fd0f5),
	.w5(32'h3a79c396),
	.w6(32'hbae5aeeb),
	.w7(32'h3a7bda66),
	.w8(32'h3a438b02),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ef597),
	.w1(32'hbb1f35f7),
	.w2(32'hbb23edd0),
	.w3(32'h3877550a),
	.w4(32'hbb08d2f8),
	.w5(32'hbb164086),
	.w6(32'hba239a24),
	.w7(32'hba81c0ae),
	.w8(32'hba7376a1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81e58),
	.w1(32'hbb21e59d),
	.w2(32'hbb245245),
	.w3(32'hbad83524),
	.w4(32'hbb12efff),
	.w5(32'hbb0ead29),
	.w6(32'hbac23ae4),
	.w7(32'hbaf27dc2),
	.w8(32'hbae111e6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf434),
	.w1(32'hba4386e7),
	.w2(32'hba640622),
	.w3(32'hba93e6b9),
	.w4(32'h3814fb02),
	.w5(32'hb9a257ee),
	.w6(32'hbaa5cffd),
	.w7(32'hbab2f78a),
	.w8(32'hb9ea151e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e82a1d),
	.w1(32'hbad6b047),
	.w2(32'hb8f2caef),
	.w3(32'hb8875559),
	.w4(32'hbb0413a1),
	.w5(32'hba71c39b),
	.w6(32'hbb369bb8),
	.w7(32'hbb06172a),
	.w8(32'hbb5f92be),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8964e5),
	.w1(32'h3a198261),
	.w2(32'h39b1f566),
	.w3(32'hb9be2937),
	.w4(32'h398d30d2),
	.w5(32'hb9732867),
	.w6(32'h3a667e40),
	.w7(32'hb9969e13),
	.w8(32'hb9448e8c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c97927),
	.w1(32'hbad474f8),
	.w2(32'hbaccb810),
	.w3(32'h37af5a97),
	.w4(32'hba8a1729),
	.w5(32'hba88e70e),
	.w6(32'hba059711),
	.w7(32'hba0b2c86),
	.w8(32'hb8d7fffd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba555f1e),
	.w1(32'h3855e2a5),
	.w2(32'h38925c1c),
	.w3(32'h394f33ba),
	.w4(32'h3a0c7aae),
	.w5(32'h38fb8f27),
	.w6(32'h39e9cc76),
	.w7(32'h39e327e8),
	.w8(32'h394ee6be),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0754a9),
	.w1(32'hb8ab70a6),
	.w2(32'h3ab04d80),
	.w3(32'h3a913e5c),
	.w4(32'h3932bde6),
	.w5(32'hba998364),
	.w6(32'h3a743b09),
	.w7(32'h3abc3900),
	.w8(32'h3a123d0d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae6439),
	.w1(32'hbae41aec),
	.w2(32'hbb17eb8e),
	.w3(32'hba5b5563),
	.w4(32'hbac4b8ae),
	.w5(32'hba45c22f),
	.w6(32'h39eb2b10),
	.w7(32'hb9cf2563),
	.w8(32'hba115761),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39525d5b),
	.w1(32'hb918ddef),
	.w2(32'hb930572b),
	.w3(32'h38598045),
	.w4(32'hb85ba7be),
	.w5(32'hb8ce1f97),
	.w6(32'hb6a9f8dd),
	.w7(32'hb85ee2f4),
	.w8(32'hb9071d28),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95da4f1),
	.w1(32'hb9659e1f),
	.w2(32'h37e641eb),
	.w3(32'h39b32dfd),
	.w4(32'hb958ac04),
	.w5(32'h39448eab),
	.w6(32'h3978246c),
	.w7(32'h3926067b),
	.w8(32'hb94d0210),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf1943),
	.w1(32'h38a406f6),
	.w2(32'h3852ed11),
	.w3(32'h36f50324),
	.w4(32'h391e7d07),
	.w5(32'h38de2e40),
	.w6(32'h38317028),
	.w7(32'hb775cacd),
	.w8(32'h385a52b7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5524f0),
	.w1(32'hb9b99605),
	.w2(32'hb9c51e2a),
	.w3(32'hba20a2e3),
	.w4(32'hb9fcda18),
	.w5(32'hb911c871),
	.w6(32'hba11918a),
	.w7(32'hb99ba990),
	.w8(32'hb9de8656),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa51e36),
	.w1(32'hb8ece7e6),
	.w2(32'hba1c9ce7),
	.w3(32'hba1d4d7a),
	.w4(32'h39fd76f4),
	.w5(32'hb97c3793),
	.w6(32'hb9cb0928),
	.w7(32'hba12164f),
	.w8(32'hba46b1c2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3220d8),
	.w1(32'hbad72957),
	.w2(32'hbb209d7a),
	.w3(32'hba0b7bfa),
	.w4(32'hba83924d),
	.w5(32'hb964e3b5),
	.w6(32'hb7825e57),
	.w7(32'hba88e170),
	.w8(32'hbaf426e8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cf0e9),
	.w1(32'hba2822e1),
	.w2(32'hb9c4f7c1),
	.w3(32'hba039470),
	.w4(32'hb70a40df),
	.w5(32'hb8eb7be7),
	.w6(32'hba410fd7),
	.w7(32'hb8e840af),
	.w8(32'h394bd056),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac55790),
	.w1(32'hba922f50),
	.w2(32'hb9b3a92f),
	.w3(32'hba7802a6),
	.w4(32'h373f05cc),
	.w5(32'h390b64d6),
	.w6(32'hba81f9cf),
	.w7(32'hba65f1e3),
	.w8(32'hb9a64254),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380754f4),
	.w1(32'hbaa84f73),
	.w2(32'hbabb947c),
	.w3(32'h39817f6e),
	.w4(32'hba5ae1f8),
	.w5(32'hba6f6865),
	.w6(32'h3a313603),
	.w7(32'hb98c6dc7),
	.w8(32'hba44cbf8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c06359),
	.w1(32'h387fe873),
	.w2(32'h39fff029),
	.w3(32'h3a32372e),
	.w4(32'h3a166800),
	.w5(32'hb988ef6c),
	.w6(32'h37e1f6cc),
	.w7(32'h39ea2773),
	.w8(32'h39b5df65),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869a3b),
	.w1(32'hba552ef4),
	.w2(32'hba0fe680),
	.w3(32'hba53857f),
	.w4(32'hb89ca770),
	.w5(32'h38c8d1c0),
	.w6(32'hb9bfc162),
	.w7(32'h39031963),
	.w8(32'hb9da4c19),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c89ff6),
	.w1(32'hb9416b92),
	.w2(32'hb90685e8),
	.w3(32'hb93758f9),
	.w4(32'h38a71eba),
	.w5(32'h377d8293),
	.w6(32'hb964f70d),
	.w7(32'h38a4f036),
	.w8(32'h38d36edb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cb393),
	.w1(32'hbaeea03a),
	.w2(32'hba735381),
	.w3(32'h3a27331d),
	.w4(32'h38e96bc5),
	.w5(32'hba0bc80f),
	.w6(32'hb96e5c80),
	.w7(32'hb8e7852f),
	.w8(32'hb93a0c8e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d44db),
	.w1(32'h39e9cf08),
	.w2(32'h391ff74c),
	.w3(32'h3a09414c),
	.w4(32'h3a8f00e9),
	.w5(32'h398bd1d2),
	.w6(32'h37c1a92a),
	.w7(32'h39e4c6c4),
	.w8(32'h3978477f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361c164a),
	.w1(32'hb6091b22),
	.w2(32'h37c111c6),
	.w3(32'h3861c0e6),
	.w4(32'h38039798),
	.w5(32'h37fdc4c1),
	.w6(32'h38524e76),
	.w7(32'h37ac36d0),
	.w8(32'h379c19d4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364143a3),
	.w1(32'hb7cfa1e0),
	.w2(32'hb6628d9f),
	.w3(32'h3796711c),
	.w4(32'h36f5a8d1),
	.w5(32'hb69b3bd9),
	.w6(32'h37c189e0),
	.w7(32'h37029571),
	.w8(32'h37b02827),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39467af2),
	.w1(32'hb9a73960),
	.w2(32'hb930a532),
	.w3(32'h39684a5c),
	.w4(32'hb82c0dd2),
	.w5(32'hb908eceb),
	.w6(32'h392cd9dd),
	.w7(32'h38a0d6f6),
	.w8(32'h3958b357),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba913b97),
	.w1(32'hb9839467),
	.w2(32'hb9dbe56b),
	.w3(32'hba1e6b85),
	.w4(32'h39a06087),
	.w5(32'h39b0e6e4),
	.w6(32'hbaa196b9),
	.w7(32'hba30d3aa),
	.w8(32'h3a12ca32),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04ec00),
	.w1(32'hbb05518c),
	.w2(32'hba90bb58),
	.w3(32'hbab7ff53),
	.w4(32'hbac3c54b),
	.w5(32'hba92ee08),
	.w6(32'hba795533),
	.w7(32'hba70323b),
	.w8(32'hba0b3d9c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37122e31),
	.w1(32'hb744168e),
	.w2(32'hb7237c37),
	.w3(32'h37ca58d1),
	.w4(32'h37092108),
	.w5(32'hb62835d5),
	.w6(32'h380689ba),
	.w7(32'h3792645c),
	.w8(32'h35f76c77),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc8108),
	.w1(32'hbadcb86e),
	.w2(32'hba9cf485),
	.w3(32'hb9bbcbc3),
	.w4(32'hba4ad472),
	.w5(32'hb9e6acc3),
	.w6(32'hb9117926),
	.w7(32'h387310dd),
	.w8(32'hba0b99c8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3adbce),
	.w1(32'h37edbff6),
	.w2(32'h394c0d95),
	.w3(32'h3938700e),
	.w4(32'h3866c811),
	.w5(32'hba14f123),
	.w6(32'h3a06953c),
	.w7(32'h3a57021c),
	.w8(32'hba185f0b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39437b15),
	.w1(32'hba87422c),
	.w2(32'hba75a92f),
	.w3(32'h3984984b),
	.w4(32'hba99e3d3),
	.w5(32'hba8c407f),
	.w6(32'h393acb88),
	.w7(32'hbad2d045),
	.w8(32'hbae0ceee),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a680d),
	.w1(32'hbae2c7b7),
	.w2(32'hba7d1c7b),
	.w3(32'hba8e5907),
	.w4(32'hba66e55c),
	.w5(32'h3a0ca7cd),
	.w6(32'hbafba969),
	.w7(32'hbb41ec9d),
	.w8(32'h38138d6c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a275e10),
	.w1(32'h39daf7a1),
	.w2(32'h394b82e0),
	.w3(32'h3a2d43f5),
	.w4(32'h3a6faead),
	.w5(32'h39f4912e),
	.w6(32'hb930344d),
	.w7(32'h38024980),
	.w8(32'h39b211f6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0ff47),
	.w1(32'h3a9efdbd),
	.w2(32'h3b0cc43d),
	.w3(32'h3b0b8b55),
	.w4(32'h3aecf42e),
	.w5(32'h3af0a958),
	.w6(32'h3b0cc588),
	.w7(32'h3ae6c693),
	.w8(32'h3af19bf0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367402),
	.w1(32'hbb1946ff),
	.w2(32'hba924a6d),
	.w3(32'hbae3d466),
	.w4(32'hba8e0547),
	.w5(32'hba08ce98),
	.w6(32'hbaf4ddcd),
	.w7(32'hb9c3ed4d),
	.w8(32'h398c763f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d067d9),
	.w1(32'h3aa2d129),
	.w2(32'h3a6d2082),
	.w3(32'h380bc911),
	.w4(32'h39094e11),
	.w5(32'hb98b5b7f),
	.w6(32'h3a82861f),
	.w7(32'hba32bad8),
	.w8(32'hb9f0b5d2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41ed2e),
	.w1(32'h3a94fbbe),
	.w2(32'h3aa9edfa),
	.w3(32'h3a23d317),
	.w4(32'h3a8c0058),
	.w5(32'h3a999a0e),
	.w6(32'h3845eb2e),
	.w7(32'h3941453b),
	.w8(32'h3a15cf49),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ea73a),
	.w1(32'hb9782438),
	.w2(32'hb901736d),
	.w3(32'h38a6012e),
	.w4(32'hb9475783),
	.w5(32'hb8b60318),
	.w6(32'h38f8c36d),
	.w7(32'hb783a1b8),
	.w8(32'hb90d663c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a1174),
	.w1(32'h381b7569),
	.w2(32'h36604342),
	.w3(32'h38ab6315),
	.w4(32'h3911a4d8),
	.w5(32'h388fcba8),
	.w6(32'hb8b09a0b),
	.w7(32'hb8163820),
	.w8(32'hb6e276e5),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac25b9e),
	.w1(32'hbae281f0),
	.w2(32'hba54de23),
	.w3(32'hbaba07b0),
	.w4(32'hba62bad0),
	.w5(32'h392d0a9f),
	.w6(32'hbabe1203),
	.w7(32'hba20c356),
	.w8(32'hb8873dd4),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3836b14a),
	.w1(32'hb8c8c961),
	.w2(32'hb905bb32),
	.w3(32'h394bf5ce),
	.w4(32'h396db2e4),
	.w5(32'h390fd5fa),
	.w6(32'h397be28b),
	.w7(32'h3933a658),
	.w8(32'h39b14964),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ae703),
	.w1(32'hba6b2272),
	.w2(32'hb981238a),
	.w3(32'hba1e105c),
	.w4(32'hb933356d),
	.w5(32'h390ab466),
	.w6(32'hba54ef7d),
	.w7(32'hb97a352e),
	.w8(32'h3a38a67b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915f0df),
	.w1(32'h3967c74b),
	.w2(32'hb8bed0a0),
	.w3(32'hb8042ecc),
	.w4(32'hb92aaa74),
	.w5(32'hb987fd20),
	.w6(32'hb8ad2fe0),
	.w7(32'hb93bb836),
	.w8(32'hb9c2d49e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83fce6),
	.w1(32'h3a9c0b86),
	.w2(32'h3aa3403e),
	.w3(32'h3b5f5eb0),
	.w4(32'h3a6f6f28),
	.w5(32'h3a8bfe4e),
	.w6(32'h3b42dbec),
	.w7(32'h3977c36e),
	.w8(32'hb93e6fc2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3ac5f),
	.w1(32'h3987cad5),
	.w2(32'h391fb038),
	.w3(32'h39aa6a46),
	.w4(32'h3993b542),
	.w5(32'h37d7af89),
	.w6(32'h39c84a5b),
	.w7(32'h39be5e3a),
	.w8(32'h38936301),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39782ad9),
	.w1(32'h384e0c84),
	.w2(32'hb85af01e),
	.w3(32'h39b02166),
	.w4(32'h38928c7d),
	.w5(32'h38577437),
	.w6(32'h3a058b68),
	.w7(32'hb6e34ee7),
	.w8(32'hb89ba972),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba696e1c),
	.w1(32'hbb03cbc5),
	.w2(32'hb9b288a5),
	.w3(32'hb989e91e),
	.w4(32'hb9d29454),
	.w5(32'h3a0410dc),
	.w6(32'hbaf47ba5),
	.w7(32'hba1f4580),
	.w8(32'h3ab1629b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59bf11),
	.w1(32'hba76e07f),
	.w2(32'h398a4568),
	.w3(32'hba3f5416),
	.w4(32'hb98093c8),
	.w5(32'h397e5f00),
	.w6(32'hbae29dbb),
	.w7(32'h3a346e59),
	.w8(32'h390b00b3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9dcb0d),
	.w1(32'h3a9fd8b4),
	.w2(32'h3a841995),
	.w3(32'h3a5bbb34),
	.w4(32'h3a356a31),
	.w5(32'h3a4f5057),
	.w6(32'h3a180938),
	.w7(32'h39f216dd),
	.w8(32'h3a03d15f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3816fa),
	.w1(32'hbb024bab),
	.w2(32'hbad4f556),
	.w3(32'hba7ab77b),
	.w4(32'hba8c3126),
	.w5(32'hbaaa7f0f),
	.w6(32'h39cfa084),
	.w7(32'hb8846dcf),
	.w8(32'hb95b6f66),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3b494),
	.w1(32'h39bb8267),
	.w2(32'hb900d9e5),
	.w3(32'h39658abd),
	.w4(32'h39527db3),
	.w5(32'h389e234c),
	.w6(32'h38be0f23),
	.w7(32'hb9cbd02e),
	.w8(32'hb94feca3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf1472),
	.w1(32'hbb27c7fe),
	.w2(32'hbad0f4ec),
	.w3(32'hb77cdbc2),
	.w4(32'hba379c81),
	.w5(32'hb83c0352),
	.w6(32'h38b7211c),
	.w7(32'hba7b761e),
	.w8(32'hb95014b5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a33175),
	.w1(32'hba0b43f3),
	.w2(32'hb9355f41),
	.w3(32'h38f225b1),
	.w4(32'hb59e714c),
	.w5(32'h3912a515),
	.w6(32'hb8e8b49a),
	.w7(32'hba314ed1),
	.w8(32'hb9f6f55d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82acd5),
	.w1(32'hbaf57f67),
	.w2(32'hba2ec54e),
	.w3(32'hbb272269),
	.w4(32'hba039775),
	.w5(32'h398ed34f),
	.w6(32'hbab7e851),
	.w7(32'h39e25b83),
	.w8(32'hb84f432d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c392ed),
	.w1(32'h396b81aa),
	.w2(32'hb8b16913),
	.w3(32'h38ce01aa),
	.w4(32'h38d99db5),
	.w5(32'hb8ac45e1),
	.w6(32'hb9f7d34b),
	.w7(32'hb8a7ddf3),
	.w8(32'h38f54de8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f6072),
	.w1(32'hba1d417a),
	.w2(32'hb9c64e75),
	.w3(32'hb94d22d0),
	.w4(32'hb970ce8b),
	.w5(32'hb9aa4d2c),
	.w6(32'hb995dea7),
	.w7(32'hba507de2),
	.w8(32'hba3cac88),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c85a21),
	.w1(32'h3747c4aa),
	.w2(32'h37a8fdee),
	.w3(32'h380d5907),
	.w4(32'h37788b17),
	.w5(32'h3724e5b1),
	.w6(32'h386ae886),
	.w7(32'h37e02037),
	.w8(32'h37c85957),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93782b1),
	.w1(32'hb5b7c0bc),
	.w2(32'h39a12269),
	.w3(32'hb9923594),
	.w4(32'h379b061e),
	.w5(32'h39d8c9ec),
	.w6(32'hb8d8dd45),
	.w7(32'h38c4ce2d),
	.w8(32'h3908d888),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989b2bd),
	.w1(32'hb903c034),
	.w2(32'hb87ab2a3),
	.w3(32'hb8c68c9f),
	.w4(32'h38c92e87),
	.w5(32'h38876939),
	.w6(32'hb8abd7b9),
	.w7(32'h3695a291),
	.w8(32'h3885be35),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58fca0),
	.w1(32'hba6dac2a),
	.w2(32'hbab8b9e9),
	.w3(32'hb9fe88e5),
	.w4(32'hba629272),
	.w5(32'hba97a68d),
	.w6(32'hba6fe0e5),
	.w7(32'hbadd1519),
	.w8(32'hbae6c6f9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67f4cda),
	.w1(32'hb7386df4),
	.w2(32'hb6aff021),
	.w3(32'hb62ac9b0),
	.w4(32'hb72d7c00),
	.w5(32'hb702ac7c),
	.w6(32'hb6a0ec11),
	.w7(32'hb69ac75d),
	.w8(32'hb5ba9964),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbcd3d),
	.w1(32'hb9f466de),
	.w2(32'hb98600c3),
	.w3(32'hb9958311),
	.w4(32'hb9745c9d),
	.w5(32'hb89549ad),
	.w6(32'hb9a73d14),
	.w7(32'hb9917ec4),
	.w8(32'hb82aa88b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9600814),
	.w1(32'hb87b6ab8),
	.w2(32'h39456fbf),
	.w3(32'hb5ba1344),
	.w4(32'h38c92393),
	.w5(32'h3984bf8b),
	.w6(32'hb9e4e973),
	.w7(32'hba060acd),
	.w8(32'hb8b29804),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2018),
	.w1(32'hb99e3521),
	.w2(32'hba1128c9),
	.w3(32'h3acc66b4),
	.w4(32'h3a8f3c06),
	.w5(32'h399eab59),
	.w6(32'h3a58f597),
	.w7(32'hb9ba9487),
	.w8(32'hba4278fb),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d7ee),
	.w1(32'h3a441dd8),
	.w2(32'hb8f2846f),
	.w3(32'hb88e1d4a),
	.w4(32'hb9a95a9b),
	.w5(32'hb94c9760),
	.w6(32'h383a6ba9),
	.w7(32'h38bd262a),
	.w8(32'h388d50ff),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca14ff),
	.w1(32'h3856acbb),
	.w2(32'hba1a5758),
	.w3(32'h3a02ee40),
	.w4(32'h3913df30),
	.w5(32'hba026702),
	.w6(32'h3a446325),
	.w7(32'h3907b352),
	.w8(32'hb9f89333),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd6a36),
	.w1(32'hbbc82104),
	.w2(32'hbb9a6399),
	.w3(32'hbbaa74fd),
	.w4(32'hbb86b147),
	.w5(32'hbb819f05),
	.w6(32'hbb55f81a),
	.w7(32'hbb191fc2),
	.w8(32'hbb60d8e9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03488),
	.w1(32'hba24f61f),
	.w2(32'hba8b6b78),
	.w3(32'hb967e464),
	.w4(32'h3a7bad0d),
	.w5(32'h3a0bcdd1),
	.w6(32'hba9b2eb9),
	.w7(32'hbadb5301),
	.w8(32'hba0ccb80),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a354abf),
	.w1(32'h39a911d1),
	.w2(32'h395e1d09),
	.w3(32'h3a38c9c7),
	.w4(32'h392f24f2),
	.w5(32'h399727cd),
	.w6(32'h3a1e7820),
	.w7(32'h39626455),
	.w8(32'hb981e2b1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d52fc7),
	.w1(32'hb7acc74c),
	.w2(32'h3533ce08),
	.w3(32'hb8044a9f),
	.w4(32'hb81e33c1),
	.w5(32'hb7e868dd),
	.w6(32'hb82982a3),
	.w7(32'hb80b01b3),
	.w8(32'hb7f8dfb4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e63821),
	.w1(32'hb9cb9bac),
	.w2(32'hb91d9528),
	.w3(32'hba27871d),
	.w4(32'hb9ee1096),
	.w5(32'hb9705492),
	.w6(32'hba45a23c),
	.w7(32'hb9ac3d56),
	.w8(32'hb8d2dd10),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eb6703),
	.w1(32'h37b8fcb1),
	.w2(32'h3785c2c8),
	.w3(32'h379c9cab),
	.w4(32'h379c7cd9),
	.w5(32'h373efcd2),
	.w6(32'h37f1b81c),
	.w7(32'h381c4c51),
	.w8(32'h38212af0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a90e7),
	.w1(32'hba24e022),
	.w2(32'hb9c50d24),
	.w3(32'h399d69e4),
	.w4(32'h38b55969),
	.w5(32'hb8dde827),
	.w6(32'h397a4ee7),
	.w7(32'h39c36676),
	.w8(32'h3756b15f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a429dbd),
	.w1(32'h3966cbae),
	.w2(32'hb9dadeef),
	.w3(32'h3a29334b),
	.w4(32'h382085b4),
	.w5(32'hb705f5b3),
	.w6(32'h3a7d9846),
	.w7(32'hb9d287f0),
	.w8(32'hba4010c0),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8ceed),
	.w1(32'hb9f58d50),
	.w2(32'hb9f3c52d),
	.w3(32'hba32d5fb),
	.w4(32'h38cde76b),
	.w5(32'hb9d724de),
	.w6(32'hba9c343a),
	.w7(32'h3724a015),
	.w8(32'h39fdedaa),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4fa91),
	.w1(32'hb995e1b5),
	.w2(32'hb894092d),
	.w3(32'hb92f782d),
	.w4(32'hb91ae506),
	.w5(32'hb7c5a168),
	.w6(32'h3831c3d5),
	.w7(32'h3899b22d),
	.w8(32'h376d85cc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92a1fa),
	.w1(32'hbb1208db),
	.w2(32'hbb1b5238),
	.w3(32'hbaa48a71),
	.w4(32'hbac9b093),
	.w5(32'hbaf78253),
	.w6(32'hba252421),
	.w7(32'hba675d73),
	.w8(32'hba9886da),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991c28),
	.w1(32'hb9c667b0),
	.w2(32'hb97ef940),
	.w3(32'h398cd32e),
	.w4(32'hb908a9ef),
	.w5(32'hb9d74274),
	.w6(32'hb985e161),
	.w7(32'hb82f2a22),
	.w8(32'hb8f9f1ff),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb48a5e64),
	.w1(32'hb705458c),
	.w2(32'h374764bc),
	.w3(32'hb74f13d8),
	.w4(32'hb77b6286),
	.w5(32'h36fa6d2b),
	.w6(32'hb69e0df5),
	.w7(32'h36f8c014),
	.w8(32'h37d24be4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e6fb1b),
	.w1(32'hb8504ee0),
	.w2(32'hba2bcd41),
	.w3(32'hb9921313),
	.w4(32'hb911bc4b),
	.w5(32'hba1c7997),
	.w6(32'hb94d4e86),
	.w7(32'h3865a5be),
	.w8(32'hb881636f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364d5468),
	.w1(32'h372d008a),
	.w2(32'h37a579d5),
	.w3(32'h368139ad),
	.w4(32'hb7588200),
	.w5(32'h36858391),
	.w6(32'h3871d76b),
	.w7(32'h381c3acc),
	.w8(32'h3818a510),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2189b8),
	.w1(32'hba35f27a),
	.w2(32'hba69e70d),
	.w3(32'hb8445f2f),
	.w4(32'h393a0610),
	.w5(32'hb7b0d643),
	.w6(32'h390bc3d2),
	.w7(32'h39899525),
	.w8(32'h383c38be),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f25d9),
	.w1(32'h3a5b6a32),
	.w2(32'h39f28e65),
	.w3(32'h3a8c4cd4),
	.w4(32'h3add308d),
	.w5(32'h3af447bc),
	.w6(32'hb815396e),
	.w7(32'h39ad1390),
	.w8(32'h3a719c08),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981316c),
	.w1(32'hb9428a8f),
	.w2(32'hba13a339),
	.w3(32'h39e05210),
	.w4(32'h39e9f0c3),
	.w5(32'hb99c6f49),
	.w6(32'h38c95a0f),
	.w7(32'h39846f5d),
	.w8(32'hb919baf7),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b9429),
	.w1(32'h399cc769),
	.w2(32'h3968297e),
	.w3(32'h3a02fd83),
	.w4(32'hb7e10e15),
	.w5(32'h3920a837),
	.w6(32'h398ad86d),
	.w7(32'hb9fe2c92),
	.w8(32'hb9baa5f5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827639),
	.w1(32'hba349c15),
	.w2(32'hba5fbb68),
	.w3(32'h38229046),
	.w4(32'h39b16523),
	.w5(32'hb972cc8d),
	.w6(32'hb9c56869),
	.w7(32'h391e9b95),
	.w8(32'h394fb47d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaeb6f),
	.w1(32'hbb0484e0),
	.w2(32'hba47f954),
	.w3(32'hbab8bf3b),
	.w4(32'hbaa675cb),
	.w5(32'hba549a5b),
	.w6(32'hbac04162),
	.w7(32'hba521d7a),
	.w8(32'hb9aa4c8f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaf4a2),
	.w1(32'hba7e522b),
	.w2(32'hba818b10),
	.w3(32'hbb114c21),
	.w4(32'hbab87686),
	.w5(32'hba658995),
	.w6(32'hbaa9334a),
	.w7(32'hbaa333d3),
	.w8(32'hbaa3da6d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3835b8b8),
	.w1(32'h3796ed55),
	.w2(32'h37d97283),
	.w3(32'h37e532b1),
	.w4(32'h378148dd),
	.w5(32'h37f3db3a),
	.w6(32'h36fbdc09),
	.w7(32'hb6ed2562),
	.w8(32'h37376723),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3702e603),
	.w1(32'h37804c5a),
	.w2(32'h3656220e),
	.w3(32'h369f75fe),
	.w4(32'hb70cc517),
	.w5(32'h35de9759),
	.w6(32'h387230ca),
	.w7(32'hb57de9cf),
	.w8(32'h36871a00),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f4df1b),
	.w1(32'hb82a917a),
	.w2(32'h3a615f94),
	.w3(32'h3ace2f65),
	.w4(32'h3a3599a1),
	.w5(32'h3a0852f0),
	.w6(32'h390c6485),
	.w7(32'h3a55cd90),
	.w8(32'h39aa6933),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fc13d),
	.w1(32'hbb15fd6f),
	.w2(32'hba544d08),
	.w3(32'hba91790a),
	.w4(32'h3a8cf3e0),
	.w5(32'h390c9627),
	.w6(32'hbaa1d132),
	.w7(32'h3b0fe162),
	.w8(32'h3a1d4818),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf8274),
	.w1(32'hb9db43fe),
	.w2(32'h3959e951),
	.w3(32'hba826f20),
	.w4(32'hb9cadaf0),
	.w5(32'h39029546),
	.w6(32'hbac441be),
	.w7(32'hb981d10f),
	.w8(32'h39c413f6),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91aec0),
	.w1(32'hb9af84aa),
	.w2(32'hba57cae7),
	.w3(32'h39c91e76),
	.w4(32'h398016c4),
	.w5(32'h3a33bcc1),
	.w6(32'h3a29831b),
	.w7(32'hba7461c7),
	.w8(32'hba213149),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967bde0),
	.w1(32'hb801d548),
	.w2(32'hb897f1b6),
	.w3(32'h34a095c7),
	.w4(32'h391eeea8),
	.w5(32'hb9446d2d),
	.w6(32'hb806e155),
	.w7(32'hb82a8dcd),
	.w8(32'hb8492b04),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c503d),
	.w1(32'hba0a58de),
	.w2(32'hb9c41899),
	.w3(32'hba538fa1),
	.w4(32'hba31ff0c),
	.w5(32'hb97f1f06),
	.w6(32'hba0a2145),
	.w7(32'hb98be4a7),
	.w8(32'hb851ba06),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6da900),
	.w1(32'h3a1440a2),
	.w2(32'h3a801921),
	.w3(32'h3b0cb403),
	.w4(32'h3a841ec8),
	.w5(32'hb8d15088),
	.w6(32'h3ab63afd),
	.w7(32'h3abfe04d),
	.w8(32'h3af0057a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165a1a),
	.w1(32'hbb7ddc47),
	.w2(32'hbb4c4b16),
	.w3(32'hbb198fb0),
	.w4(32'hbb4d743c),
	.w5(32'hbb165405),
	.w6(32'h37808713),
	.w7(32'hbb16f8ff),
	.w8(32'hbb1bc7dd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4c78a),
	.w1(32'h38024785),
	.w2(32'h397e4262),
	.w3(32'h3b0948c0),
	.w4(32'hb957badb),
	.w5(32'hba7d39b9),
	.w6(32'h3a933ea0),
	.w7(32'h3a3189eb),
	.w8(32'hba107fec),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f30c1b),
	.w1(32'h3958d60d),
	.w2(32'h39f43fe5),
	.w3(32'h397c3259),
	.w4(32'h3a4142a3),
	.w5(32'h3a50936e),
	.w6(32'hb9270e43),
	.w7(32'h393dc07b),
	.w8(32'h3a82e18d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb467584),
	.w1(32'hba5959cc),
	.w2(32'h38e78391),
	.w3(32'hbb23c743),
	.w4(32'hb943f11b),
	.w5(32'h3a59bf91),
	.w6(32'hbb3960d7),
	.w7(32'hbabebe82),
	.w8(32'h39f4c869),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f2b027),
	.w1(32'h37a58add),
	.w2(32'h37adc2c2),
	.w3(32'h37a0be25),
	.w4(32'h376820aa),
	.w5(32'h374fd760),
	.w6(32'h37e6b2d5),
	.w7(32'h3752c369),
	.w8(32'h37906511),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374a1d21),
	.w1(32'h37073d2a),
	.w2(32'h379ef77a),
	.w3(32'h36e70257),
	.w4(32'hb548f0fd),
	.w5(32'h373596e3),
	.w6(32'h376527d6),
	.w7(32'h36d7a122),
	.w8(32'h374f2fcb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385451ee),
	.w1(32'hb948a143),
	.w2(32'hb8b062af),
	.w3(32'hb8096cb3),
	.w4(32'h37be2dc1),
	.w5(32'h384b8a5a),
	.w6(32'h393f75f9),
	.w7(32'h37e0618d),
	.w8(32'hb6c5ab8a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77ecef6),
	.w1(32'hb7e8eb6f),
	.w2(32'hb7721dd8),
	.w3(32'hb7a66aba),
	.w4(32'hb7e972fe),
	.w5(32'hb7a03dcd),
	.w6(32'hb5dd735f),
	.w7(32'hb6b5cff1),
	.w8(32'h375e345f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04f7d0),
	.w1(32'h3a0644bb),
	.w2(32'h39d7f415),
	.w3(32'h3a125213),
	.w4(32'h39aa963e),
	.w5(32'h3912aca1),
	.w6(32'h39fb1e7e),
	.w7(32'h394b8bf3),
	.w8(32'hb9061aed),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2b47),
	.w1(32'hbb20e00e),
	.w2(32'h3795acbb),
	.w3(32'h38e3337a),
	.w4(32'hb7d31dbb),
	.w5(32'hba422006),
	.w6(32'hba56a6e7),
	.w7(32'hb9743fa3),
	.w8(32'h39bfbd5a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f22f52),
	.w1(32'hb94ec788),
	.w2(32'hb9a6b6f8),
	.w3(32'hb8f71815),
	.w4(32'h3910c17c),
	.w5(32'h387f463c),
	.w6(32'hb9f882bf),
	.w7(32'h3845d0ed),
	.w8(32'h382eba61),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386d564a),
	.w1(32'h3837240c),
	.w2(32'h3865b231),
	.w3(32'h3826f9b6),
	.w4(32'h38032c1d),
	.w5(32'h3816f21b),
	.w6(32'h3842be27),
	.w7(32'h37fada8c),
	.w8(32'h3841c4ca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea84fa),
	.w1(32'hba7a9ac0),
	.w2(32'hb63e5a37),
	.w3(32'h3ab00165),
	.w4(32'hba9c2544),
	.w5(32'hba85eaeb),
	.w6(32'h3aabecc4),
	.w7(32'h3948e6ca),
	.w8(32'hba532d4f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bfcdb),
	.w1(32'hba1d5f8e),
	.w2(32'hba231367),
	.w3(32'h3955dc74),
	.w4(32'h3a0ef8bb),
	.w5(32'h39b18445),
	.w6(32'h3aa15add),
	.w7(32'h3a5a7902),
	.w8(32'hb93cbc8a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810875f),
	.w1(32'h38373b09),
	.w2(32'h38330aef),
	.w3(32'hb7dd5817),
	.w4(32'h387e1944),
	.w5(32'h3875c906),
	.w6(32'h376121d4),
	.w7(32'h38869491),
	.w8(32'h38bba539),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a81f94),
	.w1(32'hbaa25c02),
	.w2(32'hba749cd7),
	.w3(32'hba072a62),
	.w4(32'hba83fff0),
	.w5(32'hba589446),
	.w6(32'h39030d96),
	.w7(32'hba1b9928),
	.w8(32'hba6290a5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38237afa),
	.w1(32'h382a9c7a),
	.w2(32'h38ddfaa8),
	.w3(32'h3896740f),
	.w4(32'h38a7816e),
	.w5(32'h38dae1f9),
	.w6(32'h38e663a0),
	.w7(32'h39228e84),
	.w8(32'h395fa009),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd8f96),
	.w1(32'h3a08c5e3),
	.w2(32'h39e97ff5),
	.w3(32'h3a10ea4c),
	.w4(32'h3a26e84d),
	.w5(32'h3a1b8f16),
	.w6(32'h39570284),
	.w7(32'h39e27568),
	.w8(32'h39f0d4bc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e2525d),
	.w1(32'hb6a2a499),
	.w2(32'h37208a06),
	.w3(32'h3828906b),
	.w4(32'h37356b98),
	.w5(32'h36d494af),
	.w6(32'h38339e29),
	.w7(32'h38112241),
	.w8(32'h37b5eb00),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c4e4bb),
	.w1(32'h3840cccb),
	.w2(32'h38752ce1),
	.w3(32'h388ba9b8),
	.w4(32'h381f019f),
	.w5(32'h3857a2dc),
	.w6(32'h389cc27d),
	.w7(32'h38521732),
	.w8(32'h388884d4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f774d),
	.w1(32'hb890d271),
	.w2(32'h3a1e718a),
	.w3(32'hba48dbcb),
	.w4(32'h3789f735),
	.w5(32'h39d8d5d1),
	.w6(32'hbaa09307),
	.w7(32'hba0390aa),
	.w8(32'h39fda4e4),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac38b32),
	.w1(32'hba0eb1a7),
	.w2(32'hba470f42),
	.w3(32'hbad9e7ca),
	.w4(32'h39ac9a03),
	.w5(32'h391e7342),
	.w6(32'hbab94e28),
	.w7(32'hba155647),
	.w8(32'hb9ec7a70),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4d57),
	.w1(32'hbb342da6),
	.w2(32'hbafc56c5),
	.w3(32'hbae3a249),
	.w4(32'hba99b034),
	.w5(32'hba7e8f85),
	.w6(32'hba62990b),
	.w7(32'hb9af3942),
	.w8(32'hba15ddf1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae002d7),
	.w1(32'hbae5d651),
	.w2(32'hba1f3458),
	.w3(32'hbaf3840f),
	.w4(32'hba654c32),
	.w5(32'h394f1eda),
	.w6(32'hbac6e4b6),
	.w7(32'hba92efa8),
	.w8(32'hba1cb69f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0439e),
	.w1(32'h39d579e5),
	.w2(32'h39d82076),
	.w3(32'h39b9cb8f),
	.w4(32'h39e2566f),
	.w5(32'h39cf2b07),
	.w6(32'h396dc8a6),
	.w7(32'h398b7505),
	.w8(32'h398cd07b),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917e8ff),
	.w1(32'h383d51d3),
	.w2(32'h370940ca),
	.w3(32'h387b5a3e),
	.w4(32'hb8f58984),
	.w5(32'hb91817ce),
	.w6(32'h37e06075),
	.w7(32'hb90eab78),
	.w8(32'hb956d0cb),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6a00c),
	.w1(32'hb8924b08),
	.w2(32'hb82ce2a9),
	.w3(32'hb870d4e7),
	.w4(32'hb8650342),
	.w5(32'hb837eb4c),
	.w6(32'hb8688870),
	.w7(32'hb882851c),
	.w8(32'hb7c43d06),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772ee13),
	.w1(32'h342281c2),
	.w2(32'hb835d061),
	.w3(32'h38994bfe),
	.w4(32'h38664254),
	.w5(32'h3748a782),
	.w6(32'h387c0ea8),
	.w7(32'h3824f0cc),
	.w8(32'hb3d4b824),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbd60c),
	.w1(32'hba213e39),
	.w2(32'hbaaf36ce),
	.w3(32'hb9c21c0a),
	.w4(32'hba20d32a),
	.w5(32'hbaae8480),
	.w6(32'hb98df900),
	.w7(32'hba4e6564),
	.w8(32'hbab46b81),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8dfcd),
	.w1(32'hb9b92736),
	.w2(32'hb8881fd2),
	.w3(32'hba184a2c),
	.w4(32'hb9eda99a),
	.w5(32'hb99e8902),
	.w6(32'hba2e6407),
	.w7(32'hba09f20d),
	.w8(32'hb9bae561),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10298),
	.w1(32'h39d54a80),
	.w2(32'hb8ccc826),
	.w3(32'h3a836cbf),
	.w4(32'h39ba4f7d),
	.w5(32'hb742e5c8),
	.w6(32'h3a1e954c),
	.w7(32'h390e54de),
	.w8(32'hb9d723de),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d94b8e),
	.w1(32'h399e13e6),
	.w2(32'hb9685734),
	.w3(32'h39e87715),
	.w4(32'hb90c29b2),
	.w5(32'hb9f58d40),
	.w6(32'h3929bd5b),
	.w7(32'hb9356215),
	.w8(32'hb94c9df1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9660652),
	.w1(32'hb8f4b9e8),
	.w2(32'hb7efefef),
	.w3(32'hb981b14b),
	.w4(32'hb910fbc6),
	.w5(32'hb88b22f0),
	.w6(32'hb97f4655),
	.w7(32'hb8b2fd28),
	.w8(32'hb82d99ed),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f43e94),
	.w1(32'hb9c559bb),
	.w2(32'hb9a78460),
	.w3(32'h382ed6fa),
	.w4(32'hba00afe7),
	.w5(32'hb9f4e2d8),
	.w6(32'h388fd46f),
	.w7(32'hb9e050c9),
	.w8(32'hb9f8541b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3825a990),
	.w1(32'h395dbd84),
	.w2(32'h39271cec),
	.w3(32'h3953355e),
	.w4(32'h39469b05),
	.w5(32'h388078d9),
	.w6(32'h39761fd0),
	.w7(32'h3920512e),
	.w8(32'h371bd30e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b91f5),
	.w1(32'hba434345),
	.w2(32'hbac4652d),
	.w3(32'hbacd9b6f),
	.w4(32'hba6a2cfd),
	.w5(32'hbabb7273),
	.w6(32'hba516bbb),
	.w7(32'hbb63824b),
	.w8(32'hbb24eb17),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364f60c9),
	.w1(32'h38f0c7c9),
	.w2(32'h392844a5),
	.w3(32'hb6ffc81f),
	.w4(32'h3858da7c),
	.w5(32'h38c72e88),
	.w6(32'h388fe8fe),
	.w7(32'h3866c956),
	.w8(32'h38b2b250),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3b59),
	.w1(32'hbabe798e),
	.w2(32'h393af866),
	.w3(32'h3978a334),
	.w4(32'h399561c4),
	.w5(32'hb8c1b43a),
	.w6(32'h39d20fc8),
	.w7(32'h3a574f6c),
	.w8(32'h3a4972cc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule