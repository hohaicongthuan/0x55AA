module layer_10_featuremap_106(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94892a9),
	.w1(32'hb9fa9bb5),
	.w2(32'h39ae0c71),
	.w3(32'hb9b27a63),
	.w4(32'h3a5b695c),
	.w5(32'h39956cca),
	.w6(32'h396eca6b),
	.w7(32'h397a6f7b),
	.w8(32'hb989d7d1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61528a),
	.w1(32'h38c68e89),
	.w2(32'hb99f7fcf),
	.w3(32'h3a4cbd5f),
	.w4(32'hba3cd643),
	.w5(32'hb9406737),
	.w6(32'hb9b01db1),
	.w7(32'hb9ad8e72),
	.w8(32'hb8a6154f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02a5ee),
	.w1(32'h37eaa7df),
	.w2(32'h38b987bc),
	.w3(32'h39970161),
	.w4(32'hb9b508a2),
	.w5(32'hb91c16cf),
	.w6(32'hb9b501f3),
	.w7(32'hb8de79a7),
	.w8(32'hb82f4501),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b4784),
	.w1(32'hbab8260a),
	.w2(32'hbab553ac),
	.w3(32'hb9ac89f3),
	.w4(32'hba80c0ef),
	.w5(32'hba739ea5),
	.w6(32'h3a153e98),
	.w7(32'h399fde8c),
	.w8(32'h3a5a39ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d4ecd),
	.w1(32'hb9585120),
	.w2(32'h390319e5),
	.w3(32'hba742f3e),
	.w4(32'hb93ccfaa),
	.w5(32'hb9068c62),
	.w6(32'hb9c8f808),
	.w7(32'hb9d993b8),
	.w8(32'hb9094dfc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372e00bd),
	.w1(32'hb9062ac5),
	.w2(32'h389de7fa),
	.w3(32'hb9221db0),
	.w4(32'hb9821a80),
	.w5(32'hb8d475cc),
	.w6(32'hb9887d11),
	.w7(32'hb8b1f3f6),
	.w8(32'hb83d5cc9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4c162),
	.w1(32'hba633109),
	.w2(32'h3aaecf91),
	.w3(32'hbb5902b6),
	.w4(32'hba21e8ad),
	.w5(32'h3b0d5980),
	.w6(32'hbac475fb),
	.w7(32'h3aa08071),
	.w8(32'h3b2cfa0f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839219),
	.w1(32'h3b4f3711),
	.w2(32'h3b2d8e8e),
	.w3(32'h3b7c709e),
	.w4(32'h3b39cc0b),
	.w5(32'h3a61e83c),
	.w6(32'h3b8f5721),
	.w7(32'h3b8dd518),
	.w8(32'h3b4ea33f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39957533),
	.w1(32'h3a80303b),
	.w2(32'h3ae5710c),
	.w3(32'h3a2f7911),
	.w4(32'h3aac2039),
	.w5(32'h3b022805),
	.w6(32'h3a9e038a),
	.w7(32'h3b0b6b3b),
	.w8(32'h3b088c25),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c27da),
	.w1(32'h3b47a584),
	.w2(32'h3a9e3395),
	.w3(32'h3ae8bbed),
	.w4(32'h3a5b546c),
	.w5(32'h39833d2c),
	.w6(32'h3b48632f),
	.w7(32'h39af81ea),
	.w8(32'h3a504915),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b007d07),
	.w1(32'hba15b8ae),
	.w2(32'hbae5acc0),
	.w3(32'h3b23efff),
	.w4(32'h39b3989c),
	.w5(32'hbab5073f),
	.w6(32'hb938100c),
	.w7(32'h39a30536),
	.w8(32'hbac9387c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43df59),
	.w1(32'hbac75d4d),
	.w2(32'h3ad0a895),
	.w3(32'hbbb5f951),
	.w4(32'hbaed726a),
	.w5(32'h3aca9985),
	.w6(32'hbaf3364e),
	.w7(32'hba801820),
	.w8(32'h3b184c91),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa43208),
	.w1(32'h3aa47186),
	.w2(32'h3a9ae1de),
	.w3(32'hba1c72c3),
	.w4(32'h39010975),
	.w5(32'h3a823d3f),
	.w6(32'hba5b35c7),
	.w7(32'h39f1aef0),
	.w8(32'h3af15ef2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38895001),
	.w1(32'h3a287311),
	.w2(32'hb9b09326),
	.w3(32'h3a59e4c3),
	.w4(32'h3a85c7a1),
	.w5(32'hb99c7daf),
	.w6(32'h3a6e9c8b),
	.w7(32'h3a3c2418),
	.w8(32'hb97b5020),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4717e),
	.w1(32'hba77e35b),
	.w2(32'hbabe130d),
	.w3(32'hba6076c1),
	.w4(32'hb9fa31da),
	.w5(32'hba942746),
	.w6(32'h39324714),
	.w7(32'hb9ce83ba),
	.w8(32'hba8f5bb6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0320e3),
	.w1(32'h3af5ae72),
	.w2(32'h392c7212),
	.w3(32'h39bd4efb),
	.w4(32'h3a813ea9),
	.w5(32'hba3cba39),
	.w6(32'h3ad9efa8),
	.w7(32'h3b00f4c7),
	.w8(32'h39a5edb2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f4d3b),
	.w1(32'hb8fae631),
	.w2(32'hb9a29593),
	.w3(32'h3989d9da),
	.w4(32'hb997e7fd),
	.w5(32'hba8dcb9b),
	.w6(32'h395511af),
	.w7(32'hb93dd4be),
	.w8(32'hbab7d2f7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950e24c),
	.w1(32'h3b31b555),
	.w2(32'h3b984b17),
	.w3(32'h3b1d3e72),
	.w4(32'h3b951fc0),
	.w5(32'h3b281e9f),
	.w6(32'h3bb19d16),
	.w7(32'h3bea591b),
	.w8(32'h3bb7444c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed7fa8),
	.w1(32'h398f1b30),
	.w2(32'h3ad0a11e),
	.w3(32'h39f9fea0),
	.w4(32'h3a94d963),
	.w5(32'h3adb32d2),
	.w6(32'h3af9babe),
	.w7(32'h3b36810e),
	.w8(32'h3b3bb9fb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387a1043),
	.w1(32'h38f32e7e),
	.w2(32'h387e7e2a),
	.w3(32'h38c6cf8a),
	.w4(32'hb7ffb0cf),
	.w5(32'h3806f1e4),
	.w6(32'hb8b49253),
	.w7(32'hb8a6116b),
	.w8(32'h37b57592),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b9079d),
	.w1(32'h372f74b8),
	.w2(32'hb88ad119),
	.w3(32'hb91259ac),
	.w4(32'h383f1a93),
	.w5(32'hb87cd92a),
	.w6(32'h392e090b),
	.w7(32'h39334cba),
	.w8(32'h398a34d0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3892fe36),
	.w1(32'hb9d93fb2),
	.w2(32'hb9a50c7c),
	.w3(32'hb9c5284f),
	.w4(32'hb98d24de),
	.w5(32'h376580f6),
	.w6(32'hba74d655),
	.w7(32'hba542c0d),
	.w8(32'hba225646),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80880d),
	.w1(32'h3b193fa4),
	.w2(32'h3c110853),
	.w3(32'h3a8fbfd4),
	.w4(32'h3ad9b6b3),
	.w5(32'h3c021be2),
	.w6(32'h3b576e3e),
	.w7(32'h3bfd0002),
	.w8(32'h3c14edda),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0401),
	.w1(32'h3ae8eaeb),
	.w2(32'h39521065),
	.w3(32'h39320ff5),
	.w4(32'hba8a4ab7),
	.w5(32'hba55011b),
	.w6(32'hb80d905e),
	.w7(32'hba153b8a),
	.w8(32'h3908fcbd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ec640),
	.w1(32'h3b0960c0),
	.w2(32'h3a7bdaf4),
	.w3(32'h37dab094),
	.w4(32'h3a13c80d),
	.w5(32'hba84c947),
	.w6(32'hba4f098b),
	.w7(32'h3abc70de),
	.w8(32'hbadf8eb8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29695f),
	.w1(32'hb9c33c74),
	.w2(32'hba7024f7),
	.w3(32'h3a57c118),
	.w4(32'hba31f1a2),
	.w5(32'hba17bdc1),
	.w6(32'h398ecd5c),
	.w7(32'hb9b53536),
	.w8(32'hb99525bd),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14e662),
	.w1(32'hb8bed7ad),
	.w2(32'hb93f2fd8),
	.w3(32'hb992cc2f),
	.w4(32'hb8fb0958),
	.w5(32'hb99c30e8),
	.w6(32'hb98339f0),
	.w7(32'hb9726958),
	.w8(32'hb9ae5b18),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39669637),
	.w1(32'hb8f52a28),
	.w2(32'hbabee2d7),
	.w3(32'hba6958f3),
	.w4(32'hbb0f8998),
	.w5(32'hbb2648db),
	.w6(32'hbaf27119),
	.w7(32'hbb2bcc6d),
	.w8(32'hbb3db432),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76b3f),
	.w1(32'hba6e0e89),
	.w2(32'hbad6febb),
	.w3(32'hb998c97e),
	.w4(32'hbaafcf46),
	.w5(32'hbb30c329),
	.w6(32'h38ba2355),
	.w7(32'hbacb8227),
	.w8(32'hbb444ed5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b150283),
	.w1(32'h3958f6b0),
	.w2(32'hbaa934fa),
	.w3(32'h399772c4),
	.w4(32'hbb3bf871),
	.w5(32'hba6730ec),
	.w6(32'hbb0691aa),
	.w7(32'hbb3b86e3),
	.w8(32'hba3b6d68),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a080fe),
	.w1(32'hb9780f51),
	.w2(32'hb9808d7f),
	.w3(32'hb8890c80),
	.w4(32'hb96200dd),
	.w5(32'hb98839a5),
	.w6(32'hb92b8653),
	.w7(32'hb936ba4a),
	.w8(32'hb950db8d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e668e),
	.w1(32'h39d8bbcd),
	.w2(32'hb964a57e),
	.w3(32'h39cad97c),
	.w4(32'h38a5f674),
	.w5(32'hba77fb0d),
	.w6(32'h3a1ae21a),
	.w7(32'hb9550180),
	.w8(32'hba97326d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9449fc0),
	.w1(32'hb9cb3c77),
	.w2(32'hba186929),
	.w3(32'hb910d91c),
	.w4(32'hba2917b8),
	.w5(32'hba7ff4c7),
	.w6(32'h37edf686),
	.w7(32'hba324409),
	.w8(32'hba253fc2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1e92e),
	.w1(32'h3a740244),
	.w2(32'h3890b899),
	.w3(32'h39d19692),
	.w4(32'h39d9c935),
	.w5(32'h3a4d3372),
	.w6(32'h39e6516b),
	.w7(32'hb7b5a344),
	.w8(32'h3a4b185c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92908ff),
	.w1(32'h3a09aef2),
	.w2(32'h399bdeed),
	.w3(32'hba3a1ab2),
	.w4(32'h38920193),
	.w5(32'h3984125f),
	.w6(32'h3a049929),
	.w7(32'h3a2466f8),
	.w8(32'h3a433c14),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994f3a3),
	.w1(32'hba04b132),
	.w2(32'h3a3986f6),
	.w3(32'h398c523a),
	.w4(32'h39941935),
	.w5(32'h3a3ed5d1),
	.w6(32'hba13bf38),
	.w7(32'h37addfc2),
	.w8(32'h3a999221),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52dab7),
	.w1(32'hbb17be16),
	.w2(32'h3b7990f9),
	.w3(32'h3a927e0c),
	.w4(32'hbb1e5789),
	.w5(32'h3a6529ae),
	.w6(32'h3ba95d18),
	.w7(32'hbb030605),
	.w8(32'h3b8f03a1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba96e8a),
	.w1(32'hba8c067d),
	.w2(32'hbb4aa77a),
	.w3(32'h3a88a0dd),
	.w4(32'hbb91cb9e),
	.w5(32'hbb4277f8),
	.w6(32'hb99cbb28),
	.w7(32'hbbac0348),
	.w8(32'hbb436490),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17dfdb),
	.w1(32'hbb5730f7),
	.w2(32'hbbacc241),
	.w3(32'hbaa4de91),
	.w4(32'hbbc30d22),
	.w5(32'hbb855616),
	.w6(32'hbb6552eb),
	.w7(32'hbbbd0586),
	.w8(32'hbb2080de),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00134a),
	.w1(32'hb98590c1),
	.w2(32'hb9ec2fa1),
	.w3(32'hba9846cf),
	.w4(32'hba793611),
	.w5(32'hba273823),
	.w6(32'hba042a3a),
	.w7(32'hba5ed649),
	.w8(32'hba1c0985),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776956),
	.w1(32'h39fd2352),
	.w2(32'h39b54eb3),
	.w3(32'h3a8d06b7),
	.w4(32'h399e0ce2),
	.w5(32'h39d7f703),
	.w6(32'h3a387233),
	.w7(32'h37fbaad5),
	.w8(32'h3986ad22),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba323974),
	.w1(32'hb94264f9),
	.w2(32'h39e30362),
	.w3(32'hba83b790),
	.w4(32'hba2594f2),
	.w5(32'h3989af26),
	.w6(32'hba83f042),
	.w7(32'h3802e355),
	.w8(32'h3a589241),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbe08a),
	.w1(32'h3983a9e7),
	.w2(32'hba62b892),
	.w3(32'hb99c7226),
	.w4(32'hb963849a),
	.w5(32'hba98c9b2),
	.w6(32'h3a882344),
	.w7(32'h38fadf83),
	.w8(32'hba811e87),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf53de),
	.w1(32'h3b7776aa),
	.w2(32'h3b92c173),
	.w3(32'h3b236892),
	.w4(32'h3a9d38c2),
	.w5(32'h3bc325a9),
	.w6(32'h3b72d8bf),
	.w7(32'h3b15056b),
	.w8(32'h3bbeb354),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61bec5),
	.w1(32'h3a7a6837),
	.w2(32'h3961141c),
	.w3(32'h3a8ee026),
	.w4(32'hbb1e33bf),
	.w5(32'hba321cbc),
	.w6(32'hb89fc33e),
	.w7(32'hbb07c292),
	.w8(32'h3a559478),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f68af),
	.w1(32'h3ad81228),
	.w2(32'h3a33a87c),
	.w3(32'hba54d557),
	.w4(32'hbb22f2a2),
	.w5(32'h3a9be075),
	.w6(32'hbac18a69),
	.w7(32'hbab57e8f),
	.w8(32'h3b328ac2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a962df3),
	.w1(32'h3a844354),
	.w2(32'h3abfcbe8),
	.w3(32'hbad1a2e5),
	.w4(32'hbafbb0cf),
	.w5(32'h3b38289a),
	.w6(32'h3a192f45),
	.w7(32'h3a256337),
	.w8(32'h3bbde9ef),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6667da),
	.w1(32'h3b1263a6),
	.w2(32'h3c0610a7),
	.w3(32'h3a51603a),
	.w4(32'h3b9091fd),
	.w5(32'h3bca9c47),
	.w6(32'h3b9bdd0d),
	.w7(32'h3c029a09),
	.w8(32'h3beb572d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a5596),
	.w1(32'h3aa9f041),
	.w2(32'h3ac0e793),
	.w3(32'h3a472877),
	.w4(32'h398f6865),
	.w5(32'h3ad7f9fb),
	.w6(32'h38d9a0f7),
	.w7(32'hb977c82c),
	.w8(32'h3af286f9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98adc15),
	.w1(32'h3a4ad16b),
	.w2(32'h3b30d978),
	.w3(32'hba6efb4c),
	.w4(32'h39d49b24),
	.w5(32'h3b61f330),
	.w6(32'hbac4ddd1),
	.w7(32'h3ab33d31),
	.w8(32'h3b616e21),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa46654),
	.w1(32'hb9163e1d),
	.w2(32'h3a07ef06),
	.w3(32'hbada3450),
	.w4(32'hba83ecc6),
	.w5(32'h39234de0),
	.w6(32'h375f590b),
	.w7(32'h38ccc77a),
	.w8(32'h393e1ae5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c1a87),
	.w1(32'h3a8628a7),
	.w2(32'h3a63a099),
	.w3(32'hb7e29111),
	.w4(32'h3a21fa47),
	.w5(32'hb717e856),
	.w6(32'h39b67a1e),
	.w7(32'h386d029a),
	.w8(32'h3aa153e9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f5b3b),
	.w1(32'h3a2493d8),
	.w2(32'h3ab32be3),
	.w3(32'h3a08ef9d),
	.w4(32'h39718116),
	.w5(32'h39e7ba60),
	.w6(32'h3a16e5e3),
	.w7(32'h3a4e8f2e),
	.w8(32'h3a2f68fe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6b3a3),
	.w1(32'h3ab4a403),
	.w2(32'h3b7285ad),
	.w3(32'hb84dd228),
	.w4(32'h3b2e4bf3),
	.w5(32'h3b3058ff),
	.w6(32'h3b533965),
	.w7(32'h3b854b78),
	.w8(32'h3b843bce),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57c5d5),
	.w1(32'h3a2a631e),
	.w2(32'h3a469c9e),
	.w3(32'h3a4265ff),
	.w4(32'h3a066129),
	.w5(32'h393d72ca),
	.w6(32'h39890d48),
	.w7(32'h39a16efa),
	.w8(32'h39794b73),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37894b32),
	.w1(32'hb87f9893),
	.w2(32'hb9f29b05),
	.w3(32'h39c33393),
	.w4(32'hb9b822f4),
	.w5(32'hba14117e),
	.w6(32'hb985d125),
	.w7(32'hba436727),
	.w8(32'hb9bf1ed7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b8bf2),
	.w1(32'hb99fe8c4),
	.w2(32'h393261e6),
	.w3(32'hb9cc97c1),
	.w4(32'hba13c726),
	.w5(32'hb9827d9f),
	.w6(32'hb9ebfbc8),
	.w7(32'hb9d8d141),
	.w8(32'hb9b9425e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7593f),
	.w1(32'hb957b8bc),
	.w2(32'h39dc27bf),
	.w3(32'hb96b5efc),
	.w4(32'h38f15f7e),
	.w5(32'h3a1973c5),
	.w6(32'hb90479f8),
	.w7(32'h39dd7818),
	.w8(32'hb9760a11),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3a762),
	.w1(32'hb9d51529),
	.w2(32'hb9818e95),
	.w3(32'hb98d6fab),
	.w4(32'hba51c75d),
	.w5(32'hb9c4a2a1),
	.w6(32'h39cd8878),
	.w7(32'h37954fb6),
	.w8(32'h39d51e0a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9978250),
	.w1(32'hba458206),
	.w2(32'hba52e383),
	.w3(32'h3a0d99fe),
	.w4(32'hb93ae2e6),
	.w5(32'hb859dc9e),
	.w6(32'h38c3af20),
	.w7(32'hb87743e6),
	.w8(32'h395c45bf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c72ff3),
	.w1(32'h3a8fcbc5),
	.w2(32'h3af56a0f),
	.w3(32'h39642c8f),
	.w4(32'h3aa848bf),
	.w5(32'h3ac07888),
	.w6(32'h3aadafe4),
	.w7(32'h3b1d43c9),
	.w8(32'h3b18a3d1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89181f),
	.w1(32'h3afb8812),
	.w2(32'h3a4f4fe8),
	.w3(32'h3b348bd7),
	.w4(32'h3aeb1d33),
	.w5(32'h3a4304e0),
	.w6(32'h3b203f8e),
	.w7(32'h3a857a00),
	.w8(32'h3a89bbd9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fc714),
	.w1(32'h39792959),
	.w2(32'h39e2e507),
	.w3(32'hb914fa74),
	.w4(32'h3a665205),
	.w5(32'h399f43b9),
	.w6(32'h39044338),
	.w7(32'hb97ae1a6),
	.w8(32'hb940cb66),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b06c0c),
	.w1(32'h3a4a28ca),
	.w2(32'h3a2cda8e),
	.w3(32'h3811000d),
	.w4(32'h3a2bb148),
	.w5(32'h3a256f09),
	.w6(32'h3a6770e2),
	.w7(32'h3a2aab3e),
	.w8(32'h3a1178cd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29d6bd),
	.w1(32'hb882b0c0),
	.w2(32'hb9f10224),
	.w3(32'h3a1336b5),
	.w4(32'hb98b0f1f),
	.w5(32'hb958c693),
	.w6(32'hb9582eb3),
	.w7(32'hb901bd96),
	.w8(32'hb8bc2981),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955cc3f),
	.w1(32'h399f0b7c),
	.w2(32'h3a01662f),
	.w3(32'h396bf7ae),
	.w4(32'h3a13cb2d),
	.w5(32'h3a048b13),
	.w6(32'h39b07202),
	.w7(32'h38e11ac3),
	.w8(32'h3873fc94),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df2e76),
	.w1(32'hba18fe58),
	.w2(32'hba8888fa),
	.w3(32'hba80d9b7),
	.w4(32'hbaada701),
	.w5(32'hbaf838a9),
	.w6(32'h3a34417f),
	.w7(32'h39812f7c),
	.w8(32'hbadb3521),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29ea66),
	.w1(32'h3b0d33c4),
	.w2(32'h3a8475f6),
	.w3(32'hb9789b3d),
	.w4(32'h398ebd78),
	.w5(32'h3a90df12),
	.w6(32'hb932165e),
	.w7(32'h3ac0ae35),
	.w8(32'h3b50e870),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a793bec),
	.w1(32'h3b21e52f),
	.w2(32'h3b767a2f),
	.w3(32'h3ae5652d),
	.w4(32'h3ab6aad6),
	.w5(32'h3afd158a),
	.w6(32'h3b333f1e),
	.w7(32'h3b5bd849),
	.w8(32'h3b8c5358),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78f91e),
	.w1(32'h3b08ffe0),
	.w2(32'h3a3b3d6c),
	.w3(32'h3abfd45e),
	.w4(32'hba6f6dcf),
	.w5(32'h3a79964d),
	.w6(32'h3a5c3296),
	.w7(32'hba972f07),
	.w8(32'h3a05b8a2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39402e9c),
	.w1(32'h39dd71e5),
	.w2(32'h3a0c05fb),
	.w3(32'hb707c9e2),
	.w4(32'h390a2897),
	.w5(32'h39874044),
	.w6(32'h398e263e),
	.w7(32'h39b80b09),
	.w8(32'h39e6e766),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0de24a),
	.w1(32'hb98574e3),
	.w2(32'hb93f7b32),
	.w3(32'h396a79a7),
	.w4(32'hb9996486),
	.w5(32'hb99572af),
	.w6(32'hb9a59e77),
	.w7(32'hb96cdbb7),
	.w8(32'hb95949b8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bef96),
	.w1(32'hb9ac9132),
	.w2(32'hb9b12dfe),
	.w3(32'hb9805efe),
	.w4(32'hb9a01996),
	.w5(32'hb9b55778),
	.w6(32'hb9bf7b43),
	.w7(32'hb9bd26e4),
	.w8(32'hb9857e35),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba319ce1),
	.w1(32'h3896cf63),
	.w2(32'h39898204),
	.w3(32'hb9e82635),
	.w4(32'h3a00dc97),
	.w5(32'h38dec52b),
	.w6(32'h3a50ae5d),
	.w7(32'h3a8ad3d8),
	.w8(32'h3a17b083),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3ec4f),
	.w1(32'h3997238b),
	.w2(32'h3a4e743a),
	.w3(32'hba449b0c),
	.w4(32'hb8ffad86),
	.w5(32'h39f75fe2),
	.w6(32'hb9bc3b1d),
	.w7(32'h3965491c),
	.w8(32'h3a86fa97),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382358c2),
	.w1(32'hb995325e),
	.w2(32'h3a9b72a8),
	.w3(32'hba467758),
	.w4(32'h3ac2fdf8),
	.w5(32'h3a8acef8),
	.w6(32'h3abf1b31),
	.w7(32'h3af2cacd),
	.w8(32'h3b1c8e9a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa52ff7),
	.w1(32'hbaea2b5e),
	.w2(32'h3b0532e9),
	.w3(32'hbac26d36),
	.w4(32'h3b4835e2),
	.w5(32'h3affc19f),
	.w6(32'h3b47bcb0),
	.w7(32'h3b7492b5),
	.w8(32'h3b5d9f6d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3bc0a),
	.w1(32'h3a932e37),
	.w2(32'h3aa00209),
	.w3(32'hba3d2557),
	.w4(32'hba21b67e),
	.w5(32'h39a63d7f),
	.w6(32'hba621b0b),
	.w7(32'hba8981ba),
	.w8(32'h39d0a0ba),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a800352),
	.w1(32'h3a80b2ee),
	.w2(32'h3a14a64c),
	.w3(32'h3a51246b),
	.w4(32'h3a0e3a69),
	.w5(32'h39fc27fe),
	.w6(32'h3aacccdd),
	.w7(32'h3ab41fe1),
	.w8(32'h3a7f2b2e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957637c),
	.w1(32'h3a375f6a),
	.w2(32'h3a29bf14),
	.w3(32'hbaa9a81a),
	.w4(32'hba974550),
	.w5(32'h3947b379),
	.w6(32'hb9d40ae8),
	.w7(32'h39c73736),
	.w8(32'h3a41ce97),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6cb72),
	.w1(32'h3a334b5d),
	.w2(32'h35e7acb2),
	.w3(32'h3a81466b),
	.w4(32'hb9380ad6),
	.w5(32'hba12e045),
	.w6(32'h3a5731fc),
	.w7(32'h38f1c941),
	.w8(32'hb9dbb9ce),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b785f),
	.w1(32'h3a003189),
	.w2(32'h3b2c1904),
	.w3(32'hb998cb4e),
	.w4(32'h3a28bc3e),
	.w5(32'h3aa6b714),
	.w6(32'h3a834ecc),
	.w7(32'h3b19a186),
	.w8(32'h3b2b57b6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395970d6),
	.w1(32'h3868627e),
	.w2(32'h38a75457),
	.w3(32'hb79d0c74),
	.w4(32'hb8d12ed8),
	.w5(32'hb794e6cd),
	.w6(32'hb8de9639),
	.w7(32'h38c9d89a),
	.w8(32'h382fadd9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f23d6),
	.w1(32'h390b0322),
	.w2(32'h3993c9ff),
	.w3(32'h38348a25),
	.w4(32'h370323c5),
	.w5(32'hb818e0c3),
	.w6(32'h373cf82e),
	.w7(32'h384ebe4f),
	.w8(32'h382b9abb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395674b1),
	.w1(32'h381c6ff1),
	.w2(32'hba39edea),
	.w3(32'hb8721303),
	.w4(32'hba0f04a5),
	.w5(32'hba2ef31c),
	.w6(32'hba80176f),
	.w7(32'hba8460e1),
	.w8(32'hba82a6e6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92133c7),
	.w1(32'hb9b4bcaa),
	.w2(32'hb8800157),
	.w3(32'hb9f3d0ec),
	.w4(32'hba198128),
	.w5(32'hba092a49),
	.w6(32'hb986e21e),
	.w7(32'hb94065f1),
	.w8(32'hb9f47c4e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a868ca4),
	.w1(32'h39e327dd),
	.w2(32'hbabdeb2d),
	.w3(32'h391899e1),
	.w4(32'hba825048),
	.w5(32'hba9da1e8),
	.w6(32'h3a3f5d24),
	.w7(32'hba8a2986),
	.w8(32'hbaa53e41),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9478813),
	.w1(32'hb7906f4e),
	.w2(32'h38d2786a),
	.w3(32'hb83f807e),
	.w4(32'h37db3dd4),
	.w5(32'h391b36e6),
	.w6(32'h3962baef),
	.w7(32'h38d3741f),
	.w8(32'h38f1eaa5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89c874),
	.w1(32'h3ab4c552),
	.w2(32'h3963d084),
	.w3(32'h357bb6e4),
	.w4(32'hb991f52f),
	.w5(32'hb88a7b37),
	.w6(32'hba02f3bc),
	.w7(32'hb9e528dd),
	.w8(32'h3a0d758d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991093f),
	.w1(32'h3a8f0164),
	.w2(32'h3b9213b2),
	.w3(32'h3b1176ea),
	.w4(32'h3b89b1ad),
	.w5(32'h3b541eda),
	.w6(32'h3bad7a16),
	.w7(32'h3bd91741),
	.w8(32'h3bb1ff45),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae81011),
	.w1(32'hb8230e88),
	.w2(32'hb8950fd2),
	.w3(32'hba166236),
	.w4(32'hbad7410e),
	.w5(32'hbad99424),
	.w6(32'hb9e5597b),
	.w7(32'hba9f7267),
	.w8(32'hbad703d2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399acf31),
	.w1(32'hba86dcfb),
	.w2(32'h3aba15e2),
	.w3(32'hba550356),
	.w4(32'hbb005cfa),
	.w5(32'h3a438b0f),
	.w6(32'h3a36420e),
	.w7(32'h3a055c24),
	.w8(32'h3ab070a2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3e52d),
	.w1(32'h39043a1c),
	.w2(32'hb966689e),
	.w3(32'hba06c798),
	.w4(32'hba934af7),
	.w5(32'hba8b538c),
	.w6(32'hb9c026ba),
	.w7(32'hba8bb640),
	.w8(32'hba2e204c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf2c5),
	.w1(32'h3acd211f),
	.w2(32'h3abee254),
	.w3(32'h3a9afbb9),
	.w4(32'h39f79a44),
	.w5(32'h3a8d1047),
	.w6(32'h3ad55609),
	.w7(32'h3adca215),
	.w8(32'h3b2b1dfc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a864462),
	.w1(32'h3aa4da73),
	.w2(32'h3a31ce21),
	.w3(32'hbabfd69e),
	.w4(32'hba807541),
	.w5(32'hba2e5d5c),
	.w6(32'hbadff59d),
	.w7(32'hba4c4c4c),
	.w8(32'hbaa651f0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5853a),
	.w1(32'h39b09aa1),
	.w2(32'hb9b4f8e8),
	.w3(32'hb9b54040),
	.w4(32'hba804c1f),
	.w5(32'hba758881),
	.w6(32'hba431676),
	.w7(32'hba99f851),
	.w8(32'hbaa1a9c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfa33f),
	.w1(32'h3ac321f9),
	.w2(32'h3b379643),
	.w3(32'h3acda6d5),
	.w4(32'h3b095d9a),
	.w5(32'h3b6ee469),
	.w6(32'h3b0da09e),
	.w7(32'h3b612834),
	.w8(32'h3b603db6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a834a),
	.w1(32'hb9f9d9ec),
	.w2(32'h3b5abb5f),
	.w3(32'hba480fc5),
	.w4(32'hb9f45b62),
	.w5(32'h3bae7c6a),
	.w6(32'h3a376e6f),
	.w7(32'h3b836447),
	.w8(32'h3c10f270),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb464ac9),
	.w1(32'hbb1670c3),
	.w2(32'h3a7ce96a),
	.w3(32'hbbac672f),
	.w4(32'hbb6af587),
	.w5(32'h3a73caba),
	.w6(32'hb9f54227),
	.w7(32'h3abcdb42),
	.w8(32'h3be7a2dd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11e741),
	.w1(32'hba73fce2),
	.w2(32'h3befa320),
	.w3(32'h3b1ebbcc),
	.w4(32'h3afb68f4),
	.w5(32'h3b5b5fdf),
	.w6(32'h3a9d5a62),
	.w7(32'h3b2237cf),
	.w8(32'h3b8b984b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01bd3b),
	.w1(32'hba8fb910),
	.w2(32'h3ab5e91d),
	.w3(32'h3b51097f),
	.w4(32'hbbc0aa87),
	.w5(32'hba3d9f92),
	.w6(32'h3b2e5b72),
	.w7(32'hbb72ab5b),
	.w8(32'h3b11fd6e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29517b),
	.w1(32'h3b1065c9),
	.w2(32'h3ac93e61),
	.w3(32'h396d7912),
	.w4(32'h3b061a03),
	.w5(32'h3b13cc8f),
	.w6(32'hbb10385c),
	.w7(32'hba5e243a),
	.w8(32'h3b18ffe4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80044),
	.w1(32'hbb42315e),
	.w2(32'h3b1e8995),
	.w3(32'hb96f8519),
	.w4(32'hbb7c7917),
	.w5(32'h3b598209),
	.w6(32'h3af58d0e),
	.w7(32'hbb0a0400),
	.w8(32'h3ba20f60),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ea644),
	.w1(32'h3a906510),
	.w2(32'h3b5819a8),
	.w3(32'hba751851),
	.w4(32'hb904d7db),
	.w5(32'h3b41f1f0),
	.w6(32'hba05c182),
	.w7(32'hb800167c),
	.w8(32'h3ba216b6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ef9c2),
	.w1(32'h3b2f2bfb),
	.w2(32'h3be13e0f),
	.w3(32'h3ad535ca),
	.w4(32'h3b15e461),
	.w5(32'h3b879943),
	.w6(32'h3b4e31da),
	.w7(32'h3af1c1ca),
	.w8(32'h3bb8ea53),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba683cdf),
	.w1(32'hba234eda),
	.w2(32'h3a6a2fa4),
	.w3(32'hbaccebf3),
	.w4(32'hbae5012a),
	.w5(32'h3ac54317),
	.w6(32'hbacb888a),
	.w7(32'hbafb2c12),
	.w8(32'h3a1efc34),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966a50a),
	.w1(32'h37d6b5fc),
	.w2(32'h39b8b327),
	.w3(32'hb92c2772),
	.w4(32'hb9a84d23),
	.w5(32'hb831c1fa),
	.w6(32'hb9921853),
	.w7(32'hb6970929),
	.w8(32'h3997c41d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95594e),
	.w1(32'h39c99afa),
	.w2(32'h3790c10d),
	.w3(32'h38c0a811),
	.w4(32'hb9a11019),
	.w5(32'hb9f2e3c3),
	.w6(32'h3a1bcc66),
	.w7(32'h39c8b02e),
	.w8(32'hb92b0394),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94647c1),
	.w1(32'hba2932ad),
	.w2(32'h39ec083a),
	.w3(32'hba520ff6),
	.w4(32'hba54df4c),
	.w5(32'h3b08d427),
	.w6(32'hb9a8a99e),
	.w7(32'hb9db6051),
	.w8(32'h3b546414),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10c571),
	.w1(32'h3a51de8f),
	.w2(32'h3adfef2b),
	.w3(32'hba0032b4),
	.w4(32'hbb354f1b),
	.w5(32'h3ae63c62),
	.w6(32'hbb338a8a),
	.w7(32'hbb358cdb),
	.w8(32'h3ab16152),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1cb29),
	.w1(32'h392fee52),
	.w2(32'h3a814689),
	.w3(32'h396c7543),
	.w4(32'hbaae6459),
	.w5(32'hb9814df2),
	.w6(32'hb9b14920),
	.w7(32'hba59d42d),
	.w8(32'hb98325e9),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4a5f),
	.w1(32'h39c6b636),
	.w2(32'h3ac1c950),
	.w3(32'h3aa84c11),
	.w4(32'h3a1d0c24),
	.w5(32'h3ac13161),
	.w6(32'h3add940c),
	.w7(32'h39d20374),
	.w8(32'h3b522918),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ea6ef),
	.w1(32'hba57c2e9),
	.w2(32'hb9e90f05),
	.w3(32'h3addd596),
	.w4(32'hba4059fc),
	.w5(32'hba7cd718),
	.w6(32'hb8daacf1),
	.w7(32'hbaeb475e),
	.w8(32'hba17d922),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b85e6),
	.w1(32'h3a4f415e),
	.w2(32'h396b81ec),
	.w3(32'h3b4332e7),
	.w4(32'hb907e9e5),
	.w5(32'hb95cfbff),
	.w6(32'h3b369662),
	.w7(32'h3b1df08c),
	.w8(32'hb9530d5d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c34ef),
	.w1(32'h393b51e4),
	.w2(32'hb9a7fdce),
	.w3(32'hb9ab9402),
	.w4(32'hba9d8af2),
	.w5(32'hba34a91a),
	.w6(32'hba1c80e4),
	.w7(32'hba98b71d),
	.w8(32'hb9d824ce),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2da83),
	.w1(32'hb99def03),
	.w2(32'hba2243c7),
	.w3(32'hb91def87),
	.w4(32'hb75c702c),
	.w5(32'hb9822264),
	.w6(32'hb92dbf29),
	.w7(32'hba076ff5),
	.w8(32'hb9f3e960),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e603b6),
	.w1(32'hb96993de),
	.w2(32'hb9d5c5af),
	.w3(32'hb9c5f54b),
	.w4(32'hb9825dac),
	.w5(32'hb9be1f9c),
	.w6(32'hb9af42f3),
	.w7(32'hb9c75de2),
	.w8(32'hb9aebd8c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e70c96),
	.w1(32'hb9a97872),
	.w2(32'hb9e82362),
	.w3(32'hb9d27167),
	.w4(32'hb94e6ed1),
	.w5(32'hb99c9996),
	.w6(32'hb9c8c7e9),
	.w7(32'hb9d28658),
	.w8(32'hb9b0b0fc),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d447b6),
	.w1(32'h389781f9),
	.w2(32'hb85875f7),
	.w3(32'hb9d07caa),
	.w4(32'h3a0ebed1),
	.w5(32'h39e7a0e4),
	.w6(32'h39874afe),
	.w7(32'h393be389),
	.w8(32'h3a16dad6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9647a1),
	.w1(32'hb8c7a699),
	.w2(32'hba81d761),
	.w3(32'h3884b40e),
	.w4(32'hbaeab808),
	.w5(32'hba4740b0),
	.w6(32'hba8d21ae),
	.w7(32'hbaa7fedc),
	.w8(32'hba489f28),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0532af),
	.w1(32'h3871b677),
	.w2(32'h3a180484),
	.w3(32'h3a050089),
	.w4(32'hb9f58334),
	.w5(32'hb894e476),
	.w6(32'h394c7ef2),
	.w7(32'hb918806c),
	.w8(32'h3a54c7eb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c3d8d5),
	.w1(32'h39920010),
	.w2(32'h3acd5cf3),
	.w3(32'hb9c4e366),
	.w4(32'h3a415582),
	.w5(32'h3a97e37d),
	.w6(32'h3a926478),
	.w7(32'h3ac7ba66),
	.w8(32'h3aeb5e33),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eee40),
	.w1(32'h38b35218),
	.w2(32'hba771a43),
	.w3(32'h3a8823b4),
	.w4(32'hba2ffc6a),
	.w5(32'hba6c7169),
	.w6(32'hba80ccf2),
	.w7(32'hba87e728),
	.w8(32'hba79295a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0040e2),
	.w1(32'h3888c5f4),
	.w2(32'h37c0cbcc),
	.w3(32'hba1335c9),
	.w4(32'h3abe522e),
	.w5(32'h3a8e7fb8),
	.w6(32'h39f7251c),
	.w7(32'h39507de3),
	.w8(32'h3a18a3cb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f38db),
	.w1(32'h3968d765),
	.w2(32'h3a861b7e),
	.w3(32'h3aa28a14),
	.w4(32'hb822962e),
	.w5(32'h3a1e006a),
	.w6(32'hb7276d03),
	.w7(32'h39c17867),
	.w8(32'h3a44ef7d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54edd8),
	.w1(32'hb8a0e50a),
	.w2(32'hb92c660b),
	.w3(32'h39ff9efb),
	.w4(32'hb8907190),
	.w5(32'hb904408a),
	.w6(32'hb915466e),
	.w7(32'hb8a74c7e),
	.w8(32'hb772c431),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78f2500),
	.w1(32'hb9d9f09a),
	.w2(32'hb977cb47),
	.w3(32'hb9e995c2),
	.w4(32'hba557768),
	.w5(32'hb924ce10),
	.w6(32'hba46f8b5),
	.w7(32'hba24dc9d),
	.w8(32'h3a3051e2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba910b71),
	.w1(32'h3a1be174),
	.w2(32'h3ae6b6f8),
	.w3(32'hba9d0096),
	.w4(32'h3a041187),
	.w5(32'h3adb6a44),
	.w6(32'h3880cd70),
	.w7(32'h3b017c54),
	.w8(32'h3b2a38b9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3790c551),
	.w1(32'h398565c5),
	.w2(32'hba480ec9),
	.w3(32'hb9cc822c),
	.w4(32'h3aa9bf6f),
	.w5(32'hb9c42caa),
	.w6(32'hb9e95000),
	.w7(32'h3b09a8f8),
	.w8(32'h3aa9096f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909c9ab),
	.w1(32'hba76f3ac),
	.w2(32'hba16ade7),
	.w3(32'h3994bc72),
	.w4(32'hb99e940d),
	.w5(32'h36e649c5),
	.w6(32'hb998bbcc),
	.w7(32'hb9a3ed6c),
	.w8(32'h3a3bd396),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3f6ea),
	.w1(32'hb899d231),
	.w2(32'hba273d9e),
	.w3(32'h3a9b5e90),
	.w4(32'h3a1a0d30),
	.w5(32'hb9941505),
	.w6(32'h39834aef),
	.w7(32'h3891ae36),
	.w8(32'h39c34fa2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994641c),
	.w1(32'hb978e3b0),
	.w2(32'hba8966d4),
	.w3(32'hb9ea0d94),
	.w4(32'h38b12f41),
	.w5(32'h3988f0a3),
	.w6(32'hb9935cc7),
	.w7(32'hb9a657a5),
	.w8(32'hba322971),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4eb30),
	.w1(32'h3b11ccdd),
	.w2(32'h3aa69bfc),
	.w3(32'h3a4a4af2),
	.w4(32'h3acb211d),
	.w5(32'h3a5d9d9b),
	.w6(32'h3aabd0f0),
	.w7(32'h3ac778f0),
	.w8(32'h3a8b99d1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee2a91),
	.w1(32'hba0174a7),
	.w2(32'hba630cbe),
	.w3(32'h3936c2de),
	.w4(32'hbad089c0),
	.w5(32'hbab3b2e0),
	.w6(32'hb9be622f),
	.w7(32'hba8597dd),
	.w8(32'hb9d804f7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c8d75),
	.w1(32'hb9ee75f7),
	.w2(32'h39a3d3ce),
	.w3(32'h3aa49376),
	.w4(32'h3ac049fe),
	.w5(32'h3a238828),
	.w6(32'h3b18993c),
	.w7(32'h3b5d21eb),
	.w8(32'h3b5f525d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b4dc0),
	.w1(32'h39b151c8),
	.w2(32'hb9e67e7c),
	.w3(32'hb9892b38),
	.w4(32'hbab2dde0),
	.w5(32'hb9266cb0),
	.w6(32'hba404ca8),
	.w7(32'hba93e52a),
	.w8(32'hb9aeb8d8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6870ec),
	.w1(32'h3ab10346),
	.w2(32'h3a969ade),
	.w3(32'hb98465ce),
	.w4(32'hb9e21668),
	.w5(32'h3a2d78a7),
	.w6(32'h3a5b1c61),
	.w7(32'h39a49042),
	.w8(32'h3aec6322),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39698023),
	.w1(32'hba866037),
	.w2(32'h3ac0460f),
	.w3(32'h3a5b747c),
	.w4(32'h3ac6a182),
	.w5(32'h3ab49122),
	.w6(32'h3a9355f5),
	.w7(32'h3b11a773),
	.w8(32'h3b33cf7e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a922cbb),
	.w1(32'h3929c8a0),
	.w2(32'hba1d6b91),
	.w3(32'h3b01da0b),
	.w4(32'hb9e21903),
	.w5(32'h39cad530),
	.w6(32'hb9d8687c),
	.w7(32'hba2dc183),
	.w8(32'h3a01f2ec),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961c4eb),
	.w1(32'h3a3833c5),
	.w2(32'h39c694cc),
	.w3(32'h3975f0b9),
	.w4(32'hba29eee6),
	.w5(32'h3a211d0f),
	.w6(32'h3afcd7ef),
	.w7(32'h3ab8f55e),
	.w8(32'h3afb2731),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74baf3),
	.w1(32'h3891344b),
	.w2(32'h3a1c3afe),
	.w3(32'h3a80c01a),
	.w4(32'h39709d64),
	.w5(32'h39dddb63),
	.w6(32'hb908e3a6),
	.w7(32'hb998318b),
	.w8(32'h39af8cf5),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3278ff),
	.w1(32'h3a64b241),
	.w2(32'hb9643fb3),
	.w3(32'h37b50d8a),
	.w4(32'hbaa2b7de),
	.w5(32'hbaa875f8),
	.w6(32'hbae8d57f),
	.w7(32'hbacd2717),
	.w8(32'hb9cc3cb4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba117b2a),
	.w1(32'hb8e7651f),
	.w2(32'hb9ba18f0),
	.w3(32'hb99d09ad),
	.w4(32'h390130e3),
	.w5(32'hba8d3f80),
	.w6(32'h3a5f1089),
	.w7(32'h3a75bd01),
	.w8(32'h3a8aefa0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c6fa7),
	.w1(32'h39b5c4ac),
	.w2(32'hb993c906),
	.w3(32'h39e507b3),
	.w4(32'h394b5086),
	.w5(32'h39811ec8),
	.w6(32'h39ce83db),
	.w7(32'h397a2803),
	.w8(32'h3a3cdea6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c069f),
	.w1(32'h39f5ea26),
	.w2(32'h3af7e503),
	.w3(32'h3a75f325),
	.w4(32'hb936d506),
	.w5(32'h39d40bd4),
	.w6(32'hb8f221e4),
	.w7(32'h3a50cb39),
	.w8(32'hb9d1157f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd15cd),
	.w1(32'hba30ffa1),
	.w2(32'hba90df25),
	.w3(32'hbab5a19f),
	.w4(32'h3951312b),
	.w5(32'h39986428),
	.w6(32'hba73a0e2),
	.w7(32'hba29aadb),
	.w8(32'h39d4e232),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1ffa7),
	.w1(32'hba51221d),
	.w2(32'h397a2ca8),
	.w3(32'h382ba2be),
	.w4(32'hbaeb9b59),
	.w5(32'hba06b8af),
	.w6(32'hba02bde7),
	.w7(32'hba923972),
	.w8(32'h3a2ff6a7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f374b),
	.w1(32'h3ac76115),
	.w2(32'h39cc35c4),
	.w3(32'hb8a7c1a5),
	.w4(32'h3a31defb),
	.w5(32'h3934874c),
	.w6(32'hb9b01475),
	.w7(32'h39330c70),
	.w8(32'h3a89f5d4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a420802),
	.w1(32'hb92383c0),
	.w2(32'hbaabc3e7),
	.w3(32'h3a6f42f6),
	.w4(32'hb9bc8cd9),
	.w5(32'hba0fb669),
	.w6(32'hba003a7e),
	.w7(32'hba553947),
	.w8(32'h38ab2c0d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f77c29),
	.w1(32'hb9dcb950),
	.w2(32'hbb4b0b1e),
	.w3(32'hba0be9db),
	.w4(32'h3a0fc428),
	.w5(32'hb994cf93),
	.w6(32'hba1f190f),
	.w7(32'hb9fbb3d6),
	.w8(32'hb9d33957),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d986f),
	.w1(32'h3ad2d796),
	.w2(32'hb8200f3c),
	.w3(32'hbb14b9f5),
	.w4(32'h3a9b5d53),
	.w5(32'h3a753406),
	.w6(32'hbaa4d593),
	.w7(32'h37f118f4),
	.w8(32'h3aff9981),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd90b8),
	.w1(32'hba817f3f),
	.w2(32'h3b1f3628),
	.w3(32'hb9f34632),
	.w4(32'hb9e6d9f7),
	.w5(32'h3ab0cb04),
	.w6(32'h3ae232ac),
	.w7(32'h3aab1afc),
	.w8(32'h3b4f4136),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b070e5f),
	.w1(32'h3a7a953a),
	.w2(32'hb9980aad),
	.w3(32'hb8588043),
	.w4(32'hbab64596),
	.w5(32'hb9eab5a2),
	.w6(32'hba1a3856),
	.w7(32'hba55b3b1),
	.w8(32'h3923a6e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb8d7b),
	.w1(32'hb9d03bac),
	.w2(32'hba314cc0),
	.w3(32'h3a903ae9),
	.w4(32'hbae3651b),
	.w5(32'h381128a9),
	.w6(32'hb9fbe54b),
	.w7(32'h3a7a600c),
	.w8(32'h3a5138ba),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b079),
	.w1(32'h3b7f362b),
	.w2(32'h3adcd62c),
	.w3(32'h3a4204ab),
	.w4(32'h3af0962e),
	.w5(32'h39a3cf2b),
	.w6(32'h3b0fd004),
	.w7(32'h3b218919),
	.w8(32'h3b801c2b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0167a5),
	.w1(32'h3a9c7086),
	.w2(32'h38e1b0ae),
	.w3(32'h3a480218),
	.w4(32'hb984845a),
	.w5(32'h3b0925f4),
	.w6(32'h3983e599),
	.w7(32'hbaa3897b),
	.w8(32'h3b0eb7a6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a381bac),
	.w1(32'hba806d15),
	.w2(32'hbab3a628),
	.w3(32'h39622b40),
	.w4(32'hbb02cea7),
	.w5(32'hbaed3a14),
	.w6(32'hba6e8915),
	.w7(32'hbaa844b4),
	.w8(32'hba9045f4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cbf02),
	.w1(32'hb95907b8),
	.w2(32'h3979cfec),
	.w3(32'hb8bd944f),
	.w4(32'hba8c2369),
	.w5(32'hb8818a17),
	.w6(32'hb8a1b915),
	.w7(32'hb852db19),
	.w8(32'hbaae74e0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44ce6e),
	.w1(32'h3819cb8f),
	.w2(32'h3a258353),
	.w3(32'hba044e23),
	.w4(32'h39be7381),
	.w5(32'h3a21bec7),
	.w6(32'h39676366),
	.w7(32'h399b73dd),
	.w8(32'h3a6305b7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce1d7b),
	.w1(32'h376d4eee),
	.w2(32'hb8cd99f2),
	.w3(32'h39a6c7bc),
	.w4(32'hb86b9f4b),
	.w5(32'h37bb86a2),
	.w6(32'hb8ffadae),
	.w7(32'hb95f0af0),
	.w8(32'h39a21dce),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c7566c),
	.w1(32'hba7a9028),
	.w2(32'h39f34d59),
	.w3(32'hb7c59add),
	.w4(32'hbad67f07),
	.w5(32'h39923f6e),
	.w6(32'hba3486eb),
	.w7(32'h3926be71),
	.w8(32'h3b18aee5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3982d98d),
	.w1(32'h3b29fc51),
	.w2(32'h3abf9dc8),
	.w3(32'h39269e49),
	.w4(32'h3ae18adf),
	.w5(32'h399750bb),
	.w6(32'h3af895da),
	.w7(32'h3986b52f),
	.w8(32'h39fa0dab),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fe4af),
	.w1(32'h39e914f4),
	.w2(32'hba7cabdf),
	.w3(32'h3b05b01b),
	.w4(32'h39a25839),
	.w5(32'hb8dace41),
	.w6(32'h39f59dbc),
	.w7(32'hba88bedd),
	.w8(32'hb90801e7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d772aa),
	.w1(32'h3a2db80b),
	.w2(32'h392f49bb),
	.w3(32'h3a7d8ebd),
	.w4(32'hb8dba77e),
	.w5(32'h383339ff),
	.w6(32'h3a78bfed),
	.w7(32'hb93156b5),
	.w8(32'h3a43a2bb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8e16c),
	.w1(32'hba9ca71f),
	.w2(32'hb9f8eadc),
	.w3(32'hbaabf8fc),
	.w4(32'hb994549e),
	.w5(32'hb82ee90a),
	.w6(32'hbae03813),
	.w7(32'h3a40a4ad),
	.w8(32'h3af21635),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9ae71),
	.w1(32'h396b524f),
	.w2(32'hba27fa59),
	.w3(32'h3a2e9636),
	.w4(32'h3a036027),
	.w5(32'h388efbc6),
	.w6(32'h39d09039),
	.w7(32'hb79a4ae3),
	.w8(32'h3a08087b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3d9dc),
	.w1(32'hb8b3042c),
	.w2(32'hb868bb80),
	.w3(32'hb9826833),
	.w4(32'hb9d4c451),
	.w5(32'hb828dd51),
	.w6(32'hb9dcb779),
	.w7(32'hb70e0855),
	.w8(32'h399fd9a6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a4db),
	.w1(32'hb95812eb),
	.w2(32'hba165b76),
	.w3(32'h3b151c78),
	.w4(32'hbaca48cb),
	.w5(32'hb98b9a65),
	.w6(32'h3abc5b7a),
	.w7(32'hbb0aa5a8),
	.w8(32'h3a07f743),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b482e),
	.w1(32'hb9e8494f),
	.w2(32'h3acc4e02),
	.w3(32'h3a2a8313),
	.w4(32'h38f450a1),
	.w5(32'h3acc19e8),
	.w6(32'h3b989815),
	.w7(32'h3b083b7d),
	.w8(32'h3b85e426),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0bb82),
	.w1(32'hba7649a5),
	.w2(32'hbaa64d85),
	.w3(32'hb9b70fc4),
	.w4(32'hba396b1b),
	.w5(32'hba5511e7),
	.w6(32'hba909f0f),
	.w7(32'hba9e2e6c),
	.w8(32'hb9f85424),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978c4b7),
	.w1(32'h39cf3d28),
	.w2(32'hba5a56eb),
	.w3(32'hb9219ea1),
	.w4(32'hbad63560),
	.w5(32'hbb18cbdd),
	.w6(32'hbaec551b),
	.w7(32'hbaee2fbc),
	.w8(32'hbb0164f7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883a7c2),
	.w1(32'hba261ec7),
	.w2(32'hba186f0b),
	.w3(32'hb7fb6516),
	.w4(32'h3a0a1965),
	.w5(32'h3a20ebee),
	.w6(32'hb8442a81),
	.w7(32'h39c49b8e),
	.w8(32'h39d74055),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1242f),
	.w1(32'hbae13b0a),
	.w2(32'hbac89281),
	.w3(32'h3ab75895),
	.w4(32'hb9f93895),
	.w5(32'hba890ac5),
	.w6(32'hbb01a0da),
	.w7(32'hbaa72d6b),
	.w8(32'hba801149),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8628fc),
	.w1(32'h3b24ce66),
	.w2(32'h3a667709),
	.w3(32'h3984ac62),
	.w4(32'h3b10e325),
	.w5(32'h3a4e681a),
	.w6(32'h3b007f3f),
	.w7(32'h3b07007a),
	.w8(32'h3ab759d8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93684b4),
	.w1(32'h3a27dc65),
	.w2(32'h3a51689e),
	.w3(32'h3982518e),
	.w4(32'hb91e6ea1),
	.w5(32'h3b17d944),
	.w6(32'h3b71def1),
	.w7(32'h3b4ee286),
	.w8(32'h3ba6214b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c2b15),
	.w1(32'h3a5d5603),
	.w2(32'h39b27534),
	.w3(32'h3ae5dbb0),
	.w4(32'h39a6b5c6),
	.w5(32'h3720c87d),
	.w6(32'h3a818182),
	.w7(32'h38bd1bcf),
	.w8(32'hbaea55fc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad68cd4),
	.w1(32'h3935339c),
	.w2(32'h393ffeb8),
	.w3(32'hb8b70e89),
	.w4(32'hb9b2b579),
	.w5(32'hb9d57f1e),
	.w6(32'h3b0c6235),
	.w7(32'hb807e4d0),
	.w8(32'h39f0fd5e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ce3da),
	.w1(32'hba214a15),
	.w2(32'hba59d485),
	.w3(32'h3a1cac20),
	.w4(32'hba2ec5b8),
	.w5(32'hba139919),
	.w6(32'hb9f40a61),
	.w7(32'hb9cd10a9),
	.w8(32'hb8d3de81),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a799a),
	.w1(32'hb9f42242),
	.w2(32'hbab0ccc1),
	.w3(32'h3950d456),
	.w4(32'hb9d19550),
	.w5(32'hba93330d),
	.w6(32'hb85eab20),
	.w7(32'hba064b8f),
	.w8(32'hb9ccfd98),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9709a44),
	.w1(32'h3a851794),
	.w2(32'h39977fc9),
	.w3(32'hba000a59),
	.w4(32'h3a6a75c6),
	.w5(32'h3ac1f86f),
	.w6(32'h3b012d5b),
	.w7(32'h38f8d2a6),
	.w8(32'h39872842),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4bcdf),
	.w1(32'h3ac61fb7),
	.w2(32'h39f1bce2),
	.w3(32'h3b089367),
	.w4(32'h39cc8a8d),
	.w5(32'h3a2f134e),
	.w6(32'h3a92dafd),
	.w7(32'h3aaf1739),
	.w8(32'h3ad60abb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a763795),
	.w1(32'hb9e7b2a1),
	.w2(32'h3a720fce),
	.w3(32'h3ac9edcb),
	.w4(32'h38af5e33),
	.w5(32'h3a07a0df),
	.w6(32'h39127ab6),
	.w7(32'h39afbc53),
	.w8(32'h38aff9c3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e5bde),
	.w1(32'h3900eb7d),
	.w2(32'h3a1b0fba),
	.w3(32'h391465ae),
	.w4(32'h38ce8657),
	.w5(32'h39d86677),
	.w6(32'hb91a20a2),
	.w7(32'h3968873f),
	.w8(32'h3a3a346e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a559271),
	.w1(32'h3a7674fe),
	.w2(32'h38148266),
	.w3(32'h3a6b6831),
	.w4(32'h3a7103d9),
	.w5(32'h3975c2af),
	.w6(32'h3accb588),
	.w7(32'h3a8cd38f),
	.w8(32'h3a8126ca),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951e0fa),
	.w1(32'hb910d4ba),
	.w2(32'h3a031ac3),
	.w3(32'hba619b35),
	.w4(32'hba45bf63),
	.w5(32'h3a4f7ab3),
	.w6(32'hbab1dd9f),
	.w7(32'h39e4d425),
	.w8(32'h3b132206),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c34f4f),
	.w1(32'h3a04ca98),
	.w2(32'h3a9a44aa),
	.w3(32'hb74bbc28),
	.w4(32'hba9d6a9f),
	.w5(32'hba817bfe),
	.w6(32'h3ab0782b),
	.w7(32'hba3c7ead),
	.w8(32'h3ad63880),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f823),
	.w1(32'h39a22bc7),
	.w2(32'hb8f93c2c),
	.w3(32'h393a5473),
	.w4(32'h3a19f4c2),
	.w5(32'h3a5cb9e4),
	.w6(32'h3908760f),
	.w7(32'h393e2983),
	.w8(32'h3a776209),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710eef1),
	.w1(32'h3b1fecee),
	.w2(32'h3b50c308),
	.w3(32'hba24b239),
	.w4(32'h3b190b05),
	.w5(32'h3bd8f432),
	.w6(32'hba9079c7),
	.w7(32'h3b75f2b3),
	.w8(32'h3be3bb86),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6166f0),
	.w1(32'h39eb1f07),
	.w2(32'hba52f409),
	.w3(32'h392bd835),
	.w4(32'hbb45ebd6),
	.w5(32'hb966763f),
	.w6(32'hba8d3351),
	.w7(32'hbb6a3561),
	.w8(32'hb92b7c2f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f9c86),
	.w1(32'hba532775),
	.w2(32'hb95adaf0),
	.w3(32'hb8926d9b),
	.w4(32'hba4b1f91),
	.w5(32'h3975d905),
	.w6(32'hba0348e5),
	.w7(32'hb9d7e1cd),
	.w8(32'h3a28ef34),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924b731),
	.w1(32'h38ee4fd4),
	.w2(32'h3aee6411),
	.w3(32'h38016f53),
	.w4(32'h395322ca),
	.w5(32'h3aa73c49),
	.w6(32'hbaa11bf4),
	.w7(32'hb8f13fb0),
	.w8(32'h3b3f470f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10beb0),
	.w1(32'h3985259c),
	.w2(32'h398259f0),
	.w3(32'h3b0b74d4),
	.w4(32'h39529af8),
	.w5(32'h3a0b24dc),
	.w6(32'hba0bb735),
	.w7(32'hba1813eb),
	.w8(32'h3a2e35e9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81906a3),
	.w1(32'hbacec042),
	.w2(32'hba94f0e4),
	.w3(32'h39c8ec98),
	.w4(32'hba797db2),
	.w5(32'hba8787eb),
	.w6(32'hbab98c6c),
	.w7(32'hba9d9a6a),
	.w8(32'hb6d7b778),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00b8b),
	.w1(32'hba243d6b),
	.w2(32'h390d5816),
	.w3(32'hbb12356d),
	.w4(32'hb9ae76c6),
	.w5(32'h3a140458),
	.w6(32'hb82915be),
	.w7(32'hba3aba1e),
	.w8(32'h3a90a456),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a9bfad),
	.w1(32'h3b05ba0b),
	.w2(32'h3a9efd3d),
	.w3(32'hba392207),
	.w4(32'h3a960d7b),
	.w5(32'h383162d7),
	.w6(32'h3ad36cc9),
	.w7(32'h3b2220f5),
	.w8(32'h3a9c5680),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e23f5),
	.w1(32'h3a9a5e63),
	.w2(32'hba097e2e),
	.w3(32'h3a0c2e6b),
	.w4(32'h39bfdf8e),
	.w5(32'hb943f2e4),
	.w6(32'hb9fbbdad),
	.w7(32'hbae8c14c),
	.w8(32'hba7611e8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990114f),
	.w1(32'h38a42fd1),
	.w2(32'hba9c47d7),
	.w3(32'h3ac09fae),
	.w4(32'hb9e4c53c),
	.w5(32'hb9ffebac),
	.w6(32'h3a220edc),
	.w7(32'h37a2ac2e),
	.w8(32'h39940b87),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dd9ea),
	.w1(32'hb9eb51fc),
	.w2(32'hba1b0644),
	.w3(32'h39f662dd),
	.w4(32'hba332717),
	.w5(32'hba06186d),
	.w6(32'h36b48346),
	.w7(32'hba48c0cb),
	.w8(32'h39862e1e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30c952),
	.w1(32'hb9c9b4e5),
	.w2(32'hba339a7b),
	.w3(32'hbaafaac8),
	.w4(32'hba12c531),
	.w5(32'hb98c699c),
	.w6(32'hba173998),
	.w7(32'hba9b1d95),
	.w8(32'hb964242a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926b17f),
	.w1(32'hb84048a6),
	.w2(32'hb892dcb4),
	.w3(32'h38fc5e73),
	.w4(32'hb930960d),
	.w5(32'h39c1618c),
	.w6(32'hb85a0c0a),
	.w7(32'hb8903606),
	.w8(32'h39ba1705),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a854b5d),
	.w1(32'h39e8ab2f),
	.w2(32'hb9d1e030),
	.w3(32'h3b018226),
	.w4(32'h3a788054),
	.w5(32'hb78ce332),
	.w6(32'h39fc075f),
	.w7(32'h389e47fb),
	.w8(32'h39b5ce97),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389614b7),
	.w1(32'h39611f58),
	.w2(32'hb994a7d8),
	.w3(32'h39cc46e9),
	.w4(32'h38ec2287),
	.w5(32'hb8a6208b),
	.w6(32'h38f389dd),
	.w7(32'hb94f40e7),
	.w8(32'h39c40f76),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a523479),
	.w1(32'hb916f8c6),
	.w2(32'h389db941),
	.w3(32'h3ab684fe),
	.w4(32'h39e7c4fd),
	.w5(32'h3a254918),
	.w6(32'h398b23d5),
	.w7(32'h398c8c47),
	.w8(32'h3a6b4079),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a464882),
	.w1(32'hba2e6030),
	.w2(32'h3a0e21bc),
	.w3(32'hb98341c4),
	.w4(32'hbb428c8f),
	.w5(32'hb98ae137),
	.w6(32'h3a79e1b7),
	.w7(32'h3a14f620),
	.w8(32'h3a587c27),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affde34),
	.w1(32'h39d359a5),
	.w2(32'h3985f70a),
	.w3(32'h3aad1264),
	.w4(32'hbac24e9e),
	.w5(32'hb9cdf1ba),
	.w6(32'hb9b8d7dc),
	.w7(32'hba7b0b7b),
	.w8(32'h39b21e5f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a49ea),
	.w1(32'hb9dc251a),
	.w2(32'h3a9b2a04),
	.w3(32'h3a0474ed),
	.w4(32'h38bfd0ef),
	.w5(32'h3ab17a26),
	.w6(32'h393442c0),
	.w7(32'h3a810ad7),
	.w8(32'h3ad18df1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acadd5f),
	.w1(32'h374e6f69),
	.w2(32'h3aa4a9e8),
	.w3(32'h3a2f6abd),
	.w4(32'hbb197232),
	.w5(32'hba9ac72f),
	.w6(32'hba8ef730),
	.w7(32'hbad004aa),
	.w8(32'hba9b2856),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2ea5a),
	.w1(32'h3acd9c83),
	.w2(32'h39b7b4f0),
	.w3(32'h3a89ec8a),
	.w4(32'h3a32483b),
	.w5(32'h3a4fc2ac),
	.w6(32'h3a4d14e8),
	.w7(32'hb8bcee45),
	.w8(32'h3a97dfb4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af20459),
	.w1(32'h3b13f85f),
	.w2(32'h39b505db),
	.w3(32'h3af56bfd),
	.w4(32'h3af13de9),
	.w5(32'hb81891b7),
	.w6(32'h3b0b4f3d),
	.w7(32'h3a35c8e9),
	.w8(32'h3a820f1d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99aed2f),
	.w1(32'hba22c8e3),
	.w2(32'hbab0aa0f),
	.w3(32'h393b860b),
	.w4(32'hb9c8da2c),
	.w5(32'hb9bd55ce),
	.w6(32'hba466731),
	.w7(32'hba83e47d),
	.w8(32'hb9435c3d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9ff8d),
	.w1(32'h3845ae86),
	.w2(32'h38859e57),
	.w3(32'hb911e317),
	.w4(32'h394bccf7),
	.w5(32'h392ad658),
	.w6(32'h399fa856),
	.w7(32'h39b9a67e),
	.w8(32'h39914024),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d47f1),
	.w1(32'hb9c43d69),
	.w2(32'hb9613a94),
	.w3(32'hba49573c),
	.w4(32'h38e32b20),
	.w5(32'h3b125aae),
	.w6(32'hbabbbfde),
	.w7(32'h39a8553d),
	.w8(32'h3b138b85),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996d583),
	.w1(32'h3b5e52df),
	.w2(32'h3b45aaa4),
	.w3(32'h3a839f56),
	.w4(32'h3aebdd9d),
	.w5(32'h3aedeb75),
	.w6(32'h3b810515),
	.w7(32'h3b802b02),
	.w8(32'h3b806002),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc8705),
	.w1(32'h3ae4880e),
	.w2(32'h3913b66b),
	.w3(32'h3aa00570),
	.w4(32'hb9c899bd),
	.w5(32'h3988e805),
	.w6(32'hb9e55ed2),
	.w7(32'h390ace46),
	.w8(32'h390f86b1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e543cb),
	.w1(32'hbae35256),
	.w2(32'h3b0a7835),
	.w3(32'hbb23f79d),
	.w4(32'hbb152c2a),
	.w5(32'h3a8b2935),
	.w6(32'hba891054),
	.w7(32'h3ab026c4),
	.w8(32'h3a2ff56f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789106a),
	.w1(32'h3964195a),
	.w2(32'hba239cba),
	.w3(32'hb7966a92),
	.w4(32'hb7d2ab49),
	.w5(32'hb995fafc),
	.w6(32'hb801ff59),
	.w7(32'hb98f70d1),
	.w8(32'h3931c49e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d759d2),
	.w1(32'h3a29135f),
	.w2(32'h38c8a223),
	.w3(32'h3a267b47),
	.w4(32'h3a44d9b3),
	.w5(32'h39fae7b8),
	.w6(32'h39c5fd33),
	.w7(32'h3a77af4d),
	.w8(32'h3a4c0017),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba2f7c),
	.w1(32'hbb4ecc0a),
	.w2(32'h3b0d62f1),
	.w3(32'hbb14f882),
	.w4(32'hbb2e495e),
	.w5(32'h3b085294),
	.w6(32'hbaee95bc),
	.w7(32'hbb2253b2),
	.w8(32'h3b553bac),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38849a15),
	.w1(32'h3aa8084a),
	.w2(32'h3aeea70e),
	.w3(32'h3ab793a5),
	.w4(32'h3b3fd798),
	.w5(32'h3ac666bc),
	.w6(32'h3b309440),
	.w7(32'h3b7349e1),
	.w8(32'h3b343548),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95bee5),
	.w1(32'hbb2574eb),
	.w2(32'h39b5cbd2),
	.w3(32'hba90d284),
	.w4(32'hb9ae25bc),
	.w5(32'h3aa623f8),
	.w6(32'h3aa08b52),
	.w7(32'h3a75a9aa),
	.w8(32'h3b590228),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926d1c),
	.w1(32'hb989ac6b),
	.w2(32'hb9aac080),
	.w3(32'h3a03c13a),
	.w4(32'hba787da2),
	.w5(32'hb9ebb8ec),
	.w6(32'hb9bd34ee),
	.w7(32'hba9eb348),
	.w8(32'h398058d8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b236ee8),
	.w1(32'h3ac4985b),
	.w2(32'hb98c0754),
	.w3(32'h3ace5013),
	.w4(32'h3978ce48),
	.w5(32'hb9682863),
	.w6(32'h3adf06d1),
	.w7(32'hb9051e85),
	.w8(32'h3aa36731),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956e480),
	.w1(32'hb99ec791),
	.w2(32'hba500350),
	.w3(32'h3961234e),
	.w4(32'h381f4f02),
	.w5(32'hb95a27a7),
	.w6(32'hb97a94b3),
	.w7(32'hb9b5ef6a),
	.w8(32'hb8a8e019),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9874e85),
	.w1(32'hba6c14c0),
	.w2(32'hb93bc725),
	.w3(32'hb7501aeb),
	.w4(32'hb9e0c0a2),
	.w5(32'hb92298ac),
	.w6(32'hb99c9c4c),
	.w7(32'hb9d34145),
	.w8(32'hb9993f7d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3d578),
	.w1(32'h396468cb),
	.w2(32'hb9efa1d4),
	.w3(32'hba36cdcd),
	.w4(32'h39851811),
	.w5(32'hba74e07e),
	.w6(32'h395c61db),
	.w7(32'hba4d3134),
	.w8(32'h3a7a5923),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d4f68),
	.w1(32'h3896e9a0),
	.w2(32'hb8ea0973),
	.w3(32'hb9e8263d),
	.w4(32'h395df3d0),
	.w5(32'h38fa05c7),
	.w6(32'h396822d8),
	.w7(32'hb8874163),
	.w8(32'h39a52f03),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9292678),
	.w1(32'hba58a72e),
	.w2(32'hba256dd5),
	.w3(32'hb9c06589),
	.w4(32'hb86794f2),
	.w5(32'h3a0a5f04),
	.w6(32'hba47298a),
	.w7(32'hb98fa150),
	.w8(32'h3a7658c2),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9392395),
	.w1(32'h3aa06cff),
	.w2(32'h3a972ad4),
	.w3(32'h392b6d68),
	.w4(32'h3a9e7c05),
	.w5(32'h3aaf14da),
	.w6(32'h3aa5288f),
	.w7(32'h3abca526),
	.w8(32'h3b3b5b14),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9faf6e),
	.w1(32'h3ab73278),
	.w2(32'hba393ab0),
	.w3(32'h3a232dcd),
	.w4(32'hba357345),
	.w5(32'hbb2fd422),
	.w6(32'h3a228197),
	.w7(32'hba7af431),
	.w8(32'h37d8294f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9183e06),
	.w1(32'h3abd5545),
	.w2(32'h3a6a1886),
	.w3(32'hbac7aeb0),
	.w4(32'h3a5364ab),
	.w5(32'h39e411db),
	.w6(32'h3aa2621b),
	.w7(32'h39403ca8),
	.w8(32'hb8891fa8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265cc5),
	.w1(32'hbabbf420),
	.w2(32'h3b59af2f),
	.w3(32'h39ff50cd),
	.w4(32'h3a8788be),
	.w5(32'h3af61088),
	.w6(32'h3b343221),
	.w7(32'h3b34e407),
	.w8(32'h3ba91bb7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd831),
	.w1(32'hb9f43c9c),
	.w2(32'h3986bb92),
	.w3(32'h39d52b8e),
	.w4(32'hb9aaa8a7),
	.w5(32'h3a153b5f),
	.w6(32'h3a036000),
	.w7(32'h3aa0e8ae),
	.w8(32'h3acfd362),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0dd93),
	.w1(32'h370967f3),
	.w2(32'hb8862c35),
	.w3(32'h3a4ee2d7),
	.w4(32'hb9588c57),
	.w5(32'hb755bd38),
	.w6(32'h38d958ea),
	.w7(32'h36c143b5),
	.w8(32'h39c038b6),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eb63e9),
	.w1(32'h3a77feec),
	.w2(32'h3aca224b),
	.w3(32'h3a5631ff),
	.w4(32'h3a452f2f),
	.w5(32'h3a8fad62),
	.w6(32'h3acf42b3),
	.w7(32'h3ad10ef0),
	.w8(32'h3b2b386c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bc54a0),
	.w1(32'hbab871a1),
	.w2(32'hbaafb5da),
	.w3(32'h37eae6be),
	.w4(32'hba664b0e),
	.w5(32'hb987b955),
	.w6(32'hbaa17e6b),
	.w7(32'hba93d0e3),
	.w8(32'hb9700045),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d9917),
	.w1(32'h37183b2e),
	.w2(32'hba26aa0e),
	.w3(32'h3903b67f),
	.w4(32'hb9588341),
	.w5(32'hb7b8a75f),
	.w6(32'hb8ac54c0),
	.w7(32'hba2c7228),
	.w8(32'h3a27112f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9622110),
	.w1(32'hb87251dd),
	.w2(32'hb95c1845),
	.w3(32'h39b681d5),
	.w4(32'hb9b4fc2a),
	.w5(32'hb92a6baf),
	.w6(32'h391010c7),
	.w7(32'hb8f0cdc0),
	.w8(32'h398421ea),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0b216),
	.w1(32'hbb00b3cf),
	.w2(32'h3801ba7a),
	.w3(32'h39a650fa),
	.w4(32'hba61e7e7),
	.w5(32'h398e3013),
	.w6(32'hbaf10b69),
	.w7(32'hba004e9a),
	.w8(32'h37c1dee4),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a3df8),
	.w1(32'h39df5b35),
	.w2(32'hba1dfd86),
	.w3(32'h39ea4459),
	.w4(32'hb9d7efe9),
	.w5(32'hb9836ade),
	.w6(32'h3a6f52ab),
	.w7(32'hb9e901d4),
	.w8(32'h37128bc3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcde41),
	.w1(32'h39d13787),
	.w2(32'h3b307873),
	.w3(32'h3a15cdbb),
	.w4(32'hb9ae7845),
	.w5(32'h3aaeb07d),
	.w6(32'h391400c7),
	.w7(32'h3abd936d),
	.w8(32'h3a1bfe57),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f17aa8),
	.w1(32'h3a67be80),
	.w2(32'h3a6855fb),
	.w3(32'h3a7863d0),
	.w4(32'h3a1352db),
	.w5(32'h3abe1b8a),
	.w6(32'h3ad0bfe6),
	.w7(32'h3aeacd0a),
	.w8(32'h3b2b94cc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab52f96),
	.w1(32'h39a30c16),
	.w2(32'h38117024),
	.w3(32'h3adb4a36),
	.w4(32'hb9454c93),
	.w5(32'hba19863c),
	.w6(32'h3abd73a4),
	.w7(32'h3a7f6d8d),
	.w8(32'h390a86af),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e082ff),
	.w1(32'hbae30252),
	.w2(32'hbabaa04b),
	.w3(32'hb98e1e67),
	.w4(32'hbac41fb8),
	.w5(32'hbab1b3fc),
	.w6(32'hba8998ea),
	.w7(32'hba986f4d),
	.w8(32'hba768d63),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba700fd0),
	.w1(32'h388ac88a),
	.w2(32'hb945ec12),
	.w3(32'hba6893e1),
	.w4(32'hb9a6d3c8),
	.w5(32'hb91f138d),
	.w6(32'h38724a83),
	.w7(32'hb6251d53),
	.w8(32'h3a0912b3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a091698),
	.w1(32'hb7dbf92f),
	.w2(32'hb7e02ef4),
	.w3(32'h3a3be33f),
	.w4(32'hb8be01e4),
	.w5(32'hb91997ed),
	.w6(32'hb935c2fc),
	.w7(32'h3964b7a3),
	.w8(32'h39b060e3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996d22c),
	.w1(32'hb888a975),
	.w2(32'h38ae63bd),
	.w3(32'h39935204),
	.w4(32'hb9c98257),
	.w5(32'h386286b5),
	.w6(32'hb944b428),
	.w7(32'hb8aaa50a),
	.w8(32'h39c9d90a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fa272),
	.w1(32'h3829db99),
	.w2(32'h38d848f5),
	.w3(32'h3591999b),
	.w4(32'h3ad7877d),
	.w5(32'h3ac15ea7),
	.w6(32'hba4e27a1),
	.w7(32'h39e320f1),
	.w8(32'h3a1c0b73),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f39ed),
	.w1(32'h399dbdce),
	.w2(32'hb9be4b51),
	.w3(32'h39f4c1f5),
	.w4(32'h39da3e45),
	.w5(32'hb8290f56),
	.w6(32'h3a0b980f),
	.w7(32'hb8c55408),
	.w8(32'h3a2a2ebe),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f22a17),
	.w1(32'hb9b3682d),
	.w2(32'hb98e2289),
	.w3(32'hba9188f2),
	.w4(32'hba52b7b2),
	.w5(32'hb94c08ed),
	.w6(32'hba39eabd),
	.w7(32'hba18699e),
	.w8(32'h39671de8),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1afefc),
	.w1(32'h3a221753),
	.w2(32'hb9844887),
	.w3(32'h3a9ee664),
	.w4(32'h3990de68),
	.w5(32'hb8a9e0b2),
	.w6(32'h37c34428),
	.w7(32'hb9942564),
	.w8(32'hba0c67a3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b9ccc),
	.w1(32'hb995c1d0),
	.w2(32'hb931721b),
	.w3(32'hb5d8c872),
	.w4(32'hba325148),
	.w5(32'hb8053550),
	.w6(32'hba42e6dc),
	.w7(32'hb9d69954),
	.w8(32'h39f3bd4b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8e1f5),
	.w1(32'hb992aadb),
	.w2(32'hbb056a7d),
	.w3(32'hb9138942),
	.w4(32'h3a8a630e),
	.w5(32'h3a0b97d4),
	.w6(32'h39813bcf),
	.w7(32'h3a1a572d),
	.w8(32'h3a9c247f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995c9fe),
	.w1(32'hb9988a3f),
	.w2(32'h3a1aa7ed),
	.w3(32'h3a0c963a),
	.w4(32'hb9acf58f),
	.w5(32'h3a24d08b),
	.w6(32'hb9389254),
	.w7(32'h3a57696f),
	.w8(32'h3add90b1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b644),
	.w1(32'h3ac6d489),
	.w2(32'h393a73eb),
	.w3(32'h3b2566d8),
	.w4(32'hb8d752ea),
	.w5(32'hba161693),
	.w6(32'h3b5f40c0),
	.w7(32'h3ad5e80f),
	.w8(32'h38881ba2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37da1152),
	.w1(32'h38b0a6aa),
	.w2(32'hb8ef66fd),
	.w3(32'h3a025aa8),
	.w4(32'h393f6783),
	.w5(32'h383f359f),
	.w6(32'h38e36961),
	.w7(32'hb93dbff1),
	.w8(32'h389770f2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe26f6),
	.w1(32'h3ad97b05),
	.w2(32'h3aaa27e4),
	.w3(32'h3aefc066),
	.w4(32'h3aae63d2),
	.w5(32'h3ab330b2),
	.w6(32'h3b4618cd),
	.w7(32'h3aac4c68),
	.w8(32'h3af6da0e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule