module layer_10_featuremap_372(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a6278),
	.w1(32'h3bd23114),
	.w2(32'h3a297ec0),
	.w3(32'h3b200b23),
	.w4(32'h3af885c6),
	.w5(32'h3c81b3d4),
	.w6(32'hbc00b779),
	.w7(32'hbb6d4c77),
	.w8(32'hbc0495f8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07408a),
	.w1(32'h3c0157dc),
	.w2(32'h3c07f7af),
	.w3(32'hba72dce5),
	.w4(32'h3b10adc5),
	.w5(32'h3c173c88),
	.w6(32'hba910149),
	.w7(32'h3bd944ef),
	.w8(32'h3c017ead),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8229a),
	.w1(32'hbb236bcc),
	.w2(32'h3b44304a),
	.w3(32'hbc2b259d),
	.w4(32'h3bd19001),
	.w5(32'h3c5f65af),
	.w6(32'h3c8bdaa3),
	.w7(32'h3c15dfc5),
	.w8(32'h39e454b3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc252e11),
	.w1(32'hbd652cbb),
	.w2(32'hbb2073db),
	.w3(32'hbc1f7e64),
	.w4(32'h3c9fe11d),
	.w5(32'hbbfdab2c),
	.w6(32'hbb41f579),
	.w7(32'h36d0ebd9),
	.w8(32'h3c143335),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2140d),
	.w1(32'hbcbb90da),
	.w2(32'h3ab6c45b),
	.w3(32'hbd68d8c0),
	.w4(32'h3b1304a6),
	.w5(32'h3aa959a4),
	.w6(32'hbc4b070a),
	.w7(32'hbab2eff8),
	.w8(32'hbd94477d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02277d),
	.w1(32'hbba88f2c),
	.w2(32'h39e4ce50),
	.w3(32'hbb803703),
	.w4(32'h3b2d5bce),
	.w5(32'h3bf81800),
	.w6(32'hbb9fbe7d),
	.w7(32'h3b700030),
	.w8(32'h3b72d9c1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12f6b9),
	.w1(32'hbc6e97a6),
	.w2(32'hbc9eb631),
	.w3(32'h3b745fb1),
	.w4(32'h3bf8584a),
	.w5(32'hbd33e19a),
	.w6(32'hbb148905),
	.w7(32'hbc497c1e),
	.w8(32'hbc05ef59),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87e57c),
	.w1(32'h390ea192),
	.w2(32'h3b8f8436),
	.w3(32'hbbc6aff5),
	.w4(32'hbc754ebb),
	.w5(32'h3cbfa26a),
	.w6(32'hbb9b8d48),
	.w7(32'h3c4df59c),
	.w8(32'h3c7dd98e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17cdea),
	.w1(32'hbc05d29e),
	.w2(32'h3c8bc181),
	.w3(32'h3c8c9bbc),
	.w4(32'h3b0ad6a8),
	.w5(32'hba4abc52),
	.w6(32'hbbdb7b89),
	.w7(32'h3b2dd361),
	.w8(32'h3b80906e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26c2f9),
	.w1(32'hbb1deae2),
	.w2(32'h3b94c733),
	.w3(32'h3bbeaca1),
	.w4(32'h3bea65b7),
	.w5(32'h3c075e3a),
	.w6(32'hbc4f17b5),
	.w7(32'h3b52db73),
	.w8(32'hba427d49),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecf4c9),
	.w1(32'h3a5b0d02),
	.w2(32'hbb43f1f9),
	.w3(32'h3c497a75),
	.w4(32'h3c6a9565),
	.w5(32'hbcbeb64c),
	.w6(32'hb840e86e),
	.w7(32'hbb419316),
	.w8(32'h3ae7759c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892f0c),
	.w1(32'hba2bdf74),
	.w2(32'hbd9f2066),
	.w3(32'h3bdc6124),
	.w4(32'hbc903203),
	.w5(32'hbca684e9),
	.w6(32'h3bd15a7a),
	.w7(32'hbc318636),
	.w8(32'hbccd794b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc019f1c),
	.w1(32'h3b25ff56),
	.w2(32'hbc4f0cdf),
	.w3(32'h3c1f7745),
	.w4(32'hba9a59aa),
	.w5(32'hbc5afc5c),
	.w6(32'h3baa2c13),
	.w7(32'hbc4ea774),
	.w8(32'hbcb4d401),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14e932),
	.w1(32'hbd25fab5),
	.w2(32'hbace2027),
	.w3(32'hbbf939ff),
	.w4(32'h3c9b22ff),
	.w5(32'hbb5cb444),
	.w6(32'hbcde3b36),
	.w7(32'h3bc076ee),
	.w8(32'h3bd929de),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a2826),
	.w1(32'h3b460824),
	.w2(32'h3baf8618),
	.w3(32'hbb1bc928),
	.w4(32'h3a4e9de0),
	.w5(32'h3c679289),
	.w6(32'hbb45a820),
	.w7(32'h3b93bd2a),
	.w8(32'h3a265968),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6073a0),
	.w1(32'hbb50c2b3),
	.w2(32'h3c0da1da),
	.w3(32'h3ce4730c),
	.w4(32'h3c8cbbeb),
	.w5(32'h3ce12d02),
	.w6(32'h3bc7c13b),
	.w7(32'h3c42e8ca),
	.w8(32'h3d298cf5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc74a68),
	.w1(32'hbc101950),
	.w2(32'hbbe27ffc),
	.w3(32'h3bf00a4d),
	.w4(32'h3ace4063),
	.w5(32'hbb11c9c7),
	.w6(32'h3a7940b5),
	.w7(32'hbb1a01f8),
	.w8(32'hbb870f9c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813836),
	.w1(32'h3c66719f),
	.w2(32'h3c5a688f),
	.w3(32'h3bdbf09c),
	.w4(32'hbb90293c),
	.w5(32'h3b61d25f),
	.w6(32'hbc0a927e),
	.w7(32'hbd7ab7e9),
	.w8(32'h3c337657),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8700b5),
	.w1(32'hbcb1421f),
	.w2(32'hbb059781),
	.w3(32'h3c243266),
	.w4(32'h39de6841),
	.w5(32'h3be25153),
	.w6(32'h3c544b7c),
	.w7(32'hbb9cb074),
	.w8(32'h3b76db36),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9284e),
	.w1(32'hbb419a6d),
	.w2(32'h3c5719b5),
	.w3(32'hbbd7fc27),
	.w4(32'h3d91188b),
	.w5(32'h3bea8fe3),
	.w6(32'hbc3fec6f),
	.w7(32'h3bdedaab),
	.w8(32'hbbc120c1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5b47),
	.w1(32'hbacb08d8),
	.w2(32'h3d1b3175),
	.w3(32'hbb236ad7),
	.w4(32'hbbcdbae2),
	.w5(32'h3b01e9c3),
	.w6(32'hbc4418e8),
	.w7(32'h3afd1a63),
	.w8(32'h3baa5b3a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beccd2d),
	.w1(32'h3c458d35),
	.w2(32'h3beeb7fa),
	.w3(32'hba6d2a8b),
	.w4(32'hbb4b8864),
	.w5(32'hbc0213de),
	.w6(32'hbce69b6f),
	.w7(32'h3b6ceb9c),
	.w8(32'h3af7a8eb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd1c5b),
	.w1(32'h3b71c645),
	.w2(32'hbd04da09),
	.w3(32'h3c70731d),
	.w4(32'h3c851d20),
	.w5(32'h3aa2c5d8),
	.w6(32'h3c99d605),
	.w7(32'hbaf06b75),
	.w8(32'hbc974cf2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85e666),
	.w1(32'h3c0436dc),
	.w2(32'h3c6401f3),
	.w3(32'h3b40d75a),
	.w4(32'hbb1abda2),
	.w5(32'h3c04c66c),
	.w6(32'hbb130293),
	.w7(32'h3b7a4b5c),
	.w8(32'h3c0d04eb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac88f4a),
	.w1(32'hbc0d3cf3),
	.w2(32'h3cf24c58),
	.w3(32'h3802afc5),
	.w4(32'h3c38132f),
	.w5(32'h3c8eb630),
	.w6(32'hbb5c67c3),
	.w7(32'h3b9ac698),
	.w8(32'h3c821ffa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaec325),
	.w1(32'hbbc39681),
	.w2(32'hbb2286bd),
	.w3(32'hbb8e120e),
	.w4(32'hbc0dfeb7),
	.w5(32'hb967434e),
	.w6(32'h3b454976),
	.w7(32'h3bb865e9),
	.w8(32'hbb7888ee),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90a459),
	.w1(32'hbbe87ef3),
	.w2(32'hbb8a10b8),
	.w3(32'h3bf77c7d),
	.w4(32'h3a216501),
	.w5(32'hbae7a210),
	.w6(32'h3bbbfc28),
	.w7(32'h3b3e9eb9),
	.w8(32'hbbf1af51),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa11f6e),
	.w1(32'hbcd2bc25),
	.w2(32'hbbf3abf2),
	.w3(32'hbc22cf87),
	.w4(32'hbcbb0b9c),
	.w5(32'h3d222442),
	.w6(32'h3c23bfc9),
	.w7(32'hbbf547b9),
	.w8(32'h3b7f9306),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84fc03),
	.w1(32'hbb22ee0f),
	.w2(32'hbd50ac33),
	.w3(32'h3c2fbf30),
	.w4(32'hbba46d75),
	.w5(32'h3ba93aa3),
	.w6(32'h3bace4a4),
	.w7(32'h3a578092),
	.w8(32'h3b4dd414),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c158e26),
	.w1(32'h3b0913bf),
	.w2(32'h3c9b442f),
	.w3(32'hbbf3e60c),
	.w4(32'hbddb30f4),
	.w5(32'hbcccf43c),
	.w6(32'hbbe97191),
	.w7(32'hbbdcbbdd),
	.w8(32'h3c1d533f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31a3d0),
	.w1(32'hbae47ee6),
	.w2(32'h3d242e19),
	.w3(32'hbbdc372f),
	.w4(32'h3b6731e4),
	.w5(32'h3b22943d),
	.w6(32'h3b92799e),
	.w7(32'h3b9bcc76),
	.w8(32'hbb2eb3c0),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f455),
	.w1(32'hbb4c76cc),
	.w2(32'h3bac6e5f),
	.w3(32'h3c54b324),
	.w4(32'h3b9c441c),
	.w5(32'h3c3deece),
	.w6(32'h3a84fcf2),
	.w7(32'hbcd2cfc6),
	.w8(32'hbd137371),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c055dd2),
	.w1(32'hbc33d893),
	.w2(32'h3bf61065),
	.w3(32'h3bd0c2c3),
	.w4(32'h3babb133),
	.w5(32'h3b7e02ab),
	.w6(32'h3ac67159),
	.w7(32'hba72b55c),
	.w8(32'h3c8bab2f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b907),
	.w1(32'h3d143c1c),
	.w2(32'h3c18bed9),
	.w3(32'h3be491d6),
	.w4(32'h3c26ec40),
	.w5(32'h3c754ed1),
	.w6(32'h3a40c5c7),
	.w7(32'h3b37e135),
	.w8(32'h3abb9d3d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205ff1),
	.w1(32'h3b49bf42),
	.w2(32'hbbb167df),
	.w3(32'hbc21539a),
	.w4(32'hbbd960aa),
	.w5(32'h3bf6c92d),
	.w6(32'hba85a62d),
	.w7(32'h3b0934a4),
	.w8(32'h3b0b968f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7ff33),
	.w1(32'h3be12711),
	.w2(32'hbca4abf8),
	.w3(32'hbc2e28a1),
	.w4(32'hbbaa7ab8),
	.w5(32'hbc615cba),
	.w6(32'h3b465cf0),
	.w7(32'hbbfc453e),
	.w8(32'hbba45e0c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa817d),
	.w1(32'h3d40e6f5),
	.w2(32'hbc216356),
	.w3(32'h3d13e940),
	.w4(32'h3d41bfa8),
	.w5(32'h3c23bfcf),
	.w6(32'h3d342b9c),
	.w7(32'h3ca5051f),
	.w8(32'hbd011047),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190554),
	.w1(32'h3b270650),
	.w2(32'h3bc3c238),
	.w3(32'hbc2d8b7f),
	.w4(32'hbc439e5d),
	.w5(32'h3bc1d700),
	.w6(32'hbc3c8b83),
	.w7(32'hbc1a5f31),
	.w8(32'h3ca84e05),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8da9a8),
	.w1(32'hbc8cadb0),
	.w2(32'h3bc39820),
	.w3(32'hbcfcb60e),
	.w4(32'hbcf36597),
	.w5(32'hbc88ae98),
	.w6(32'hbc7823b7),
	.w7(32'hbd18888c),
	.w8(32'hbc3d80ee),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6408e6),
	.w1(32'h3b93100a),
	.w2(32'h3a3f1f29),
	.w3(32'h3aac0782),
	.w4(32'hbb816624),
	.w5(32'hb910de46),
	.w6(32'h3caa2592),
	.w7(32'h3b581d87),
	.w8(32'hbcd1ef9e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba564a40),
	.w1(32'hbbbbe0f5),
	.w2(32'h38fb05e1),
	.w3(32'hbc8da86e),
	.w4(32'hbc0f6916),
	.w5(32'h3c4783f4),
	.w6(32'h3a8be003),
	.w7(32'h3b53b08f),
	.w8(32'h3b0bb682),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a9e9),
	.w1(32'hbc8b53b7),
	.w2(32'h3c725ed8),
	.w3(32'hba7dcae8),
	.w4(32'h3d5f1f9f),
	.w5(32'hbc4e2107),
	.w6(32'h3afeefb2),
	.w7(32'hbb29b6f8),
	.w8(32'h3bb7200a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83de08),
	.w1(32'hbbf7cca5),
	.w2(32'hbbddc733),
	.w3(32'hbbb6735a),
	.w4(32'hbc9d3fd5),
	.w5(32'h3b5f19c6),
	.w6(32'h3a174566),
	.w7(32'hbb7ea400),
	.w8(32'hb991285e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae17671),
	.w1(32'hbc7bb5d1),
	.w2(32'h3c9264cf),
	.w3(32'h3b9c3b8b),
	.w4(32'h3a1f5b63),
	.w5(32'h3be56564),
	.w6(32'hbaf9a9fb),
	.w7(32'hbc55fed9),
	.w8(32'h3b3955e7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e0098),
	.w1(32'hbcabffc8),
	.w2(32'h3c05e0ad),
	.w3(32'hbae998b2),
	.w4(32'hb9438873),
	.w5(32'h3c9abad0),
	.w6(32'hbabbd17e),
	.w7(32'hbba1ea3d),
	.w8(32'h3bcb7a6e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28b802),
	.w1(32'h3c072903),
	.w2(32'h3c56ae0d),
	.w3(32'hba31dd80),
	.w4(32'h3c0292a7),
	.w5(32'h3c62cc36),
	.w6(32'hbc533098),
	.w7(32'h3c1ffa40),
	.w8(32'h3c22eb32),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55df3d),
	.w1(32'h3ba52d20),
	.w2(32'h3bf6e2f2),
	.w3(32'hbc2f8108),
	.w4(32'h3b740ab8),
	.w5(32'h3b058829),
	.w6(32'hbb0f31bf),
	.w7(32'h3be6be98),
	.w8(32'h3c264f71),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c804229),
	.w1(32'hba493679),
	.w2(32'hbc92580a),
	.w3(32'h3c13ce01),
	.w4(32'h3c673846),
	.w5(32'hbc0f17a6),
	.w6(32'hbcc777dc),
	.w7(32'h3c5b1fe6),
	.w8(32'hbcc5f910),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba40ce),
	.w1(32'h3c6fb628),
	.w2(32'h3b94dd64),
	.w3(32'hbc75fd8d),
	.w4(32'h3a835011),
	.w5(32'h3b30641d),
	.w6(32'h3acf8fef),
	.w7(32'hbbe4a999),
	.w8(32'h3b2c3940),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc988641),
	.w1(32'h3c4eb13b),
	.w2(32'hba2b72d2),
	.w3(32'hbc7299b6),
	.w4(32'hbb6c09bb),
	.w5(32'hbc550934),
	.w6(32'h3c2d3ef0),
	.w7(32'hbaddbe1f),
	.w8(32'hbb6bff45),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b4fc8),
	.w1(32'h37e454d0),
	.w2(32'h3badb8fc),
	.w3(32'h3acba70e),
	.w4(32'h3b35527a),
	.w5(32'h39e160f7),
	.w6(32'hbc2a6f50),
	.w7(32'hbaabd979),
	.w8(32'h3b40f6a5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52d7d),
	.w1(32'h3c3077e0),
	.w2(32'h3c1f48d6),
	.w3(32'hbd695216),
	.w4(32'hbd118d2e),
	.w5(32'hb9c7ce0b),
	.w6(32'h3a7015b1),
	.w7(32'hba82a04b),
	.w8(32'hbb63308c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82e485),
	.w1(32'hba7aad45),
	.w2(32'hb63f3405),
	.w3(32'hba40e626),
	.w4(32'hbb97206a),
	.w5(32'h3c3ed89f),
	.w6(32'hbb4f21ee),
	.w7(32'h3a74dff2),
	.w8(32'h3c77bbf9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e896f),
	.w1(32'h3c16c4e7),
	.w2(32'h39d586d8),
	.w3(32'hba49a802),
	.w4(32'h3b4c22b3),
	.w5(32'hbb4a4d3d),
	.w6(32'h3c9d3e37),
	.w7(32'hbbab4447),
	.w8(32'hbc4ba68e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb422),
	.w1(32'hba940aa2),
	.w2(32'hbbdb5041),
	.w3(32'h3adfb1d9),
	.w4(32'hbc75641c),
	.w5(32'hbcee3c03),
	.w6(32'hbb39b978),
	.w7(32'hbaf00bbc),
	.w8(32'hba8ccea7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47a592),
	.w1(32'h3bd5fbfc),
	.w2(32'h3acd9ac9),
	.w3(32'hbb914125),
	.w4(32'hbb875b51),
	.w5(32'h3bbccd00),
	.w6(32'h3be5ab73),
	.w7(32'hb9cdfa5e),
	.w8(32'h3acfebb1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1e55e),
	.w1(32'h3b9ee7d6),
	.w2(32'hb981a546),
	.w3(32'h3cba0c00),
	.w4(32'h3afdb955),
	.w5(32'hbc5249ff),
	.w6(32'hbbec9f14),
	.w7(32'hbaf0d64d),
	.w8(32'hbb0d3b35),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0772c8),
	.w1(32'h3bae23a3),
	.w2(32'hbb560309),
	.w3(32'h3c83e964),
	.w4(32'hbba8b191),
	.w5(32'h3a0a3d24),
	.w6(32'hbb802523),
	.w7(32'hbb7aeea0),
	.w8(32'h3c865293),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf32fa1),
	.w1(32'hba197107),
	.w2(32'h3b874c49),
	.w3(32'h3c28eb70),
	.w4(32'h3b22d14c),
	.w5(32'h3bacb0c1),
	.w6(32'hbc240bac),
	.w7(32'hbcae9b8d),
	.w8(32'hbb2ad13d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c162d20),
	.w1(32'h3b127e86),
	.w2(32'hbace66d3),
	.w3(32'h3c5dc0d5),
	.w4(32'h3b0f2cfc),
	.w5(32'h37ccef63),
	.w6(32'hbbda2fe6),
	.w7(32'hbbe3100a),
	.w8(32'h3a3ee409),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9245cc),
	.w1(32'h3b802d2e),
	.w2(32'h3ac64a22),
	.w3(32'h3b0ba716),
	.w4(32'h3bc3d237),
	.w5(32'h39d97110),
	.w6(32'hbccb9c4c),
	.w7(32'h3bed4374),
	.w8(32'h3ac89c8b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d67d),
	.w1(32'hbab2ee16),
	.w2(32'h3c2c4a29),
	.w3(32'hbb554dc9),
	.w4(32'h3ada12bf),
	.w5(32'h3c176133),
	.w6(32'hbc48af85),
	.w7(32'h393166b7),
	.w8(32'h3c956774),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77737a),
	.w1(32'h3bb7ae46),
	.w2(32'hb9084367),
	.w3(32'hbb9a6654),
	.w4(32'hbb7e83f3),
	.w5(32'h3c2cb578),
	.w6(32'h3bac3904),
	.w7(32'h3b71e4ad),
	.w8(32'h3b44ae02),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62afe2),
	.w1(32'hbd29105c),
	.w2(32'h3bc4accc),
	.w3(32'hb9d1d4c7),
	.w4(32'h3b5cfa7a),
	.w5(32'hbc188f51),
	.w6(32'h3b5b6b62),
	.w7(32'hbb93d5ff),
	.w8(32'hbb9c78fe),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb304e4),
	.w1(32'h3b2d5f62),
	.w2(32'hbacbf40f),
	.w3(32'hbbe94faf),
	.w4(32'hbab0f308),
	.w5(32'h3b112672),
	.w6(32'hbba847d4),
	.w7(32'h3acf887b),
	.w8(32'h3a5f9176),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3ec68),
	.w1(32'hbc5257b7),
	.w2(32'h3b1770fe),
	.w3(32'h3c081fe0),
	.w4(32'h3b96b5a2),
	.w5(32'hbb81715d),
	.w6(32'hbae8008b),
	.w7(32'hbbe920d3),
	.w8(32'hbcb6a11a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd73aa8),
	.w1(32'h3bba6f14),
	.w2(32'h3a753344),
	.w3(32'h3bb173f4),
	.w4(32'h3bfadeb6),
	.w5(32'h3c7c1175),
	.w6(32'h3c892f08),
	.w7(32'h3b534f3e),
	.w8(32'h3c8824b6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa1ad9),
	.w1(32'h3b149e7d),
	.w2(32'hbbf8d699),
	.w3(32'h3b2137a2),
	.w4(32'hb9fabbca),
	.w5(32'h3a98dec0),
	.w6(32'hbc0469a9),
	.w7(32'h3c373dc6),
	.w8(32'h3c98157b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf02861),
	.w1(32'hbd3e544b),
	.w2(32'h3c8e42ce),
	.w3(32'h3b4cac2a),
	.w4(32'h39a5c538),
	.w5(32'h3bd011cc),
	.w6(32'h3a673be3),
	.w7(32'h3b20bb47),
	.w8(32'h3c661232),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8682e1),
	.w1(32'h3c1f82a8),
	.w2(32'hbba91334),
	.w3(32'hbb498a90),
	.w4(32'hbc52623c),
	.w5(32'h3b9884f5),
	.w6(32'h3b8dec97),
	.w7(32'hbc376864),
	.w8(32'h3c70837c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb67aad),
	.w1(32'hbb2043e3),
	.w2(32'hbc4ddb02),
	.w3(32'hba88ab18),
	.w4(32'h3c20ab80),
	.w5(32'h3c049f52),
	.w6(32'h3c13064e),
	.w7(32'hbc689dd0),
	.w8(32'h3c43ab25),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a48b4),
	.w1(32'hb9f08a6d),
	.w2(32'hbb247e70),
	.w3(32'hbb5fe726),
	.w4(32'h3bb19b98),
	.w5(32'h3b4d7cad),
	.w6(32'hbbe5c414),
	.w7(32'h3b49f16f),
	.w8(32'hbbf69c8d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef36b3),
	.w1(32'h3bc98d9e),
	.w2(32'h3aa11b63),
	.w3(32'hbbed193a),
	.w4(32'hbbd64381),
	.w5(32'h3ce7c8d0),
	.w6(32'hbb113fe7),
	.w7(32'hbbe3350b),
	.w8(32'h3b304a4f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bc030),
	.w1(32'h3aa5b2f0),
	.w2(32'hbc033ae8),
	.w3(32'hbc5c3cdf),
	.w4(32'h3bf30c60),
	.w5(32'hbb292bb3),
	.w6(32'h3c239879),
	.w7(32'hbb940c41),
	.w8(32'h3c8fbb5a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccd9dc),
	.w1(32'hb9ad9332),
	.w2(32'h39906159),
	.w3(32'hbc0aa52e),
	.w4(32'h3ce289ab),
	.w5(32'hbbf4ca47),
	.w6(32'hbd129c01),
	.w7(32'hba77495c),
	.w8(32'h3ca594e4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b835223),
	.w1(32'h3b803968),
	.w2(32'hbd047aa7),
	.w3(32'h3c60aac2),
	.w4(32'h3bc31d9c),
	.w5(32'hba861db1),
	.w6(32'h3cc7d650),
	.w7(32'h39396d96),
	.w8(32'hbc37e2f2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45ac90),
	.w1(32'hbccbcaf0),
	.w2(32'h3bb07822),
	.w3(32'h3c7a34a6),
	.w4(32'hbbf6c5c3),
	.w5(32'h3c10bfbb),
	.w6(32'h3cbed80a),
	.w7(32'h3bd0c87b),
	.w8(32'h3c364e61),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c541799),
	.w1(32'h3b3fdc96),
	.w2(32'h3c8475c8),
	.w3(32'h3c3ef6ae),
	.w4(32'h3b9f625d),
	.w5(32'h3c44ca8c),
	.w6(32'h3ba4c054),
	.w7(32'hbce0dba2),
	.w8(32'h3cc9fb53),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad32b8d),
	.w1(32'h3b61bb38),
	.w2(32'hbb755d26),
	.w3(32'h3abb20f6),
	.w4(32'h3b968914),
	.w5(32'h3b0393d9),
	.w6(32'h3c9b98d5),
	.w7(32'hbb7082c7),
	.w8(32'h3bfa7aa5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35f3b8),
	.w1(32'h3b9f70ef),
	.w2(32'hbc755808),
	.w3(32'hb9dae7de),
	.w4(32'hbbee0dcf),
	.w5(32'h3c73f569),
	.w6(32'h3be61bf8),
	.w7(32'h3d8c3376),
	.w8(32'h3b16c44b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8247c06),
	.w1(32'hbbd7e22d),
	.w2(32'h3bb960b0),
	.w3(32'hbb9243c2),
	.w4(32'hbc5444a4),
	.w5(32'h3c9dcc52),
	.w6(32'hba489beb),
	.w7(32'hbb902394),
	.w8(32'h3b1f571c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc3ca5),
	.w1(32'h3cf5f668),
	.w2(32'hbbb4131a),
	.w3(32'h3c528782),
	.w4(32'hbaee6641),
	.w5(32'h3c11c5b4),
	.w6(32'hbabdef76),
	.w7(32'hba1528fc),
	.w8(32'h3c463dae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f40f1),
	.w1(32'hbc5e8ff1),
	.w2(32'h3b7dc437),
	.w3(32'h3b731988),
	.w4(32'h3c8a9464),
	.w5(32'hbbcd877d),
	.w6(32'h3b165e3c),
	.w7(32'hbc0e7c5d),
	.w8(32'hbb60f795),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb8a9),
	.w1(32'h3c337b24),
	.w2(32'h3b429305),
	.w3(32'h3aa2719f),
	.w4(32'h3b30f127),
	.w5(32'hba33eff9),
	.w6(32'h3b9c05a0),
	.w7(32'h3bc22814),
	.w8(32'hb71a4f0c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe67cad),
	.w1(32'h3b99edd1),
	.w2(32'hbcc65667),
	.w3(32'h3b0fa1c2),
	.w4(32'h3c28f9eb),
	.w5(32'h3b11fc06),
	.w6(32'hbc605a41),
	.w7(32'h3c2e4a30),
	.w8(32'h3b08a79f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08cd56),
	.w1(32'h3b7486c1),
	.w2(32'h3c09a150),
	.w3(32'h399cac4c),
	.w4(32'hbba5dfc4),
	.w5(32'hbada61f1),
	.w6(32'hbc2bd005),
	.w7(32'hbb8296cd),
	.w8(32'hbb417013),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881f181),
	.w1(32'h3cbf500e),
	.w2(32'h3c1676c1),
	.w3(32'h3b22e88a),
	.w4(32'h39f25c07),
	.w5(32'h3c8e3327),
	.w6(32'h3c02ed32),
	.w7(32'h3c841c58),
	.w8(32'h3c4a6a89),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc558190),
	.w1(32'hbb80b692),
	.w2(32'h3b82641f),
	.w3(32'h3b68c0ce),
	.w4(32'hbc7e380b),
	.w5(32'hbbb8e99b),
	.w6(32'h3b9eba23),
	.w7(32'h3b088294),
	.w8(32'h3c6dc9bf),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca08718),
	.w1(32'h3c39d9c9),
	.w2(32'h3bce04c4),
	.w3(32'hb9bebbd7),
	.w4(32'h3bf5206b),
	.w5(32'h3c2c7b00),
	.w6(32'h3c564d76),
	.w7(32'hbbab5a76),
	.w8(32'h3be5fc99),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91cda6),
	.w1(32'h3c400ba6),
	.w2(32'hbc75f906),
	.w3(32'h3b57fde1),
	.w4(32'hbc2c90b3),
	.w5(32'h3c29ded9),
	.w6(32'h3c4a176f),
	.w7(32'hbc2c5daf),
	.w8(32'h3c40cdc9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81e969),
	.w1(32'hb9c955f7),
	.w2(32'hbc174cae),
	.w3(32'hbc038ef1),
	.w4(32'hbc887cb0),
	.w5(32'hbb132f3c),
	.w6(32'hbc81a612),
	.w7(32'hbc0fe2d8),
	.w8(32'hbb0d320d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86d0cb),
	.w1(32'hbc04f924),
	.w2(32'h3aa73d5b),
	.w3(32'h3c7dc807),
	.w4(32'h3bfeb218),
	.w5(32'hbc356120),
	.w6(32'h3ca5fd74),
	.w7(32'h3c15b558),
	.w8(32'hbc02e911),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe070e),
	.w1(32'h3b198b8e),
	.w2(32'h3bcd8583),
	.w3(32'hbc0726bf),
	.w4(32'hbbecf092),
	.w5(32'hbbab8f79),
	.w6(32'hbca07edd),
	.w7(32'hbc958c69),
	.w8(32'hb830bebc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f4590),
	.w1(32'hbc3748c8),
	.w2(32'hbb854846),
	.w3(32'h3c21f4f3),
	.w4(32'h3ca1cfbc),
	.w5(32'h3bca7c2c),
	.w6(32'h3bbe3ed7),
	.w7(32'h3cad0b23),
	.w8(32'h3ceff309),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc221b30),
	.w1(32'hbb4d97a6),
	.w2(32'h3b12e64a),
	.w3(32'h3c14e47a),
	.w4(32'h3c8c2712),
	.w5(32'h3b95df00),
	.w6(32'h3b21e8b0),
	.w7(32'h3c650512),
	.w8(32'h3c715df8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e5075),
	.w1(32'hbb20aa51),
	.w2(32'h3b3d11d1),
	.w3(32'hbb8c8d76),
	.w4(32'hbc2ff4c6),
	.w5(32'h3b3b3c43),
	.w6(32'hbb3182fa),
	.w7(32'hbc126af3),
	.w8(32'h3c5cd2a4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b407872),
	.w1(32'h3c3af655),
	.w2(32'h3b857411),
	.w3(32'h3c1beec0),
	.w4(32'h3c55aa97),
	.w5(32'hbc04c959),
	.w6(32'hbc0fe632),
	.w7(32'h3c031135),
	.w8(32'hb9b40a28),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cc363),
	.w1(32'h3c654d62),
	.w2(32'h3c31d7c3),
	.w3(32'h3be9b46f),
	.w4(32'h3bdec256),
	.w5(32'h3b93b9d1),
	.w6(32'hbb83d7d5),
	.w7(32'hb791ae5a),
	.w8(32'hbb68ffbc),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f0bc9),
	.w1(32'hbc306fad),
	.w2(32'hbc025bcc),
	.w3(32'hbc89020b),
	.w4(32'hba956926),
	.w5(32'hbc3e0cd3),
	.w6(32'h3bd158c5),
	.w7(32'hbce8b6f7),
	.w8(32'hbbbb7967),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c12d2),
	.w1(32'h3cc32200),
	.w2(32'hbbc6e90b),
	.w3(32'h3b2e0eb1),
	.w4(32'h3cea2f61),
	.w5(32'hbba54474),
	.w6(32'h3ce2f773),
	.w7(32'h3cd3567e),
	.w8(32'h3a879fc7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8bfae),
	.w1(32'hbbd3c22f),
	.w2(32'h3c5aab44),
	.w3(32'hbc881cb0),
	.w4(32'hbc54a53a),
	.w5(32'h3c3a4c57),
	.w6(32'hbbc404d2),
	.w7(32'hbc9f1e4f),
	.w8(32'h3ca80ddd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba57fa1),
	.w1(32'h3b8763b7),
	.w2(32'h3ca7062e),
	.w3(32'h3b723ae7),
	.w4(32'h3cbd610a),
	.w5(32'h3bd33a3d),
	.w6(32'h3a98564e),
	.w7(32'h3add6089),
	.w8(32'h3c49af8a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c849da3),
	.w1(32'h3c6d8331),
	.w2(32'hbc598748),
	.w3(32'h3cac08ef),
	.w4(32'h3c5158d9),
	.w5(32'hbb90bc08),
	.w6(32'h3ca7db8f),
	.w7(32'hbc011769),
	.w8(32'hbc65f57c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966d947),
	.w1(32'h3af57abc),
	.w2(32'h3c5a0cb6),
	.w3(32'hba3bceaa),
	.w4(32'h3ac52275),
	.w5(32'hbb470183),
	.w6(32'hbb1d9673),
	.w7(32'h3c17cce8),
	.w8(32'h3ce0e668),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f0c2),
	.w1(32'h3cbb0de4),
	.w2(32'h3aef15dd),
	.w3(32'h3c274180),
	.w4(32'h3d0c5e7b),
	.w5(32'h3bece5e6),
	.w6(32'h3c4ff07a),
	.w7(32'h3cd1642f),
	.w8(32'hbc57f66f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c222192),
	.w1(32'hbb9d9347),
	.w2(32'hbc5320c0),
	.w3(32'hbbf91627),
	.w4(32'hbc99b150),
	.w5(32'hbc86b4a2),
	.w6(32'hbb1251fb),
	.w7(32'hbc37c376),
	.w8(32'hbc2d23ba),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e43ab),
	.w1(32'h3c1c46ae),
	.w2(32'h3c59211e),
	.w3(32'h3c23a82b),
	.w4(32'hb92a41c6),
	.w5(32'h3a4c5638),
	.w6(32'hbbe9e089),
	.w7(32'h3abb46f3),
	.w8(32'h38a9d6a5),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135e85),
	.w1(32'h3b75ccf0),
	.w2(32'h3ba6d21b),
	.w3(32'hbb594a60),
	.w4(32'h3c0bd2de),
	.w5(32'h3bfd5ced),
	.w6(32'hbc2d0c1c),
	.w7(32'h3b52b16e),
	.w8(32'hbb6b41a1),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce225a4),
	.w1(32'hbc2c829f),
	.w2(32'h3bcae34a),
	.w3(32'h3c9b5aae),
	.w4(32'hbbac4c9f),
	.w5(32'hbc4e62f9),
	.w6(32'h3c99fe1d),
	.w7(32'hbc3fd6ac),
	.w8(32'hbbf8413c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d8992),
	.w1(32'hbac8ed6f),
	.w2(32'h3b89ee1e),
	.w3(32'hbc057a2a),
	.w4(32'hbba85e56),
	.w5(32'h3c8a0795),
	.w6(32'h3bb21ba9),
	.w7(32'h3b9af261),
	.w8(32'h3c28471f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb2b6),
	.w1(32'hbc09f553),
	.w2(32'hbc33aae3),
	.w3(32'hbcacdb51),
	.w4(32'hbca1907f),
	.w5(32'hbce2387e),
	.w6(32'h3be238e5),
	.w7(32'hbbfb8604),
	.w8(32'h39b28a75),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9863b5),
	.w1(32'h3b766c00),
	.w2(32'hbb60c29c),
	.w3(32'h3b4745bd),
	.w4(32'h37a55206),
	.w5(32'h3c17642b),
	.w6(32'hbb016ab3),
	.w7(32'h3bcb8ae7),
	.w8(32'h3bb924ad),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94e932),
	.w1(32'h3c7ef728),
	.w2(32'h3bec42f8),
	.w3(32'h3c46fc24),
	.w4(32'h3c99967e),
	.w5(32'h3b59dcff),
	.w6(32'hbbf78b5d),
	.w7(32'h3c011582),
	.w8(32'hbb0f6eff),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bcc0b),
	.w1(32'hbbdccedf),
	.w2(32'h3c28355d),
	.w3(32'hbbab04e4),
	.w4(32'h3d36ee86),
	.w5(32'h3caaf81d),
	.w6(32'hbbbdf2b4),
	.w7(32'h3c04d54a),
	.w8(32'h3c9dadf2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be042b2),
	.w1(32'h3a9c1056),
	.w2(32'hb9655344),
	.w3(32'hbacfeca8),
	.w4(32'hbbf81e8a),
	.w5(32'hbbeb9bf4),
	.w6(32'hbaccb319),
	.w7(32'h3c139390),
	.w8(32'hbbe2c58c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9910b4),
	.w1(32'hbb7408bb),
	.w2(32'h3977f170),
	.w3(32'hbba72fe1),
	.w4(32'h3bb8327a),
	.w5(32'hbb23ee6d),
	.w6(32'hbb95fd20),
	.w7(32'h3aadbb7e),
	.w8(32'h3b819b57),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8489d22),
	.w1(32'h3b8d9351),
	.w2(32'h3c04dde3),
	.w3(32'h3be3118f),
	.w4(32'h3ce292e5),
	.w5(32'h3cbb1d7b),
	.w6(32'hba3dd5d1),
	.w7(32'h3b8dd163),
	.w8(32'h3d083a16),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc820ac),
	.w1(32'h3c590dd0),
	.w2(32'hbbc489f4),
	.w3(32'hbc8661e6),
	.w4(32'h39a6ebe7),
	.w5(32'h39d44c1d),
	.w6(32'h3c4cbc4a),
	.w7(32'h3a39610e),
	.w8(32'hbaf3b63e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb39d11),
	.w1(32'hbc6db682),
	.w2(32'h3bd12a72),
	.w3(32'hb792d60e),
	.w4(32'h3c083abe),
	.w5(32'h3b975668),
	.w6(32'h3a91380f),
	.w7(32'hb950fe48),
	.w8(32'h3c5da465),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfcacf8),
	.w1(32'h3be3d370),
	.w2(32'h3b4b4543),
	.w3(32'hbbf12375),
	.w4(32'hbc3c2ad5),
	.w5(32'h3bd5a592),
	.w6(32'hbb836a21),
	.w7(32'h3cf34b25),
	.w8(32'hbb13a588),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9204),
	.w1(32'hbbdf2407),
	.w2(32'hbc800f8a),
	.w3(32'hbc1b613d),
	.w4(32'h3bbf64da),
	.w5(32'hbc957f30),
	.w6(32'h3c42c855),
	.w7(32'h3c8670c8),
	.w8(32'hbb08fde2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a2cbd),
	.w1(32'hbc09c913),
	.w2(32'hbc6abd3f),
	.w3(32'hbb5b1986),
	.w4(32'h3cd0b8ae),
	.w5(32'hbbdc9173),
	.w6(32'h3c8edeba),
	.w7(32'hbb23c912),
	.w8(32'h3a47ca83),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ad626),
	.w1(32'h3bd3afa7),
	.w2(32'h3cb17e72),
	.w3(32'h3bf7eb6a),
	.w4(32'h3c9c6977),
	.w5(32'hbb271d88),
	.w6(32'hbc8438de),
	.w7(32'h3be6c766),
	.w8(32'h3cf2de73),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffb12a),
	.w1(32'hbc807945),
	.w2(32'hbbdbedfa),
	.w3(32'hbae98152),
	.w4(32'hbca2cf00),
	.w5(32'hbbe57ba8),
	.w6(32'hbbaa2b5a),
	.w7(32'h3b0b175e),
	.w8(32'hbafa0c6c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1acbe3),
	.w1(32'h3c0027a7),
	.w2(32'hbc35eb6c),
	.w3(32'h3c22e6e4),
	.w4(32'h39ed669c),
	.w5(32'h3c3de931),
	.w6(32'hbb906907),
	.w7(32'hbb62cb88),
	.w8(32'h3be139ce),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ff31),
	.w1(32'hb9ca81a0),
	.w2(32'h3c9bf774),
	.w3(32'hbbbe8b9f),
	.w4(32'hbb898331),
	.w5(32'hbc57ac65),
	.w6(32'hbb10d3ca),
	.w7(32'h3c3d15bb),
	.w8(32'hbb8ef05e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c535f),
	.w1(32'hbc34ca3e),
	.w2(32'h3bed0153),
	.w3(32'h3c38a8b0),
	.w4(32'hba881f3a),
	.w5(32'hbc996524),
	.w6(32'hbb5e3100),
	.w7(32'hbce68178),
	.w8(32'hb92f765c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be64cdb),
	.w1(32'hbcba9c76),
	.w2(32'hbcac694c),
	.w3(32'h3c18c494),
	.w4(32'h3bff4e03),
	.w5(32'hbc7d7aea),
	.w6(32'h3b004de7),
	.w7(32'hbbe0b499),
	.w8(32'hbc046aba),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf51a02),
	.w1(32'h3b2970c0),
	.w2(32'h3b61454f),
	.w3(32'h3c738af6),
	.w4(32'h3c732ef3),
	.w5(32'h3c23a475),
	.w6(32'h3c2b80d2),
	.w7(32'hbc1e114e),
	.w8(32'h3ae88d57),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb72da8),
	.w1(32'h3c7e4c50),
	.w2(32'hbb10f35e),
	.w3(32'h3aaf2852),
	.w4(32'h3b191662),
	.w5(32'hbbd396c0),
	.w6(32'h3ad0d53f),
	.w7(32'hba853a81),
	.w8(32'h3ab1eab8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a7880),
	.w1(32'h3b83dd95),
	.w2(32'h3a4942d6),
	.w3(32'hbcd851d3),
	.w4(32'hbb7427ec),
	.w5(32'h3cd82c9f),
	.w6(32'hbb6ec987),
	.w7(32'h3c212967),
	.w8(32'h3c98aeae),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9144),
	.w1(32'h3bbb3ec6),
	.w2(32'h3b9fd495),
	.w3(32'h3ad7f328),
	.w4(32'h3cb655c8),
	.w5(32'hb9bd2b67),
	.w6(32'h3b6f0898),
	.w7(32'h3c05f9f6),
	.w8(32'h3b55e332),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fd9b0),
	.w1(32'h3ab7eaad),
	.w2(32'h3c13cc69),
	.w3(32'hba9bbafb),
	.w4(32'h3b8c58ac),
	.w5(32'h3cf51de0),
	.w6(32'h39c4f256),
	.w7(32'hbbdb52d9),
	.w8(32'h3c8296c0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836bd9),
	.w1(32'hbbde134e),
	.w2(32'hbbc65358),
	.w3(32'h3c0a2d0f),
	.w4(32'h3c94e2bf),
	.w5(32'h3cbcc063),
	.w6(32'h3b320d5d),
	.w7(32'h3c265cfc),
	.w8(32'hbb556dcb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccee3d9),
	.w1(32'hbbb4b407),
	.w2(32'hbcdb6343),
	.w3(32'h3c4eda61),
	.w4(32'hbb244438),
	.w5(32'h39aa8f09),
	.w6(32'h3af7627f),
	.w7(32'h3aa94254),
	.w8(32'h3af33652),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a6e6c),
	.w1(32'h3bb8167a),
	.w2(32'h3b45b114),
	.w3(32'hbc04556b),
	.w4(32'hbc15d0cc),
	.w5(32'h3b8f0dd3),
	.w6(32'hbb7f1464),
	.w7(32'h3b062318),
	.w8(32'h3b965fe7),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cb34a),
	.w1(32'hbba14ad5),
	.w2(32'hbb861b63),
	.w3(32'h3ba8b582),
	.w4(32'h3c127a76),
	.w5(32'h3c9a0dd6),
	.w6(32'h3c5945ca),
	.w7(32'h3bbf71b7),
	.w8(32'h3b0a20bd),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18493f),
	.w1(32'h3c341d12),
	.w2(32'hbc261485),
	.w3(32'h3b535535),
	.w4(32'h3c4d1655),
	.w5(32'hbc1c77a3),
	.w6(32'h3bfdbfab),
	.w7(32'h3bab2cf1),
	.w8(32'hbc912267),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca01800),
	.w1(32'h3c63442a),
	.w2(32'h3c88f906),
	.w3(32'h3c04d79e),
	.w4(32'h3cd14cd3),
	.w5(32'h3ca1481b),
	.w6(32'hbc8173d7),
	.w7(32'hbaaeaa49),
	.w8(32'h3c743f58),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d51ad),
	.w1(32'hbb18b476),
	.w2(32'h3adb099b),
	.w3(32'h3c62217f),
	.w4(32'h3c16cf18),
	.w5(32'h3ad396d7),
	.w6(32'hbb92499a),
	.w7(32'h3acea56d),
	.w8(32'h3bd06c20),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2420d5),
	.w1(32'h3ad07487),
	.w2(32'h3b58ab59),
	.w3(32'h3c258067),
	.w4(32'hbc395d4f),
	.w5(32'hba88f01d),
	.w6(32'hbc68f846),
	.w7(32'h3c4016d2),
	.w8(32'h3b128f62),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c3024),
	.w1(32'hbc5055e0),
	.w2(32'h3c862b23),
	.w3(32'hbd0cdfca),
	.w4(32'hbd82c80f),
	.w5(32'hbc987b08),
	.w6(32'h3b1f0bac),
	.w7(32'hbce362c1),
	.w8(32'h3cadca0c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61c61b),
	.w1(32'h3a8f8e5e),
	.w2(32'h3b8f7bf6),
	.w3(32'h3b984098),
	.w4(32'h3c40436a),
	.w5(32'h3caf86e5),
	.w6(32'hba168d42),
	.w7(32'h3c3147d5),
	.w8(32'hbc4d02b5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cba38db),
	.w1(32'h3b9dcb50),
	.w2(32'hbbb8042b),
	.w3(32'hbbd70523),
	.w4(32'hba305838),
	.w5(32'hbb6040c9),
	.w6(32'h3aeaa4cd),
	.w7(32'hbc03449f),
	.w8(32'h3c60dcad),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc86dc6),
	.w1(32'hbc356a6b),
	.w2(32'h3c70e7bf),
	.w3(32'hbbcfe908),
	.w4(32'hbb4de90d),
	.w5(32'hbb5a4abf),
	.w6(32'h3c37cf66),
	.w7(32'hba9da87a),
	.w8(32'hbbd40edd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340a4a),
	.w1(32'h3c2a7899),
	.w2(32'hbce8ef46),
	.w3(32'hb93c3f2d),
	.w4(32'hbcc3ef0d),
	.w5(32'hbc620dd7),
	.w6(32'hbbb2eee4),
	.w7(32'h3d290cf1),
	.w8(32'hb944eb0b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f08b),
	.w1(32'hb911eaff),
	.w2(32'hbb2531cf),
	.w3(32'hbb9d7b6d),
	.w4(32'h3c2edaa8),
	.w5(32'h3c89a457),
	.w6(32'hbbf3b223),
	.w7(32'hbbd06b27),
	.w8(32'h3bea9bfb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12219d),
	.w1(32'hbb5a71ca),
	.w2(32'h3b8d63ab),
	.w3(32'hbb6d367a),
	.w4(32'h3ca7a88b),
	.w5(32'h3b0274f0),
	.w6(32'hbabb9dbc),
	.w7(32'hbcc09095),
	.w8(32'h3bba751d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d83f),
	.w1(32'hbcda2618),
	.w2(32'h3a890bf8),
	.w3(32'hbc3e0d57),
	.w4(32'hbc7b0570),
	.w5(32'h3bc812ba),
	.w6(32'hbab7cbcb),
	.w7(32'h3b51a770),
	.w8(32'hbc1efb03),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c741d03),
	.w1(32'hbb3db239),
	.w2(32'hbc7702a1),
	.w3(32'h3b92f71a),
	.w4(32'hbb3a02c4),
	.w5(32'hbb0b536f),
	.w6(32'h3c765183),
	.w7(32'hbb627595),
	.w8(32'h3c5e1a8a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe2044),
	.w1(32'h3c647c37),
	.w2(32'h3c21e4d4),
	.w3(32'hbae0cb83),
	.w4(32'hbbcc36dd),
	.w5(32'hbbc6e2bf),
	.w6(32'h3bcac5a1),
	.w7(32'h3cc8b3e6),
	.w8(32'hbcbfde0f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c907758),
	.w1(32'h3c60b24d),
	.w2(32'hbca7856d),
	.w3(32'h3c758bd9),
	.w4(32'hba30786b),
	.w5(32'hbba25a82),
	.w6(32'hbb939fbb),
	.w7(32'h3be4d010),
	.w8(32'hbcf4bcd3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a23ab),
	.w1(32'h3bf5e209),
	.w2(32'h3aa0d33e),
	.w3(32'hbc6bdb15),
	.w4(32'hbb368703),
	.w5(32'hbbb7cac6),
	.w6(32'hbc7f69eb),
	.w7(32'hbd0c8f05),
	.w8(32'hb91714ac),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a524c6b),
	.w1(32'h3a6e3d70),
	.w2(32'h3add0116),
	.w3(32'hbc4ddcaa),
	.w4(32'hb9f6cbcc),
	.w5(32'h3b7649c0),
	.w6(32'h3c30986d),
	.w7(32'h3a9c9d96),
	.w8(32'h3c31008c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e7ae0),
	.w1(32'hbb22ce96),
	.w2(32'hbc28d269),
	.w3(32'h3b699e0f),
	.w4(32'h3c91d1c2),
	.w5(32'hbc2c432d),
	.w6(32'hbc39c788),
	.w7(32'hbc02ab1e),
	.w8(32'h3acbbde4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9f6be),
	.w1(32'h3af6d2f5),
	.w2(32'h3c5cf091),
	.w3(32'h3ba55737),
	.w4(32'hbc3c86f8),
	.w5(32'hbb75f720),
	.w6(32'hbb98d2f6),
	.w7(32'h3c812964),
	.w8(32'h3c8a8cd6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d3791),
	.w1(32'h3a5af3f3),
	.w2(32'h3be7f6be),
	.w3(32'hbc012b6f),
	.w4(32'h38b75119),
	.w5(32'h3ac4340c),
	.w6(32'h3a41c8d7),
	.w7(32'h3c0c37f3),
	.w8(32'h3c8c5db7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe8729),
	.w1(32'h3c44e272),
	.w2(32'hba0b1e50),
	.w3(32'h3b123f8d),
	.w4(32'hbaeff865),
	.w5(32'h3ba2c03c),
	.w6(32'hbc383cc0),
	.w7(32'h3b2b434c),
	.w8(32'h3c0e25a3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce013f),
	.w1(32'hbb1e2fb8),
	.w2(32'hbb071af4),
	.w3(32'hbc432293),
	.w4(32'h3c102b78),
	.w5(32'hba978e41),
	.w6(32'hbac48d10),
	.w7(32'hbd076cc6),
	.w8(32'hbc1f28e5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2bb335),
	.w1(32'h3bb37c09),
	.w2(32'hbc89391c),
	.w3(32'hbb96b890),
	.w4(32'h392aa385),
	.w5(32'hbc32ac03),
	.w6(32'h3c299326),
	.w7(32'hbacd5e1c),
	.w8(32'h3ce356c9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae910e8),
	.w1(32'h3c135c12),
	.w2(32'hbbd63220),
	.w3(32'hbbba1dd5),
	.w4(32'hbcaaf506),
	.w5(32'hbc970aad),
	.w6(32'h3c328635),
	.w7(32'hbbf2d2bc),
	.w8(32'hbbd3c1eb),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a8b5c),
	.w1(32'h3a3e6691),
	.w2(32'hbb1712bf),
	.w3(32'h3b0d4e95),
	.w4(32'hbc2d77f8),
	.w5(32'hbc101aca),
	.w6(32'h3ac6f1c0),
	.w7(32'hbca13102),
	.w8(32'hbc8fd730),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59b3b),
	.w1(32'hbb4cb87e),
	.w2(32'h3bcb44aa),
	.w3(32'hbca0d7af),
	.w4(32'h3cb22d2f),
	.w5(32'hbbc5d35e),
	.w6(32'h3ad37e1e),
	.w7(32'hbc465f52),
	.w8(32'h3b141abf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6da61e),
	.w1(32'hbb81b12f),
	.w2(32'hbb3ef5f1),
	.w3(32'hbccbea33),
	.w4(32'h3c99ea97),
	.w5(32'h3abb123c),
	.w6(32'hbc596938),
	.w7(32'hbb2990e6),
	.w8(32'h3c440beb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b8022),
	.w1(32'hbbf2acb6),
	.w2(32'hbbb331f0),
	.w3(32'h3bbf9dba),
	.w4(32'hbb5d13f4),
	.w5(32'h3c2798f8),
	.w6(32'h3ba5da8e),
	.w7(32'hbadcef28),
	.w8(32'hbc6a130c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207403),
	.w1(32'h3b78df67),
	.w2(32'h3ca674c6),
	.w3(32'hbba4ee50),
	.w4(32'h3b80cac4),
	.w5(32'hbb36967f),
	.w6(32'hbcbbc692),
	.w7(32'h3b7abb84),
	.w8(32'hb91761d0),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d30f8),
	.w1(32'h3b525779),
	.w2(32'hbd27c0ec),
	.w3(32'h3c17df80),
	.w4(32'h3c588f7c),
	.w5(32'hbc2f5dcb),
	.w6(32'hbc033a7f),
	.w7(32'h3b950378),
	.w8(32'hbaf4a5e0),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf6d27),
	.w1(32'hbb63425f),
	.w2(32'h3c503c61),
	.w3(32'hbcdc3816),
	.w4(32'hbbf3fd80),
	.w5(32'hba26e1ad),
	.w6(32'hbc0f4dca),
	.w7(32'h3b217ac6),
	.w8(32'h3c9af130),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c403b4a),
	.w1(32'hb95fc2dc),
	.w2(32'h3ad68cc0),
	.w3(32'h3c2fe2eb),
	.w4(32'hbb914907),
	.w5(32'hbb516f13),
	.w6(32'h3cdaaba5),
	.w7(32'hba45c693),
	.w8(32'h3a008710),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba892b9f),
	.w1(32'h3b807d87),
	.w2(32'h3b70a811),
	.w3(32'h3b94c953),
	.w4(32'h3b4f0ac5),
	.w5(32'hbb8db9f6),
	.w6(32'h3b8353b3),
	.w7(32'h3b1cfb14),
	.w8(32'h3ca8bfa1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd91e6a),
	.w1(32'h3c64e032),
	.w2(32'h3be101b0),
	.w3(32'hbb9a0d17),
	.w4(32'h3b0b26b9),
	.w5(32'h3c01af83),
	.w6(32'hba5a293f),
	.w7(32'h3b0a83aa),
	.w8(32'hbcfbc21e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a641611),
	.w1(32'hbb002482),
	.w2(32'h3b91e54c),
	.w3(32'h3c0a5aa7),
	.w4(32'h3b0791d1),
	.w5(32'hbafd8a96),
	.w6(32'h3c5e2db4),
	.w7(32'h3b918dac),
	.w8(32'h3b21ef3a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93f2b6),
	.w1(32'hbc0cd20f),
	.w2(32'h3c0facc0),
	.w3(32'h3b08b1e7),
	.w4(32'hb9925322),
	.w5(32'h3c572a36),
	.w6(32'h3bec9c13),
	.w7(32'h3be3851d),
	.w8(32'h3c217ac4),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc68eb),
	.w1(32'hba82ffd8),
	.w2(32'h3b3514dc),
	.w3(32'h3c02af82),
	.w4(32'h3b66299d),
	.w5(32'h3c39e830),
	.w6(32'h3c28e41e),
	.w7(32'h3c31c17e),
	.w8(32'h395efca9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd082c6a),
	.w1(32'h3ad031be),
	.w2(32'h3ace8325),
	.w3(32'h3c925281),
	.w4(32'h3c0932d1),
	.w5(32'hbb30061c),
	.w6(32'hb9beba19),
	.w7(32'hbbdb376d),
	.w8(32'hbb371105),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc254280),
	.w1(32'hbabc0aba),
	.w2(32'h3c1b702f),
	.w3(32'hbb06c3d0),
	.w4(32'hba62fc41),
	.w5(32'hbb13f93b),
	.w6(32'h3b1df316),
	.w7(32'h3ca43174),
	.w8(32'h3bfa81da),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42e12f),
	.w1(32'hbbf2e333),
	.w2(32'h3bf3a35f),
	.w3(32'hbaab071f),
	.w4(32'h3c3ef038),
	.w5(32'h3c4f0bba),
	.w6(32'h3b0ec248),
	.w7(32'h3bd2dbaa),
	.w8(32'h3bc0b767),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40f684),
	.w1(32'h3bd288af),
	.w2(32'hbb8f3964),
	.w3(32'hbd0de133),
	.w4(32'hbc154d75),
	.w5(32'hbbfeb3b4),
	.w6(32'h3c53341d),
	.w7(32'hbcb65112),
	.w8(32'hbc337b2e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09194a),
	.w1(32'hb9dcc541),
	.w2(32'h3c2f817f),
	.w3(32'h3b53e391),
	.w4(32'hbb5f646c),
	.w5(32'h3bdd6604),
	.w6(32'hbb25f04b),
	.w7(32'h3a82d89d),
	.w8(32'hba9a1540),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd91f81),
	.w1(32'h3c605c7c),
	.w2(32'hbc6d55c5),
	.w3(32'h3b9e1dd8),
	.w4(32'h3c133b5a),
	.w5(32'h3ace7f69),
	.w6(32'h3b27163d),
	.w7(32'hbbb2c80f),
	.w8(32'hbbd420cc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f4d10),
	.w1(32'hbbb11830),
	.w2(32'h3c1446b2),
	.w3(32'h3c246451),
	.w4(32'h3bb79e45),
	.w5(32'h3c8a1de2),
	.w6(32'h3c830ca1),
	.w7(32'hb9cfd436),
	.w8(32'h3c819bd7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4ecd),
	.w1(32'h3c03c268),
	.w2(32'h3c045e01),
	.w3(32'hbc90d859),
	.w4(32'h3c98d765),
	.w5(32'hbaa809b1),
	.w6(32'hbb80cae4),
	.w7(32'hbb3b791d),
	.w8(32'hbaebc441),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab405d4),
	.w1(32'hbb274fc4),
	.w2(32'h3b2e300e),
	.w3(32'hbbed7aa1),
	.w4(32'h3abe2ba8),
	.w5(32'h3beb83e0),
	.w6(32'h394daa05),
	.w7(32'h3b0c04cf),
	.w8(32'h3c1879dc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801e6c),
	.w1(32'hba841427),
	.w2(32'hbcd00c47),
	.w3(32'h3a0f33b0),
	.w4(32'h3a552677),
	.w5(32'h3a999b76),
	.w6(32'hbc39bb87),
	.w7(32'h3bc81e7c),
	.w8(32'hbc82ffd1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08c9ad),
	.w1(32'h3c1227a7),
	.w2(32'h3c29ba79),
	.w3(32'h3c111aa2),
	.w4(32'h3c0bfcee),
	.w5(32'h3be27226),
	.w6(32'hbc5ca437),
	.w7(32'h3c23629a),
	.w8(32'hbc15a60d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e6b2),
	.w1(32'h3c6475e5),
	.w2(32'hbc4d2c3c),
	.w3(32'hba125175),
	.w4(32'h3c17b1d3),
	.w5(32'hbb6abaee),
	.w6(32'h3c20a0ef),
	.w7(32'h3bc7b41d),
	.w8(32'hbc6048a2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f1015),
	.w1(32'hbb125c8b),
	.w2(32'h3b0ef748),
	.w3(32'hba65e2fd),
	.w4(32'hba9621e4),
	.w5(32'h3ba05a58),
	.w6(32'hbb4feaea),
	.w7(32'hbcfa3526),
	.w8(32'hbb2943e3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8db6f0),
	.w1(32'hbbd65a2d),
	.w2(32'h3983536a),
	.w3(32'h3b438193),
	.w4(32'h3c55e70f),
	.w5(32'hbc1c3484),
	.w6(32'h3c0aba6b),
	.w7(32'h3a237fed),
	.w8(32'h3bcddc00),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d50b7ce),
	.w1(32'h3c30ba8a),
	.w2(32'h3cae1441),
	.w3(32'h3bb9f734),
	.w4(32'h3baef9f8),
	.w5(32'h3b55ba2e),
	.w6(32'h3cfd314d),
	.w7(32'h3c4090f2),
	.w8(32'h3cb573c9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17ccb4),
	.w1(32'h3ad18b27),
	.w2(32'hbab54b17),
	.w3(32'hbbe65727),
	.w4(32'hba1d953d),
	.w5(32'hbbfe9b38),
	.w6(32'hbb8e2b2f),
	.w7(32'hbbbb702a),
	.w8(32'hbc5eeb20),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37763d),
	.w1(32'h3ba409cb),
	.w2(32'hb95f3f6f),
	.w3(32'hbceaec43),
	.w4(32'h3bb1aab3),
	.w5(32'hbb4c0d8a),
	.w6(32'h3bcc09bf),
	.w7(32'hbb1f9664),
	.w8(32'h3bf5486a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beafa24),
	.w1(32'hbd057cab),
	.w2(32'hbc62ea22),
	.w3(32'hbb1d94aa),
	.w4(32'hbbb133d7),
	.w5(32'h3b9d6a8a),
	.w6(32'h3b70bd9b),
	.w7(32'hba8a0b04),
	.w8(32'hbc1d951d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe79f10),
	.w1(32'hbb70423d),
	.w2(32'h3b48b2bf),
	.w3(32'hba183150),
	.w4(32'hbb7f40cc),
	.w5(32'h35cd55df),
	.w6(32'h3af3a751),
	.w7(32'hbb5f497c),
	.w8(32'h3aed6a79),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba615c9),
	.w1(32'hbc5994fc),
	.w2(32'hbbe846ba),
	.w3(32'h3c1117ec),
	.w4(32'h3cc8a31c),
	.w5(32'hbb9d8c43),
	.w6(32'h3bd5ac76),
	.w7(32'hbbabda66),
	.w8(32'hbb741078),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3778),
	.w1(32'h3b0da1da),
	.w2(32'h3b9fc03e),
	.w3(32'h3bd0a6e7),
	.w4(32'h397720b1),
	.w5(32'h3ad36ef3),
	.w6(32'h3be5754b),
	.w7(32'hbb85dcd2),
	.w8(32'h3b920852),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf5d93),
	.w1(32'h3c47db65),
	.w2(32'h3c9b0736),
	.w3(32'h3c4502bb),
	.w4(32'h3b531d10),
	.w5(32'h3c566f6b),
	.w6(32'h3b194710),
	.w7(32'h3ab5e7a3),
	.w8(32'h3ba888da),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf12a02),
	.w1(32'hbb7fc625),
	.w2(32'hbc02b79d),
	.w3(32'h3b58f323),
	.w4(32'hbb82dd8a),
	.w5(32'h3b84a8a9),
	.w6(32'hb992b708),
	.w7(32'h3b83d563),
	.w8(32'h3bada431),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58c020),
	.w1(32'h3b0549b8),
	.w2(32'hbc498abf),
	.w3(32'h3a9edd4f),
	.w4(32'hbb1b6217),
	.w5(32'hbb8c50d4),
	.w6(32'h3c071d0a),
	.w7(32'h3acdd7a6),
	.w8(32'h3b7a20b0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124ff4),
	.w1(32'h3cbf1258),
	.w2(32'hbbc169fc),
	.w3(32'hbb75b610),
	.w4(32'h3b8c3ad7),
	.w5(32'hbb874958),
	.w6(32'h3c717b6d),
	.w7(32'h3b252bf6),
	.w8(32'h3c9e7913),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83dad9),
	.w1(32'hbbc71566),
	.w2(32'h3af6a0af),
	.w3(32'hbc3ccb9f),
	.w4(32'hbc9242dc),
	.w5(32'hbb10da1d),
	.w6(32'h3922201f),
	.w7(32'h3a9bde73),
	.w8(32'hbba51345),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc568103),
	.w1(32'hbbb0c902),
	.w2(32'h3b0e58c6),
	.w3(32'h3b27db5b),
	.w4(32'h3cb88c72),
	.w5(32'h3c776b09),
	.w6(32'h3afe5337),
	.w7(32'hbb15b297),
	.w8(32'h3bd5ac31),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7a74a),
	.w1(32'h38cf7a10),
	.w2(32'hbcc535aa),
	.w3(32'h3d014b21),
	.w4(32'h3a99724b),
	.w5(32'h3c79c639),
	.w6(32'hbbab60b6),
	.w7(32'hbb834f4c),
	.w8(32'hbb012f9c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84c7d),
	.w1(32'h3c8c2a36),
	.w2(32'hbbe6f253),
	.w3(32'hbb3f6863),
	.w4(32'hbb8f6665),
	.w5(32'hbab272b6),
	.w6(32'h3bccfac0),
	.w7(32'h3bc08b7c),
	.w8(32'h3b44d8ed),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3990e9),
	.w1(32'hbd01458d),
	.w2(32'h3cbd9a7c),
	.w3(32'h3aa813df),
	.w4(32'h3bbe080e),
	.w5(32'hbb48e8ce),
	.w6(32'hbc5c94c3),
	.w7(32'h3be161a6),
	.w8(32'h3be566c2),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099234),
	.w1(32'h3c706d20),
	.w2(32'hba2b57c8),
	.w3(32'h3bb0fc05),
	.w4(32'hbc49777c),
	.w5(32'h38e498d2),
	.w6(32'h3cc69753),
	.w7(32'h3b51287b),
	.w8(32'h3c614fc5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bd1f7),
	.w1(32'hbb8290e4),
	.w2(32'hbc81f461),
	.w3(32'h3b33432d),
	.w4(32'hb945d3b5),
	.w5(32'h3d01124b),
	.w6(32'h3c13e9d1),
	.w7(32'hbc0c3a74),
	.w8(32'h3acbec8e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09371b),
	.w1(32'hbbec5dfb),
	.w2(32'h3cabc962),
	.w3(32'hbc51a0a8),
	.w4(32'hbc21bbf8),
	.w5(32'h3bef8483),
	.w6(32'h3c163628),
	.w7(32'h3bb7aced),
	.w8(32'h3bfc08ed),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30fc61),
	.w1(32'hbbaebfa0),
	.w2(32'h3c09e96e),
	.w3(32'hbaa4d212),
	.w4(32'hbc55248c),
	.w5(32'h3b413e66),
	.w6(32'hbc87f47f),
	.w7(32'h3c0f865e),
	.w8(32'h3c227625),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63b069),
	.w1(32'h3c8fc4e6),
	.w2(32'h3a54fad9),
	.w3(32'h39f2ea05),
	.w4(32'h3a7b4f5e),
	.w5(32'h3b8f48e4),
	.w6(32'hbcb2a02a),
	.w7(32'h3baa47c0),
	.w8(32'h3a896716),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b209678),
	.w1(32'hbc0df24a),
	.w2(32'hba8d8500),
	.w3(32'h3b794d91),
	.w4(32'h3c1bc19d),
	.w5(32'h3b98fb1f),
	.w6(32'hbaedf545),
	.w7(32'hbb2b09b4),
	.w8(32'hbbaecd48),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8dc61),
	.w1(32'h3c0bf1f7),
	.w2(32'hb991a17f),
	.w3(32'h3b6807ab),
	.w4(32'h3a4502e3),
	.w5(32'h3bba4add),
	.w6(32'hbc569fd7),
	.w7(32'hbbe4ebbd),
	.w8(32'hbb35428d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc327603),
	.w1(32'hbc495148),
	.w2(32'h3bca4e82),
	.w3(32'hbb1b2945),
	.w4(32'hbbaa0393),
	.w5(32'h3c438b47),
	.w6(32'hbbb0f727),
	.w7(32'hbbc94020),
	.w8(32'hbd129ec3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72daf1),
	.w1(32'hbc8cc689),
	.w2(32'h3c6374a6),
	.w3(32'hbb907d5c),
	.w4(32'h3b16b1f6),
	.w5(32'h3c9c7fb7),
	.w6(32'h3bfadefc),
	.w7(32'hbb4ac9ae),
	.w8(32'h3ba5d136),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7237c8),
	.w1(32'hbc9cf688),
	.w2(32'h3c84d25c),
	.w3(32'h3c8d5f46),
	.w4(32'h3bb6376a),
	.w5(32'h3c37f7c6),
	.w6(32'hbaf7c326),
	.w7(32'h3b624364),
	.w8(32'h3c33c6be),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4983f5),
	.w1(32'h3d1ad1b0),
	.w2(32'hbb5ae81d),
	.w3(32'h39ae7041),
	.w4(32'h3bff60dc),
	.w5(32'hbb5ca2c9),
	.w6(32'h3c9eba07),
	.w7(32'h3b142247),
	.w8(32'hbaa8e7cd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f750a),
	.w1(32'h3a9a8cfd),
	.w2(32'h3b29dcd8),
	.w3(32'h3b5a4890),
	.w4(32'h3bebc604),
	.w5(32'hba9516be),
	.w6(32'hbcb1d129),
	.w7(32'hb7d48de6),
	.w8(32'hbb6608f3),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06368c),
	.w1(32'hbc1e97ac),
	.w2(32'h3b9daf17),
	.w3(32'h398d47e8),
	.w4(32'h3c2c71a7),
	.w5(32'h3accb945),
	.w6(32'hbd093403),
	.w7(32'h3b9d27bc),
	.w8(32'h3c4648be),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce6ac),
	.w1(32'hbc066b7c),
	.w2(32'hbd3d0a11),
	.w3(32'h3a18b677),
	.w4(32'hbc021fb4),
	.w5(32'hbd330bea),
	.w6(32'h3c77d71b),
	.w7(32'hbb7349da),
	.w8(32'hbd66a877),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6e98),
	.w1(32'hbb143150),
	.w2(32'h3a8cefbd),
	.w3(32'h3b868736),
	.w4(32'hbcad8e7b),
	.w5(32'hbcb2b149),
	.w6(32'h3c865c49),
	.w7(32'h3b3bec92),
	.w8(32'h3b23a75a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c339d77),
	.w1(32'h3c2facef),
	.w2(32'h3ba87aa9),
	.w3(32'h3cedac4c),
	.w4(32'hbb5f6e57),
	.w5(32'h3b65fe00),
	.w6(32'hbb3d0e0c),
	.w7(32'hbb97269c),
	.w8(32'hbba76f96),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434f19),
	.w1(32'h3b8ef3e3),
	.w2(32'h3bf3a8fc),
	.w3(32'hbcd19a67),
	.w4(32'h3cb6fbb6),
	.w5(32'h3aa96c9a),
	.w6(32'hbbd0c0d6),
	.w7(32'h3a364175),
	.w8(32'hbbf8e8bd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c962e0b),
	.w1(32'hb950368d),
	.w2(32'h3b58f870),
	.w3(32'h3ce651e8),
	.w4(32'hb9070589),
	.w5(32'h3b69287e),
	.w6(32'h3a815f77),
	.w7(32'h3c220284),
	.w8(32'h3d03ab45),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dfd34),
	.w1(32'h3babe85f),
	.w2(32'h3c88d3a8),
	.w3(32'h3cacfe2e),
	.w4(32'h3b18ad1f),
	.w5(32'h3c5b9816),
	.w6(32'hbc4eda4a),
	.w7(32'hbbe59436),
	.w8(32'h3ab4499d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bd094),
	.w1(32'h3c21377f),
	.w2(32'hbc6b1031),
	.w3(32'h3c6d2af9),
	.w4(32'h3b13b6f6),
	.w5(32'hbafcdb77),
	.w6(32'hb9e2454b),
	.w7(32'h3b427e56),
	.w8(32'hbc4d8e15),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf856b4),
	.w1(32'h3a13fe53),
	.w2(32'h3b9a8c4e),
	.w3(32'h3a9353e4),
	.w4(32'hbbca4cbd),
	.w5(32'hbc1fa802),
	.w6(32'h3bf8742d),
	.w7(32'h3c103a35),
	.w8(32'hbc190e1e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca52125),
	.w1(32'h3c0c90e0),
	.w2(32'hbc663818),
	.w3(32'hbc01ccf6),
	.w4(32'h3bcad685),
	.w5(32'hbc1b5cfb),
	.w6(32'h3c45bdd4),
	.w7(32'h3c6b1850),
	.w8(32'hbb8399fd),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3c24f),
	.w1(32'hba2b0e49),
	.w2(32'h3c9a0c31),
	.w3(32'hbb94311e),
	.w4(32'hbc5ec49e),
	.w5(32'h3be0e025),
	.w6(32'h3bb91591),
	.w7(32'hbbe547a5),
	.w8(32'h3c8d42aa),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4498),
	.w1(32'hbb3bb3dd),
	.w2(32'hbb677c95),
	.w3(32'h3c488b8b),
	.w4(32'hbac45416),
	.w5(32'hbbc7c625),
	.w6(32'h3b3128ea),
	.w7(32'h3b66556d),
	.w8(32'h3c168625),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadf542),
	.w1(32'h3c8c97da),
	.w2(32'hba0084c2),
	.w3(32'h3ae6e151),
	.w4(32'h3bc5938c),
	.w5(32'h3bd21305),
	.w6(32'hb986b17f),
	.w7(32'h3c22ba44),
	.w8(32'hba1a12c9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02ea9c),
	.w1(32'hbb079f7b),
	.w2(32'h3b9644ba),
	.w3(32'hba910aaa),
	.w4(32'h3aab35d7),
	.w5(32'hbc912f7b),
	.w6(32'hbc25ff3e),
	.w7(32'h3bc72f08),
	.w8(32'h3bc5e33a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43566),
	.w1(32'h3bbda85e),
	.w2(32'hbc9d7fe6),
	.w3(32'h3c2570ea),
	.w4(32'hba233693),
	.w5(32'hbbb51351),
	.w6(32'h3c9ccfee),
	.w7(32'hba2f2c81),
	.w8(32'hbd4cf7cd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e0f31),
	.w1(32'hbb0125bb),
	.w2(32'hbccc2a91),
	.w3(32'h3c3504e2),
	.w4(32'h3c92268c),
	.w5(32'h3b10a743),
	.w6(32'hbc2b2f4d),
	.w7(32'hbbd856fd),
	.w8(32'hbc1f66e8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1d1e),
	.w1(32'hbb029c59),
	.w2(32'hbb248f98),
	.w3(32'hbb81c2f0),
	.w4(32'hbc357acc),
	.w5(32'hbbe8abfe),
	.w6(32'hbbfbdfd0),
	.w7(32'hbc05fe51),
	.w8(32'hbcd5a56c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985159),
	.w1(32'h3aa6ac90),
	.w2(32'h3b0ca14b),
	.w3(32'h3b6619fa),
	.w4(32'hbbfff1db),
	.w5(32'h3c10393b),
	.w6(32'h3bee317a),
	.w7(32'hbb2d3017),
	.w8(32'hbc0ae9cd),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2ade),
	.w1(32'h3bf52907),
	.w2(32'hbb613b95),
	.w3(32'h3b770ce7),
	.w4(32'h3c072ef3),
	.w5(32'h3b3f206c),
	.w6(32'hbb2dd076),
	.w7(32'h3c42aa8c),
	.w8(32'h3ad8fd65),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf651d9),
	.w1(32'h3bc6a0e1),
	.w2(32'h3ba9b4fa),
	.w3(32'h3b85c9b6),
	.w4(32'hbc03adac),
	.w5(32'hbc1a16e3),
	.w6(32'h3b35fdad),
	.w7(32'h3bcffa86),
	.w8(32'hbc63d1f7),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccb6e1),
	.w1(32'h371bb391),
	.w2(32'h3be1ddef),
	.w3(32'hb7956284),
	.w4(32'h3ae427e4),
	.w5(32'hbd09d1c6),
	.w6(32'hbd1100df),
	.w7(32'h3b8b58ae),
	.w8(32'h3b68e3a0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3101f2),
	.w1(32'hbc696837),
	.w2(32'h3a3e5a53),
	.w3(32'h3bb3a06f),
	.w4(32'h3bb41e33),
	.w5(32'h3bbb44a2),
	.w6(32'h3befbcd7),
	.w7(32'h3a33415a),
	.w8(32'h3b0b0f90),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e992d),
	.w1(32'h3c139965),
	.w2(32'h3c199e30),
	.w3(32'h3b250d5c),
	.w4(32'h3a09a990),
	.w5(32'hbb93aa79),
	.w6(32'h3a80eed4),
	.w7(32'h3b522323),
	.w8(32'h3c422663),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc4e32),
	.w1(32'hbb9568a8),
	.w2(32'h3bbb4cce),
	.w3(32'h3bda14c4),
	.w4(32'h3a325105),
	.w5(32'hba644304),
	.w6(32'hbbba1081),
	.w7(32'hbcab3c00),
	.w8(32'h3b3229e1),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344ba9),
	.w1(32'h3a1d4b3c),
	.w2(32'hbc1fb9e8),
	.w3(32'h3bb7c074),
	.w4(32'hbb6ce688),
	.w5(32'h392dba4b),
	.w6(32'h3ab5da5d),
	.w7(32'hbccd0804),
	.w8(32'hbbcf18fc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43b99),
	.w1(32'hbcb46cdc),
	.w2(32'hbc06d9c2),
	.w3(32'h3b9d6e72),
	.w4(32'h3af7baee),
	.w5(32'h3be380f4),
	.w6(32'h3a7ef156),
	.w7(32'hbcd99961),
	.w8(32'h3b0eec2e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24b10e),
	.w1(32'hba443edf),
	.w2(32'h3c0718f5),
	.w3(32'hbb507ea3),
	.w4(32'hbacac9f6),
	.w5(32'h3c403167),
	.w6(32'hbb708ce7),
	.w7(32'h3bb868fb),
	.w8(32'h3ba6f88f),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82cf34),
	.w1(32'h3c6893fe),
	.w2(32'hbbff9a9a),
	.w3(32'hbbe584ea),
	.w4(32'hbcdc073b),
	.w5(32'h3bfa5e21),
	.w6(32'h3c42c5e2),
	.w7(32'h3c991d13),
	.w8(32'h3c525140),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a91c5a),
	.w1(32'h3a0b2b8d),
	.w2(32'h3b89bd13),
	.w3(32'h3b01dc2b),
	.w4(32'hbbc3d735),
	.w5(32'h3be0daa2),
	.w6(32'h3b5ef753),
	.w7(32'h3c3ef227),
	.w8(32'h3b63590e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2549c4),
	.w1(32'hb96c8f7f),
	.w2(32'h3b087692),
	.w3(32'h3ac5b854),
	.w4(32'hbae5a61c),
	.w5(32'h3c21e79d),
	.w6(32'h3c13c44a),
	.w7(32'h3ba8eb4c),
	.w8(32'h3bb6e289),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b7245),
	.w1(32'h3c3c8ad7),
	.w2(32'h3a69c17d),
	.w3(32'hbc5b8208),
	.w4(32'h3b9e8459),
	.w5(32'h3cafbba7),
	.w6(32'h3bebd679),
	.w7(32'h3cc51e83),
	.w8(32'h3c1f6d61),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadcf51),
	.w1(32'h3b922966),
	.w2(32'h399bfce1),
	.w3(32'h3bfd4df3),
	.w4(32'hbb94a808),
	.w5(32'hbb99c745),
	.w6(32'h38c06620),
	.w7(32'hbbb999b7),
	.w8(32'h3b5f9029),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcee15c),
	.w1(32'h3c6ecb62),
	.w2(32'hbb2734a2),
	.w3(32'hba8a2b29),
	.w4(32'h3aedc6ba),
	.w5(32'hbcda8254),
	.w6(32'hbb869cda),
	.w7(32'hbc9f2369),
	.w8(32'h3b3b35a0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61aff7),
	.w1(32'h3bb30351),
	.w2(32'h3b0ee699),
	.w3(32'h3ad1d6b9),
	.w4(32'h3c481168),
	.w5(32'h3b99410f),
	.w6(32'h3bf14233),
	.w7(32'h3bbb6ca4),
	.w8(32'h3aa60e2c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d8665),
	.w1(32'h3ce3d0c8),
	.w2(32'h3ba51451),
	.w3(32'h3b12f458),
	.w4(32'hbcc100fd),
	.w5(32'h3bf846a8),
	.w6(32'hbab01e0e),
	.w7(32'hbc06302e),
	.w8(32'h39867b81),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c896688),
	.w1(32'h3b8d4c6f),
	.w2(32'h3b7e29b7),
	.w3(32'hbc9a46c9),
	.w4(32'h3c385e5b),
	.w5(32'hbc7c7f77),
	.w6(32'hbb7d106b),
	.w7(32'h3baa7b80),
	.w8(32'hbcb120e2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951a3e),
	.w1(32'h3b39ec32),
	.w2(32'h3b3bfd4c),
	.w3(32'hbc38d0ac),
	.w4(32'hbc0bd3fc),
	.w5(32'h3a8f85e9),
	.w6(32'h3a2b253d),
	.w7(32'hbbafc6e7),
	.w8(32'h3c23deba),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadd460),
	.w1(32'hbcbb0f40),
	.w2(32'h3c974037),
	.w3(32'h3cbaa704),
	.w4(32'h3c23ccba),
	.w5(32'h3cd4c19d),
	.w6(32'h3c882613),
	.w7(32'h3d0403ca),
	.w8(32'h3c8b73d3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bece9af),
	.w1(32'hb9207775),
	.w2(32'hbbf73a69),
	.w3(32'hba8f57ae),
	.w4(32'hbb0722e2),
	.w5(32'hbc0a5627),
	.w6(32'h3b6637e0),
	.w7(32'hbc44b983),
	.w8(32'h3c1d7edb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53dbdf),
	.w1(32'hb909cabc),
	.w2(32'h3bb6e3a1),
	.w3(32'h3ca76d57),
	.w4(32'h3c00052e),
	.w5(32'hbba25373),
	.w6(32'hbb7f5095),
	.w7(32'hbbfa556b),
	.w8(32'hbb69e880),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule