module layer_10_featuremap_332(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa76825),
	.w1(32'h3b236fe0),
	.w2(32'hba9f0e51),
	.w3(32'h3c0cdf7b),
	.w4(32'h3a950ff3),
	.w5(32'hbbb00681),
	.w6(32'h3bc7136f),
	.w7(32'hbbc847b0),
	.w8(32'hbb3278a1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3881f0),
	.w1(32'hbc3f28cd),
	.w2(32'hbc050654),
	.w3(32'hbc79e16d),
	.w4(32'hbc55d98a),
	.w5(32'hbab020cc),
	.w6(32'hbba7c9cf),
	.w7(32'hbb9fb657),
	.w8(32'hbaf4a4e0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc284777),
	.w1(32'hbb6ea457),
	.w2(32'hba86f7e5),
	.w3(32'h3b9dd155),
	.w4(32'h3bdd4e12),
	.w5(32'hbb1cb19b),
	.w6(32'h3b3b8bd4),
	.w7(32'h3ba8b818),
	.w8(32'hbb164584),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59b11d),
	.w1(32'hbc2e8ba3),
	.w2(32'hbc0d3987),
	.w3(32'hbb7fd1bd),
	.w4(32'hbb788d3e),
	.w5(32'hbb4c1d3c),
	.w6(32'hbba36ec3),
	.w7(32'hbb6b250b),
	.w8(32'hbb642e4b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3223a),
	.w1(32'hba35f328),
	.w2(32'hbb54eb44),
	.w3(32'h3b36fff6),
	.w4(32'h3b67442b),
	.w5(32'h3b53228c),
	.w6(32'h3b2f4df8),
	.w7(32'h3b8cda5a),
	.w8(32'hbb0e206e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d7941),
	.w1(32'h3b582a0c),
	.w2(32'h3b0c7c47),
	.w3(32'h3ac1066b),
	.w4(32'h3ad91629),
	.w5(32'hbb87568f),
	.w6(32'h3a0d36e9),
	.w7(32'h3a4a1e83),
	.w8(32'hbb2a2d16),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86c3b0),
	.w1(32'hbc90bfd8),
	.w2(32'hbc8b47bc),
	.w3(32'hbc4b00e9),
	.w4(32'hbc34d74c),
	.w5(32'h3b8afaa0),
	.w6(32'hbc51fe4f),
	.w7(32'hbbd2fe6a),
	.w8(32'h3b009809),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07e522),
	.w1(32'h3c7d1cba),
	.w2(32'h3cd2c417),
	.w3(32'h3c926586),
	.w4(32'h3cb02a19),
	.w5(32'h3c420b4a),
	.w6(32'h3c9a9719),
	.w7(32'h3900069d),
	.w8(32'hbbd5fa69),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7204b0),
	.w1(32'h3b728265),
	.w2(32'h3b2ac201),
	.w3(32'h39d66554),
	.w4(32'hb8af55cd),
	.w5(32'h3bceae33),
	.w6(32'hbb3ef65d),
	.w7(32'hbb4dcaae),
	.w8(32'h3b0a4971),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf8116),
	.w1(32'h3beaee9b),
	.w2(32'h3bd25934),
	.w3(32'h3b733235),
	.w4(32'h3b4ed35f),
	.w5(32'h3ba31e42),
	.w6(32'hba78d30f),
	.w7(32'hba8d043e),
	.w8(32'hba9c380c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c2f3),
	.w1(32'hbb1c6c12),
	.w2(32'h3a231a18),
	.w3(32'hbbac8348),
	.w4(32'hba84da41),
	.w5(32'h3b0861d0),
	.w6(32'hbbbcced0),
	.w7(32'h387ca317),
	.w8(32'h3b6012c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38e051),
	.w1(32'hbc5e6068),
	.w2(32'hbc007f25),
	.w3(32'h3b9d88ee),
	.w4(32'hbb8109d0),
	.w5(32'hbb34eabc),
	.w6(32'hbbee0fad),
	.w7(32'h3b608493),
	.w8(32'hbb1dbaf6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71bb99),
	.w1(32'h3c86332d),
	.w2(32'h3c06c552),
	.w3(32'h3c4ed982),
	.w4(32'h3b8119f3),
	.w5(32'h3b294d80),
	.w6(32'h3c165a59),
	.w7(32'hbb1b5c58),
	.w8(32'h398796f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc63f),
	.w1(32'h3bdc860d),
	.w2(32'h3c040f9e),
	.w3(32'h3b0fc05d),
	.w4(32'h3b3f6e23),
	.w5(32'h39eacab4),
	.w6(32'h3b857a74),
	.w7(32'h3ae4ae60),
	.w8(32'hba723739),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038f3b),
	.w1(32'hbbd73f21),
	.w2(32'hbbbc6059),
	.w3(32'hbc42b8af),
	.w4(32'hbc210789),
	.w5(32'hbb5d0004),
	.w6(32'hbb3decbe),
	.w7(32'hbba6724f),
	.w8(32'h36d274d1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36463c),
	.w1(32'h3b9988f2),
	.w2(32'h3b24a541),
	.w3(32'h38056f0e),
	.w4(32'hba879e1d),
	.w5(32'h3b352a0c),
	.w6(32'hbae5f5b5),
	.w7(32'h3abd7913),
	.w8(32'h3adef642),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46b21d),
	.w1(32'h3b16bb73),
	.w2(32'h395100c7),
	.w3(32'h3b953c2e),
	.w4(32'hba88ac68),
	.w5(32'h39aa95d5),
	.w6(32'h3c19acec),
	.w7(32'h3b214401),
	.w8(32'hbb0e4037),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84bf96),
	.w1(32'h3bfec700),
	.w2(32'h3be51f3b),
	.w3(32'hbb5fe3df),
	.w4(32'h3b50e3e6),
	.w5(32'h3bc44d47),
	.w6(32'hbc054d80),
	.w7(32'hbbeca1fe),
	.w8(32'hba34285f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9308d),
	.w1(32'hba965371),
	.w2(32'hb931bda1),
	.w3(32'hbab024d7),
	.w4(32'h3b693306),
	.w5(32'h3b183238),
	.w6(32'hbbc36e80),
	.w7(32'hbbab3ef8),
	.w8(32'h3ab90b29),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61079c),
	.w1(32'h3b906101),
	.w2(32'hbb438cce),
	.w3(32'hbb208c7f),
	.w4(32'hbb8fface),
	.w5(32'h3ba78c41),
	.w6(32'hb91f70a4),
	.w7(32'hbbaf9e50),
	.w8(32'h3bea2352),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60033c),
	.w1(32'hbadbe186),
	.w2(32'hbbb1d1c4),
	.w3(32'h3b0d3ec6),
	.w4(32'hb9bf98d7),
	.w5(32'h3bd6a026),
	.w6(32'h3a1cbe2a),
	.w7(32'hbba4c15d),
	.w8(32'h3bcc2460),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba11581),
	.w1(32'hbacb3a45),
	.w2(32'hbba4c743),
	.w3(32'h3ae0f837),
	.w4(32'hba4b3d1f),
	.w5(32'hb926b817),
	.w6(32'h3a9c33cb),
	.w7(32'hbb0aad91),
	.w8(32'hba50683a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b876277),
	.w1(32'h3bb41cf0),
	.w2(32'h3b37a70f),
	.w3(32'hbaac9958),
	.w4(32'hbc742205),
	.w5(32'hbb27ca1f),
	.w6(32'hbbbaa8ca),
	.w7(32'hbc2821f2),
	.w8(32'hbc853170),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7343cb),
	.w1(32'h3a37cf9c),
	.w2(32'h3bb30d1e),
	.w3(32'hbb9731fa),
	.w4(32'hbbc5a82c),
	.w5(32'hbb905760),
	.w6(32'hbbdf1a8a),
	.w7(32'hbbd396dc),
	.w8(32'hbc0ae141),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21a792),
	.w1(32'hbc6565b1),
	.w2(32'hbc17703b),
	.w3(32'hbc1f0a26),
	.w4(32'hbbdc9395),
	.w5(32'hbc1a767c),
	.w6(32'hbbe6890b),
	.w7(32'hbb9b03f3),
	.w8(32'hbc08b34a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a065dd8),
	.w1(32'h3b7f001e),
	.w2(32'h3a895c77),
	.w3(32'h394dbfdf),
	.w4(32'hb987691e),
	.w5(32'hbb92c7ff),
	.w6(32'h3c0d1244),
	.w7(32'h3b9c906d),
	.w8(32'hbb8b12a4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2de012),
	.w1(32'h39f3cee1),
	.w2(32'hb803cabe),
	.w3(32'hbabb334c),
	.w4(32'hba0f35a7),
	.w5(32'h3bb20376),
	.w6(32'h3b4cdb1b),
	.w7(32'hb88ea9cf),
	.w8(32'h3ba997de),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980d87a),
	.w1(32'h3c9b3988),
	.w2(32'hbc709080),
	.w3(32'h3c015cce),
	.w4(32'h3c8771bb),
	.w5(32'hbbf6ffa1),
	.w6(32'h3c7a42ca),
	.w7(32'h3c52ea07),
	.w8(32'hbb5b5fe1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0aa9),
	.w1(32'hbbe71f29),
	.w2(32'hbc0b6a99),
	.w3(32'hbb18f86c),
	.w4(32'hbb8d769a),
	.w5(32'h3a946bd5),
	.w6(32'hbb3cd62e),
	.w7(32'hbb94ce7d),
	.w8(32'h3bcbd1d1),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb7be3),
	.w1(32'hbc31bacd),
	.w2(32'hbc560dd0),
	.w3(32'hbc3753e8),
	.w4(32'h3a688732),
	.w5(32'hbc205f45),
	.w6(32'h397d5ad9),
	.w7(32'hbad55e37),
	.w8(32'hbc048d76),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd26af4),
	.w1(32'h3be70612),
	.w2(32'h3ab2e88a),
	.w3(32'h3ace0f3a),
	.w4(32'hb92f36ee),
	.w5(32'h3b47177e),
	.w6(32'h3a5e5757),
	.w7(32'h3b7a7267),
	.w8(32'hb9ade4dd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8409f5),
	.w1(32'hbb0d9576),
	.w2(32'hbac2ded9),
	.w3(32'h3c45d932),
	.w4(32'h3bed542b),
	.w5(32'hbb3d2c28),
	.w6(32'h3a4c306c),
	.w7(32'h3a97412e),
	.w8(32'hbaefe4c5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8825ea),
	.w1(32'h394b4b4f),
	.w2(32'h3973aa4a),
	.w3(32'h3b17e6dd),
	.w4(32'hbb75a9ea),
	.w5(32'h3ab54ea1),
	.w6(32'h3a1ee5b7),
	.w7(32'hbbf59e2d),
	.w8(32'hbbc7985c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb876f05),
	.w1(32'hbb6f1889),
	.w2(32'hbb71b00a),
	.w3(32'hbaf9a3d1),
	.w4(32'hbbc87ab0),
	.w5(32'hbb4c386e),
	.w6(32'hbb37c29d),
	.w7(32'hbb2eb05b),
	.w8(32'hbb9e6448),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5a1e),
	.w1(32'hbb345afe),
	.w2(32'hbba1e79b),
	.w3(32'hbb31d32b),
	.w4(32'hbac5135f),
	.w5(32'hbb1f4a5c),
	.w6(32'hbbb44e3f),
	.w7(32'hbbb13171),
	.w8(32'hbba2b40d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8c277),
	.w1(32'hbbfbcba5),
	.w2(32'hbb21e327),
	.w3(32'h3af9a471),
	.w4(32'hbb9f0222),
	.w5(32'hb7722592),
	.w6(32'hbb57f3b2),
	.w7(32'hbc04ca63),
	.w8(32'hbbe2fc7d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dbb8c),
	.w1(32'hbc92273e),
	.w2(32'h3c9ed29a),
	.w3(32'h3c61c6e3),
	.w4(32'hbcff21b9),
	.w5(32'hbcc40ae6),
	.w6(32'h3b388502),
	.w7(32'hbcef6536),
	.w8(32'hbc90eceb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6eaa3d),
	.w1(32'hbc874b52),
	.w2(32'hbc7e747b),
	.w3(32'hbc247168),
	.w4(32'hbbf80ed7),
	.w5(32'hbcd6487d),
	.w6(32'hbb1c27e6),
	.w7(32'hbc4adb22),
	.w8(32'hbc82eb2d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77e595),
	.w1(32'hbc52649a),
	.w2(32'hbcd3f56f),
	.w3(32'hbbbb3b5d),
	.w4(32'h3b4cea4c),
	.w5(32'hbc15a804),
	.w6(32'h3b1f972c),
	.w7(32'h3c47573b),
	.w8(32'h3bc5b5b3),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade09b1),
	.w1(32'hbc1f4454),
	.w2(32'hbbfeb1b8),
	.w3(32'hbbce849c),
	.w4(32'hbb8c6f3d),
	.w5(32'hbb7cdef7),
	.w6(32'hbc2eab36),
	.w7(32'hbc1bb9a9),
	.w8(32'hbb68064f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba885c89),
	.w1(32'h3bd2729d),
	.w2(32'h3b035d64),
	.w3(32'h3b15b9b5),
	.w4(32'hb93c959b),
	.w5(32'h3b6921b2),
	.w6(32'h3b585ebc),
	.w7(32'hba0f1c14),
	.w8(32'h3bcb548e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6689e),
	.w1(32'h3b9adfd5),
	.w2(32'h3b0aefcb),
	.w3(32'h3a1a900d),
	.w4(32'hb9c5f05c),
	.w5(32'h371c5ba2),
	.w6(32'h3c1c2a6d),
	.w7(32'h3bb48c72),
	.w8(32'hbaf76803),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff64c3),
	.w1(32'h3aa35104),
	.w2(32'h3bddf29e),
	.w3(32'hba8b33b7),
	.w4(32'h3bed10e8),
	.w5(32'hbb9b73ac),
	.w6(32'hbbbeedee),
	.w7(32'h3a8e7f5f),
	.w8(32'hbbb5ca12),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50938e),
	.w1(32'h3c01ea20),
	.w2(32'h3bceeb6d),
	.w3(32'hbb368320),
	.w4(32'hbb0a655c),
	.w5(32'h3ba52e78),
	.w6(32'hba8e0e41),
	.w7(32'h3b4d5adb),
	.w8(32'h3bea6663),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af94bdf),
	.w1(32'hbb4a2df6),
	.w2(32'hb9ec32f2),
	.w3(32'hbbea0f4a),
	.w4(32'hbc2918ad),
	.w5(32'hba05799a),
	.w6(32'hbb4145be),
	.w7(32'hbc091646),
	.w8(32'hb9b30292),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c899b68),
	.w1(32'h3c8eb32e),
	.w2(32'h3bebc7b1),
	.w3(32'h3c4cf2f8),
	.w4(32'h3af3668a),
	.w5(32'hbc0e641d),
	.w6(32'h3cc6f7c6),
	.w7(32'h3c02946b),
	.w8(32'hbc90d8d4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6138bf),
	.w1(32'hba416ec3),
	.w2(32'hbb701048),
	.w3(32'hbbeb54b5),
	.w4(32'hbc0c5eee),
	.w5(32'h3952e326),
	.w6(32'hbb305cef),
	.w7(32'hbb98dd9c),
	.w8(32'hbad93007),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb11d6c),
	.w1(32'h3aacd1be),
	.w2(32'h3bf7904b),
	.w3(32'h3c44bc5e),
	.w4(32'h3ac230c5),
	.w5(32'h3b0c04d0),
	.w6(32'hbb96c179),
	.w7(32'hbc8d760e),
	.w8(32'hbb9ff7c4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff2818),
	.w1(32'h3a95c42a),
	.w2(32'h3b1b14dc),
	.w3(32'hbaca70ab),
	.w4(32'hbb19174c),
	.w5(32'h39de886a),
	.w6(32'hbb7cf405),
	.w7(32'hbb06daba),
	.w8(32'h3b68734e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d4d9),
	.w1(32'h3a91138d),
	.w2(32'hbb620eae),
	.w3(32'hbae2f30e),
	.w4(32'hbb80cc03),
	.w5(32'hbb19082b),
	.w6(32'h3b285158),
	.w7(32'hbb5b262a),
	.w8(32'hbb03de5e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae48013),
	.w1(32'h3b9b18f6),
	.w2(32'hba949669),
	.w3(32'h3bf63002),
	.w4(32'h3a074ec1),
	.w5(32'hbb0f5511),
	.w6(32'h3bde0aee),
	.w7(32'h3ad96954),
	.w8(32'hbb8dbb09),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae743fe),
	.w1(32'hb732237f),
	.w2(32'h3a628ce4),
	.w3(32'hbbaf917e),
	.w4(32'hbb40a75e),
	.w5(32'hbb2bdbb7),
	.w6(32'hbbc1a75b),
	.w7(32'hbae3a9f3),
	.w8(32'hbc099e11),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8284df),
	.w1(32'hbae5852e),
	.w2(32'h3a9e652b),
	.w3(32'hbb92e24a),
	.w4(32'hba9ef6da),
	.w5(32'h3bbdb2c7),
	.w6(32'hbad72b91),
	.w7(32'h3b080fdb),
	.w8(32'h3c3e031a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d6696),
	.w1(32'h3b34f182),
	.w2(32'h3c502876),
	.w3(32'hb9c4d75a),
	.w4(32'h3c2d52f0),
	.w5(32'hb99029af),
	.w6(32'hbb559696),
	.w7(32'h3b0edf34),
	.w8(32'h3b0c39e9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5c644),
	.w1(32'h3ba7424b),
	.w2(32'hba842d56),
	.w3(32'hb772c9d5),
	.w4(32'hbab02949),
	.w5(32'hbad7c3cc),
	.w6(32'hb829ec33),
	.w7(32'hbb7fc346),
	.w8(32'hbbce1628),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e9ed7),
	.w1(32'hbb101448),
	.w2(32'hba9e3800),
	.w3(32'hbba9aded),
	.w4(32'hbb0d9e7b),
	.w5(32'h3abd4750),
	.w6(32'hbb64f90f),
	.w7(32'hbb8655d7),
	.w8(32'h3a719931),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4e191),
	.w1(32'h3b6054b1),
	.w2(32'h3b1c9816),
	.w3(32'h3b8ac64f),
	.w4(32'h3ac0a129),
	.w5(32'h3bfde675),
	.w6(32'h3b0227c3),
	.w7(32'h38e76df3),
	.w8(32'h3bfb6fc5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a2f9),
	.w1(32'hbaedaabc),
	.w2(32'h3ae5d69c),
	.w3(32'hbafa8d33),
	.w4(32'h3aa4e5ef),
	.w5(32'hbadd367e),
	.w6(32'h39231aff),
	.w7(32'h387e2db2),
	.w8(32'h3a35d5dd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d1873),
	.w1(32'hbab24850),
	.w2(32'hbba73861),
	.w3(32'hbb20ee92),
	.w4(32'hbbad4e14),
	.w5(32'hbc31056f),
	.w6(32'h3a210f37),
	.w7(32'hbb6a93ef),
	.w8(32'hbc3246c6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50c55),
	.w1(32'hb96d5202),
	.w2(32'h3c1116bf),
	.w3(32'hba4c0350),
	.w4(32'h3c081762),
	.w5(32'hbb0ba23e),
	.w6(32'h3b3faff3),
	.w7(32'h3c9c5391),
	.w8(32'hbb375b4f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad80975),
	.w1(32'h3ad6fa5e),
	.w2(32'hbb06f325),
	.w3(32'h3a1faf38),
	.w4(32'h3b0333e3),
	.w5(32'h3b850be2),
	.w6(32'h3af1beda),
	.w7(32'h3b499896),
	.w8(32'h3c325d53),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03c13c),
	.w1(32'h3cd2cee1),
	.w2(32'h3bef6754),
	.w3(32'hbbaab176),
	.w4(32'h3bf61809),
	.w5(32'h3ad6dae6),
	.w6(32'h3c43f020),
	.w7(32'h3c9b0fa6),
	.w8(32'hba840025),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b1128),
	.w1(32'hbbbd223e),
	.w2(32'hbbf053f0),
	.w3(32'hb99f8590),
	.w4(32'hbac52bac),
	.w5(32'hbacaa483),
	.w6(32'hbb8657a3),
	.w7(32'hbb7f64a8),
	.w8(32'hbadce143),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f6d57),
	.w1(32'hba9736e3),
	.w2(32'hb9f5ab15),
	.w3(32'hbb6b30a0),
	.w4(32'hbb01bd4a),
	.w5(32'hba830fd0),
	.w6(32'hba9693f4),
	.w7(32'hbb56c206),
	.w8(32'h3a918ec5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd7016),
	.w1(32'hbaac3607),
	.w2(32'hba82129e),
	.w3(32'hbc08d750),
	.w4(32'hbbcb38c4),
	.w5(32'hbb9c79c0),
	.w6(32'hbb64574c),
	.w7(32'hbb9ad48f),
	.w8(32'hbbfd1500),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00c346),
	.w1(32'hbb0ff992),
	.w2(32'hbb14bfa9),
	.w3(32'hbb8e67e8),
	.w4(32'hb7f5145d),
	.w5(32'h3b3a7721),
	.w6(32'hbc02ed27),
	.w7(32'hba7a38c5),
	.w8(32'h398bd982),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc910940),
	.w1(32'h3c282505),
	.w2(32'h3ba41798),
	.w3(32'hbbfacd1b),
	.w4(32'h3c378673),
	.w5(32'hbc1b30bc),
	.w6(32'hbc5cdb93),
	.w7(32'h3bb76938),
	.w8(32'h3bf08f4d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bd33e),
	.w1(32'h3b983e79),
	.w2(32'h3bc4b12c),
	.w3(32'hba452c47),
	.w4(32'h3b457870),
	.w5(32'h3c4855ed),
	.w6(32'h39802cb0),
	.w7(32'hbc01c8de),
	.w8(32'hbc2a3b72),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fff2),
	.w1(32'h3c7f4934),
	.w2(32'h3bedd8fd),
	.w3(32'hba631f7b),
	.w4(32'hbb593f4b),
	.w5(32'h3af34d14),
	.w6(32'h3bb39ec4),
	.w7(32'hbb090a48),
	.w8(32'hbc240197),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ca99),
	.w1(32'hbc8995ad),
	.w2(32'hbc747122),
	.w3(32'hbca44011),
	.w4(32'hbca27048),
	.w5(32'hbcbd398a),
	.w6(32'hbc2b5c55),
	.w7(32'hbc875310),
	.w8(32'hbc9eb8e3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bca02),
	.w1(32'h3aa384a3),
	.w2(32'h3bab3c0f),
	.w3(32'h3a14781f),
	.w4(32'h3bae9b31),
	.w5(32'h3b02b524),
	.w6(32'h3a4f31a1),
	.w7(32'h3bb69eb2),
	.w8(32'h3b8c2e8b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924c45b),
	.w1(32'hbbf6655a),
	.w2(32'hbbaf7c32),
	.w3(32'h3b581082),
	.w4(32'hbb61caea),
	.w5(32'hbb61d976),
	.w6(32'h368f8b52),
	.w7(32'hbb87c45f),
	.w8(32'hbbacfe25),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc162ba5),
	.w1(32'hbb73f415),
	.w2(32'h3b908a08),
	.w3(32'hb8de74ea),
	.w4(32'h3b1babda),
	.w5(32'h3b5feaf8),
	.w6(32'hb92c2f7a),
	.w7(32'h3ac2314a),
	.w8(32'h3b32f1b3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42578a),
	.w1(32'h3ba13191),
	.w2(32'h3a956d1c),
	.w3(32'h39ff3310),
	.w4(32'hba8c87c2),
	.w5(32'h3bdb2890),
	.w6(32'h3a3d2efd),
	.w7(32'h3acd4f81),
	.w8(32'h3b16b4be),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeae7e8),
	.w1(32'h3ac55d3a),
	.w2(32'h3bc2f5b6),
	.w3(32'hbad8fcf2),
	.w4(32'h3bd69d9f),
	.w5(32'h3b0583a9),
	.w6(32'hbb55e770),
	.w7(32'h3b8b81b2),
	.w8(32'hba261eab),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c5ed),
	.w1(32'h39a4e496),
	.w2(32'h3af89a81),
	.w3(32'h3bbcefcc),
	.w4(32'hba94e41b),
	.w5(32'hbc0e87d0),
	.w6(32'hbb816c70),
	.w7(32'hbbef9b6d),
	.w8(32'hbc186e8b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7513d),
	.w1(32'hbb140727),
	.w2(32'h3c2c8d06),
	.w3(32'h3bddadc8),
	.w4(32'hba4f902b),
	.w5(32'hbb0eb40b),
	.w6(32'hbb0cd8f8),
	.w7(32'hbc1fe9b0),
	.w8(32'hbbccb8e7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e74b),
	.w1(32'hbc15250d),
	.w2(32'hbc21c0ff),
	.w3(32'hbc02c7f2),
	.w4(32'hbc22e95b),
	.w5(32'hbc09ef2d),
	.w6(32'hbc00d2a9),
	.w7(32'hbc305bc9),
	.w8(32'hbc41df99),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d372c),
	.w1(32'h3ba19404),
	.w2(32'h3c047dec),
	.w3(32'hba9a8ad3),
	.w4(32'h3ae73c62),
	.w5(32'h3c095ea1),
	.w6(32'hbadd2986),
	.w7(32'h3ab08489),
	.w8(32'h3b95ffd8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc5621),
	.w1(32'h3b21e9d3),
	.w2(32'h3b6636b8),
	.w3(32'hbb6dec09),
	.w4(32'hbbec2f81),
	.w5(32'h37c4c9c2),
	.w6(32'hbba87d42),
	.w7(32'hbb4a95d6),
	.w8(32'h3bf113e9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68d5a4),
	.w1(32'hbbca53b8),
	.w2(32'hbb98ccd2),
	.w3(32'hba8db417),
	.w4(32'h3a8da4d7),
	.w5(32'hbb82d561),
	.w6(32'hbc39944c),
	.w7(32'hbc081d9f),
	.w8(32'hbbade770),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a622f42),
	.w1(32'h3b42b4c6),
	.w2(32'h3b99187e),
	.w3(32'h3a6a4723),
	.w4(32'hbac2dafb),
	.w5(32'h3b54884b),
	.w6(32'hbb602ed8),
	.w7(32'hbb984b23),
	.w8(32'hb9788791),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2fc5f),
	.w1(32'hbb2f9fc4),
	.w2(32'hbb56d6ca),
	.w3(32'hbb33e426),
	.w4(32'hbb26ffa2),
	.w5(32'hb9130df2),
	.w6(32'hb8d1722e),
	.w7(32'hbaa400d2),
	.w8(32'hbb0858a6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c36a9),
	.w1(32'hbc1701e5),
	.w2(32'hba0e1c6d),
	.w3(32'hbc010d25),
	.w4(32'h3b1ab67d),
	.w5(32'h3b4caa4b),
	.w6(32'hbbcac074),
	.w7(32'h3a80e416),
	.w8(32'h3ae2c566),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13e440),
	.w1(32'hbb37c3d6),
	.w2(32'hbb694697),
	.w3(32'hbaf45a4d),
	.w4(32'hbb23678a),
	.w5(32'h3ad60da8),
	.w6(32'hbaa93ef5),
	.w7(32'hbac5e96f),
	.w8(32'hba0e7ba2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ca44b),
	.w1(32'h3c122536),
	.w2(32'h3bc68ab5),
	.w3(32'h3b9e2608),
	.w4(32'h3bb20241),
	.w5(32'hbb817c6b),
	.w6(32'h3c1aedb0),
	.w7(32'h3c88d683),
	.w8(32'hb904ad21),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb673c4),
	.w1(32'hbbdec366),
	.w2(32'hbaaa5b5c),
	.w3(32'hbbd599f2),
	.w4(32'hb9fd7a77),
	.w5(32'hbc36b98f),
	.w6(32'hbab37076),
	.w7(32'h3a2c4de8),
	.w8(32'hbc346830),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba8158),
	.w1(32'hba927e6e),
	.w2(32'hbb34d664),
	.w3(32'hbb1f8c48),
	.w4(32'hbb5d2131),
	.w5(32'hbb3ff91f),
	.w6(32'hbb269016),
	.w7(32'hbaed7c12),
	.w8(32'hbb179ba6),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8a83),
	.w1(32'h3ab67e40),
	.w2(32'hbb334f01),
	.w3(32'hbbd4ee34),
	.w4(32'hbc45d529),
	.w5(32'hb7a88fca),
	.w6(32'hbb007e15),
	.w7(32'hbc62ec76),
	.w8(32'hbbbd0b42),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386f4c46),
	.w1(32'hbb0db38c),
	.w2(32'h3c10d9ad),
	.w3(32'hbb9a8d15),
	.w4(32'h3bcc0e4e),
	.w5(32'h3c2aca27),
	.w6(32'hbbeb7ca9),
	.w7(32'hbb017702),
	.w8(32'h3bc56977),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97fde),
	.w1(32'hbbad099b),
	.w2(32'hbc1d510a),
	.w3(32'h3b4db69b),
	.w4(32'hbb391c55),
	.w5(32'hbbf6e7e5),
	.w6(32'hb9253d48),
	.w7(32'hb9a60687),
	.w8(32'hbb5456ba),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b6884),
	.w1(32'h3ae8765c),
	.w2(32'hbad51b8c),
	.w3(32'h3ad47bc0),
	.w4(32'hbca65203),
	.w5(32'hbc96daae),
	.w6(32'hbb8a5f2f),
	.w7(32'hbc54ba18),
	.w8(32'h392bea4b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707868),
	.w1(32'hbc555e61),
	.w2(32'hbc245e94),
	.w3(32'hbc0470ed),
	.w4(32'hbc446cdb),
	.w5(32'hba98cf78),
	.w6(32'hbb1ea9d7),
	.w7(32'hbbfa33db),
	.w8(32'hbbc3f5a8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc026e55),
	.w1(32'h3c2bd093),
	.w2(32'h3c805f17),
	.w3(32'hb9038ba4),
	.w4(32'h3c2ea5e8),
	.w5(32'h3ca0cdec),
	.w6(32'hbbad9537),
	.w7(32'hbb2aef7f),
	.w8(32'h3c4c6b17),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaae31a),
	.w1(32'hbc01ab05),
	.w2(32'hbb12872b),
	.w3(32'hbafd61bd),
	.w4(32'hbbf6cf37),
	.w5(32'hbc1e7473),
	.w6(32'hbbf956e3),
	.w7(32'hbc3192dd),
	.w8(32'hbc041a69),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc406d2c),
	.w1(32'hbc3d73ce),
	.w2(32'hbb77e9f7),
	.w3(32'hbaaa6b55),
	.w4(32'h3be616a2),
	.w5(32'hbc74a480),
	.w6(32'hbb7d40d3),
	.w7(32'hbae82771),
	.w8(32'hbc149370),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817079),
	.w1(32'hbb7fca2e),
	.w2(32'hbb9650fa),
	.w3(32'hbbb2a1d2),
	.w4(32'hbbbc6396),
	.w5(32'h3a1539cd),
	.w6(32'hbb9e659e),
	.w7(32'hbb50e0bb),
	.w8(32'h3a9a2977),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44e3c1),
	.w1(32'h3c0c52d5),
	.w2(32'h3bc52475),
	.w3(32'h3a5a59fa),
	.w4(32'hbae2e58f),
	.w5(32'h3b61e0b0),
	.w6(32'hba4432b8),
	.w7(32'hbbbb213f),
	.w8(32'h3ad6c784),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b8e52),
	.w1(32'hbaf7a24b),
	.w2(32'hbbb6218d),
	.w3(32'hbb8bf138),
	.w4(32'hbc242b05),
	.w5(32'hbc958c17),
	.w6(32'hbc3b6919),
	.w7(32'hbc667a7b),
	.w8(32'hbc47af6d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf8873),
	.w1(32'hbb3fe961),
	.w2(32'h3c247db1),
	.w3(32'h3ca9be18),
	.w4(32'hbcc8a81e),
	.w5(32'hbb1144ab),
	.w6(32'h3befd3bb),
	.w7(32'hbc9d4ae2),
	.w8(32'hbc81a295),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe806cb),
	.w1(32'hbc81943b),
	.w2(32'hbc11a2ae),
	.w3(32'hbc09fa37),
	.w4(32'hbc089af5),
	.w5(32'hbc329026),
	.w6(32'hbbe3a352),
	.w7(32'hbbf85544),
	.w8(32'hbc40769b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad0304),
	.w1(32'hbc1ca2b9),
	.w2(32'hbb482b67),
	.w3(32'hbc2158a5),
	.w4(32'hbc396996),
	.w5(32'hbc286aeb),
	.w6(32'hbc534606),
	.w7(32'hbc46b492),
	.w8(32'hbc35656f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4e2a8),
	.w1(32'hbc54e2e5),
	.w2(32'hbb395d69),
	.w3(32'hbadd80db),
	.w4(32'hbcfdf510),
	.w5(32'hbc8924ef),
	.w6(32'hbc22d9d1),
	.w7(32'hbcdbcbdf),
	.w8(32'hbc071b3d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb410d3a),
	.w1(32'hbb0a54d7),
	.w2(32'hbb5cebfb),
	.w3(32'h3a41dffc),
	.w4(32'hbb335f06),
	.w5(32'h3a77f8d6),
	.w6(32'h3b0a3de2),
	.w7(32'hbb6a3817),
	.w8(32'h390bd0b6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf07ec),
	.w1(32'hbb9e9d75),
	.w2(32'h3c096582),
	.w3(32'h3c3e137f),
	.w4(32'hbb855092),
	.w5(32'hbc081653),
	.w6(32'hbb5708c7),
	.w7(32'hbd12dc3b),
	.w8(32'hbcb78287),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0ee2),
	.w1(32'hbb9ca99c),
	.w2(32'h381ee950),
	.w3(32'h3bc6faff),
	.w4(32'hba70321a),
	.w5(32'hbb847e35),
	.w6(32'h3b9fbb92),
	.w7(32'hb95f6127),
	.w8(32'hbaa359e8),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb856231f),
	.w1(32'hbb07141d),
	.w2(32'hba57200c),
	.w3(32'hba256cfd),
	.w4(32'hbb19c272),
	.w5(32'hbb5807c2),
	.w6(32'hba4ef6d0),
	.w7(32'hbb2dd279),
	.w8(32'hbb045ac3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24037f),
	.w1(32'hb9d9ffb3),
	.w2(32'hbaba29a5),
	.w3(32'hbb97e25c),
	.w4(32'hbb68bc81),
	.w5(32'hbb772e4b),
	.w6(32'hbb435c1d),
	.w7(32'hbb03af1c),
	.w8(32'hbb695fe7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b043f05),
	.w1(32'h3b7afa2e),
	.w2(32'h3b2da335),
	.w3(32'h39d7dcf2),
	.w4(32'hba2fa0c6),
	.w5(32'h3c07cb9f),
	.w6(32'h3b007b02),
	.w7(32'hbaf3c27c),
	.w8(32'h3ba68cff),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc793aa),
	.w1(32'h39daddd4),
	.w2(32'h3b3200fa),
	.w3(32'hba8aa247),
	.w4(32'h3a98a6e5),
	.w5(32'h3ac17e63),
	.w6(32'hbbdad693),
	.w7(32'hbb4445e6),
	.w8(32'hbb2fa794),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68ca95),
	.w1(32'h3c2538e0),
	.w2(32'h3bd66961),
	.w3(32'h39991799),
	.w4(32'h3b71c0cd),
	.w5(32'hbb5c704b),
	.w6(32'h3c5220de),
	.w7(32'h3c2c09d4),
	.w8(32'h3b230c0c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e1535),
	.w1(32'hba9f366c),
	.w2(32'hbb2c2f9c),
	.w3(32'hbb7c35fe),
	.w4(32'hba3c31ae),
	.w5(32'h3b5e9e2b),
	.w6(32'hbb9bf155),
	.w7(32'hbb065dbb),
	.w8(32'hba01ebeb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a03fd),
	.w1(32'hbc1910df),
	.w2(32'hbbe3c6e8),
	.w3(32'h3bda854c),
	.w4(32'h3aa26e57),
	.w5(32'hbbab182d),
	.w6(32'hbc08a7b8),
	.w7(32'hbc831660),
	.w8(32'hbcd6a6e3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376b6d),
	.w1(32'h3bfe6206),
	.w2(32'h3be82f74),
	.w3(32'h3b3d570f),
	.w4(32'hb9efd2fc),
	.w5(32'h3b3151b1),
	.w6(32'hbaf04ce1),
	.w7(32'h3bc54eb9),
	.w8(32'h3b8f8a86),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6302e),
	.w1(32'h3b1021b1),
	.w2(32'h3bcf66b2),
	.w3(32'hbb0dcc03),
	.w4(32'hbaf2e595),
	.w5(32'hba25d7a0),
	.w6(32'hbb5e6214),
	.w7(32'hbb57d09b),
	.w8(32'hba8cd9c8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d9bde),
	.w1(32'h39af83ba),
	.w2(32'h3aaca144),
	.w3(32'hbabf8754),
	.w4(32'h3ac09627),
	.w5(32'hbb1c750a),
	.w6(32'hbb26db57),
	.w7(32'hba4f54f4),
	.w8(32'hbaae5416),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb766a46),
	.w1(32'hbb7962dc),
	.w2(32'hbb68d91d),
	.w3(32'h3a8534ac),
	.w4(32'hbb5e7cf3),
	.w5(32'hbacd8633),
	.w6(32'h3a894f6f),
	.w7(32'hbb59d403),
	.w8(32'hbb72b9e2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c01af),
	.w1(32'h3a4acf16),
	.w2(32'h3b1cce0a),
	.w3(32'hbb0695c4),
	.w4(32'h3b02f3a1),
	.w5(32'hbaa5a42f),
	.w6(32'hba4d1154),
	.w7(32'h3b02e222),
	.w8(32'hba1467bd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7df859),
	.w1(32'hbb06b65a),
	.w2(32'hbb619d87),
	.w3(32'h390c20e3),
	.w4(32'hbb3c935e),
	.w5(32'hbbb0bab4),
	.w6(32'h3b00bd15),
	.w7(32'hba9cead3),
	.w8(32'hbb70dea8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ea6b),
	.w1(32'hbb0dc539),
	.w2(32'hbb435f2c),
	.w3(32'hbbabb5b5),
	.w4(32'hbc035d98),
	.w5(32'hba8bad84),
	.w6(32'hbc13b499),
	.w7(32'hbc4ac233),
	.w8(32'hbbbda6d1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc15b5),
	.w1(32'hbb90e0d3),
	.w2(32'hbb5b0de4),
	.w3(32'h3b0155bd),
	.w4(32'h3aae0df1),
	.w5(32'h3bd36be8),
	.w6(32'hbb5ca50b),
	.w7(32'hbb4f0ddf),
	.w8(32'h3afe5f9a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe32661),
	.w1(32'hbad5de55),
	.w2(32'h3ad4e44f),
	.w3(32'h3bc29a72),
	.w4(32'h3a23861d),
	.w5(32'hbbc26e97),
	.w6(32'hbbba5450),
	.w7(32'h391c710f),
	.w8(32'hbbd2208f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3774eb7f),
	.w1(32'hbbc99935),
	.w2(32'hbb638106),
	.w3(32'hbc31b03b),
	.w4(32'h3b29a865),
	.w5(32'hba421eb0),
	.w6(32'hbbb34925),
	.w7(32'h3b7fb5e6),
	.w8(32'h3b693b03),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21d2b5),
	.w1(32'h3bee8bf3),
	.w2(32'h3c2149cc),
	.w3(32'h3b5de1e2),
	.w4(32'h3b60927f),
	.w5(32'hba2a1a36),
	.w6(32'hbb157488),
	.w7(32'h3bfb4d7b),
	.w8(32'hbb1393e6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e710),
	.w1(32'h3b6e5d6a),
	.w2(32'h3c09c85a),
	.w3(32'hbb454cc4),
	.w4(32'h3a4738e3),
	.w5(32'h3b0709c6),
	.w6(32'hbb9f2418),
	.w7(32'h3b593f81),
	.w8(32'h3a9a3ca0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c241366),
	.w1(32'h3b31d047),
	.w2(32'h3b341050),
	.w3(32'hb9fbba40),
	.w4(32'hbb28c5e2),
	.w5(32'h3b0847d5),
	.w6(32'hbb0d6fa0),
	.w7(32'hbad9574d),
	.w8(32'h3aaadf4e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7a0b7),
	.w1(32'h3b97e54d),
	.w2(32'h3bfddc98),
	.w3(32'h3b0a1f81),
	.w4(32'h3b80aafc),
	.w5(32'hbb883257),
	.w6(32'hbb4f19ca),
	.w7(32'h3acd7c10),
	.w8(32'h391e7362),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcbea2),
	.w1(32'hba0dc29b),
	.w2(32'hb98277ea),
	.w3(32'h3ac61afb),
	.w4(32'h3b5a9017),
	.w5(32'h3cbb4259),
	.w6(32'hbc2c991f),
	.w7(32'hbc9d3cea),
	.w8(32'hbc7a4f7a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b737819),
	.w1(32'h3bca6726),
	.w2(32'h3be9978e),
	.w3(32'h3b26cbe3),
	.w4(32'h3c809ecf),
	.w5(32'h3c3f4e77),
	.w6(32'hbc7ddd2d),
	.w7(32'hba8ed28d),
	.w8(32'h3c29d111),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b8130),
	.w1(32'h3c0ab80b),
	.w2(32'h3c34e9c6),
	.w3(32'h3a0bbd1b),
	.w4(32'h3b8a27fe),
	.w5(32'hbb17cfed),
	.w6(32'hbc102516),
	.w7(32'h3b60012f),
	.w8(32'hbb757263),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8342a3),
	.w1(32'hb8065ef1),
	.w2(32'h3ad71ea2),
	.w3(32'h3a30510d),
	.w4(32'h3ac20ff8),
	.w5(32'h38dd773c),
	.w6(32'hbb48fa0f),
	.w7(32'hbbed0967),
	.w8(32'hbb90ff7b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab020eb),
	.w1(32'hb96c8a6f),
	.w2(32'hbaa74786),
	.w3(32'hbaa7e553),
	.w4(32'hbaddcf1d),
	.w5(32'hbc24bd93),
	.w6(32'h3959c381),
	.w7(32'hba902509),
	.w8(32'hbbdfc4a1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03dca7),
	.w1(32'hbb303bb3),
	.w2(32'hbb9fbcf2),
	.w3(32'hbbec6c9d),
	.w4(32'hbbac9c50),
	.w5(32'h3bbd6dde),
	.w6(32'hbbe7f34f),
	.w7(32'hbbbda30c),
	.w8(32'h3a93bac3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8864fe),
	.w1(32'hbad02208),
	.w2(32'h3b18ad1d),
	.w3(32'hbbc2db5b),
	.w4(32'h3b0b9471),
	.w5(32'hbc0664d4),
	.w6(32'hbc225595),
	.w7(32'h38efe353),
	.w8(32'hbc002e9f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb363548),
	.w1(32'hbb0ec9e7),
	.w2(32'h3b923b7f),
	.w3(32'hbb358c57),
	.w4(32'hbb4138aa),
	.w5(32'hbc1dd4ed),
	.w6(32'hbc5c3050),
	.w7(32'hbb8eda1e),
	.w8(32'hbb6e1e33),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39e412),
	.w1(32'hbc39a041),
	.w2(32'hbc4f49d4),
	.w3(32'hbb7945a7),
	.w4(32'hbbb265c6),
	.w5(32'hbab92f10),
	.w6(32'h3b68d6b7),
	.w7(32'hbc0142ae),
	.w8(32'hbad12b8b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b917aa7),
	.w1(32'h3b04fe81),
	.w2(32'h3ba7f182),
	.w3(32'h3b75aba9),
	.w4(32'hba71032b),
	.w5(32'h3b25c61b),
	.w6(32'hbb9abc06),
	.w7(32'h3aaa9033),
	.w8(32'hba954caa),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d0f23),
	.w1(32'hbba98936),
	.w2(32'h3ae4ee43),
	.w3(32'h3b372945),
	.w4(32'hbbd9bee5),
	.w5(32'hbbc90fad),
	.w6(32'hbc0d261f),
	.w7(32'hbc0d9f4f),
	.w8(32'hbb8d2ba2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b492d4d),
	.w1(32'hbb7bd148),
	.w2(32'hbae424b1),
	.w3(32'h3a3e5634),
	.w4(32'hbae55522),
	.w5(32'hbab67a80),
	.w6(32'hbbade2e7),
	.w7(32'hbc137b70),
	.w8(32'hbc444c62),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2abf82),
	.w1(32'hbaad0ba9),
	.w2(32'h3affb459),
	.w3(32'h3aa78fb2),
	.w4(32'h394e81b2),
	.w5(32'h3bfd3ed7),
	.w6(32'hbbb0d3b7),
	.w7(32'hbb8db857),
	.w8(32'h3c1fa156),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66be6d),
	.w1(32'h3afb579e),
	.w2(32'h3b095c60),
	.w3(32'h3a79a48f),
	.w4(32'hbb932ca3),
	.w5(32'h3b47eb81),
	.w6(32'hbb4b67af),
	.w7(32'hbbc7aa0e),
	.w8(32'h3ab85540),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeecc97),
	.w1(32'hbc4e956c),
	.w2(32'hbcae7073),
	.w3(32'hbc467434),
	.w4(32'hbb9c0cd2),
	.w5(32'hbbc3d3d8),
	.w6(32'hbc0d3185),
	.w7(32'hbb76d3c1),
	.w8(32'hbb82ce4b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4393fd),
	.w1(32'h3acfd79f),
	.w2(32'h3bb289f0),
	.w3(32'hbaa59f56),
	.w4(32'hbaf1609e),
	.w5(32'hbaad84a7),
	.w6(32'h3b9ef708),
	.w7(32'hbb3cce4d),
	.w8(32'hbb7e9884),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abff133),
	.w1(32'hb9140a54),
	.w2(32'h3bdf2759),
	.w3(32'h3b89b538),
	.w4(32'h3b2760cb),
	.w5(32'hbb42a11c),
	.w6(32'hbb24f427),
	.w7(32'h3aa19cda),
	.w8(32'hbb916474),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79afb1),
	.w1(32'hbb268f1f),
	.w2(32'hb9916586),
	.w3(32'hbaff0241),
	.w4(32'h3b67501c),
	.w5(32'hbb27bb30),
	.w6(32'hbc060606),
	.w7(32'hba3e7ef7),
	.w8(32'hbb87d140),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e52a8a),
	.w1(32'hbb2d04cb),
	.w2(32'hbb4569a8),
	.w3(32'h39ba14e1),
	.w4(32'hbac7d3ca),
	.w5(32'hbaee65dd),
	.w6(32'hbb8047a1),
	.w7(32'hbbae5549),
	.w8(32'hba2701a5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb490f78),
	.w1(32'hbbe20c27),
	.w2(32'hbaca3795),
	.w3(32'hbb5734b8),
	.w4(32'hbb86c5e8),
	.w5(32'hbbd51b31),
	.w6(32'h3a99a068),
	.w7(32'hbbdd2349),
	.w8(32'hbb9c2963),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c650368),
	.w1(32'h3c0bb747),
	.w2(32'h3b5ef830),
	.w3(32'h3ada92de),
	.w4(32'h3b6ba443),
	.w5(32'h3b5edfb7),
	.w6(32'hbb1002c7),
	.w7(32'hbaefe319),
	.w8(32'h3afb9059),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa72f7),
	.w1(32'h3b97a41c),
	.w2(32'h3baf0d36),
	.w3(32'h3bd1587e),
	.w4(32'h3a9f7f64),
	.w5(32'hb9e81651),
	.w6(32'hba373a94),
	.w7(32'h3a3905db),
	.w8(32'hba25efba),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41eaa0),
	.w1(32'h3b218211),
	.w2(32'h3a2219f3),
	.w3(32'hba7a9e4a),
	.w4(32'hbab768d2),
	.w5(32'h3b1803ca),
	.w6(32'hb980dae3),
	.w7(32'hbb864f80),
	.w8(32'h3b8ddbfc),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c87e6),
	.w1(32'hb9da9aef),
	.w2(32'hbad41080),
	.w3(32'hbb720b4e),
	.w4(32'hbb80a497),
	.w5(32'hb9e4c349),
	.w6(32'hbba8eed9),
	.w7(32'hbbd3697a),
	.w8(32'h3a835b7c),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e533),
	.w1(32'hbbc54d1e),
	.w2(32'h3c0118a1),
	.w3(32'h3ba913d0),
	.w4(32'hbc220f0a),
	.w5(32'hbc14746a),
	.w6(32'hbbbb51e3),
	.w7(32'hbc8035fa),
	.w8(32'hbbc33ff2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f415),
	.w1(32'h3bb343a0),
	.w2(32'hbc5101f2),
	.w3(32'hbbfc4ab8),
	.w4(32'hba2ac96a),
	.w5(32'hbc95e688),
	.w6(32'hbbab9e09),
	.w7(32'hbab551a5),
	.w8(32'hbc00b0cc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20ecf1),
	.w1(32'hbb230285),
	.w2(32'hba2ea1eb),
	.w3(32'hbbc9dee9),
	.w4(32'h39207f78),
	.w5(32'hbb7e0e3f),
	.w6(32'h3a008816),
	.w7(32'h3a97e369),
	.w8(32'hbb662503),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2bcc5),
	.w1(32'hbb167065),
	.w2(32'hbb042a55),
	.w3(32'hbb1788e7),
	.w4(32'hbae4101d),
	.w5(32'h3b578ca3),
	.w6(32'hbae44b7c),
	.w7(32'hba921d6c),
	.w8(32'h3a9bb13d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8524),
	.w1(32'h3b4e2d88),
	.w2(32'h3baaacad),
	.w3(32'h3b6f9941),
	.w4(32'h3b828525),
	.w5(32'hbb85a4b5),
	.w6(32'hbbef6f85),
	.w7(32'hbac18069),
	.w8(32'hbc0cb8a2),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb553ddc),
	.w1(32'hbb84352e),
	.w2(32'h3a84a141),
	.w3(32'hbc257835),
	.w4(32'hbc364e6c),
	.w5(32'h39c5fd84),
	.w6(32'hbc1e691f),
	.w7(32'hbbfb1a0f),
	.w8(32'hbacbcfa4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92810e),
	.w1(32'hbb552363),
	.w2(32'hbb126eb5),
	.w3(32'hbab76c4a),
	.w4(32'h3abfd6d4),
	.w5(32'hbb86c3b7),
	.w6(32'hba5e0b73),
	.w7(32'h3b1e9c05),
	.w8(32'h3943a5fc),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac93021),
	.w1(32'h3b158651),
	.w2(32'h3aae4dde),
	.w3(32'h3a60100c),
	.w4(32'hbb737e6e),
	.w5(32'h3a06dd46),
	.w6(32'hbb6be125),
	.w7(32'hbae5cc37),
	.w8(32'hbab3e81b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac19d23),
	.w1(32'hba2a6db9),
	.w2(32'hbb3fd7a4),
	.w3(32'h3b23712b),
	.w4(32'hbb615302),
	.w5(32'hbb64f750),
	.w6(32'hba1574ed),
	.w7(32'hbb3ab7b7),
	.w8(32'hbb4209bf),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a55e9e),
	.w1(32'h3b68bfc3),
	.w2(32'h3b63086f),
	.w3(32'hba1506be),
	.w4(32'hbb3a0e1d),
	.w5(32'h3a32cb1d),
	.w6(32'hbbc21425),
	.w7(32'hbbb73cab),
	.w8(32'hbb765102),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ad6d1),
	.w1(32'hbb5be670),
	.w2(32'hb8fb3d4e),
	.w3(32'hbb8d35f1),
	.w4(32'hbb4d3da9),
	.w5(32'h3a5f2833),
	.w6(32'hbbd10509),
	.w7(32'h3aa9cb5c),
	.w8(32'h3b690e42),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2290c),
	.w1(32'hba9ef158),
	.w2(32'hbbb6b0bf),
	.w3(32'hbb8af9d9),
	.w4(32'hbbc3b675),
	.w5(32'hbbdc9423),
	.w6(32'hbb8e76ff),
	.w7(32'hbbe0778a),
	.w8(32'hbbc0f723),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00768e),
	.w1(32'h3af6c13c),
	.w2(32'h3ac22bab),
	.w3(32'h3abf802a),
	.w4(32'hba9af50b),
	.w5(32'h3aa8c036),
	.w6(32'h3af36a47),
	.w7(32'h3aa1277f),
	.w8(32'h3b650678),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f3645),
	.w1(32'hbb5d10d4),
	.w2(32'hbb8e85d7),
	.w3(32'hbb1accae),
	.w4(32'h3b8adf95),
	.w5(32'h3b737cd5),
	.w6(32'hbb89dcb3),
	.w7(32'h3b771c61),
	.w8(32'h3b3be8aa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b266a80),
	.w1(32'hbb3913a8),
	.w2(32'h3b3c7cf7),
	.w3(32'hbb647755),
	.w4(32'h3b9b215a),
	.w5(32'h39374ad9),
	.w6(32'hbbd0faa7),
	.w7(32'h3b42bcee),
	.w8(32'h3b9a2910),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d354a5),
	.w1(32'h3c0f3b38),
	.w2(32'h3c06c20e),
	.w3(32'hba4cfb55),
	.w4(32'h3a4d07c7),
	.w5(32'h3b7b7862),
	.w6(32'hbb3c13a2),
	.w7(32'hbb0a04e5),
	.w8(32'h3ac89cdf),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9cec),
	.w1(32'hbb018a6f),
	.w2(32'hbb738556),
	.w3(32'hbc007486),
	.w4(32'hbb79b882),
	.w5(32'h3b65cb23),
	.w6(32'hbb82ff7c),
	.w7(32'hbc046c2d),
	.w8(32'hba9eee6f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae05b10),
	.w1(32'hbba16c18),
	.w2(32'h3b1ae674),
	.w3(32'h3c2d3611),
	.w4(32'h3b62d8f6),
	.w5(32'h3be6f7ca),
	.w6(32'h3a467414),
	.w7(32'hbbfb22be),
	.w8(32'hbbf93753),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f96346),
	.w1(32'hba138c71),
	.w2(32'hba179d32),
	.w3(32'hb92793a7),
	.w4(32'h38eb963b),
	.w5(32'h3b52c6d3),
	.w6(32'h399ffe70),
	.w7(32'hba59511c),
	.w8(32'hba0252a3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0681b1),
	.w1(32'hbaedae40),
	.w2(32'h3aac9e93),
	.w3(32'hba6a719f),
	.w4(32'hba8e7413),
	.w5(32'hbbd1ae93),
	.w6(32'h39c47c38),
	.w7(32'hbb83208a),
	.w8(32'hbbf46383),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cd41fa),
	.w1(32'h3bdf31cc),
	.w2(32'h3b40f2d4),
	.w3(32'hbbca99b0),
	.w4(32'h3b669ead),
	.w5(32'hbb3efc3d),
	.w6(32'hbb944d62),
	.w7(32'h3b397fce),
	.w8(32'h3a226297),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c011446),
	.w1(32'h3bd65bda),
	.w2(32'h3a2f025b),
	.w3(32'hbb11c494),
	.w4(32'h3a48b726),
	.w5(32'h3ba467ce),
	.w6(32'hbb870b29),
	.w7(32'hbb108b44),
	.w8(32'h39437d45),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac53fed),
	.w1(32'h3bb9b71f),
	.w2(32'h3b30d8cf),
	.w3(32'h3a209602),
	.w4(32'h3b173cb0),
	.w5(32'hb98a4140),
	.w6(32'h3a846d7c),
	.w7(32'hbb80e8fc),
	.w8(32'h398f5c76),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981d431),
	.w1(32'h3bb76e5c),
	.w2(32'h3b9bc301),
	.w3(32'hba922482),
	.w4(32'hb9fb7f12),
	.w5(32'h3c079eff),
	.w6(32'hbb87e615),
	.w7(32'hbba19b3f),
	.w8(32'h3bd2dac2),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c1cea),
	.w1(32'h3b38d38c),
	.w2(32'h3b152160),
	.w3(32'h3b8a13db),
	.w4(32'h3b07c21e),
	.w5(32'h3b195769),
	.w6(32'h3b177df4),
	.w7(32'h3a8305c7),
	.w8(32'hba958720),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a58d),
	.w1(32'h3b45dd6d),
	.w2(32'h3be65499),
	.w3(32'hbb556a6f),
	.w4(32'h37b0772c),
	.w5(32'h3b1cbd06),
	.w6(32'hbc3a90d5),
	.w7(32'hbb2b4750),
	.w8(32'h3b0fbdf2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb941193f),
	.w1(32'h3a8e7060),
	.w2(32'h3b4436de),
	.w3(32'h3ae4835a),
	.w4(32'h396b1efd),
	.w5(32'hbb948692),
	.w6(32'h3b070b97),
	.w7(32'h3a103ed5),
	.w8(32'hbb6055f1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08b51),
	.w1(32'hb9a723af),
	.w2(32'hba42a99a),
	.w3(32'hba61fff0),
	.w4(32'h39cc5fce),
	.w5(32'hbb36a87a),
	.w6(32'hba8d2ab9),
	.w7(32'hb786674e),
	.w8(32'hbb4e2ab6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa936e),
	.w1(32'h3980c5aa),
	.w2(32'hbb092328),
	.w3(32'hbb94b6c1),
	.w4(32'hbafdd312),
	.w5(32'hbb596f10),
	.w6(32'hb957e9be),
	.w7(32'h3a87102d),
	.w8(32'h3a92f121),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03c57),
	.w1(32'hbbdc8115),
	.w2(32'hbb3a0236),
	.w3(32'h3b38ee07),
	.w4(32'h3bac68f8),
	.w5(32'h3c307cdf),
	.w6(32'hbc115b1d),
	.w7(32'hbb0406eb),
	.w8(32'h398f36ad),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17f87d),
	.w1(32'h39e1d1d1),
	.w2(32'hbb2078ac),
	.w3(32'h3acf4d8b),
	.w4(32'h3b33db37),
	.w5(32'h3a9129c7),
	.w6(32'hba8961d7),
	.w7(32'h3aec700f),
	.w8(32'h3b63b544),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad575),
	.w1(32'h3b2d1804),
	.w2(32'hbb161a0c),
	.w3(32'hbb7c1c31),
	.w4(32'hbb488f52),
	.w5(32'h3a60e3c3),
	.w6(32'hba440506),
	.w7(32'hbb380954),
	.w8(32'hbb779776),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba089dc1),
	.w1(32'hbbe7abb9),
	.w2(32'hbbfcd195),
	.w3(32'hbb1cdab5),
	.w4(32'hbbc37305),
	.w5(32'hbb5fd268),
	.w6(32'hbbf25fa9),
	.w7(32'hbbbd5370),
	.w8(32'hbb7f0b97),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2cb55),
	.w1(32'hbbdf71b9),
	.w2(32'hbb073e87),
	.w3(32'h3b06eac8),
	.w4(32'hbbce3c02),
	.w5(32'hba8428ef),
	.w6(32'h3b0463b9),
	.w7(32'hbad90392),
	.w8(32'hbbfe3346),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d2ac8),
	.w1(32'hbc51c57d),
	.w2(32'hbb8013ab),
	.w3(32'hb99f5373),
	.w4(32'hbc7eabc0),
	.w5(32'hbb98424b),
	.w6(32'hbbe8ae9c),
	.w7(32'hbc954ee1),
	.w8(32'hbb9044e4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f11ae8),
	.w1(32'hb95e97f5),
	.w2(32'h3b4feb7b),
	.w3(32'h3a955984),
	.w4(32'h3af2d01c),
	.w5(32'hbba24ba0),
	.w6(32'hba03b54f),
	.w7(32'h3aef74c9),
	.w8(32'hba767128),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c624dd1),
	.w1(32'h3c816d44),
	.w2(32'hbb8b1a04),
	.w3(32'h3a7e3ad2),
	.w4(32'hbb601ab0),
	.w5(32'h3c397da2),
	.w6(32'h3b859edb),
	.w7(32'hbc294717),
	.w8(32'h3b3a8474),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cd5c9),
	.w1(32'h3bd0dbb5),
	.w2(32'hbc01b24a),
	.w3(32'hbc1dfb76),
	.w4(32'hbbcc91ef),
	.w5(32'hbcaaa655),
	.w6(32'hbbc87541),
	.w7(32'hbbb2b1d0),
	.w8(32'hbbdd9fbb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97bf15),
	.w1(32'h3b0ef60e),
	.w2(32'h3bb3a41a),
	.w3(32'hbb202523),
	.w4(32'hba6705b2),
	.w5(32'hbbcd8132),
	.w6(32'hbb2d1274),
	.w7(32'hba9eea1d),
	.w8(32'hba84f2df),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b793b53),
	.w1(32'h3a90e3be),
	.w2(32'hbad70f78),
	.w3(32'hb7d22669),
	.w4(32'hba6d74a9),
	.w5(32'h39418300),
	.w6(32'hbb6f01f8),
	.w7(32'hbb32c7c1),
	.w8(32'h3b4d9eab),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2c689),
	.w1(32'hbac6cd52),
	.w2(32'hbb872ef2),
	.w3(32'hbb13ddc2),
	.w4(32'hbba059da),
	.w5(32'hbb380a31),
	.w6(32'hbb118b9e),
	.w7(32'hbb33fb30),
	.w8(32'h39a54b49),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b1c99),
	.w1(32'hbb1fd276),
	.w2(32'hbb3fad11),
	.w3(32'hbb699079),
	.w4(32'hbb91620e),
	.w5(32'hbb1274e6),
	.w6(32'hbb96b742),
	.w7(32'hbac98937),
	.w8(32'h3a875985),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab75487),
	.w1(32'hbbf00985),
	.w2(32'hbba932cd),
	.w3(32'hbab00518),
	.w4(32'hbb6c261d),
	.w5(32'hbaa624d8),
	.w6(32'hbbcbe924),
	.w7(32'hbbbe9b8a),
	.w8(32'hbb98b083),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe92e0),
	.w1(32'hbbc8144f),
	.w2(32'hbbc35705),
	.w3(32'hbb5258f9),
	.w4(32'hba86130e),
	.w5(32'hba21dff4),
	.w6(32'hbb23cad3),
	.w7(32'hbbbf89ed),
	.w8(32'h38e19c14),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b417614),
	.w1(32'h3af875bc),
	.w2(32'h3b34af98),
	.w3(32'hbb2f1d5b),
	.w4(32'hbbc3ca9c),
	.w5(32'hbba0dcdb),
	.w6(32'h3a930c0a),
	.w7(32'hbbd41ec1),
	.w8(32'hbb163d1f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8646be),
	.w1(32'hbb228aaa),
	.w2(32'hbb85a28a),
	.w3(32'hbb238e41),
	.w4(32'hbaecd7a1),
	.w5(32'h3b9f0321),
	.w6(32'hbb285e46),
	.w7(32'hbba2788f),
	.w8(32'h3b1c696a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081636),
	.w1(32'h3c611ade),
	.w2(32'h3bf8adf6),
	.w3(32'h3c1b9032),
	.w4(32'h3b6136ec),
	.w5(32'h3b1788f4),
	.w6(32'h3c20edc1),
	.w7(32'hbae936cb),
	.w8(32'h39cc5c6d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5159),
	.w1(32'hb904b9de),
	.w2(32'h3a0bcfe0),
	.w3(32'h3b5c9cfa),
	.w4(32'hbb3d00f6),
	.w5(32'hbba9363a),
	.w6(32'h3b475480),
	.w7(32'hbb5ff59f),
	.w8(32'h3b00441f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ad53b),
	.w1(32'hb9d9bd3f),
	.w2(32'hbc3850b4),
	.w3(32'hbb8de1fe),
	.w4(32'h3a671719),
	.w5(32'hbbca28fa),
	.w6(32'hbbab4fed),
	.w7(32'hbbbe6327),
	.w8(32'hb9049bb6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaf5d7),
	.w1(32'h39c94a86),
	.w2(32'h3b7fec35),
	.w3(32'h3a90041f),
	.w4(32'h38f55560),
	.w5(32'h3bfa298a),
	.w6(32'hbaf2641e),
	.w7(32'hb9cff913),
	.w8(32'h3ba3aa89),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19180b),
	.w1(32'h3c042fc6),
	.w2(32'h3ba83c7f),
	.w3(32'hbb62d27f),
	.w4(32'h3adbcbcc),
	.w5(32'hba177d2f),
	.w6(32'h3adb0748),
	.w7(32'h3b3182ce),
	.w8(32'hbbc10dc5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb17b4),
	.w1(32'h3899e95b),
	.w2(32'h3b3e3323),
	.w3(32'hbadd9c69),
	.w4(32'h3b978eac),
	.w5(32'h3b4a8ad5),
	.w6(32'hbbcc0e9e),
	.w7(32'hbb163fba),
	.w8(32'hba5bbaff),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40341b),
	.w1(32'hbb7b4c30),
	.w2(32'hbbc870df),
	.w3(32'hbbd471af),
	.w4(32'hbbc8f349),
	.w5(32'hbc4d8792),
	.w6(32'hbbb443f0),
	.w7(32'hbbc39598),
	.w8(32'hbc096271),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85e7bb),
	.w1(32'hbb558065),
	.w2(32'hbad88f39),
	.w3(32'hbb4f2d57),
	.w4(32'hbb335696),
	.w5(32'hbb943a62),
	.w6(32'hbba3400f),
	.w7(32'hbbb8f0fc),
	.w8(32'hbbf6a522),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1103e),
	.w1(32'hbab34dad),
	.w2(32'hbaa9df4d),
	.w3(32'hb9edabec),
	.w4(32'hbaaeab49),
	.w5(32'h3a85dc5e),
	.w6(32'h3ac84d38),
	.w7(32'hba9f40be),
	.w8(32'hba230273),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc167ef),
	.w1(32'hb7218fb3),
	.w2(32'hbb7fa33f),
	.w3(32'hbbf9cbab),
	.w4(32'hbbc740b3),
	.w5(32'hbc08989b),
	.w6(32'hbbbe2c1a),
	.w7(32'hbbda3b5d),
	.w8(32'hbc56175f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713e41),
	.w1(32'h3bbcaab3),
	.w2(32'h3c16fb26),
	.w3(32'hbb233252),
	.w4(32'h3bce390e),
	.w5(32'h3c1ff62b),
	.w6(32'hbc024b28),
	.w7(32'hb9831a90),
	.w8(32'h3c4069e9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f9d9d),
	.w1(32'h3be02d31),
	.w2(32'hb89bd63c),
	.w3(32'h3c107c52),
	.w4(32'h3b029303),
	.w5(32'h3aebc610),
	.w6(32'h3c4db7dc),
	.w7(32'hbb464ef9),
	.w8(32'hbbd064b6),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78a740),
	.w1(32'h3a8e8416),
	.w2(32'h3b304313),
	.w3(32'h3acaab2e),
	.w4(32'h3a92b4fc),
	.w5(32'hbafe8aa1),
	.w6(32'hbb3b88d7),
	.w7(32'h380e75bb),
	.w8(32'hb942e7aa),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80cefa),
	.w1(32'h3acd93ed),
	.w2(32'hba9d9f28),
	.w3(32'hbb5b3504),
	.w4(32'hbab36817),
	.w5(32'hbbcc29ed),
	.w6(32'hbb757c0f),
	.w7(32'hba96cad5),
	.w8(32'hbb09b505),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bfc54),
	.w1(32'hbbe3990a),
	.w2(32'hbb7aa094),
	.w3(32'h399acc4a),
	.w4(32'hbbf5a171),
	.w5(32'h3c09840d),
	.w6(32'hbba7e8dd),
	.w7(32'hbcc4e6be),
	.w8(32'hbc4d6ba5),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37302f),
	.w1(32'hba62271f),
	.w2(32'h3b2f6312),
	.w3(32'hb9d04420),
	.w4(32'hbba27f8a),
	.w5(32'hb9451efe),
	.w6(32'hbbd34a4b),
	.w7(32'hbc1505c9),
	.w8(32'hbc05a56e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb209d2),
	.w1(32'h3b248550),
	.w2(32'h3b6f2f08),
	.w3(32'hbba674ce),
	.w4(32'hbbc6044e),
	.w5(32'hbb0533c2),
	.w6(32'hbc46ebfa),
	.w7(32'hbc34c1dc),
	.w8(32'hbc30e604),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02b863),
	.w1(32'hbc27688f),
	.w2(32'hbc2bce03),
	.w3(32'h3b1c6ad5),
	.w4(32'hbc783a70),
	.w5(32'hbcd8d9f9),
	.w6(32'hbc1dd7b7),
	.w7(32'hbc2294f1),
	.w8(32'hb9c8aa0f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78d3d),
	.w1(32'h3b88967c),
	.w2(32'h3abce676),
	.w3(32'hbb91ae29),
	.w4(32'hbb22e238),
	.w5(32'h3abb0d62),
	.w6(32'hbbc4e6d8),
	.w7(32'hbb1d7153),
	.w8(32'hbae2508c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620e18),
	.w1(32'hba5875fb),
	.w2(32'h3bce743d),
	.w3(32'hba506746),
	.w4(32'h3b3f7791),
	.w5(32'h3baa8b9e),
	.w6(32'hbb963375),
	.w7(32'h3931cc9e),
	.w8(32'h3b3eeea6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18af57),
	.w1(32'hbc97fc10),
	.w2(32'h3a14da31),
	.w3(32'h3c974ff5),
	.w4(32'hbbb29cd2),
	.w5(32'h3c2b9a88),
	.w6(32'h39a618ae),
	.w7(32'hbbbaf689),
	.w8(32'hbb285f54),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40b717),
	.w1(32'h3c2d4cce),
	.w2(32'h3bd24292),
	.w3(32'h3bbb1b0e),
	.w4(32'h3b8d4d13),
	.w5(32'hbb9bd341),
	.w6(32'h3a8edf4e),
	.w7(32'hbbbc3077),
	.w8(32'hbc076eea),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8b2e),
	.w1(32'hbc83e45e),
	.w2(32'hbba31976),
	.w3(32'h3baeb497),
	.w4(32'hbc972082),
	.w5(32'hbb66eb25),
	.w6(32'hb91f04da),
	.w7(32'hbca49975),
	.w8(32'hbc134ab9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceaf36),
	.w1(32'hbc471b81),
	.w2(32'hbc098d48),
	.w3(32'hbba084eb),
	.w4(32'hbbd37127),
	.w5(32'hbc160ac1),
	.w6(32'hbc2765b3),
	.w7(32'hbba335cf),
	.w8(32'hbbf63d31),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadfe1d),
	.w1(32'hbc26d599),
	.w2(32'hbc3e6901),
	.w3(32'hbc1cbb21),
	.w4(32'hbc26980e),
	.w5(32'hbc1917ba),
	.w6(32'hbb45618c),
	.w7(32'hbbaf41f3),
	.w8(32'hbb5b4e4a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf892f1),
	.w1(32'h3a9be059),
	.w2(32'h3b0c4848),
	.w3(32'hbab88245),
	.w4(32'h3b97890e),
	.w5(32'h3b03bc37),
	.w6(32'hbb9c7abb),
	.w7(32'h3b02a7e5),
	.w8(32'h3b007445),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd864b),
	.w1(32'hba5d10f8),
	.w2(32'hba8194e4),
	.w3(32'h3b523df4),
	.w4(32'h3b4d0b78),
	.w5(32'h3bb0544b),
	.w6(32'h39436718),
	.w7(32'hbb1f9850),
	.w8(32'h3bbe2c52),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11a3ab),
	.w1(32'h3bff8f42),
	.w2(32'h39cd42f0),
	.w3(32'h3c05b1ce),
	.w4(32'h3b23a137),
	.w5(32'hbae85171),
	.w6(32'h3b9bd3f2),
	.w7(32'hbb90b819),
	.w8(32'hbaa0f7eb),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b92e),
	.w1(32'hbb36f913),
	.w2(32'hbb8c05e2),
	.w3(32'hbb4311bc),
	.w4(32'hbb58d000),
	.w5(32'hb8a0a594),
	.w6(32'hbb1be569),
	.w7(32'hbaf50bcf),
	.w8(32'hbab7ba90),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba157585),
	.w1(32'hbb95fac5),
	.w2(32'h3a139276),
	.w3(32'hb8802913),
	.w4(32'h3aa5a57f),
	.w5(32'h3b2aea2b),
	.w6(32'hbb9fc142),
	.w7(32'hbb00874b),
	.w8(32'hba459302),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b8e38),
	.w1(32'h3b7e9c65),
	.w2(32'h3bd021b4),
	.w3(32'hbbbc5b10),
	.w4(32'hbbc3caac),
	.w5(32'h3bba0590),
	.w6(32'hbbf9f86e),
	.w7(32'hbb9828f1),
	.w8(32'hbb1d797c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72729d),
	.w1(32'h39d5a1b8),
	.w2(32'h3bc56948),
	.w3(32'hbb8e0e75),
	.w4(32'hb89e312f),
	.w5(32'hbad12816),
	.w6(32'hbbeeec32),
	.w7(32'hbb877f84),
	.w8(32'hbaea2254),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20bd9f),
	.w1(32'h39c0821c),
	.w2(32'hba72a3f1),
	.w3(32'hbadb2764),
	.w4(32'hbac869c2),
	.w5(32'h3a21f0a9),
	.w6(32'hba84e086),
	.w7(32'h3b039caa),
	.w8(32'hb7191fe9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3097d5),
	.w1(32'hbc5f039b),
	.w2(32'h3b84b575),
	.w3(32'h3c81cf1c),
	.w4(32'hbc80af1c),
	.w5(32'hbbd7d9b0),
	.w6(32'h3b405e38),
	.w7(32'hbca8d1fb),
	.w8(32'hbc068927),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afda0b9),
	.w1(32'h3ade910f),
	.w2(32'h3acef22d),
	.w3(32'hbb7a9834),
	.w4(32'hbb6624c7),
	.w5(32'h3babea90),
	.w6(32'hbb9b0ffb),
	.w7(32'hbad56d38),
	.w8(32'hbb1fa24e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4a3b4),
	.w1(32'hbba4eed3),
	.w2(32'hbb2a96e1),
	.w3(32'h3a23b800),
	.w4(32'hba539d70),
	.w5(32'hba020f2a),
	.w6(32'hbc03f9cf),
	.w7(32'hbbada7ef),
	.w8(32'h3b054a74),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b053694),
	.w1(32'h3acda529),
	.w2(32'h3a97058e),
	.w3(32'h3b361329),
	.w4(32'h3aca0a32),
	.w5(32'hba9a31ff),
	.w6(32'hbafb2a68),
	.w7(32'hb9a3d56b),
	.w8(32'h3a17d989),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642b22),
	.w1(32'hbb2c9fae),
	.w2(32'hbb347452),
	.w3(32'hbb342bb6),
	.w4(32'hbbc8352b),
	.w5(32'h3b4bdafe),
	.w6(32'h3a9b13de),
	.w7(32'h39dac0e4),
	.w8(32'h3ac848ea),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b325315),
	.w1(32'h3bfe86d3),
	.w2(32'h3bf3c785),
	.w3(32'h3b8b7be8),
	.w4(32'h3aa83972),
	.w5(32'h38cb4236),
	.w6(32'h3b745455),
	.w7(32'h3a864d58),
	.w8(32'h39bdb9d3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3eb9c),
	.w1(32'h3b17e9a7),
	.w2(32'h3b7210fb),
	.w3(32'hbb039016),
	.w4(32'h373789b2),
	.w5(32'h39c6b696),
	.w6(32'hbb246c59),
	.w7(32'h39ea084e),
	.w8(32'h3b8a3179),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f1de9),
	.w1(32'h3a401571),
	.w2(32'h3bb7c05e),
	.w3(32'hbaad7208),
	.w4(32'hbb2067d0),
	.w5(32'hbad09ef7),
	.w6(32'h3ac97bdc),
	.w7(32'h3b8245ed),
	.w8(32'hbb5a260a),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96c953),
	.w1(32'hbbd5ca22),
	.w2(32'hbbf311e5),
	.w3(32'hb8c15648),
	.w4(32'hbba55507),
	.w5(32'hbb762619),
	.w6(32'hb8bda1ff),
	.w7(32'hba9b27ce),
	.w8(32'hbbc44f0c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba992a0),
	.w1(32'h3af604e7),
	.w2(32'h3b84a7cf),
	.w3(32'hbbd0fd0f),
	.w4(32'hbbaa7641),
	.w5(32'hbba63ff2),
	.w6(32'hbbfce12e),
	.w7(32'hbb024671),
	.w8(32'h3ae5c162),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995e36),
	.w1(32'h3b49768e),
	.w2(32'h3ba85cc4),
	.w3(32'hbaf05e02),
	.w4(32'hb9c0d42a),
	.w5(32'h3b37548c),
	.w6(32'hbaa37ea0),
	.w7(32'hbb44de70),
	.w8(32'h3ab108e0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b809238),
	.w1(32'h3c07f73b),
	.w2(32'h3b7d0f51),
	.w3(32'hb8eba6bb),
	.w4(32'h3b013580),
	.w5(32'hbae9f825),
	.w6(32'hba5e1a4a),
	.w7(32'hb94ecdd5),
	.w8(32'h3aaaebcf),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db21b),
	.w1(32'hbab793a0),
	.w2(32'hbba81ae4),
	.w3(32'hbb8dec4c),
	.w4(32'hba7ce0e3),
	.w5(32'h3acd4b6c),
	.w6(32'hbb757da7),
	.w7(32'hbbbdcb76),
	.w8(32'hba9925af),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a69c2),
	.w1(32'hbb6592ce),
	.w2(32'hbb1b4fee),
	.w3(32'hba99567c),
	.w4(32'hbad01267),
	.w5(32'h3bb35de6),
	.w6(32'hbb18a367),
	.w7(32'hbabecb75),
	.w8(32'h3b781591),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c035be7),
	.w1(32'h3c037aa2),
	.w2(32'h3be81169),
	.w3(32'h3b944a43),
	.w4(32'h3be48aed),
	.w5(32'h3b9c1316),
	.w6(32'h3a810f95),
	.w7(32'h3b09669d),
	.w8(32'hbb2ce06a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b667),
	.w1(32'hbb702e48),
	.w2(32'hbb88df29),
	.w3(32'h3b5c9a10),
	.w4(32'h3a250f46),
	.w5(32'hbb2c0539),
	.w6(32'hbae30b22),
	.w7(32'hbaa387e4),
	.w8(32'hbb875699),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33a395),
	.w1(32'h3b7e19c7),
	.w2(32'h3bcba7e2),
	.w3(32'hbbda7d51),
	.w4(32'h3b94d71e),
	.w5(32'h3c24e8e3),
	.w6(32'hbc2d2286),
	.w7(32'hbb2ca065),
	.w8(32'h3b2d8e40),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1410f0),
	.w1(32'hbb4873ca),
	.w2(32'h3b0d7342),
	.w3(32'h3b2a8f7e),
	.w4(32'h3b815b78),
	.w5(32'h39166d08),
	.w6(32'hbbc6d3bf),
	.w7(32'h38fe5678),
	.w8(32'h39b512be),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15055b),
	.w1(32'hb9d5ab70),
	.w2(32'hbb0bd985),
	.w3(32'hbb15df35),
	.w4(32'hbb34e03e),
	.w5(32'hbb0544ec),
	.w6(32'h3ac30423),
	.w7(32'h3a75e04a),
	.w8(32'hba81c3e4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39313440),
	.w1(32'h39250889),
	.w2(32'hbb383be7),
	.w3(32'h3b858d26),
	.w4(32'h3b0e08a1),
	.w5(32'hbb93baf0),
	.w6(32'h3b0be32e),
	.w7(32'h3af5691a),
	.w8(32'h3bb79608),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae14d79),
	.w1(32'hba9ef691),
	.w2(32'hb98fffcf),
	.w3(32'hbba1629d),
	.w4(32'hbc22be50),
	.w5(32'h37453bec),
	.w6(32'h3baa89c2),
	.w7(32'h3a508a7c),
	.w8(32'h3b82df2a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa247e4),
	.w1(32'h3aaa57c7),
	.w2(32'hba27836d),
	.w3(32'h3a3df498),
	.w4(32'hbb1e5d9b),
	.w5(32'h3b39d352),
	.w6(32'h3b2b6354),
	.w7(32'hbab6871f),
	.w8(32'hb9892c37),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1525a3),
	.w1(32'h3b91f6ee),
	.w2(32'h3b37d6f4),
	.w3(32'h3a9826a9),
	.w4(32'hbb154db8),
	.w5(32'hbb431c75),
	.w6(32'hbaef6325),
	.w7(32'hbb705c79),
	.w8(32'hbb120b57),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4196d3),
	.w1(32'h3c8f6d5a),
	.w2(32'h3c6a0c4d),
	.w3(32'hbc25db03),
	.w4(32'h3c3ead0e),
	.w5(32'h3c225aa4),
	.w6(32'hbc420fb1),
	.w7(32'h3bc8bcc7),
	.w8(32'h3b583c06),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a7083),
	.w1(32'h3b2d49ed),
	.w2(32'h3a88293f),
	.w3(32'h3a8eee45),
	.w4(32'h3a9fb3df),
	.w5(32'h3b07be37),
	.w6(32'hba887dbc),
	.w7(32'hbb1154a3),
	.w8(32'h39cbfc4e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38c39),
	.w1(32'hbbc1d507),
	.w2(32'hbb45e449),
	.w3(32'h39b67725),
	.w4(32'hbb591f35),
	.w5(32'hbc0c9de9),
	.w6(32'hbc079452),
	.w7(32'hbc850e07),
	.w8(32'hbc80821a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule