module layer_10_featuremap_21(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b209a8f),
	.w1(32'hbbc8dee1),
	.w2(32'h3b912030),
	.w3(32'hbb305320),
	.w4(32'hbc8775e1),
	.w5(32'hbb0d7a21),
	.w6(32'hb9d7202c),
	.w7(32'hbc3f6c6a),
	.w8(32'h3bc07f1f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70ddbe),
	.w1(32'h3c1e1d39),
	.w2(32'hbc044637),
	.w3(32'hba2796c4),
	.w4(32'hbc175ae7),
	.w5(32'h3c126d15),
	.w6(32'h3af26084),
	.w7(32'hbb286419),
	.w8(32'hbabcb616),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8532d0),
	.w1(32'hbb7e9d48),
	.w2(32'hbb427472),
	.w3(32'h3c4b91af),
	.w4(32'h3c1f90e6),
	.w5(32'hbbbd0353),
	.w6(32'h3b70b634),
	.w7(32'h3b1bf42b),
	.w8(32'hbb47936f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4bcb0),
	.w1(32'hbb0c4588),
	.w2(32'hbcb7eddd),
	.w3(32'hbc288925),
	.w4(32'h3adc7018),
	.w5(32'hbbd135e0),
	.w6(32'hbb03a11a),
	.w7(32'hbb0c4fe2),
	.w8(32'hbbb32209),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc766c8),
	.w1(32'hbca460d1),
	.w2(32'hbb2c3ae0),
	.w3(32'h3a5e7e1d),
	.w4(32'hbbbf5ac9),
	.w5(32'h3b8d8810),
	.w6(32'hbacb5f2f),
	.w7(32'h389c9749),
	.w8(32'h3b79e2fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf92b19),
	.w1(32'hbb7982cc),
	.w2(32'hbb9ffc54),
	.w3(32'hbb8e98ae),
	.w4(32'hbb942d51),
	.w5(32'hba929f6b),
	.w6(32'hbc2166ca),
	.w7(32'hbaadd484),
	.w8(32'hbb247613),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776863),
	.w1(32'hbba0678b),
	.w2(32'hbcca2e53),
	.w3(32'h3a56b42c),
	.w4(32'h3b4d2421),
	.w5(32'hbc53fe51),
	.w6(32'h3a459914),
	.w7(32'hbc114300),
	.w8(32'hbc487267),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860027),
	.w1(32'hbb88f2ae),
	.w2(32'h3c3f8da5),
	.w3(32'hbbe383c9),
	.w4(32'hbb2224c9),
	.w5(32'h3bdf3b91),
	.w6(32'h3aa44ca8),
	.w7(32'hbb0fcaf9),
	.w8(32'hbb60351a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1cfed),
	.w1(32'h3c1adc73),
	.w2(32'hbb8ce252),
	.w3(32'h3a27058b),
	.w4(32'hbb600f39),
	.w5(32'h389b865c),
	.w6(32'hbc1fdea7),
	.w7(32'hbc3bbd78),
	.w8(32'h3b3114b3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb687297),
	.w1(32'hbbc8edab),
	.w2(32'hbb5c23d3),
	.w3(32'h3b545866),
	.w4(32'h3b57a3a9),
	.w5(32'hbaf652cb),
	.w6(32'h3bf4dfdf),
	.w7(32'h3c006952),
	.w8(32'hbb725b39),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3215b),
	.w1(32'hb8092559),
	.w2(32'h3bc6574d),
	.w3(32'hbafa3b7d),
	.w4(32'hbb36b8d8),
	.w5(32'h3b0c3feb),
	.w6(32'hbb74eba7),
	.w7(32'hbb5aa8c8),
	.w8(32'h3a556ff5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6136a),
	.w1(32'hbb7a1092),
	.w2(32'hbc1a8fa9),
	.w3(32'h3ba74d25),
	.w4(32'h3b835c48),
	.w5(32'hbbca954e),
	.w6(32'hbb716714),
	.w7(32'hbbc4b88e),
	.w8(32'hbbbf5ac8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac457df),
	.w1(32'hba03666e),
	.w2(32'hbc0f6505),
	.w3(32'hbb6729ca),
	.w4(32'hbae2b23e),
	.w5(32'hbb0c839b),
	.w6(32'hbba94027),
	.w7(32'hbba03929),
	.w8(32'hbb8d1917),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d738a),
	.w1(32'hbb1bf3d8),
	.w2(32'h3c83c09a),
	.w3(32'hbc1d73b9),
	.w4(32'h3a14e5f1),
	.w5(32'hbc5758af),
	.w6(32'hbb882502),
	.w7(32'hbb2b80a1),
	.w8(32'hbc7de235),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf9172),
	.w1(32'h3c6e280a),
	.w2(32'hbc9aeeca),
	.w3(32'hbc6de54f),
	.w4(32'hbb9f0057),
	.w5(32'hba665b9a),
	.w6(32'hbc9c0593),
	.w7(32'hbc5681e1),
	.w8(32'h3c47ca10),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd066bfc),
	.w1(32'hbcdc764a),
	.w2(32'h3894065f),
	.w3(32'hbc63306d),
	.w4(32'hbc04c648),
	.w5(32'h3ab87bce),
	.w6(32'h3c48124f),
	.w7(32'h3b777477),
	.w8(32'h3b7fa24d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2275de),
	.w1(32'hbab27823),
	.w2(32'h3b845c62),
	.w3(32'h38e607ed),
	.w4(32'hba976812),
	.w5(32'hbb616482),
	.w6(32'h39cb3544),
	.w7(32'hb8cc7d1a),
	.w8(32'hbc52db97),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6b6c6),
	.w1(32'h3ae7b621),
	.w2(32'h3b489f16),
	.w3(32'hbb9b057d),
	.w4(32'hbaf49e36),
	.w5(32'h3bb230b8),
	.w6(32'hbc8567ff),
	.w7(32'hbc9d7684),
	.w8(32'h3ab17bcb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92dc28),
	.w1(32'hbb94b8c9),
	.w2(32'hbbdd9321),
	.w3(32'hbb035a6c),
	.w4(32'hbb13d6ea),
	.w5(32'hbb5c89ba),
	.w6(32'hbb9f921e),
	.w7(32'hbbb5d8c7),
	.w8(32'hbbd58029),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29a92f),
	.w1(32'h3bf327be),
	.w2(32'h3c679a38),
	.w3(32'hbbc1a561),
	.w4(32'hbb10921e),
	.w5(32'h3c1b404e),
	.w6(32'hbc5708f0),
	.w7(32'hbc5ba5e4),
	.w8(32'h388084a7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c429bed),
	.w1(32'h3c16c032),
	.w2(32'hbb34fcbe),
	.w3(32'h3a3a8526),
	.w4(32'hbbbecc94),
	.w5(32'h3ab4f42d),
	.w6(32'hbb879699),
	.w7(32'hbb8e1c32),
	.w8(32'hbbd9f909),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6082fe),
	.w1(32'h38ce0a74),
	.w2(32'hbc6899b1),
	.w3(32'hbbe66be1),
	.w4(32'hbbbc5eaf),
	.w5(32'h3b2bfa75),
	.w6(32'hbc3e35e7),
	.w7(32'hbc25e648),
	.w8(32'h3c36b38a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9850a0),
	.w1(32'hbc14241f),
	.w2(32'h3b19a944),
	.w3(32'h3b8878a7),
	.w4(32'h3b797e07),
	.w5(32'h3ba71837),
	.w6(32'h3c14022d),
	.w7(32'h3b9b9f9a),
	.w8(32'hbb02d4c6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76b8ae),
	.w1(32'h3b928d90),
	.w2(32'h3b8ef943),
	.w3(32'h3b63a1c7),
	.w4(32'h3beeb050),
	.w5(32'hbb600f73),
	.w6(32'hba1ea78f),
	.w7(32'h3b3db667),
	.w8(32'hba99b18a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb396c9),
	.w1(32'h3adefd41),
	.w2(32'hbaf891f0),
	.w3(32'hbb9d1bf3),
	.w4(32'h3938d4f5),
	.w5(32'hbc2ca8ec),
	.w6(32'h3a5196af),
	.w7(32'hba553ebf),
	.w8(32'hbc679d70),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb922c88),
	.w1(32'hb9375f68),
	.w2(32'h3bb75d33),
	.w3(32'hbbe98cbb),
	.w4(32'hbc3372e4),
	.w5(32'h3a0abdff),
	.w6(32'hbc8a3e5e),
	.w7(32'hbc5556e9),
	.w8(32'hbc20fd8c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d8f9a),
	.w1(32'h3c05cea0),
	.w2(32'h3a9660c2),
	.w3(32'h3a92a507),
	.w4(32'h3b43f839),
	.w5(32'hba81a1f5),
	.w6(32'hbb596e80),
	.w7(32'hbae54282),
	.w8(32'h3a8a2f27),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6edb),
	.w1(32'h3bacb227),
	.w2(32'hbc2e796f),
	.w3(32'hba04ed84),
	.w4(32'h3a77eb20),
	.w5(32'h3b3abc97),
	.w6(32'h3b2bcace),
	.w7(32'h3bfc08d1),
	.w8(32'h3c4f53ab),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e574),
	.w1(32'hbc888ce3),
	.w2(32'h3c213fb2),
	.w3(32'hbb033ce7),
	.w4(32'hbb664f55),
	.w5(32'h3b98100d),
	.w6(32'hba02638a),
	.w7(32'hbbda8bce),
	.w8(32'h3ab4bd28),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50064f),
	.w1(32'hbb3e9b1d),
	.w2(32'h3b812160),
	.w3(32'hbb838085),
	.w4(32'hbb947825),
	.w5(32'h390ff1e5),
	.w6(32'hba323fb8),
	.w7(32'h3b2c8b89),
	.w8(32'hb9ecc46f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05c95b),
	.w1(32'hbb89b5e2),
	.w2(32'h3a1fd6b5),
	.w3(32'hbb60741f),
	.w4(32'hbb5a2b54),
	.w5(32'h3b53d661),
	.w6(32'h3aefe278),
	.w7(32'h3b0bf5d0),
	.w8(32'h3b06a4fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f139),
	.w1(32'hbb87f2af),
	.w2(32'hbae18baa),
	.w3(32'h3b40fd84),
	.w4(32'h3b900f6e),
	.w5(32'h3bd5f134),
	.w6(32'h3c5f3339),
	.w7(32'h3c08d0c6),
	.w8(32'h3c95782d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38213f),
	.w1(32'hbbad3255),
	.w2(32'hbbb69ead),
	.w3(32'h3c439bcf),
	.w4(32'h3bda0a4b),
	.w5(32'hbb3fc3b5),
	.w6(32'h3c4e4f7f),
	.w7(32'h3c264ce7),
	.w8(32'h3a9a6675),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49dfb6),
	.w1(32'hbbb157ad),
	.w2(32'h3b6cb1b2),
	.w3(32'hbbf4e763),
	.w4(32'hbbc67979),
	.w5(32'hbc1c890f),
	.w6(32'h38ed0062),
	.w7(32'h3b794afb),
	.w8(32'hbc212bab),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8612e1),
	.w1(32'hbc1f711f),
	.w2(32'hbb786992),
	.w3(32'hbbcbcea7),
	.w4(32'hbbd1f4bd),
	.w5(32'hbb647f61),
	.w6(32'hbbc98da9),
	.w7(32'hbb8d04e6),
	.w8(32'hbade26db),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8abec1),
	.w1(32'hba57d833),
	.w2(32'hbc181ef3),
	.w3(32'hbb263c1e),
	.w4(32'hbb25d1f0),
	.w5(32'h3bd3b0d4),
	.w6(32'hbbcb7b58),
	.w7(32'hbbb87ec6),
	.w8(32'hb9b385c7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c292975),
	.w1(32'hb8de6ea1),
	.w2(32'hbc63449f),
	.w3(32'h3b04f19e),
	.w4(32'hbb789580),
	.w5(32'hbb7492df),
	.w6(32'hbad1f6ff),
	.w7(32'h3b21200c),
	.w8(32'hbc0e7e09),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4adc),
	.w1(32'hbbc58d23),
	.w2(32'h3c379758),
	.w3(32'hbb87a33b),
	.w4(32'hbbb82321),
	.w5(32'h398cb592),
	.w6(32'hbaa60175),
	.w7(32'h3b820e99),
	.w8(32'hbc1c852f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14623d),
	.w1(32'h39b78149),
	.w2(32'hbc77eb09),
	.w3(32'hbc4c3046),
	.w4(32'hbc679641),
	.w5(32'hbbd5ff39),
	.w6(32'hbc3696f3),
	.w7(32'hbc8bd195),
	.w8(32'hb9a02a3f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce2c58),
	.w1(32'hbc0b836a),
	.w2(32'h3b9075ec),
	.w3(32'hbc08d369),
	.w4(32'h3b34b4fa),
	.w5(32'h3a4081f4),
	.w6(32'h3aa3564e),
	.w7(32'h3b9ccaca),
	.w8(32'hbc6ca799),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a712576),
	.w1(32'h3a761d95),
	.w2(32'h3be6c722),
	.w3(32'hbbdd2de8),
	.w4(32'hbb71d4d6),
	.w5(32'h3bccc62d),
	.w6(32'hbc8755fe),
	.w7(32'hbc3f85bd),
	.w8(32'h3c1d6439),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf415ea),
	.w1(32'hba81d20f),
	.w2(32'hbb961020),
	.w3(32'h3c4db958),
	.w4(32'h3b60affb),
	.w5(32'h3af97933),
	.w6(32'h3b659729),
	.w7(32'h3bac1644),
	.w8(32'h3ba0bb3d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95dda7),
	.w1(32'hbb1b83e9),
	.w2(32'hbc28276c),
	.w3(32'hba22fb13),
	.w4(32'h3bd09e95),
	.w5(32'hbb65cc79),
	.w6(32'h3bdfebc3),
	.w7(32'h3b05de27),
	.w8(32'hba758276),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dc3f3),
	.w1(32'hbca69792),
	.w2(32'h3a35635b),
	.w3(32'hbbd7a029),
	.w4(32'hbbf20755),
	.w5(32'h3b2d9fd0),
	.w6(32'hbb2c0e37),
	.w7(32'hbb7aaf65),
	.w8(32'hbbbe3ebb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2212d0),
	.w1(32'h3a4d7003),
	.w2(32'h3baa159e),
	.w3(32'hbb7c98a3),
	.w4(32'h3a9ebfc8),
	.w5(32'hbb4036a3),
	.w6(32'hbbbcf8f2),
	.w7(32'hbc8ac020),
	.w8(32'hbb7b2aad),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed17e2),
	.w1(32'h3b1f2bdb),
	.w2(32'h3b262437),
	.w3(32'hbbacb8f2),
	.w4(32'hbb30e50d),
	.w5(32'h3c0efab3),
	.w6(32'hbbdc5b5c),
	.w7(32'hbc48810f),
	.w8(32'hbb63378b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba747268),
	.w1(32'hbc138e10),
	.w2(32'hba94a4c7),
	.w3(32'hbb4190b7),
	.w4(32'hbbbaa734),
	.w5(32'h3c15c60c),
	.w6(32'hbb629425),
	.w7(32'hba1fb57d),
	.w8(32'hba030161),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22a57a),
	.w1(32'hbce59185),
	.w2(32'hbc3fa7e7),
	.w3(32'h3b41412a),
	.w4(32'h3c88738e),
	.w5(32'h3a8ddb14),
	.w6(32'h3b0816f6),
	.w7(32'h3c85c783),
	.w8(32'h3b333020),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc3627),
	.w1(32'hbbcd0650),
	.w2(32'hbb70df3e),
	.w3(32'h3b7e11e5),
	.w4(32'h3b9cabc5),
	.w5(32'hbc176112),
	.w6(32'h3ba7b538),
	.w7(32'h3b9a09a8),
	.w8(32'hbbeac58f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb1aa),
	.w1(32'hbb2c1db8),
	.w2(32'hbbb78a1d),
	.w3(32'hbbd2f214),
	.w4(32'hbb830261),
	.w5(32'hbad30059),
	.w6(32'hbc14625a),
	.w7(32'hbc99ef33),
	.w8(32'h3b263e4e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f17d58),
	.w1(32'h3a9c46b3),
	.w2(32'h3ab88578),
	.w3(32'hbaee7ac8),
	.w4(32'hba008bd7),
	.w5(32'h3bf77904),
	.w6(32'h3b5ba644),
	.w7(32'h3a77a48f),
	.w8(32'h3ca17e3b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba912f6c),
	.w1(32'hbc123185),
	.w2(32'h3a5487ed),
	.w3(32'h3c09286c),
	.w4(32'h3b780138),
	.w5(32'hbb002eb2),
	.w6(32'h3cd20363),
	.w7(32'h3c651f8a),
	.w8(32'h3b3371d7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8c060),
	.w1(32'h3a42cf5b),
	.w2(32'h3c1ff855),
	.w3(32'h37bf9a33),
	.w4(32'h3a71153c),
	.w5(32'hb9e89c29),
	.w6(32'h3ba041dc),
	.w7(32'hb9bc478e),
	.w8(32'h3af40e7c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6457e),
	.w1(32'h3c4d55bc),
	.w2(32'hbbd9f89e),
	.w3(32'h3c12cea3),
	.w4(32'h3bedbbf3),
	.w5(32'hbbf9a77b),
	.w6(32'h3cbb6815),
	.w7(32'h3c91f561),
	.w8(32'hbbbeb31f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ac61f),
	.w1(32'h3ba0e6a8),
	.w2(32'hbb2cf3dc),
	.w3(32'hbbad6141),
	.w4(32'h3c3c7412),
	.w5(32'hbb6032fe),
	.w6(32'hbbe90711),
	.w7(32'hbaccb1be),
	.w8(32'hbb48e517),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77bf6e),
	.w1(32'hbb20398e),
	.w2(32'h39bbb4bc),
	.w3(32'hbbf7b287),
	.w4(32'hbaca6dfc),
	.w5(32'hbb4bf475),
	.w6(32'hbbecdf4d),
	.w7(32'hbc03d014),
	.w8(32'h3b7f5e42),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1273a),
	.w1(32'hb99dbf46),
	.w2(32'hbcaa4627),
	.w3(32'hb9e8c0d5),
	.w4(32'hb80aa27e),
	.w5(32'hbba3ae10),
	.w6(32'hbbed38bf),
	.w7(32'hbaca6912),
	.w8(32'hbc719626),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4f66e),
	.w1(32'hbcdfd744),
	.w2(32'hbb2eb232),
	.w3(32'hbbddb65e),
	.w4(32'hbb145820),
	.w5(32'hbbaa785a),
	.w6(32'hbc958ad7),
	.w7(32'hbbb54484),
	.w8(32'h3c9ab30a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeedbfe),
	.w1(32'hbbdd581c),
	.w2(32'hbcbbe8bf),
	.w3(32'hbb6cc41a),
	.w4(32'hbb797459),
	.w5(32'hbca90146),
	.w6(32'h3cc63397),
	.w7(32'h3caebded),
	.w8(32'hbc9d8bd2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd055dd3),
	.w1(32'hbceebe0d),
	.w2(32'hbc620e16),
	.w3(32'hbcf68eb5),
	.w4(32'hbce84436),
	.w5(32'hbad7a0b7),
	.w6(32'hbccd2608),
	.w7(32'hbc983cb3),
	.w8(32'h3b5a298b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7bede),
	.w1(32'hbc91ca6c),
	.w2(32'hb975442d),
	.w3(32'h3abe0df9),
	.w4(32'h3b02e5e5),
	.w5(32'hbb9d64ae),
	.w6(32'h3c74d328),
	.w7(32'h3bf103ef),
	.w8(32'hbb22c056),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee7e26),
	.w1(32'hbc20c01d),
	.w2(32'hbbf61004),
	.w3(32'hbbff4636),
	.w4(32'hbae2a1e2),
	.w5(32'h3ac6166e),
	.w6(32'h3ac2d2a3),
	.w7(32'hbb903ce0),
	.w8(32'h3b908984),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb247631),
	.w1(32'hbb4bd046),
	.w2(32'h3b118ec2),
	.w3(32'hbab585ca),
	.w4(32'h39d38644),
	.w5(32'hbb88a4ff),
	.w6(32'hbb59cb94),
	.w7(32'h3b5cc056),
	.w8(32'h3b0aa371),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e68f0),
	.w1(32'hbaadc5c2),
	.w2(32'hbb78cc6c),
	.w3(32'hbb8f3845),
	.w4(32'hbb7d2470),
	.w5(32'h3b2e5ea4),
	.w6(32'h3afe6404),
	.w7(32'hb8b26947),
	.w8(32'hb8cb56e2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3986b97b),
	.w1(32'h3a893ec7),
	.w2(32'h3c847e75),
	.w3(32'h3b83ca65),
	.w4(32'h3bd2c13e),
	.w5(32'h3be6b0f0),
	.w6(32'h3c11ae38),
	.w7(32'hba87a594),
	.w8(32'h3c527c37),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb38945),
	.w1(32'h3c8b18cc),
	.w2(32'hbaa028e3),
	.w3(32'h3c3cd302),
	.w4(32'h3c155929),
	.w5(32'h3ae53000),
	.w6(32'h3cc0e1ef),
	.w7(32'h3cafa2f8),
	.w8(32'h3b8ddb2f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91b015),
	.w1(32'hbc952051),
	.w2(32'hbc3614a4),
	.w3(32'h39a5fbcf),
	.w4(32'hbbf37733),
	.w5(32'h39d00de1),
	.w6(32'h3bf12f74),
	.w7(32'h3ba337a8),
	.w8(32'h3c0ee2eb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500003),
	.w1(32'h3a2ffa94),
	.w2(32'h39ee2010),
	.w3(32'h3ad6a152),
	.w4(32'h3bed89bd),
	.w5(32'h3b06ae01),
	.w6(32'h3a8a6b12),
	.w7(32'h3a6f2156),
	.w8(32'h3b306257),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f0ff2),
	.w1(32'hbb9aec84),
	.w2(32'h3c0727a1),
	.w3(32'hbb56b6a7),
	.w4(32'h3b70c984),
	.w5(32'h3bcec77d),
	.w6(32'hbbf727e8),
	.w7(32'hba94a748),
	.w8(32'hbb200d4b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b8d8f),
	.w1(32'h3c83680b),
	.w2(32'h3b735580),
	.w3(32'h3bc3c1aa),
	.w4(32'h3ba500af),
	.w5(32'h3c3050d1),
	.w6(32'hbbea15e9),
	.w7(32'hbba12478),
	.w8(32'h3b55310f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc4aaab),
	.w1(32'hbc987771),
	.w2(32'hbbf6ac40),
	.w3(32'h3a8b286f),
	.w4(32'h3bc97ac4),
	.w5(32'hbb39ea81),
	.w6(32'h3ba0a084),
	.w7(32'h3a67aa33),
	.w8(32'h3abb6b95),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb529cb4),
	.w1(32'hbb1950a3),
	.w2(32'hba5aff37),
	.w3(32'hbb1884b7),
	.w4(32'h3b55aa22),
	.w5(32'hbaa9e0fa),
	.w6(32'h3b61b2ef),
	.w7(32'h3c1dd427),
	.w8(32'hbae5c60c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab54ef),
	.w1(32'hbbd5fa54),
	.w2(32'h3a21f74f),
	.w3(32'h3bed3de6),
	.w4(32'hba310f78),
	.w5(32'h39e0f693),
	.w6(32'h3a8ab230),
	.w7(32'h3b821186),
	.w8(32'hbb9c9722),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc47bf8),
	.w1(32'hbbdd5013),
	.w2(32'hbabdbca8),
	.w3(32'hba0a003b),
	.w4(32'h39b0e3fb),
	.w5(32'h3651d640),
	.w6(32'h3b54df88),
	.w7(32'hbaabea94),
	.w8(32'hba232f9b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aa88c),
	.w1(32'hbbb671a0),
	.w2(32'hbc477f01),
	.w3(32'hbb6d71ef),
	.w4(32'hbb21b97e),
	.w5(32'hbb222441),
	.w6(32'hbbe03920),
	.w7(32'hbb85de94),
	.w8(32'h39f8f3e3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7488d4),
	.w1(32'hbc894d2d),
	.w2(32'hbbd651da),
	.w3(32'hbb8263e2),
	.w4(32'hbb65a4c0),
	.w5(32'h3b6239e2),
	.w6(32'hb98e9f1a),
	.w7(32'h3b175cde),
	.w8(32'h3b461f50),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3f22f),
	.w1(32'hbc205625),
	.w2(32'hbc0471b4),
	.w3(32'h3b5ec111),
	.w4(32'hb8cd3177),
	.w5(32'h3b4d520c),
	.w6(32'h3bf86d4d),
	.w7(32'h3bafebd1),
	.w8(32'hba00828c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90df1b),
	.w1(32'h39aa2771),
	.w2(32'h3a75196e),
	.w3(32'hbc28060f),
	.w4(32'hbbe34559),
	.w5(32'hbb7a4d85),
	.w6(32'hbb46ed0b),
	.w7(32'h390d47d5),
	.w8(32'hbc02e9b0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb091491),
	.w1(32'hbb0c15fd),
	.w2(32'hb971e01a),
	.w3(32'hbb3cc934),
	.w4(32'h3c169f64),
	.w5(32'h3b029e38),
	.w6(32'hbb990a8d),
	.w7(32'h3b4bfe85),
	.w8(32'h3a8627d5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c440ab2),
	.w1(32'hbb8f79b5),
	.w2(32'hbc0a0b37),
	.w3(32'h3bb8c362),
	.w4(32'hbb816b10),
	.w5(32'h3bd404e7),
	.w6(32'h3b0f4a6e),
	.w7(32'h3b18037b),
	.w8(32'hba981dab),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d3f2),
	.w1(32'hbc2a0753),
	.w2(32'hbaffd2fa),
	.w3(32'h3ba98a54),
	.w4(32'h3c254bf9),
	.w5(32'h3b4e7745),
	.w6(32'hbb2b49b7),
	.w7(32'h3b98f5a8),
	.w8(32'h3ba310e5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea8c57),
	.w1(32'hbbdb0b66),
	.w2(32'h3b5b0531),
	.w3(32'hbb353ed1),
	.w4(32'hbb85ce8f),
	.w5(32'h3bc3d38b),
	.w6(32'h3b28d7c1),
	.w7(32'hba85dabc),
	.w8(32'h3bbfe7a0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7589dd),
	.w1(32'h3b0078de),
	.w2(32'hbb3f409e),
	.w3(32'h3aa685dd),
	.w4(32'hba9953db),
	.w5(32'hbb049577),
	.w6(32'h3a96075e),
	.w7(32'hbbdc4a53),
	.w8(32'hbb90c87b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03bcb2),
	.w1(32'hbafb87ca),
	.w2(32'hbb80d94c),
	.w3(32'hba638066),
	.w4(32'h3b9430c4),
	.w5(32'hbaba159b),
	.w6(32'hbbdeed3c),
	.w7(32'hbc0bca9a),
	.w8(32'h395fdd02),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba934408),
	.w1(32'h3a9b79a0),
	.w2(32'hbbd9b545),
	.w3(32'h3b99b75f),
	.w4(32'h3abe5705),
	.w5(32'h3bd09d0a),
	.w6(32'hb9fc5a29),
	.w7(32'h3bbdd821),
	.w8(32'hbb9427a6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9f83),
	.w1(32'h3c040034),
	.w2(32'hba171582),
	.w3(32'hbba299ae),
	.w4(32'h3bc578a2),
	.w5(32'h3b8ac1a8),
	.w6(32'hbbdd1ae9),
	.w7(32'h3a05915d),
	.w8(32'h39f91737),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbd27),
	.w1(32'hbade5dd9),
	.w2(32'h3bf33d9e),
	.w3(32'h3996b3f7),
	.w4(32'hbafcea9b),
	.w5(32'h3aa10781),
	.w6(32'h3b8cb4a4),
	.w7(32'h3a609453),
	.w8(32'hbb528f5e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea17cf),
	.w1(32'h3b7c6fa5),
	.w2(32'hbc1ef070),
	.w3(32'h3b56a648),
	.w4(32'h3b404047),
	.w5(32'hba42f322),
	.w6(32'hb9c8d317),
	.w7(32'hb9e44ab7),
	.w8(32'h3a6fb534),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67117b),
	.w1(32'h3b259b67),
	.w2(32'hbc11ff0a),
	.w3(32'h3c03faa9),
	.w4(32'h3c130d36),
	.w5(32'hbb7993f4),
	.w6(32'h3b882f9b),
	.w7(32'h3b8721df),
	.w8(32'hbbfcad38),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc227de8),
	.w1(32'hbc480b99),
	.w2(32'h3c8d1254),
	.w3(32'hbc0c33f2),
	.w4(32'hbb137312),
	.w5(32'h3c5af154),
	.w6(32'hbc1e52db),
	.w7(32'hbbf1615d),
	.w8(32'h3c797acd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d04ee2c),
	.w1(32'h3cd66615),
	.w2(32'hbb174c74),
	.w3(32'h3c809673),
	.w4(32'h3c8c178c),
	.w5(32'h3b8a461f),
	.w6(32'h3d0d37c2),
	.w7(32'h3cfbef8a),
	.w8(32'h3c599e8d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21f38e),
	.w1(32'hbc4c322c),
	.w2(32'hbb935d34),
	.w3(32'h3becd8e0),
	.w4(32'h3a8e2f1d),
	.w5(32'hbc17da3a),
	.w6(32'h3c9846fb),
	.w7(32'h3c0d579d),
	.w8(32'hbc1f8e82),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cf52a),
	.w1(32'h3bff074a),
	.w2(32'hb9f2631d),
	.w3(32'hbba30618),
	.w4(32'hbb64945e),
	.w5(32'h39f7b07a),
	.w6(32'hbc14d11d),
	.w7(32'hbc05b1cb),
	.w8(32'hbb87b4da),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d76be),
	.w1(32'hbc2fd138),
	.w2(32'hbadb3b28),
	.w3(32'h3b193dda),
	.w4(32'h3b06a6aa),
	.w5(32'hba1e9b92),
	.w6(32'h384f5ab8),
	.w7(32'hba011f4c),
	.w8(32'h3aeb990e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072d91),
	.w1(32'hbbd5dd40),
	.w2(32'h3b5ae1dc),
	.w3(32'hbb22d5cb),
	.w4(32'hbb03a2bb),
	.w5(32'hbaefbd98),
	.w6(32'h3b17f9a9),
	.w7(32'hbb164678),
	.w8(32'h3b6e7cee),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45a904),
	.w1(32'h3c14c93f),
	.w2(32'h3bcb7998),
	.w3(32'hbadff1d4),
	.w4(32'hbb447aa6),
	.w5(32'hb9fa7357),
	.w6(32'h398a1350),
	.w7(32'h3b813067),
	.w8(32'h3b2bc43b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb719825),
	.w1(32'hbb77fcbe),
	.w2(32'h3a200fae),
	.w3(32'hba6aaccf),
	.w4(32'hbb532532),
	.w5(32'h3bb9d241),
	.w6(32'hbc2b6393),
	.w7(32'hbb0d94a8),
	.w8(32'h395b40d4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f409f),
	.w1(32'hbbfb633d),
	.w2(32'hbc2f850f),
	.w3(32'hb9358663),
	.w4(32'h3b79ebf4),
	.w5(32'h3b7d3452),
	.w6(32'h3aa83a54),
	.w7(32'hbb426a1f),
	.w8(32'h3b1cc615),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38c878),
	.w1(32'hbc994c57),
	.w2(32'hbbbd7640),
	.w3(32'h3b11fd98),
	.w4(32'hbc05b4ce),
	.w5(32'hbba54aab),
	.w6(32'h3a6f3393),
	.w7(32'h3b17da9f),
	.w8(32'hbb7267b9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5703a),
	.w1(32'hbb49b3a8),
	.w2(32'hb9bc2278),
	.w3(32'hbc1b9c84),
	.w4(32'hba88d50f),
	.w5(32'h3bc3bdc6),
	.w6(32'hbc42846c),
	.w7(32'hbbf503ea),
	.w8(32'hbc2781d9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e008c),
	.w1(32'hbb654609),
	.w2(32'h3b1ca0aa),
	.w3(32'hbbc9bc16),
	.w4(32'hbb1b407b),
	.w5(32'hba7a3bf5),
	.w6(32'hbb709299),
	.w7(32'hbba94852),
	.w8(32'hbb566a39),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1964d2),
	.w1(32'hb948a95c),
	.w2(32'h3bcd2bc8),
	.w3(32'hbbb301d2),
	.w4(32'h3a35e942),
	.w5(32'hbac66fb1),
	.w6(32'hbb6ca41d),
	.w7(32'hba6d1ed1),
	.w8(32'hbc35cef0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc77f8),
	.w1(32'hbc26d83a),
	.w2(32'hbbef3ec9),
	.w3(32'hbc52322d),
	.w4(32'hbc4fbf25),
	.w5(32'h3b7c64cf),
	.w6(32'hbbeb3801),
	.w7(32'hbbe944f1),
	.w8(32'h3c122a40),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c080f51),
	.w1(32'h3c6ff83a),
	.w2(32'hbb3550ff),
	.w3(32'h3c1489d5),
	.w4(32'h3c2bc1e2),
	.w5(32'hbc3ef43e),
	.w6(32'h3ca0967f),
	.w7(32'h3c867ec1),
	.w8(32'hbb63c25c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6661c),
	.w1(32'h3a6eaf0e),
	.w2(32'hbb45b28c),
	.w3(32'hbbbd9975),
	.w4(32'h3b7a7851),
	.w5(32'h3c0733fb),
	.w6(32'hbb57baf0),
	.w7(32'hb8eb1385),
	.w8(32'hbbfee326),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf252f8),
	.w1(32'hbc1f6dc7),
	.w2(32'hbc446b52),
	.w3(32'hbbd028f8),
	.w4(32'h3a6d4d4d),
	.w5(32'hba735712),
	.w6(32'hbba854ac),
	.w7(32'hbb843907),
	.w8(32'hbbd6c3fa),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d972),
	.w1(32'hbb86cf05),
	.w2(32'hbad362b8),
	.w3(32'h39bf6819),
	.w4(32'h3be855ae),
	.w5(32'hbabcc4dc),
	.w6(32'hbb440e39),
	.w7(32'h3b95fc29),
	.w8(32'hbad30e9a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62e4bc),
	.w1(32'hbc3115d2),
	.w2(32'hbb297cc9),
	.w3(32'hbbf1e241),
	.w4(32'hbae52f7e),
	.w5(32'hbb36e0b0),
	.w6(32'hbb9fb4d9),
	.w7(32'hbb54d388),
	.w8(32'hbaa10b0d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f3835),
	.w1(32'hbba93bde),
	.w2(32'hbb9e8921),
	.w3(32'h3b1f3702),
	.w4(32'h3afd76be),
	.w5(32'hbb830885),
	.w6(32'hbb914d2f),
	.w7(32'h3b6e5ed1),
	.w8(32'hbbd38a3a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce66e8),
	.w1(32'hbb10104e),
	.w2(32'h3a52d65e),
	.w3(32'hbb2e3d18),
	.w4(32'hbb9d485c),
	.w5(32'hbbb8757e),
	.w6(32'hbc156fc6),
	.w7(32'hbb805694),
	.w8(32'hbb5e957b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac96616),
	.w1(32'hbbbc9a16),
	.w2(32'h3b228d3f),
	.w3(32'hbbf53e0a),
	.w4(32'hbaa76408),
	.w5(32'hbbf62771),
	.w6(32'hbb43dfaa),
	.w7(32'h3a3e519d),
	.w8(32'hbbd4f63f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941ccc),
	.w1(32'hba87bdbd),
	.w2(32'hbbb4fd1e),
	.w3(32'h3b724908),
	.w4(32'h3b0bf0e8),
	.w5(32'h3a4fdefd),
	.w6(32'h3b5c36dc),
	.w7(32'h3c60199c),
	.w8(32'h3be8ed74),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0d68),
	.w1(32'h3b2bf4b2),
	.w2(32'hbc43a63a),
	.w3(32'h3b8d3164),
	.w4(32'hbb0957c3),
	.w5(32'hba710f95),
	.w6(32'h3b02813f),
	.w7(32'hba77c0c2),
	.w8(32'hbbf02237),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb441a1),
	.w1(32'hbcc55d7a),
	.w2(32'hbc24daec),
	.w3(32'h3afda915),
	.w4(32'hbb991c97),
	.w5(32'hbb1a127a),
	.w6(32'hbc0107b9),
	.w7(32'hbb07ab19),
	.w8(32'h3bc13e0e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d469e),
	.w1(32'hbcd7ade6),
	.w2(32'hbc3de48f),
	.w3(32'hbc28b11b),
	.w4(32'hbc89d21f),
	.w5(32'hbc6bf00d),
	.w6(32'hbb57d796),
	.w7(32'hbb5bb069),
	.w8(32'hbc9fc0a8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90e3f0),
	.w1(32'hbc914c92),
	.w2(32'h3cfbedf8),
	.w3(32'hbcbb1808),
	.w4(32'hbcc53b1e),
	.w5(32'h3c2d46fb),
	.w6(32'hbcd5ff5f),
	.w7(32'hbccd2f35),
	.w8(32'h3cf00930),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3e56ca),
	.w1(32'h3d392ac1),
	.w2(32'hbc5ef780),
	.w3(32'h3cd39cd1),
	.w4(32'h3ced0cab),
	.w5(32'hbc9e449b),
	.w6(32'h3d6a3a60),
	.w7(32'h3d5034f5),
	.w8(32'hbcbf4983),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a6ef6),
	.w1(32'hbcb634f3),
	.w2(32'hbc01443d),
	.w3(32'hbcc533a3),
	.w4(32'hbcd324f5),
	.w5(32'h3b58986d),
	.w6(32'hbcd4e10d),
	.w7(32'hbcbedbe2),
	.w8(32'hbbf50420),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09bda2),
	.w1(32'hbb8062b1),
	.w2(32'h3abbc0cd),
	.w3(32'h3b912729),
	.w4(32'h3b29c85d),
	.w5(32'hbb2e80a8),
	.w6(32'h3c0c8359),
	.w7(32'h3abde380),
	.w8(32'hba4cc259),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54a3da),
	.w1(32'h3b382cc6),
	.w2(32'h3a6a621d),
	.w3(32'hbb079f11),
	.w4(32'hbbbc5df6),
	.w5(32'hbaac019b),
	.w6(32'hbb6778d3),
	.w7(32'h3ae2858c),
	.w8(32'h39633828),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabed251),
	.w1(32'hbb4fe9c2),
	.w2(32'h3b3d754a),
	.w3(32'hbc13dec4),
	.w4(32'hbb3be1b7),
	.w5(32'h3b19b0b5),
	.w6(32'h3ab0841d),
	.w7(32'hbb08b30c),
	.w8(32'hbac25107),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af85bba),
	.w1(32'hbb264c32),
	.w2(32'hbaf59835),
	.w3(32'hb9bd1c11),
	.w4(32'hbaa44cc0),
	.w5(32'h3a2a6d20),
	.w6(32'hbb146640),
	.w7(32'hbb59e678),
	.w8(32'hbb5c0611),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c02c2),
	.w1(32'h3b4d032e),
	.w2(32'h3b7364f3),
	.w3(32'hb9b9dc8f),
	.w4(32'h3a2117f2),
	.w5(32'h3b993a9d),
	.w6(32'hbbad0133),
	.w7(32'hbb5dc077),
	.w8(32'h3c3ba23e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc7c40),
	.w1(32'hbb9a597b),
	.w2(32'hbc5c6ffc),
	.w3(32'hba5b990d),
	.w4(32'h3be448b4),
	.w5(32'hbbaf7b37),
	.w6(32'h3c7f849f),
	.w7(32'h3c0481cc),
	.w8(32'hbc41df2c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6876d9),
	.w1(32'hbc7db6b5),
	.w2(32'hbc15421a),
	.w3(32'hbc39774b),
	.w4(32'hbc176d01),
	.w5(32'hbb62f2df),
	.w6(32'hbc92828e),
	.w7(32'hbc805141),
	.w8(32'h3b2968e8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b5ba1),
	.w1(32'hbbd56b3b),
	.w2(32'hbba93006),
	.w3(32'hbb42c2f0),
	.w4(32'h3ba4f734),
	.w5(32'hbad26869),
	.w6(32'h3c401215),
	.w7(32'h3a41a665),
	.w8(32'h3bbd96ba),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9e1e),
	.w1(32'hbbc477a2),
	.w2(32'hbb82e76d),
	.w3(32'h3bb9cbbd),
	.w4(32'hbad8154f),
	.w5(32'hbba79eed),
	.w6(32'h3a1063cd),
	.w7(32'hbb8e8dc8),
	.w8(32'hbb810376),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf71bdb),
	.w1(32'h3be96242),
	.w2(32'hbc2d502d),
	.w3(32'h3b2f33f4),
	.w4(32'hbac1b1ea),
	.w5(32'hbaa97b18),
	.w6(32'hbbcd6bc0),
	.w7(32'hbc1a29e4),
	.w8(32'hbbff8f4a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc308a26),
	.w1(32'hbc8b99b1),
	.w2(32'hbba2e07d),
	.w3(32'hbadf5f8f),
	.w4(32'hbb9ecb41),
	.w5(32'hbba0b4fe),
	.w6(32'h3bca0455),
	.w7(32'hbc3d7721),
	.w8(32'hbb784964),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8a926),
	.w1(32'hbbb69598),
	.w2(32'hba839169),
	.w3(32'hbbc48125),
	.w4(32'hbb83ef78),
	.w5(32'h3b798c8c),
	.w6(32'hba2d2f11),
	.w7(32'h3bbe8eb1),
	.w8(32'h3baae155),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd94ce9),
	.w1(32'h3bd2dc68),
	.w2(32'hba4cbd93),
	.w3(32'h3c56958a),
	.w4(32'h3bcc238d),
	.w5(32'h3bcb3127),
	.w6(32'h38b91085),
	.w7(32'h3b1ce0e0),
	.w8(32'h3bd156aa),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e6d5),
	.w1(32'hb981363e),
	.w2(32'hbc530da1),
	.w3(32'h3b27a0a8),
	.w4(32'h3bc65990),
	.w5(32'hbc9624d4),
	.w6(32'hb92f3c49),
	.w7(32'hbb8554fe),
	.w8(32'hbcde8caa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf54d),
	.w1(32'hba9ab031),
	.w2(32'h3b91c1f0),
	.w3(32'hbc3125a4),
	.w4(32'hbc12ae89),
	.w5(32'h3bc4b63a),
	.w6(32'hbccaef9a),
	.w7(32'hbcbc18e3),
	.w8(32'h3a8f6deb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce51c7),
	.w1(32'h3b281e71),
	.w2(32'h3bd1b230),
	.w3(32'h3bd50d98),
	.w4(32'h38f29a0e),
	.w5(32'h3bf92066),
	.w6(32'hbb447b82),
	.w7(32'hbbfd1c2b),
	.w8(32'h3bb4f280),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0db513),
	.w1(32'hbbd6ef91),
	.w2(32'hbc3e5916),
	.w3(32'h3b1501ef),
	.w4(32'hb73ebaea),
	.w5(32'hbc7bc307),
	.w6(32'hb96e17c2),
	.w7(32'hbb4fa183),
	.w8(32'hbc064df6),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a91e8),
	.w1(32'hbc08b8f5),
	.w2(32'h3c037874),
	.w3(32'hbca06c17),
	.w4(32'hbc8eec4e),
	.w5(32'hbabb6c37),
	.w6(32'hbbddbb62),
	.w7(32'hba837c31),
	.w8(32'hbbbe65a1),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50d44d),
	.w1(32'hba2c4e98),
	.w2(32'h3bc44a4d),
	.w3(32'h3be38867),
	.w4(32'h3c170e29),
	.w5(32'h3ad8a27f),
	.w6(32'h3c5d84c2),
	.w7(32'h3c8450bb),
	.w8(32'h3bf34304),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0672ce),
	.w1(32'h3b54d60c),
	.w2(32'hbb79eea4),
	.w3(32'h3bd2eafc),
	.w4(32'h3b504121),
	.w5(32'h3a7a8704),
	.w6(32'h3bbae4be),
	.w7(32'h3bdf40d8),
	.w8(32'h3b087f70),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cb35a),
	.w1(32'h3b3ec349),
	.w2(32'h3a0dfc5d),
	.w3(32'h3a4a19e4),
	.w4(32'hbabbc960),
	.w5(32'h3a891bbb),
	.w6(32'hba6f3f60),
	.w7(32'hbaaef9f9),
	.w8(32'hb9c78f6f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ab416),
	.w1(32'hbc12cb78),
	.w2(32'hbbcad742),
	.w3(32'hbb1ccbaf),
	.w4(32'hbb210696),
	.w5(32'hba06badb),
	.w6(32'h3bcce21a),
	.w7(32'hbbb449a2),
	.w8(32'hbb575b5a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbceff),
	.w1(32'hbb7c8a0c),
	.w2(32'hbba7a46e),
	.w3(32'hba7ed8e7),
	.w4(32'h3b1aaa02),
	.w5(32'hb8eb4f12),
	.w6(32'hbbb6f0f6),
	.w7(32'hbb9b2f00),
	.w8(32'hbb8a0a34),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71f87),
	.w1(32'h3a807289),
	.w2(32'h3c9b95da),
	.w3(32'h3bbdd695),
	.w4(32'h3ba0d0f3),
	.w5(32'h3c6c4512),
	.w6(32'h3babc2f2),
	.w7(32'hbb79bd31),
	.w8(32'h3ce04841),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23dd04),
	.w1(32'h3c9e1771),
	.w2(32'hbc2fcbc8),
	.w3(32'h3c7601bf),
	.w4(32'h3c89c39b),
	.w5(32'hbc4ccc84),
	.w6(32'h3ceb9472),
	.w7(32'h3cdf3a0a),
	.w8(32'hbc811c3b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaaaf5b),
	.w1(32'hbcbbbc1d),
	.w2(32'h3a850cf5),
	.w3(32'hbc92d74b),
	.w4(32'hbc8c62ce),
	.w5(32'h3ba8e315),
	.w6(32'hbc83a67c),
	.w7(32'hbc61d866),
	.w8(32'h3b92538b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2b55e),
	.w1(32'h388838a4),
	.w2(32'h3b06c373),
	.w3(32'h3bae188b),
	.w4(32'h3ae26688),
	.w5(32'hbb2cf197),
	.w6(32'h3bb55489),
	.w7(32'h3aedd843),
	.w8(32'h3c5ce872),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10865f),
	.w1(32'hbbeeb83b),
	.w2(32'hbb5e4bb3),
	.w3(32'h3b550bcf),
	.w4(32'hbb6e565a),
	.w5(32'hbb0fcb60),
	.w6(32'h3ccd9c21),
	.w7(32'h3cae240a),
	.w8(32'hba953083),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c56d8),
	.w1(32'hba7de421),
	.w2(32'h3b83f88d),
	.w3(32'hbbbe86eb),
	.w4(32'hbba6b599),
	.w5(32'h3beac9ee),
	.w6(32'hbb85cfb4),
	.w7(32'hbb62788f),
	.w8(32'h3c388837),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd10d7),
	.w1(32'h3b3ac81a),
	.w2(32'hbb96234f),
	.w3(32'h3bbf26ae),
	.w4(32'h3c7c1e92),
	.w5(32'hb5813bca),
	.w6(32'h3c516f95),
	.w7(32'h3c8d4d1b),
	.w8(32'h3b4eb6cf),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1eb4c),
	.w1(32'hbb50a247),
	.w2(32'hbb1dfb62),
	.w3(32'h3a7260ba),
	.w4(32'h39f52a74),
	.w5(32'h3bbc93a1),
	.w6(32'h3bb31c93),
	.w7(32'h3ad66a7e),
	.w8(32'h3b0f2c5e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1efa29),
	.w1(32'hbc3ecf5a),
	.w2(32'hbc61b0cc),
	.w3(32'hbbb5ef5e),
	.w4(32'hbb46af40),
	.w5(32'hba18dd81),
	.w6(32'h3accb34b),
	.w7(32'hbb1b5cdf),
	.w8(32'hbb5e9283),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b2b51),
	.w1(32'hbba17bee),
	.w2(32'h3b87dfaa),
	.w3(32'hb976f803),
	.w4(32'h3b033bf4),
	.w5(32'h3b66c099),
	.w6(32'hbbd9ce12),
	.w7(32'hba90f8b1),
	.w8(32'h3a1da444),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f2381),
	.w1(32'h3ab95d7e),
	.w2(32'hbc3c30c2),
	.w3(32'h3a87223f),
	.w4(32'h3ad382fb),
	.w5(32'hb9d9baeb),
	.w6(32'h3b0fd0a5),
	.w7(32'h3b8b410e),
	.w8(32'hbb8e70d0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f87b0),
	.w1(32'h3c10fd00),
	.w2(32'h3b73ea0e),
	.w3(32'h3adc4861),
	.w4(32'h3b924372),
	.w5(32'hbbc9b020),
	.w6(32'hbba782e5),
	.w7(32'h39f5b5eb),
	.w8(32'h3b870b62),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7eb742),
	.w1(32'hba929779),
	.w2(32'hba85b809),
	.w3(32'h3a5c4673),
	.w4(32'hba642c1f),
	.w5(32'hbab2867b),
	.w6(32'h3b7bd5bc),
	.w7(32'hbb8c81fc),
	.w8(32'hbbaa736b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b400fda),
	.w1(32'h3ace1713),
	.w2(32'h387726d2),
	.w3(32'h3b089e7c),
	.w4(32'hb824b186),
	.w5(32'h3a160bcd),
	.w6(32'hbb0864d2),
	.w7(32'h3b61b239),
	.w8(32'hb9ed8906),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a79c5),
	.w1(32'h3ac8c5b2),
	.w2(32'h3bd70c7c),
	.w3(32'hba414e36),
	.w4(32'h3a8136e8),
	.w5(32'hbbdf45ba),
	.w6(32'hbacd315f),
	.w7(32'hb9d72e6c),
	.w8(32'hbc60bb71),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc839be4),
	.w1(32'h3bc0b207),
	.w2(32'h3c846e74),
	.w3(32'hbc5283fe),
	.w4(32'h3c91b5f2),
	.w5(32'h3cf7f5a3),
	.w6(32'h3bf6a23f),
	.w7(32'h3c4889a0),
	.w8(32'h3cad7fbf),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d034e65),
	.w1(32'hbcac402a),
	.w2(32'h3a717318),
	.w3(32'h3c8f1690),
	.w4(32'hbc32c790),
	.w5(32'hb9c72b5d),
	.w6(32'hbc4db32a),
	.w7(32'h3c31a625),
	.w8(32'hb9033385),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b0a62),
	.w1(32'hbb5c089b),
	.w2(32'hbb910ec1),
	.w3(32'hbb398758),
	.w4(32'hbba63c0a),
	.w5(32'h3b44a8c9),
	.w6(32'hba636dc0),
	.w7(32'hbb39f312),
	.w8(32'h3bb57445),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4260f1),
	.w1(32'hbc94d788),
	.w2(32'h3ac0ba2a),
	.w3(32'hbbfd03c3),
	.w4(32'hbc689cbf),
	.w5(32'h3c2df18a),
	.w6(32'hbc855666),
	.w7(32'hbbe0f52f),
	.w8(32'h3c13794d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21c6fa),
	.w1(32'hbbe0d9f4),
	.w2(32'hba760e14),
	.w3(32'h3bf22fda),
	.w4(32'hbc1ba9be),
	.w5(32'hb991e609),
	.w6(32'hbc95b69f),
	.w7(32'hbc2ce203),
	.w8(32'h3a179fc2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2ff12),
	.w1(32'h3a49a386),
	.w2(32'hbcaba9d6),
	.w3(32'hbb270366),
	.w4(32'hba7bfc8f),
	.w5(32'hbc919b86),
	.w6(32'h3b65e51e),
	.w7(32'h3ad6fd8f),
	.w8(32'h3ba517d2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecdf09),
	.w1(32'h3b6904a0),
	.w2(32'h3c184483),
	.w3(32'h3c9609f0),
	.w4(32'h3b961818),
	.w5(32'h3bb2ab53),
	.w6(32'h3ad02f3f),
	.w7(32'hbc218724),
	.w8(32'h3a7224d0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af51deb),
	.w1(32'h3aac1490),
	.w2(32'h3ce8452b),
	.w3(32'hba4edfa6),
	.w4(32'h3aa715cc),
	.w5(32'h3be08f52),
	.w6(32'h3ab6bc20),
	.w7(32'h39384f98),
	.w8(32'hbcd3fc3f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79e612),
	.w1(32'hbbc19638),
	.w2(32'hbbe6db6a),
	.w3(32'hbc866026),
	.w4(32'h3c8bfc15),
	.w5(32'hbba9fab7),
	.w6(32'h3c65f1e2),
	.w7(32'h3ca0f814),
	.w8(32'hbb86439a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00cb4a),
	.w1(32'hbb765a3d),
	.w2(32'h3c88241e),
	.w3(32'hbbd59bb5),
	.w4(32'hbb544327),
	.w5(32'hbb933bcd),
	.w6(32'h385735b4),
	.w7(32'hbc0881ba),
	.w8(32'hbc33be7e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc040f),
	.w1(32'hbc30a517),
	.w2(32'hbbd708d1),
	.w3(32'hbd0fe14e),
	.w4(32'h3a3fc26b),
	.w5(32'hbbc54d91),
	.w6(32'hbbccebdc),
	.w7(32'h3ca9b318),
	.w8(32'hbb9d7de4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc450cda),
	.w1(32'h3b17e336),
	.w2(32'h3bd3598b),
	.w3(32'hbc8cf4ef),
	.w4(32'h3c0ad312),
	.w5(32'h3bbb3dba),
	.w6(32'h3c0712f8),
	.w7(32'h3bcb5a7c),
	.w8(32'hba0ce616),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1753bb),
	.w1(32'hbaa5069a),
	.w2(32'hbaeb4c78),
	.w3(32'h3b9989b7),
	.w4(32'h3a81e75c),
	.w5(32'hbb815bbc),
	.w6(32'hbc57d293),
	.w7(32'hbb3c91e4),
	.w8(32'hbbfda345),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbb2c3),
	.w1(32'hbbb9b233),
	.w2(32'h3c050f7d),
	.w3(32'hbbbc1f47),
	.w4(32'hbbb3842f),
	.w5(32'h3c539121),
	.w6(32'hbc1f1d53),
	.w7(32'hbbbd3ae5),
	.w8(32'h3ba3bbf5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b737a),
	.w1(32'h3b2b610d),
	.w2(32'hba24e91f),
	.w3(32'hbc19adb8),
	.w4(32'hbc2973c0),
	.w5(32'hbb0e20fa),
	.w6(32'hbc08481e),
	.w7(32'h3bd2332a),
	.w8(32'hbb740a04),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72ca91),
	.w1(32'hbb9fb798),
	.w2(32'hbca92f60),
	.w3(32'hbb2511e2),
	.w4(32'hbadbfff7),
	.w5(32'h3b835af2),
	.w6(32'hbb3e53d7),
	.w7(32'hbac5cbb5),
	.w8(32'h3c80b634),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8781),
	.w1(32'h3c3cf1f9),
	.w2(32'hbbf948ca),
	.w3(32'h3ce91b89),
	.w4(32'hbc754a51),
	.w5(32'h3c9268dd),
	.w6(32'hbbb67e1c),
	.w7(32'hbcb69638),
	.w8(32'hbaf7c49f),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36ce36),
	.w1(32'hbc46cd35),
	.w2(32'h3c1fbd62),
	.w3(32'h3ad08f3f),
	.w4(32'hbcaae459),
	.w5(32'h3ce75fcc),
	.w6(32'hbccd93fb),
	.w7(32'h3c1b6240),
	.w8(32'h3c45b536),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b85a),
	.w1(32'h396636c4),
	.w2(32'hbc130595),
	.w3(32'h3bbcc8bc),
	.w4(32'hbc1f63a2),
	.w5(32'h3c1726c3),
	.w6(32'hbca076e7),
	.w7(32'hbabbabd3),
	.w8(32'h3c94fcef),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c668b91),
	.w1(32'h3aa05087),
	.w2(32'hb8afa84e),
	.w3(32'h3cde4224),
	.w4(32'hbc95ad79),
	.w5(32'h3aba8209),
	.w6(32'hbb79866f),
	.w7(32'hbc1ba47f),
	.w8(32'hb891b4f3),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0bccd),
	.w1(32'hbba48584),
	.w2(32'hbc44723b),
	.w3(32'hbaa72331),
	.w4(32'hba62e25a),
	.w5(32'hbc38f516),
	.w6(32'hbb3d89b7),
	.w7(32'h39658dd6),
	.w8(32'hbbe3daed),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6730),
	.w1(32'hbc81ffd7),
	.w2(32'h3c0219d0),
	.w3(32'hbc7afe76),
	.w4(32'hbc8c5a2d),
	.w5(32'hbb849993),
	.w6(32'hbc7eed8d),
	.w7(32'hbbcbe3df),
	.w8(32'h3bbebeef),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2464),
	.w1(32'h3bc3248b),
	.w2(32'hba9b89ee),
	.w3(32'h3c8628da),
	.w4(32'h3c3f083c),
	.w5(32'h3c94c082),
	.w6(32'h3c6df804),
	.w7(32'h3baf684a),
	.w8(32'h3b131e92),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c772473),
	.w1(32'h3b81f021),
	.w2(32'hbc1f9b99),
	.w3(32'h3bab040b),
	.w4(32'h3c712831),
	.w5(32'hbaae4d99),
	.w6(32'hbbe96a56),
	.w7(32'h3ccb8e7c),
	.w8(32'h3c0cfe39),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabafbb7),
	.w1(32'h3aea96b3),
	.w2(32'h3a88f13d),
	.w3(32'h3cb33d76),
	.w4(32'h3bf8fc57),
	.w5(32'hbb87a5e7),
	.w6(32'h3c790ae5),
	.w7(32'h3c46aa16),
	.w8(32'h3c379782),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c341451),
	.w1(32'h3c625f12),
	.w2(32'h3c830885),
	.w3(32'h3c2164ec),
	.w4(32'h3c027c41),
	.w5(32'hbbdfcce2),
	.w6(32'h3bbcfa7e),
	.w7(32'h3bf24719),
	.w8(32'hbb67c4a3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84915c5),
	.w1(32'hbb3b90f6),
	.w2(32'hbc062b42),
	.w3(32'hbce0fa9e),
	.w4(32'h3c11853c),
	.w5(32'hbbfad65d),
	.w6(32'h3c984ca8),
	.w7(32'h3c01119c),
	.w8(32'h3c9321da),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34286a),
	.w1(32'h3c4d458c),
	.w2(32'h3bbf929c),
	.w3(32'h3b439bf7),
	.w4(32'hbc22f666),
	.w5(32'h3b16d0b2),
	.w6(32'hb9d5dd08),
	.w7(32'hbca372df),
	.w8(32'hbc47fd71),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9e83),
	.w1(32'hbbdd80ae),
	.w2(32'hbc05d53e),
	.w3(32'hbcb47a0d),
	.w4(32'h3b9064d6),
	.w5(32'hbb9900f8),
	.w6(32'hbc549e9b),
	.w7(32'h3c21edb4),
	.w8(32'hbb43a86f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4138b),
	.w1(32'h3a90df31),
	.w2(32'hbb43396a),
	.w3(32'h3b1d2daa),
	.w4(32'hbba72fe6),
	.w5(32'h3a159546),
	.w6(32'hbb7bf0c6),
	.w7(32'hbb90ecbe),
	.w8(32'hbbf3e4e0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393254f3),
	.w1(32'h3c2a5a37),
	.w2(32'hba7d45dd),
	.w3(32'hba7c2795),
	.w4(32'h3c200637),
	.w5(32'hba01ca93),
	.w6(32'h3ae9510d),
	.w7(32'h3bffb5ac),
	.w8(32'hbbdc60b0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3302bd),
	.w1(32'hbc0b6de1),
	.w2(32'hbc87b425),
	.w3(32'hbb8c18a1),
	.w4(32'hba693bba),
	.w5(32'h3b02ce6a),
	.w6(32'hbaa7fb66),
	.w7(32'h3b6e152d),
	.w8(32'hb87559b8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70dce6),
	.w1(32'hbc64f998),
	.w2(32'h3bbfe713),
	.w3(32'hbbbc5cf2),
	.w4(32'hbc349185),
	.w5(32'h3b17a91a),
	.w6(32'hbc37bb8a),
	.w7(32'h39192aa0),
	.w8(32'hbc2d7252),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58430f),
	.w1(32'hbc0532c1),
	.w2(32'hbbe0ed69),
	.w3(32'hbc9e77cb),
	.w4(32'hbcb12162),
	.w5(32'h3aadf918),
	.w6(32'hbd0d096d),
	.w7(32'hbba7da91),
	.w8(32'hbb4e0fc0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb04466),
	.w1(32'hbaeb3975),
	.w2(32'hbb6c6df4),
	.w3(32'h3968b153),
	.w4(32'hbaa9c506),
	.w5(32'hbb984657),
	.w6(32'h3a45bf8a),
	.w7(32'h3c0c61f4),
	.w8(32'hbc3715e8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4767f),
	.w1(32'hbaf295ae),
	.w2(32'h3c41ff93),
	.w3(32'hbba41570),
	.w4(32'h3c2581b8),
	.w5(32'h3c4d891d),
	.w6(32'hbb2b807e),
	.w7(32'h3c151e2f),
	.w8(32'h3aa59d6f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54be5),
	.w1(32'h3ba30f48),
	.w2(32'hbb3ad299),
	.w3(32'h3b9a705c),
	.w4(32'h3b44c295),
	.w5(32'hbbb50499),
	.w6(32'hbc432b95),
	.w7(32'h3b224331),
	.w8(32'h3b092acf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc1f1a),
	.w1(32'hbad19856),
	.w2(32'hbbf165e7),
	.w3(32'hbba976ee),
	.w4(32'hbaa0701b),
	.w5(32'hbbc60e91),
	.w6(32'hbb43c68b),
	.w7(32'hbba1ef9a),
	.w8(32'hbc1c4f57),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e023b),
	.w1(32'hba918d31),
	.w2(32'hba0fdb6b),
	.w3(32'h376dcb3f),
	.w4(32'h3a903eba),
	.w5(32'h3b7ba971),
	.w6(32'hbaefa21c),
	.w7(32'hbb99f5d9),
	.w8(32'hbb71e528),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13b319),
	.w1(32'h3c0694ac),
	.w2(32'h3ab9e0b2),
	.w3(32'h3c13134e),
	.w4(32'hbb3c8402),
	.w5(32'hbbc27fbf),
	.w6(32'h3b0f339f),
	.w7(32'h3c002a33),
	.w8(32'hbb22d65e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b11fa),
	.w1(32'h3b776bfb),
	.w2(32'hbb91d5b3),
	.w3(32'h3b6aab73),
	.w4(32'h3b870104),
	.w5(32'hbbb1e65c),
	.w6(32'h3c171758),
	.w7(32'hbaf24818),
	.w8(32'hbba65932),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d61e0),
	.w1(32'hbb842756),
	.w2(32'hbc70e4cd),
	.w3(32'hbbcfe4e9),
	.w4(32'hbb6c8769),
	.w5(32'hbc0f6e52),
	.w6(32'hbc034403),
	.w7(32'hbbd5924d),
	.w8(32'hbc111a61),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97991),
	.w1(32'h3a39a10e),
	.w2(32'h3b517d5b),
	.w3(32'hba11e9e6),
	.w4(32'h3bce8e97),
	.w5(32'hbb68f4c0),
	.w6(32'hba68b687),
	.w7(32'h3c1fd2bf),
	.w8(32'hbb309908),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dfb1a),
	.w1(32'h3b267c81),
	.w2(32'h3c438a97),
	.w3(32'hbc20f5ba),
	.w4(32'h3bc02e3e),
	.w5(32'h3c32dd84),
	.w6(32'hbb92e1b9),
	.w7(32'h3c11495b),
	.w8(32'h3acc7afa),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64486a),
	.w1(32'h3ba64899),
	.w2(32'h39313565),
	.w3(32'h3b46a536),
	.w4(32'hbc3fc986),
	.w5(32'hbbe39610),
	.w6(32'hbc77be84),
	.w7(32'hbb264ea4),
	.w8(32'h3aff1505),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aaa2f),
	.w1(32'hbc0a604d),
	.w2(32'h3a108b13),
	.w3(32'hbc1fd521),
	.w4(32'h3b5c1b1c),
	.w5(32'hbae723f7),
	.w6(32'hbc11436f),
	.w7(32'hbb0c9a0c),
	.w8(32'hbb83c3dd),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56279b),
	.w1(32'hbb8f7588),
	.w2(32'hbbd178c1),
	.w3(32'hbbce2838),
	.w4(32'hbb82f546),
	.w5(32'h3aff25f2),
	.w6(32'hbbe79591),
	.w7(32'hbbd3bdbf),
	.w8(32'h3ad38fa6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cb9a5),
	.w1(32'hbb735e34),
	.w2(32'h382fbef4),
	.w3(32'h3b9053b7),
	.w4(32'hbc0bd415),
	.w5(32'hbb79ec7e),
	.w6(32'hbba55bb7),
	.w7(32'hb916d37c),
	.w8(32'hbba0363e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc41572),
	.w1(32'hbc03ce03),
	.w2(32'hbadaf547),
	.w3(32'hbbb8a042),
	.w4(32'hbc0e3342),
	.w5(32'h3bb812a0),
	.w6(32'hbb503911),
	.w7(32'hbbbbcb32),
	.w8(32'hbbd5665b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07db7a),
	.w1(32'hbb9bdcf8),
	.w2(32'hbbdb0511),
	.w3(32'hbbdd584d),
	.w4(32'hbc2b0695),
	.w5(32'h3aef72a5),
	.w6(32'hbb59bf48),
	.w7(32'h3bb6f364),
	.w8(32'hbbaf6edc),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188cbd),
	.w1(32'hbc045831),
	.w2(32'h3b9887b3),
	.w3(32'hbca57834),
	.w4(32'hbc5975cf),
	.w5(32'h388e0b4e),
	.w6(32'hbcdce828),
	.w7(32'hb9a29024),
	.w8(32'h3a8a73da),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b5ada),
	.w1(32'hbb0b1ba4),
	.w2(32'hbc2d551f),
	.w3(32'hbb9a86c2),
	.w4(32'hba175869),
	.w5(32'hbb039d4e),
	.w6(32'h3a33f8e3),
	.w7(32'h3b64963a),
	.w8(32'h3b6ff831),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ea60b),
	.w1(32'h3a790b7e),
	.w2(32'h3a3805e4),
	.w3(32'h3c0b8ca4),
	.w4(32'h3bb04c0c),
	.w5(32'h3a25677e),
	.w6(32'h3b752cb4),
	.w7(32'hbaec780b),
	.w8(32'hbac09c87),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e5263),
	.w1(32'h3aedc6d0),
	.w2(32'h3c882d4f),
	.w3(32'h3ad77a7e),
	.w4(32'h3b15168b),
	.w5(32'h3be489a9),
	.w6(32'h3b485a16),
	.w7(32'h3b381f8d),
	.w8(32'hbcad331a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1e4ea),
	.w1(32'h3b885467),
	.w2(32'h3c3539ff),
	.w3(32'hbc4b66f4),
	.w4(32'h3ccb6404),
	.w5(32'h3c8e5460),
	.w6(32'h3cc11d60),
	.w7(32'h3cc86505),
	.w8(32'h3bd89a45),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c971244),
	.w1(32'h3b080c5c),
	.w2(32'h3ba038a5),
	.w3(32'h3c31bcf7),
	.w4(32'hbcd754aa),
	.w5(32'h3c803a57),
	.w6(32'hbc467578),
	.w7(32'hbbf8c0aa),
	.w8(32'h3a6cd7c8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c657ef8),
	.w1(32'h3bed4040),
	.w2(32'h3c06aca5),
	.w3(32'h3c11ae81),
	.w4(32'h3bd00745),
	.w5(32'h3b2c0ae8),
	.w6(32'hb79b312a),
	.w7(32'h3a2bbc9a),
	.w8(32'hbc22982f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dd7d2),
	.w1(32'h3b22c379),
	.w2(32'h3935d3cf),
	.w3(32'hbbec46a4),
	.w4(32'h3c800612),
	.w5(32'hbbc911dc),
	.w6(32'h3ccdb0ad),
	.w7(32'h3c024760),
	.w8(32'hbb8a9e27),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a970557),
	.w1(32'hbc45d170),
	.w2(32'hbcbc4556),
	.w3(32'hbb313214),
	.w4(32'h3a5d5aeb),
	.w5(32'hbc4c67c4),
	.w6(32'h3c18a3a0),
	.w7(32'h3c1d2c62),
	.w8(32'hbb6784c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe91de6),
	.w1(32'hbbc4071e),
	.w2(32'h3b114d8e),
	.w3(32'hbb8f209b),
	.w4(32'hbbc9d4b8),
	.w5(32'h3c75308d),
	.w6(32'hbbbc830a),
	.w7(32'hbb97d551),
	.w8(32'h3ca4f2eb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24b213),
	.w1(32'h3c871ed6),
	.w2(32'hbc33f01e),
	.w3(32'h3cd6c344),
	.w4(32'h3c8b4e1f),
	.w5(32'h3b0cb6a7),
	.w6(32'h3ce19f66),
	.w7(32'hbb0365f6),
	.w8(32'h3c3c24d7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab0786),
	.w1(32'h3c0ac41b),
	.w2(32'hbbecf463),
	.w3(32'h3be72a12),
	.w4(32'hbb09a9cf),
	.w5(32'hba84d5b1),
	.w6(32'h3baded56),
	.w7(32'hbc27c06d),
	.w8(32'hbb591145),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8877c),
	.w1(32'h3b521e5d),
	.w2(32'hbad50916),
	.w3(32'h3bfc440e),
	.w4(32'hbbeeda54),
	.w5(32'h3c3066f6),
	.w6(32'hbbd7cb28),
	.w7(32'hbc8f2f16),
	.w8(32'h3bb19cff),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149919),
	.w1(32'h3c154cef),
	.w2(32'hba53cc1b),
	.w3(32'h3c45e474),
	.w4(32'h3c4a8481),
	.w5(32'h3b2253e0),
	.w6(32'h3c1f84d7),
	.w7(32'h3acc6d3e),
	.w8(32'hbb849c01),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03383e),
	.w1(32'hb9bf5336),
	.w2(32'h3ba2eab4),
	.w3(32'hba7009e1),
	.w4(32'hbb8163da),
	.w5(32'h3a093547),
	.w6(32'hbb704602),
	.w7(32'hbb68b329),
	.w8(32'hba39f132),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac32fcb),
	.w1(32'h3b9b8cac),
	.w2(32'h3ba76857),
	.w3(32'h3b043c42),
	.w4(32'h3a84b1dd),
	.w5(32'hbbd5b91b),
	.w6(32'h3a8edc35),
	.w7(32'h3ba937a0),
	.w8(32'hba874b88),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb679e82),
	.w1(32'h3bbc53e7),
	.w2(32'h3cd90e76),
	.w3(32'hba9a7c89),
	.w4(32'hbbb18345),
	.w5(32'h3d797185),
	.w6(32'hbb98c58e),
	.w7(32'h39aaf71b),
	.w8(32'h3d2091fe),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d55efb2),
	.w1(32'h3bb1587f),
	.w2(32'hbbfb42a2),
	.w3(32'h3d6b09c4),
	.w4(32'hbce428b3),
	.w5(32'h3c114b8d),
	.w6(32'hbc65873e),
	.w7(32'hbc0be6f2),
	.w8(32'h3ab2ef13),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6727dd),
	.w1(32'hbb50b537),
	.w2(32'h3b8adef2),
	.w3(32'h3ae6b863),
	.w4(32'hbb28bcdb),
	.w5(32'h3c9538af),
	.w6(32'hbb1fa502),
	.w7(32'h3b8af40e),
	.w8(32'h3c02576d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82033d),
	.w1(32'h3b2407fa),
	.w2(32'hbc0e4757),
	.w3(32'hba9ac49b),
	.w4(32'hba5dc949),
	.w5(32'h3bbf27b1),
	.w6(32'hbb7e95c8),
	.w7(32'h3bc702c8),
	.w8(32'h3bf3cb14),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5b4ae),
	.w1(32'h3c3f0e7c),
	.w2(32'hba91a8c5),
	.w3(32'h3c4b2c52),
	.w4(32'h3c7ee41e),
	.w5(32'h3a3a032a),
	.w6(32'h3c943576),
	.w7(32'h3c1e0644),
	.w8(32'h3a876158),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a3d6b),
	.w1(32'hbbd2153c),
	.w2(32'h3bd631bb),
	.w3(32'h3bc77b73),
	.w4(32'hbbcc0641),
	.w5(32'h3c593dea),
	.w6(32'hbbe6c9a7),
	.w7(32'hbc86a5d3),
	.w8(32'h3b6265bf),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc88e98),
	.w1(32'hbbbedeca),
	.w2(32'h3be67d2e),
	.w3(32'h39f6f247),
	.w4(32'hbbb253e1),
	.w5(32'h3c648cd5),
	.w6(32'hbb91e532),
	.w7(32'h3c5d6841),
	.w8(32'hbbe4cedc),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f8b38),
	.w1(32'h3aa31161),
	.w2(32'hba485678),
	.w3(32'h3b8a24e9),
	.w4(32'hbc1a8a8b),
	.w5(32'hbb8a5761),
	.w6(32'hbc11767f),
	.w7(32'h3b8217aa),
	.w8(32'hbc14ef41),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67c090),
	.w1(32'h3a2cb88e),
	.w2(32'hbca75650),
	.w3(32'hbc76c383),
	.w4(32'h3c1f09d8),
	.w5(32'hb9312b43),
	.w6(32'hba88056e),
	.w7(32'h3c025fed),
	.w8(32'h3ba62156),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963307c),
	.w1(32'h3b1f48d4),
	.w2(32'hbb4c844e),
	.w3(32'h3bcc602a),
	.w4(32'h3a8ccc0d),
	.w5(32'h3bc750c3),
	.w6(32'h3b257771),
	.w7(32'hbc0ad89b),
	.w8(32'h3b51e944),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba94186),
	.w1(32'h3c54de32),
	.w2(32'h3971f369),
	.w3(32'h3c55c8d8),
	.w4(32'h3c062bc3),
	.w5(32'hbb833430),
	.w6(32'h3bb5cae0),
	.w7(32'h3b7433f4),
	.w8(32'hbbefb973),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2ccfa),
	.w1(32'h3b7748d2),
	.w2(32'h3998cbbd),
	.w3(32'hbbb1ddff),
	.w4(32'h3ca2cb49),
	.w5(32'h397e848a),
	.w6(32'h3c2fa98d),
	.w7(32'h3c78dfef),
	.w8(32'h3b04af00),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036abb),
	.w1(32'h3bcedcc9),
	.w2(32'h3bf47be8),
	.w3(32'hbb272403),
	.w4(32'h3c413312),
	.w5(32'h3c174ab0),
	.w6(32'h3c2998f4),
	.w7(32'h3c3f97f6),
	.w8(32'h3bc79178),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030971),
	.w1(32'hbc304114),
	.w2(32'h3b405fc8),
	.w3(32'hbc05fd2d),
	.w4(32'hbb9e6e6c),
	.w5(32'h3c47075b),
	.w6(32'hbc465008),
	.w7(32'h3c1f8144),
	.w8(32'hbb929bec),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb270),
	.w1(32'h3b2973db),
	.w2(32'hbb479f95),
	.w3(32'h398bddee),
	.w4(32'h3b67d29d),
	.w5(32'hbbf2b33f),
	.w6(32'hbb956ee8),
	.w7(32'h3b2c998c),
	.w8(32'hbbc11b1f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20368),
	.w1(32'hbc0bb329),
	.w2(32'hbc10ad49),
	.w3(32'hbc5d8bf1),
	.w4(32'hbc93da94),
	.w5(32'h3b56a1f2),
	.w6(32'hbcb06592),
	.w7(32'hbbe076e5),
	.w8(32'hb89b2318),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4d6e2),
	.w1(32'hbc3dac71),
	.w2(32'hbbdc7dca),
	.w3(32'hbc3d4565),
	.w4(32'hbc37db05),
	.w5(32'hba08a92d),
	.w6(32'hbc48cce6),
	.w7(32'h3ac79ded),
	.w8(32'hbc30ab49),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca5a4),
	.w1(32'hbc2aef3e),
	.w2(32'hbc6fb009),
	.w3(32'hbbf69031),
	.w4(32'hbbb528f2),
	.w5(32'hbc7f5a62),
	.w6(32'hbc2e749e),
	.w7(32'hbb8773ad),
	.w8(32'h3a7698b7),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98511c),
	.w1(32'h3b91a823),
	.w2(32'h39d51681),
	.w3(32'hbb798fb5),
	.w4(32'h3c07ddeb),
	.w5(32'h3c12e09d),
	.w6(32'h3c594cb2),
	.w7(32'h3c430ed9),
	.w8(32'hba8d5e9e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f20ee),
	.w1(32'hbc74e1ab),
	.w2(32'hbb2f4a8d),
	.w3(32'hbc1c4fb5),
	.w4(32'hbcd9e70c),
	.w5(32'h3bec70d2),
	.w6(32'hbcc96e5b),
	.w7(32'h3ad01fde),
	.w8(32'h3c2851ee),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7816d4),
	.w1(32'h3ab1c90d),
	.w2(32'h3b614ecf),
	.w3(32'hbb181f37),
	.w4(32'hbc1c0689),
	.w5(32'hbbf13e0f),
	.w6(32'hbc19a6ea),
	.w7(32'hb995ae0c),
	.w8(32'hbbcd02ba),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba929646),
	.w1(32'h3b16098c),
	.w2(32'hbbdf8550),
	.w3(32'hbbcc748e),
	.w4(32'h3c08e817),
	.w5(32'hbc04efc0),
	.w6(32'hbb2b3f89),
	.w7(32'h3c07249c),
	.w8(32'h3b9fb9b5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d7d8a),
	.w1(32'hbb396ecb),
	.w2(32'hb87bf8e2),
	.w3(32'hbb8e1d3e),
	.w4(32'hba828af5),
	.w5(32'hba9d2457),
	.w6(32'h3a9aba6b),
	.w7(32'h3b6ed62b),
	.w8(32'hbb7206e1),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33d405),
	.w1(32'h39197591),
	.w2(32'h3c634041),
	.w3(32'hba457153),
	.w4(32'h3b919e0d),
	.w5(32'h3b893d1a),
	.w6(32'h3b43d06e),
	.w7(32'h3ba21b06),
	.w8(32'h3c036aa2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad01607),
	.w1(32'h3b01b13c),
	.w2(32'h3c6773bc),
	.w3(32'h3c20eda1),
	.w4(32'h3bb37da8),
	.w5(32'h3c077877),
	.w6(32'h3c221f2b),
	.w7(32'h3b483093),
	.w8(32'h3b93da0a),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12b303),
	.w1(32'hbb6d28d1),
	.w2(32'hbbaeee25),
	.w3(32'hbb31452f),
	.w4(32'hbaaefdfd),
	.w5(32'h3b46cd53),
	.w6(32'hbc28c7f2),
	.w7(32'h3bbdf0f0),
	.w8(32'h3ba4d7e6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b131123),
	.w1(32'h39e80731),
	.w2(32'hb9c115ba),
	.w3(32'h3c0740b5),
	.w4(32'hbbb25c8f),
	.w5(32'hbb024cae),
	.w6(32'hbb5717e2),
	.w7(32'h3b919984),
	.w8(32'hbb25be14),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5e5f9),
	.w1(32'hbb6fd25b),
	.w2(32'hbb00eca5),
	.w3(32'hbbaff435),
	.w4(32'hbb33ec69),
	.w5(32'hba75e4d5),
	.w6(32'hbb5c3275),
	.w7(32'hbb127c45),
	.w8(32'h3a3013f0),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff7718),
	.w1(32'hbb916937),
	.w2(32'h3bdb4d9b),
	.w3(32'hba15404a),
	.w4(32'hbc06fc56),
	.w5(32'h3ba183b2),
	.w6(32'hbbb491fb),
	.w7(32'hbb27f4b8),
	.w8(32'h3bbd8acb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213680),
	.w1(32'h3b79f37e),
	.w2(32'hbbee8686),
	.w3(32'hba081b00),
	.w4(32'h3b8b6484),
	.w5(32'hbbc4e2ed),
	.w6(32'hba416dab),
	.w7(32'h3c64043a),
	.w8(32'hbb92957e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c2d1),
	.w1(32'h3af09e0b),
	.w2(32'h3b6a68ed),
	.w3(32'hbac39fb3),
	.w4(32'h3b9ee969),
	.w5(32'hbaa07deb),
	.w6(32'h3bbc1fb4),
	.w7(32'h3befadfa),
	.w8(32'h3c5390ca),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b9f6),
	.w1(32'h3c0f011e),
	.w2(32'h3ba5f6ab),
	.w3(32'h3c8b2028),
	.w4(32'h3cb347b4),
	.w5(32'hb9a16894),
	.w6(32'h3cf6b504),
	.w7(32'h3bb7ee1d),
	.w8(32'h3b6cef7b),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31a70b),
	.w1(32'hbbb38208),
	.w2(32'h3b9997be),
	.w3(32'h3bfae61d),
	.w4(32'hbc3ca97e),
	.w5(32'h3b992f55),
	.w6(32'hbc5edcb9),
	.w7(32'h384b252f),
	.w8(32'hbbd6d665),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47b14f),
	.w1(32'hbb0e5479),
	.w2(32'h3c9fd03b),
	.w3(32'h3b61f29c),
	.w4(32'hbc1e2ddf),
	.w5(32'h3d01c3df),
	.w6(32'hbc82897c),
	.w7(32'hbbac753f),
	.w8(32'hbc03998d),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule