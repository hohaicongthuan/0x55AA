module layer_10_featuremap_108(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e4432),
	.w1(32'hbb9a0b4f),
	.w2(32'h3b3c656f),
	.w3(32'hb810f40f),
	.w4(32'h3a9d5b13),
	.w5(32'h3be9bbf0),
	.w6(32'h3a78a631),
	.w7(32'h3b093a8e),
	.w8(32'h3a179d69),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a7a2),
	.w1(32'h39fa3ac1),
	.w2(32'h3aa83791),
	.w3(32'h39eb9838),
	.w4(32'hba93765a),
	.w5(32'hba8e0c21),
	.w6(32'h39d9c072),
	.w7(32'h39c56d1d),
	.w8(32'hb9c5a761),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce4814),
	.w1(32'h3b0781cb),
	.w2(32'h3b48afee),
	.w3(32'hba925bd1),
	.w4(32'hb9b6340e),
	.w5(32'h3afa9861),
	.w6(32'hba8d8c3f),
	.w7(32'hba8614aa),
	.w8(32'hbabd944b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add7423),
	.w1(32'h3a833f2a),
	.w2(32'hbac4bdb9),
	.w3(32'hb91f821c),
	.w4(32'hbbf64bf3),
	.w5(32'hbc0620a2),
	.w6(32'hbb615a5a),
	.w7(32'hbb8499aa),
	.w8(32'hbb0f9262),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad142fd),
	.w1(32'h3a04534b),
	.w2(32'h3b31f33e),
	.w3(32'hbbe20a86),
	.w4(32'h3a400c26),
	.w5(32'h39da337c),
	.w6(32'hb984aebc),
	.w7(32'hba457e83),
	.w8(32'hb9897aa7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3328a0),
	.w1(32'h3a5ab896),
	.w2(32'h37b03b20),
	.w3(32'h3b22a7cc),
	.w4(32'hbaea9a00),
	.w5(32'hbb2ee714),
	.w6(32'h3ac28880),
	.w7(32'h3a7a2f9c),
	.w8(32'h3aca1b8b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2fab),
	.w1(32'h39930aa7),
	.w2(32'h3ab332fd),
	.w3(32'h3a351067),
	.w4(32'hbb007378),
	.w5(32'hba45c2e7),
	.w6(32'h3a2fbee1),
	.w7(32'h38a1e085),
	.w8(32'h394d0398),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d113),
	.w1(32'h39983e88),
	.w2(32'hb99e44e2),
	.w3(32'hbb2551c1),
	.w4(32'hb9f4115a),
	.w5(32'hb9c8d37a),
	.w6(32'hb935205e),
	.w7(32'hbb118f81),
	.w8(32'h380fe41a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4a408),
	.w1(32'hba5d19d7),
	.w2(32'h39f1aa44),
	.w3(32'h399446e7),
	.w4(32'hbaaf77d6),
	.w5(32'hb9e060ad),
	.w6(32'h3a6749a7),
	.w7(32'h39d74a96),
	.w8(32'h3a921923),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8b7ac),
	.w1(32'hba46dcc8),
	.w2(32'hbaeb3cf5),
	.w3(32'hba603d7e),
	.w4(32'hb8269bb0),
	.w5(32'hba685de9),
	.w6(32'h3acb184d),
	.w7(32'hba3a3638),
	.w8(32'h3a4c9197),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8003cce),
	.w1(32'h3b302465),
	.w2(32'h3b538ce9),
	.w3(32'hba3cede5),
	.w4(32'hba57c603),
	.w5(32'h3ac1586a),
	.w6(32'hbb9a3d68),
	.w7(32'hbab881d0),
	.w8(32'hbb47d126),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b570ab9),
	.w1(32'h3ae8f392),
	.w2(32'hbb1a357f),
	.w3(32'hb96719f1),
	.w4(32'hb9e9bf9e),
	.w5(32'hbb731016),
	.w6(32'h3b98580e),
	.w7(32'h3b1c423d),
	.w8(32'h3ba247f0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cc405),
	.w1(32'hbb53fc34),
	.w2(32'hbaf26d6b),
	.w3(32'hbac93cc4),
	.w4(32'hbb1fd42b),
	.w5(32'hbb00d66a),
	.w6(32'hbaa43f53),
	.w7(32'hbb12ae9d),
	.w8(32'hbad2fd2a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f2389),
	.w1(32'h3b86f653),
	.w2(32'h3a400b6f),
	.w3(32'hba66de30),
	.w4(32'h3b26071b),
	.w5(32'h37b1d2c9),
	.w6(32'h3b87258a),
	.w7(32'h3ab68a3a),
	.w8(32'h3b2229e2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52cef1),
	.w1(32'h3a8ccf2c),
	.w2(32'hba061110),
	.w3(32'h3b0ac56d),
	.w4(32'hbacdecae),
	.w5(32'hbb146d36),
	.w6(32'h38a0b0a6),
	.w7(32'h3b2ab58a),
	.w8(32'h3b85fec0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be40a),
	.w1(32'hb9e75e46),
	.w2(32'h3abeb388),
	.w3(32'h3a9a2ae0),
	.w4(32'hbacffa2e),
	.w5(32'hbb033dd1),
	.w6(32'h3a90fed2),
	.w7(32'h3a9bba2f),
	.w8(32'h3aca8efa),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d7867),
	.w1(32'hbaa321d7),
	.w2(32'hba1fb434),
	.w3(32'hbad04e55),
	.w4(32'h3c60c64e),
	.w5(32'h3c637287),
	.w6(32'hbac8db32),
	.w7(32'hba9cc7a4),
	.w8(32'hbabb1968),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ccb6b),
	.w1(32'h3a7c349f),
	.w2(32'h3ae326de),
	.w3(32'h3c415e2f),
	.w4(32'hbaaa9003),
	.w5(32'h3b14c559),
	.w6(32'hba7bb464),
	.w7(32'hbaf144f0),
	.w8(32'hba315482),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886fa6d),
	.w1(32'hbb0e88fe),
	.w2(32'hb92566d2),
	.w3(32'hba9f70d8),
	.w4(32'hbb3a59bd),
	.w5(32'hb7c1da7f),
	.w6(32'hbaeacc03),
	.w7(32'hbb0e9201),
	.w8(32'hba748fdf),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919090a),
	.w1(32'hb8f96bf8),
	.w2(32'h3ab48bfe),
	.w3(32'hbac9452c),
	.w4(32'hbac680d5),
	.w5(32'hb9c5b934),
	.w6(32'h3a923051),
	.w7(32'h3a245549),
	.w8(32'h3a9aa79a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d80b9),
	.w1(32'hbab9aa61),
	.w2(32'hbb876633),
	.w3(32'hbab6fc2a),
	.w4(32'hbb41c9fd),
	.w5(32'hbb83d3cd),
	.w6(32'hba027339),
	.w7(32'hbb0dddba),
	.w8(32'hba851551),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb905569f),
	.w1(32'h3b11fafb),
	.w2(32'h3a7cfb29),
	.w3(32'hbb2d1282),
	.w4(32'hbc00e3af),
	.w5(32'hbb8e015b),
	.w6(32'hbb2aafcc),
	.w7(32'h39c35659),
	.w8(32'hba456aa6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfa5f0),
	.w1(32'h3c8d49e9),
	.w2(32'h3c68c14e),
	.w3(32'hbc182985),
	.w4(32'hbb49923e),
	.w5(32'h3ac132a2),
	.w6(32'hbbbd2e22),
	.w7(32'hbb4bab81),
	.w8(32'hbb8083cb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c999f97),
	.w1(32'h396b2307),
	.w2(32'hb9911675),
	.w3(32'hba2c296f),
	.w4(32'h398a7628),
	.w5(32'hbaad1f1c),
	.w6(32'h3b0f5067),
	.w7(32'h3a414962),
	.w8(32'h3a674070),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9a492),
	.w1(32'hbb5e868a),
	.w2(32'hbac60d80),
	.w3(32'hb99e5d0e),
	.w4(32'hb9a571c8),
	.w5(32'hba388fea),
	.w6(32'hbb177a09),
	.w7(32'hbb3e7100),
	.w8(32'hbb4095e5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66c56f),
	.w1(32'h3b961c15),
	.w2(32'h3b873fe1),
	.w3(32'h3a239dd0),
	.w4(32'h3be75e94),
	.w5(32'h3bf3a34f),
	.w6(32'h3b4a0745),
	.w7(32'h3bbed768),
	.w8(32'h3a1d5622),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee40c8),
	.w1(32'hb8163888),
	.w2(32'h3a1ca04e),
	.w3(32'h3bd7eac1),
	.w4(32'hba8f4a78),
	.w5(32'hbab51a2b),
	.w6(32'h3a974aa1),
	.w7(32'h3a622eef),
	.w8(32'h3a3be9d0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8f52e),
	.w1(32'h392a2dba),
	.w2(32'h3b916742),
	.w3(32'hba1ede9d),
	.w4(32'hba5a8b75),
	.w5(32'hbaf8652c),
	.w6(32'h3a32678b),
	.w7(32'h37a6b516),
	.w8(32'h39fe76b6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e8cf6),
	.w1(32'hba583e8b),
	.w2(32'hbb1adc93),
	.w3(32'hba2835f4),
	.w4(32'h3adcf141),
	.w5(32'h3b0187b7),
	.w6(32'hbacee972),
	.w7(32'hbb6abe12),
	.w8(32'hbb2c61b2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa107f1),
	.w1(32'hbb8a7850),
	.w2(32'hbb9d8d10),
	.w3(32'h3b3115e9),
	.w4(32'h3c61ecff),
	.w5(32'h3c4da2ad),
	.w6(32'h3929d051),
	.w7(32'hbaa0feaf),
	.w8(32'hbb4324e2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c8b1),
	.w1(32'hbac115eb),
	.w2(32'hbb1c82f4),
	.w3(32'h3c57811f),
	.w4(32'hbae7468e),
	.w5(32'hbb03f772),
	.w6(32'hba02469c),
	.w7(32'hbadb994f),
	.w8(32'hb92a5797),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a59e4),
	.w1(32'hb899a8cf),
	.w2(32'hb920a47a),
	.w3(32'hbaa26352),
	.w4(32'hbaa490c1),
	.w5(32'hbad68d1e),
	.w6(32'h39ca6260),
	.w7(32'hba2d10c5),
	.w8(32'hba23704a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aa418),
	.w1(32'hbaaa4e56),
	.w2(32'h3a3bc1e2),
	.w3(32'hba96762a),
	.w4(32'hbb1ac5d8),
	.w5(32'h3b1a6e90),
	.w6(32'hba397d71),
	.w7(32'hbb1d2f72),
	.w8(32'hbabc661f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d3b9e),
	.w1(32'hbb7ab110),
	.w2(32'hbb362461),
	.w3(32'hb9a13402),
	.w4(32'hbaea26b5),
	.w5(32'hbbab4163),
	.w6(32'hbb3eb6d4),
	.w7(32'hbb3a4ce2),
	.w8(32'hbb180dbf),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c79262),
	.w1(32'hba9e6804),
	.w2(32'hbb067bad),
	.w3(32'hbb81e9ef),
	.w4(32'hbae756d2),
	.w5(32'hbacbb3c2),
	.w6(32'hb9fde4dd),
	.w7(32'hbb04354b),
	.w8(32'hba824096),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae31f1b),
	.w1(32'h3966eaa7),
	.w2(32'h389f9a32),
	.w3(32'hbb09b94a),
	.w4(32'hbaf57a85),
	.w5(32'hbab975b8),
	.w6(32'h3a89e22f),
	.w7(32'h3a03e0fc),
	.w8(32'h3aaf9147),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad64287),
	.w1(32'hba63168b),
	.w2(32'h3a0c8889),
	.w3(32'hba43612d),
	.w4(32'hbb4f3643),
	.w5(32'hbadb8d56),
	.w6(32'hbb47367b),
	.w7(32'hbb4cd21a),
	.w8(32'hbb861d79),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f26c2),
	.w1(32'h3a9c15c1),
	.w2(32'h3ac45bc3),
	.w3(32'hb6fe1304),
	.w4(32'h3a2f64ff),
	.w5(32'h380631d9),
	.w6(32'h3b07a15a),
	.w7(32'h3aa0c69d),
	.w8(32'hb94595dc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b44ba7),
	.w1(32'h3aa23c8a),
	.w2(32'h3a9ca17a),
	.w3(32'h3986c244),
	.w4(32'h39cf2f11),
	.w5(32'hba65196a),
	.w6(32'h3b6bf805),
	.w7(32'h3b3d4f1f),
	.w8(32'h3b08d8d1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dcffa),
	.w1(32'h3a17405e),
	.w2(32'h3a7432b6),
	.w3(32'h3a0f8f75),
	.w4(32'hb8d37198),
	.w5(32'hb9e8e885),
	.w6(32'h3a88463d),
	.w7(32'h39dac126),
	.w8(32'hb9e4f238),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f5670),
	.w1(32'hbba47488),
	.w2(32'hbbcaeea3),
	.w3(32'hb9f453a9),
	.w4(32'h3bd44445),
	.w5(32'h3bcd8880),
	.w6(32'hb9b1c83e),
	.w7(32'h3a91cb2a),
	.w8(32'hbb4aa784),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4a240),
	.w1(32'h3a11ac7c),
	.w2(32'h3ab7d1e4),
	.w3(32'h3b891215),
	.w4(32'hbaf26038),
	.w5(32'hbaea8849),
	.w6(32'hba931ff9),
	.w7(32'h39bfd81d),
	.w8(32'h3af2b88c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c63423),
	.w1(32'hba232fd2),
	.w2(32'h384f0607),
	.w3(32'hbaf4f6b2),
	.w4(32'hbab64055),
	.w5(32'hbaa7e8b1),
	.w6(32'hba00bf8f),
	.w7(32'hba8e3f5f),
	.w8(32'hbad821e6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada2ac0),
	.w1(32'h3b345ba4),
	.w2(32'h3989666c),
	.w3(32'hbb38b7c8),
	.w4(32'h3b4193b6),
	.w5(32'h3a53e08b),
	.w6(32'h3b879038),
	.w7(32'h3ac8e4cc),
	.w8(32'h3b404193),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb4205),
	.w1(32'h3b116ae3),
	.w2(32'h3b7d8fb0),
	.w3(32'h3b0534da),
	.w4(32'h3909d488),
	.w5(32'hba771142),
	.w6(32'h3b0f52ff),
	.w7(32'h3a28e2db),
	.w8(32'h3a98718d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b807cdf),
	.w1(32'h39de4813),
	.w2(32'h3b167678),
	.w3(32'hbaadce77),
	.w4(32'hbaf32957),
	.w5(32'hbb2e73d6),
	.w6(32'h39c2049d),
	.w7(32'hba49e84a),
	.w8(32'h3a4a1c58),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a228af5),
	.w1(32'hb9774235),
	.w2(32'hbb97c78b),
	.w3(32'hbb0b2662),
	.w4(32'hbb2ceee0),
	.w5(32'hbbbd9060),
	.w6(32'hba7b1edd),
	.w7(32'h3b4dbf04),
	.w8(32'h3aa674fb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbad9a8),
	.w1(32'hbb4f1d80),
	.w2(32'hbb0d50a1),
	.w3(32'hbb9c9bfb),
	.w4(32'h3a63aacd),
	.w5(32'h3bab987d),
	.w6(32'hbbec6722),
	.w7(32'hbc21418c),
	.w8(32'hbbfecd5b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adefda6),
	.w1(32'h398bd529),
	.w2(32'h3a9a6da4),
	.w3(32'h3b6bfd53),
	.w4(32'hbac4ea74),
	.w5(32'hba24498d),
	.w6(32'h3a86abdc),
	.w7(32'h39c6ebd8),
	.w8(32'hba57b5c7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc7694),
	.w1(32'h3aa7a266),
	.w2(32'h3a299809),
	.w3(32'hbacef434),
	.w4(32'h399c2c29),
	.w5(32'hba2d1b14),
	.w6(32'h3aae5b34),
	.w7(32'h3a0f5195),
	.w8(32'h3a8be5cb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e74a4),
	.w1(32'h3abe1fe3),
	.w2(32'hb8662d8d),
	.w3(32'h3968fb25),
	.w4(32'h3aee85d7),
	.w5(32'h3aab6575),
	.w6(32'h3a2ed04e),
	.w7(32'h3a87fefb),
	.w8(32'h3ac90005),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998fa7f),
	.w1(32'h3b70bfce),
	.w2(32'h3c260d3d),
	.w3(32'hb896bfad),
	.w4(32'h39c1c3c3),
	.w5(32'h3a885a4f),
	.w6(32'h3b48215b),
	.w7(32'h3b90dc94),
	.w8(32'h3b0ff3ec),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cacb7),
	.w1(32'hb96ab277),
	.w2(32'h3a6aeed8),
	.w3(32'hbb7aa311),
	.w4(32'hbb1df7a3),
	.w5(32'hbb5da750),
	.w6(32'h3a0f0944),
	.w7(32'h3a342912),
	.w8(32'h37cc5869),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99e7e1),
	.w1(32'hbaba2192),
	.w2(32'h3882cf9b),
	.w3(32'hbb78fa56),
	.w4(32'hbad3da23),
	.w5(32'h3a849a65),
	.w6(32'hbb107350),
	.w7(32'hbb386141),
	.w8(32'hbb1bb6da),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7d71a),
	.w1(32'hba876e25),
	.w2(32'hba9806d3),
	.w3(32'h3a8d49f4),
	.w4(32'hba49e0d1),
	.w5(32'h3a0771ee),
	.w6(32'h392ce195),
	.w7(32'h39fdad59),
	.w8(32'hbb0683fe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b2bee),
	.w1(32'hbbc0d02e),
	.w2(32'hbb9c3e8a),
	.w3(32'hba3e5918),
	.w4(32'hbb1ee871),
	.w5(32'hba0bdfa1),
	.w6(32'hb947e8b4),
	.w7(32'h3a0702ba),
	.w8(32'h3a52e4dd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37c27),
	.w1(32'hb9651e8d),
	.w2(32'h3a35b29b),
	.w3(32'hbb4ebe33),
	.w4(32'hb98aef5d),
	.w5(32'hbaec52e5),
	.w6(32'hb8fb0317),
	.w7(32'hba1c1396),
	.w8(32'hb80aabd5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a040df7),
	.w1(32'hba3bfb9b),
	.w2(32'h3b08f469),
	.w3(32'hbab455ac),
	.w4(32'h3a8ac14e),
	.w5(32'h3b083cde),
	.w6(32'h3a803578),
	.w7(32'h3b18fa98),
	.w8(32'h3b379091),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ebc99),
	.w1(32'h3a41e65d),
	.w2(32'h3aa85acd),
	.w3(32'h3a14e548),
	.w4(32'hba84aefd),
	.w5(32'hba252bb4),
	.w6(32'h3a6e8672),
	.w7(32'hb7e210c9),
	.w8(32'h39ed7889),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cd4346),
	.w1(32'h3ab7eda6),
	.w2(32'h3ab80f2a),
	.w3(32'hbabb35e6),
	.w4(32'hb96ba933),
	.w5(32'hb99ef9e1),
	.w6(32'h3aed768f),
	.w7(32'h3aa88019),
	.w8(32'h3af77109),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e69764),
	.w1(32'h39cdb684),
	.w2(32'h3b09e5dd),
	.w3(32'hbac002d5),
	.w4(32'hba858024),
	.w5(32'h394a51b8),
	.w6(32'hba2ce4ca),
	.w7(32'hba15d9ed),
	.w8(32'hb8a10b56),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d73e81),
	.w1(32'h37b6f5da),
	.w2(32'h3a77196c),
	.w3(32'hbad2a4d6),
	.w4(32'hba9fccf8),
	.w5(32'hb92c2ce1),
	.w6(32'hba39cad0),
	.w7(32'hbaa1dfb8),
	.w8(32'hb809fa50),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b0109),
	.w1(32'hba0138f2),
	.w2(32'h3b29e5fe),
	.w3(32'hba966516),
	.w4(32'h3898c515),
	.w5(32'h3b682b7c),
	.w6(32'h3873e510),
	.w7(32'hbb7ac96d),
	.w8(32'hbb248cb8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3599),
	.w1(32'h3af8f0a3),
	.w2(32'h3a091acb),
	.w3(32'hbb6f7b91),
	.w4(32'h3ab70804),
	.w5(32'h39a11de6),
	.w6(32'h3b444dbd),
	.w7(32'h3aac1a15),
	.w8(32'h3afafa48),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a891a2b),
	.w1(32'hba7a7f68),
	.w2(32'h3a1c41a9),
	.w3(32'h3a3528ed),
	.w4(32'hbb3f480c),
	.w5(32'hba03e8e2),
	.w6(32'hba2aabdb),
	.w7(32'hb8d914e8),
	.w8(32'h3a1eb303),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6edc6d),
	.w1(32'hb9af6ca4),
	.w2(32'h39ba1178),
	.w3(32'hba4eef17),
	.w4(32'hbab59085),
	.w5(32'hbac511d2),
	.w6(32'hba7a222b),
	.w7(32'hbb31f760),
	.w8(32'hba9f795e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba941aad),
	.w1(32'hbadf0759),
	.w2(32'hb982a40d),
	.w3(32'hbac2efd2),
	.w4(32'h3bde52b2),
	.w5(32'h3be5bdaa),
	.w6(32'hba620cc6),
	.w7(32'h3a91ece1),
	.w8(32'hba79fe89),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd9ead),
	.w1(32'h3c0b5c99),
	.w2(32'h3b3e4edb),
	.w3(32'h3b612028),
	.w4(32'h3bd7ef33),
	.w5(32'h3bbdde31),
	.w6(32'hba770f2e),
	.w7(32'hba3340d2),
	.w8(32'hbbc08c4e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda4cab),
	.w1(32'h3a351350),
	.w2(32'h3a7e56a7),
	.w3(32'h3adaa9e2),
	.w4(32'hb9b42ec4),
	.w5(32'h389bf195),
	.w6(32'h3a536fd5),
	.w7(32'h3af0392d),
	.w8(32'h3aea06f9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abf8e9),
	.w1(32'hbaa239e2),
	.w2(32'hba51f398),
	.w3(32'hb9d27fae),
	.w4(32'h3a9c4619),
	.w5(32'hba1bde7a),
	.w6(32'h3a96f1a8),
	.w7(32'h3a1490a0),
	.w8(32'h3964e56f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0346f7),
	.w1(32'h3aacbb19),
	.w2(32'h3abfbe03),
	.w3(32'h3b349f66),
	.w4(32'hb91fa9a1),
	.w5(32'h38ac257b),
	.w6(32'h3a0a3517),
	.w7(32'hba0ec9a1),
	.w8(32'hb891135f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5d0c3),
	.w1(32'h3a9a3fb9),
	.w2(32'h3a86c38e),
	.w3(32'hba16c8ee),
	.w4(32'hb6c91d52),
	.w5(32'hb9c60b37),
	.w6(32'h3adf28de),
	.w7(32'h3b07de7a),
	.w8(32'h3b1e2bd2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d8cf),
	.w1(32'h3a969052),
	.w2(32'h3a9d0ea6),
	.w3(32'h39533271),
	.w4(32'hba010ec2),
	.w5(32'hb7864e46),
	.w6(32'h3ada2ea9),
	.w7(32'h3ac04921),
	.w8(32'h3adef9cc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86cb12),
	.w1(32'h391a4a74),
	.w2(32'hba3cfce3),
	.w3(32'hba178417),
	.w4(32'hbacc3a08),
	.w5(32'hbace6fca),
	.w6(32'hb8f71741),
	.w7(32'hbab475a3),
	.w8(32'hba3a5bad),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe42e),
	.w1(32'hba0f63e7),
	.w2(32'h3abf45d4),
	.w3(32'hbabf005c),
	.w4(32'hbaf4f5e3),
	.w5(32'hba89183b),
	.w6(32'h39312a75),
	.w7(32'hb9f75022),
	.w8(32'h390d7091),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2581f8),
	.w1(32'h391391fb),
	.w2(32'hbbb4b470),
	.w3(32'hbade1ca6),
	.w4(32'hbb17be45),
	.w5(32'hba955ace),
	.w6(32'h39f4702a),
	.w7(32'h3b294f07),
	.w8(32'hb8326343),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc490570),
	.w1(32'h3a0d2920),
	.w2(32'h39b665f8),
	.w3(32'hbb17ee7f),
	.w4(32'hba0e248c),
	.w5(32'hb9c95711),
	.w6(32'hb8d2015f),
	.w7(32'hbad70bba),
	.w8(32'hb9a86b18),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f7d0a),
	.w1(32'hbb1dfac8),
	.w2(32'hb8776049),
	.w3(32'h39cae362),
	.w4(32'hbb38fb25),
	.w5(32'hba94e4b5),
	.w6(32'hbb0de132),
	.w7(32'hbb609f1c),
	.w8(32'hbafb98a2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6cac85),
	.w1(32'h3a7d40f7),
	.w2(32'hbb47357a),
	.w3(32'hbaba2b98),
	.w4(32'h3938239a),
	.w5(32'h3af45329),
	.w6(32'h3a0e6acc),
	.w7(32'h3abd272d),
	.w8(32'hba4c0987),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e0356),
	.w1(32'hbb4ea883),
	.w2(32'hbba049dd),
	.w3(32'h3b42909b),
	.w4(32'hbb2beffb),
	.w5(32'hbb723f0a),
	.w6(32'hbaf13535),
	.w7(32'hbb82baa2),
	.w8(32'hbaa78cbc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f7acf),
	.w1(32'hba970f83),
	.w2(32'hbb4af037),
	.w3(32'hbb0ef802),
	.w4(32'hbaf93357),
	.w5(32'hbb2dbdea),
	.w6(32'hba51d561),
	.w7(32'hba5ec495),
	.w8(32'hbb53d5b0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6547dc),
	.w1(32'hbab2af5d),
	.w2(32'h3a55ea62),
	.w3(32'hbbb15675),
	.w4(32'hbb24571a),
	.w5(32'hba9e6563),
	.w6(32'hba72f38e),
	.w7(32'hbac60ec0),
	.w8(32'hb954e66f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396abdfa),
	.w1(32'hba3807af),
	.w2(32'h394a4d03),
	.w3(32'hbaa2751e),
	.w4(32'h3a16d0e8),
	.w5(32'h3aaa24d7),
	.w6(32'hba831e69),
	.w7(32'hbac3a916),
	.w8(32'hbae074e3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a4620),
	.w1(32'h38446c1d),
	.w2(32'h3ae337f4),
	.w3(32'h3a6d2c00),
	.w4(32'hbaa08139),
	.w5(32'hb9a1a963),
	.w6(32'h3a8e3c1d),
	.w7(32'hb9dadb6a),
	.w8(32'h3919d71e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86a71d),
	.w1(32'h3b1a2a2c),
	.w2(32'h3ac52173),
	.w3(32'hb9ce0ad5),
	.w4(32'hbb75d3d8),
	.w5(32'hbb0d025b),
	.w6(32'hbb37f889),
	.w7(32'hbbac1bf9),
	.w8(32'hbb92f17b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac9d4e),
	.w1(32'hb930eb5d),
	.w2(32'h3ad62dc5),
	.w3(32'hbac1df68),
	.w4(32'h3af5cf63),
	.w5(32'h3aecdfaf),
	.w6(32'hba62b734),
	.w7(32'hba4ad478),
	.w8(32'hbaa61407),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b9c87),
	.w1(32'hbabcb38e),
	.w2(32'hbb40c7c0),
	.w3(32'h3b568b38),
	.w4(32'h3b84e8b0),
	.w5(32'h3b056456),
	.w6(32'h3a0a9be2),
	.w7(32'hb8487e73),
	.w8(32'hba28e411),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2dd5),
	.w1(32'hbae7d848),
	.w2(32'hbb24d720),
	.w3(32'hb9875f4e),
	.w4(32'hbab38d82),
	.w5(32'hbafb0712),
	.w6(32'hba2a48c4),
	.w7(32'hbadb87cb),
	.w8(32'hba46e009),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ad3a3),
	.w1(32'hba1d71af),
	.w2(32'h38f2ddc5),
	.w3(32'hb8849c6c),
	.w4(32'hb8e598db),
	.w5(32'hb9a12449),
	.w6(32'h3a9d6649),
	.w7(32'h3a7a5bc2),
	.w8(32'hbacd29fd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fecbc),
	.w1(32'hbb187a0b),
	.w2(32'hbb2dcd4d),
	.w3(32'hbb7fbf66),
	.w4(32'hbb7b6d9d),
	.w5(32'hbad9890e),
	.w6(32'hbb954f85),
	.w7(32'hbbaeef7b),
	.w8(32'hbaeda6d3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e1e6c),
	.w1(32'h3a89da33),
	.w2(32'hba149459),
	.w3(32'hbb15e9a6),
	.w4(32'hba9bedf4),
	.w5(32'hbb149c9f),
	.w6(32'h38b5d8c4),
	.w7(32'hbaaa9e5c),
	.w8(32'hba78848a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78cf96),
	.w1(32'h3a56c3ab),
	.w2(32'h3a40347f),
	.w3(32'hba9f05b8),
	.w4(32'hb963f4f1),
	.w5(32'h3a15174e),
	.w6(32'h390b96cb),
	.w7(32'hba8563c9),
	.w8(32'h3a385955),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbf3c7),
	.w1(32'hba9fe870),
	.w2(32'hba9f49bc),
	.w3(32'h3a63ad62),
	.w4(32'hbb4f879a),
	.w5(32'hbb40c1b2),
	.w6(32'hba4fddf6),
	.w7(32'hbaaa6aba),
	.w8(32'hbb28c718),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9701d8a),
	.w1(32'hbae36238),
	.w2(32'hbb64311c),
	.w3(32'hbabf292c),
	.w4(32'hbb19f7e6),
	.w5(32'hbb278ec1),
	.w6(32'hb97b426f),
	.w7(32'h3a52e3ee),
	.w8(32'h381d7c46),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeef9df),
	.w1(32'h3b675571),
	.w2(32'h3b904f85),
	.w3(32'hbb0958cd),
	.w4(32'h3a4a634f),
	.w5(32'h3aab5e1c),
	.w6(32'h3aab6817),
	.w7(32'h3aa0fe62),
	.w8(32'h379644c9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5862ab),
	.w1(32'hbb3de119),
	.w2(32'hbbd30ffb),
	.w3(32'h3a566a23),
	.w4(32'hb99773c4),
	.w5(32'h38381c99),
	.w6(32'h3b410b6f),
	.w7(32'h3af517e3),
	.w8(32'h3adb7849),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbc5ea),
	.w1(32'h3bd013d3),
	.w2(32'h3bb97815),
	.w3(32'h3b0f3e05),
	.w4(32'hbbbdcb86),
	.w5(32'hbb3db1f9),
	.w6(32'hbb4dd080),
	.w7(32'hba2c8b3d),
	.w8(32'hbb884444),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfb218),
	.w1(32'h3a47a982),
	.w2(32'h3b1a37df),
	.w3(32'hbba3e473),
	.w4(32'h3a6208a8),
	.w5(32'h3b29149b),
	.w6(32'h3ab4123f),
	.w7(32'hb9e8d7eb),
	.w8(32'hbaaf3610),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b092f48),
	.w1(32'h39cf6ca7),
	.w2(32'h3ae408db),
	.w3(32'h3a64c208),
	.w4(32'hba9bf24f),
	.w5(32'hbaa76f76),
	.w6(32'h3a80eaac),
	.w7(32'h39e53b22),
	.w8(32'h39282b9a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a050733),
	.w1(32'hbb936c17),
	.w2(32'hbb533075),
	.w3(32'hbb8286e4),
	.w4(32'hbba3b170),
	.w5(32'hbb75a68c),
	.w6(32'hbbe54ffe),
	.w7(32'hbbdd9c85),
	.w8(32'hbbe36b1e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2282af),
	.w1(32'h3a607453),
	.w2(32'h3b30f022),
	.w3(32'h3ac2e09d),
	.w4(32'h3b611f52),
	.w5(32'h3acad15a),
	.w6(32'h3a0883ac),
	.w7(32'h3b378afa),
	.w8(32'hba41a485),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39948018),
	.w1(32'hb95dc850),
	.w2(32'hbb7194ee),
	.w3(32'hba4ee1f2),
	.w4(32'h3a97a114),
	.w5(32'hbb3b4481),
	.w6(32'h3ab69bf9),
	.w7(32'h3acd67f8),
	.w8(32'h3ab0c96b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3245c),
	.w1(32'h3b85533e),
	.w2(32'hb9121cba),
	.w3(32'h3ba2e322),
	.w4(32'h3ad64b7f),
	.w5(32'hb9abda7b),
	.w6(32'h3b56ab47),
	.w7(32'h3a0f2ae2),
	.w8(32'h3b093d9c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f4c2c),
	.w1(32'h3a9aeda7),
	.w2(32'h3a35d20b),
	.w3(32'h3ac756bc),
	.w4(32'hbabe95ff),
	.w5(32'hbb035570),
	.w6(32'h3a8ac840),
	.w7(32'h3b0bb1fd),
	.w8(32'h3b0c927a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d635),
	.w1(32'hba1ba9cb),
	.w2(32'hbad26fbc),
	.w3(32'hbb13d860),
	.w4(32'hba56a22f),
	.w5(32'hbaebf9d3),
	.w6(32'hba476945),
	.w7(32'hbb0192d0),
	.w8(32'hbabcec32),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0689e2),
	.w1(32'hbad8dd6f),
	.w2(32'hba966881),
	.w3(32'h3ae298e0),
	.w4(32'hbb2da40e),
	.w5(32'hbb508dce),
	.w6(32'h3a9d0a50),
	.w7(32'h3970ca5b),
	.w8(32'hba21495f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3719d63d),
	.w1(32'h3b34861c),
	.w2(32'h3b69fbb5),
	.w3(32'hbaec4fa2),
	.w4(32'hbb1c81de),
	.w5(32'hb9d752b6),
	.w6(32'hb8be31fd),
	.w7(32'hb9bc075d),
	.w8(32'hba34cef0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30079d),
	.w1(32'h3ac2acfe),
	.w2(32'hba5a28fa),
	.w3(32'hbaeaf0c7),
	.w4(32'hbadd7e8d),
	.w5(32'hbb086fc3),
	.w6(32'hba537a97),
	.w7(32'hbb098b86),
	.w8(32'hba1f4721),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcec52),
	.w1(32'h3a830c4c),
	.w2(32'hba950d74),
	.w3(32'hba9c0681),
	.w4(32'h39d64c1d),
	.w5(32'hba94afd1),
	.w6(32'h3ae12e3b),
	.w7(32'h38c5bbac),
	.w8(32'h3a2c7bad),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ab2a),
	.w1(32'h3b07d521),
	.w2(32'h3aceffa6),
	.w3(32'h3accbffb),
	.w4(32'hba9791b9),
	.w5(32'hba152c66),
	.w6(32'h3b6e820c),
	.w7(32'h3b1f0e1a),
	.w8(32'h3b262177),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b85b),
	.w1(32'h3ade6348),
	.w2(32'h3b4353af),
	.w3(32'h3a115c5b),
	.w4(32'hba7c5552),
	.w5(32'hbad0bd6c),
	.w6(32'h3b305037),
	.w7(32'h3b0aed3b),
	.w8(32'h3a8eb6a5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adea6e3),
	.w1(32'h3a1e8fe2),
	.w2(32'h3bae7e3c),
	.w3(32'hba9cb394),
	.w4(32'hb8be171e),
	.w5(32'h3b8fe54c),
	.w6(32'h3b0380c3),
	.w7(32'h3a5b0529),
	.w8(32'hba9d0e3e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acd82f),
	.w1(32'h39e070f3),
	.w2(32'h3b31f895),
	.w3(32'hbb2c7b8a),
	.w4(32'hbb056370),
	.w5(32'hba4c5271),
	.w6(32'hb96e07e1),
	.w7(32'h3754cf2d),
	.w8(32'h3acc54a5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae42b2),
	.w1(32'h39dacdca),
	.w2(32'h38b26935),
	.w3(32'hbaf63f2c),
	.w4(32'hba8b3a83),
	.w5(32'hb9dcd0c1),
	.w6(32'hba6e1876),
	.w7(32'h3a23bb02),
	.w8(32'h3b3435cc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e04659),
	.w1(32'hbb3ddd51),
	.w2(32'hbb403207),
	.w3(32'hbaa5f3a7),
	.w4(32'hbb8ac05b),
	.w5(32'hbb8e6f7f),
	.w6(32'hbacd14aa),
	.w7(32'hbb67bd50),
	.w8(32'hbb83bee0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572642),
	.w1(32'h3b262d0b),
	.w2(32'hb90b353f),
	.w3(32'hbb9fc26e),
	.w4(32'h3a442e64),
	.w5(32'hba30ad37),
	.w6(32'h3b211d63),
	.w7(32'h3a02c196),
	.w8(32'h3ad464f1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228dc7),
	.w1(32'h3a445f38),
	.w2(32'h39101c76),
	.w3(32'h3a9580f1),
	.w4(32'h38edb098),
	.w5(32'hb8b6552a),
	.w6(32'h3aa8f3ec),
	.w7(32'h3a07aea9),
	.w8(32'h3a7e0111),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1759f),
	.w1(32'h3a58d27c),
	.w2(32'hb9e8e488),
	.w3(32'h3a2e9589),
	.w4(32'hb9fb5596),
	.w5(32'hba1b02b0),
	.w6(32'h3ad53b11),
	.w7(32'h39cbf9a9),
	.w8(32'h3a900b4d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92af67),
	.w1(32'h3ae10687),
	.w2(32'h3b3a5d4a),
	.w3(32'h3a115929),
	.w4(32'hbb295acd),
	.w5(32'hbaa2ef56),
	.w6(32'h3abf2876),
	.w7(32'h3a88c6ba),
	.w8(32'h3b38bcce),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1def),
	.w1(32'hbb126ec4),
	.w2(32'h3944c10d),
	.w3(32'hb9e43777),
	.w4(32'hbb2b51df),
	.w5(32'h3978a5f2),
	.w6(32'hba92bc0b),
	.w7(32'hba97ae42),
	.w8(32'hba694186),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01048d),
	.w1(32'h3ad9fefa),
	.w2(32'h3b5832c1),
	.w3(32'hbb7ab4a1),
	.w4(32'hbb015bb7),
	.w5(32'hbb420e01),
	.w6(32'h3874dd82),
	.w7(32'h3a63aa6d),
	.w8(32'h3b2b50a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ca864),
	.w1(32'h39b15274),
	.w2(32'h3b09b115),
	.w3(32'hbacf706a),
	.w4(32'hbabf0ecb),
	.w5(32'hba188cbe),
	.w6(32'h3aaea6a7),
	.w7(32'h3a7714b3),
	.w8(32'h3acf8501),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d677),
	.w1(32'h3a7ae418),
	.w2(32'hb9bc3b9a),
	.w3(32'h3923a6fd),
	.w4(32'hb939d04d),
	.w5(32'hbb280fef),
	.w6(32'h3b214c43),
	.w7(32'h3a7186ab),
	.w8(32'h3785ed44),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8030f),
	.w1(32'hbac7c2bc),
	.w2(32'hbad04b63),
	.w3(32'hb986d35a),
	.w4(32'hbab290b6),
	.w5(32'hbaf1eade),
	.w6(32'hb98cab2f),
	.w7(32'h3a76e0bc),
	.w8(32'h3b36f36d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80bdb7),
	.w1(32'hbac2bdc8),
	.w2(32'hbb377503),
	.w3(32'hbb0c494c),
	.w4(32'hbb5517ce),
	.w5(32'hbb5f3a3f),
	.w6(32'hb95e67f6),
	.w7(32'h391682c9),
	.w8(32'h39552cab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a146849),
	.w1(32'hbacc7ae0),
	.w2(32'hbb67c564),
	.w3(32'hbb1d3c1d),
	.w4(32'hbb1bfe2e),
	.w5(32'hbb6837c2),
	.w6(32'hb9c16537),
	.w7(32'hbb101df0),
	.w8(32'hb928cecf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e3f9b),
	.w1(32'h3b9085cc),
	.w2(32'h39ca2f75),
	.w3(32'hbad4b470),
	.w4(32'h3b8b528f),
	.w5(32'h3bdb3e40),
	.w6(32'hbb82286a),
	.w7(32'hbc588fcb),
	.w8(32'hbb8e3909),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b6129),
	.w1(32'h3ae7f7b7),
	.w2(32'h3bbc2ff6),
	.w3(32'hbb2ba35a),
	.w4(32'h3a6cc217),
	.w5(32'h3c0ba27e),
	.w6(32'hbb84f87c),
	.w7(32'hbc1b550e),
	.w8(32'hbbb5a0e8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a036440),
	.w1(32'h3b94c392),
	.w2(32'h3cdd3b5f),
	.w3(32'hbacabda7),
	.w4(32'hbbb77eaf),
	.w5(32'h3b3a4bf9),
	.w6(32'h3c27f407),
	.w7(32'h3b32662e),
	.w8(32'hbc02d468),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb136261),
	.w1(32'hbb8c108f),
	.w2(32'h3a82908e),
	.w3(32'h3b73c0e0),
	.w4(32'hbb689b2a),
	.w5(32'hbc00d661),
	.w6(32'h3b7992fd),
	.w7(32'h3c85a6f8),
	.w8(32'h3b84a164),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a883f03),
	.w1(32'hbc225267),
	.w2(32'hbc1208fa),
	.w3(32'hbb5ca7e0),
	.w4(32'h3a2373b0),
	.w5(32'hbb478517),
	.w6(32'hbb8f3b17),
	.w7(32'h3bfaad81),
	.w8(32'h3b2e32fb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf67453),
	.w1(32'hbc6792d3),
	.w2(32'hbc4f3012),
	.w3(32'hba607461),
	.w4(32'hba84dee0),
	.w5(32'h3b39d3a6),
	.w6(32'h3a07d7b4),
	.w7(32'hbb9ebbc9),
	.w8(32'h3ba851c8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b8e0b),
	.w1(32'hbb1294f5),
	.w2(32'hbc30bf89),
	.w3(32'h3b81b4b7),
	.w4(32'h3bd94652),
	.w5(32'h3ac50af3),
	.w6(32'hbc0ed59c),
	.w7(32'hbc4df1e4),
	.w8(32'h3a48ccbf),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cc3c4),
	.w1(32'h3b5ec97c),
	.w2(32'h3bbf4712),
	.w3(32'hbc00067d),
	.w4(32'hb9c1df7f),
	.w5(32'h3bf0f31b),
	.w6(32'h3a3cc53f),
	.w7(32'hbb10d4d9),
	.w8(32'hb96136fd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ef4c5),
	.w1(32'hbc092a35),
	.w2(32'hbb089c5f),
	.w3(32'hbbbcb0c0),
	.w4(32'hbbbf5c53),
	.w5(32'hbc222f1c),
	.w6(32'h3a5cb272),
	.w7(32'h3c681f39),
	.w8(32'h3b4c2f9d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b3513),
	.w1(32'h3b4d8a2d),
	.w2(32'h3b5a6de9),
	.w3(32'hbba1b68c),
	.w4(32'h3b9487bb),
	.w5(32'h3c55234c),
	.w6(32'hbbd11a2b),
	.w7(32'hbc928cfd),
	.w8(32'hbc1e25d0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a133),
	.w1(32'h3b8f9eea),
	.w2(32'h3b813b16),
	.w3(32'h3ab36d79),
	.w4(32'h3a5719fa),
	.w5(32'h3b8d6e26),
	.w6(32'hbb614466),
	.w7(32'hbbd635f0),
	.w8(32'hbb1fe25d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af1a71),
	.w1(32'hbc5b5337),
	.w2(32'hbc580b5a),
	.w3(32'hba6e52ee),
	.w4(32'hbc0799c5),
	.w5(32'hbc920366),
	.w6(32'h3c30e0a5),
	.w7(32'h3d0eea9b),
	.w8(32'h3c5ed7a0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca4b1),
	.w1(32'hbcff6e64),
	.w2(32'hbd0fd813),
	.w3(32'hbbbbf008),
	.w4(32'hbb535ef1),
	.w5(32'hbb75a162),
	.w6(32'hbbab81cb),
	.w7(32'hba897508),
	.w8(32'h3a6938df),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf0a033),
	.w1(32'hbb9d6ef5),
	.w2(32'hbc02c361),
	.w3(32'hbb42961e),
	.w4(32'hbbd1f441),
	.w5(32'hbbf5bbbf),
	.w6(32'hbbf77702),
	.w7(32'hbc4d41df),
	.w8(32'hbbb082ce),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc129753),
	.w1(32'hbb539a75),
	.w2(32'hbb96c286),
	.w3(32'hbbcede2f),
	.w4(32'hbb100a33),
	.w5(32'hb8afca20),
	.w6(32'hbbacdb85),
	.w7(32'hbc0e20ad),
	.w8(32'hbb9dc212),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947727),
	.w1(32'h3be88b78),
	.w2(32'h3b13c99e),
	.w3(32'hbb3fec4a),
	.w4(32'h3c1e88a0),
	.w5(32'h3cc84c18),
	.w6(32'hbbb4006c),
	.w7(32'hbcdfc3ca),
	.w8(32'hbc91c451),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84481b),
	.w1(32'h3a3e56fb),
	.w2(32'h3bb8ac0b),
	.w3(32'h3c1a6ec4),
	.w4(32'h3bdf154e),
	.w5(32'h3b160b7c),
	.w6(32'hba8522bc),
	.w7(32'hbbacb7f7),
	.w8(32'h3b863321),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc316a5f),
	.w1(32'h3b890ed8),
	.w2(32'h3b381bbd),
	.w3(32'hbb5fd97c),
	.w4(32'hbb80ac23),
	.w5(32'h3a6b9cac),
	.w6(32'hbb0facee),
	.w7(32'hbbf0570a),
	.w8(32'hbb8f75eb),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce2486),
	.w1(32'hbb34ca2c),
	.w2(32'h3bd23c3b),
	.w3(32'hbb9fba86),
	.w4(32'hbb16fc6e),
	.w5(32'h3b82c097),
	.w6(32'hbb7a75ae),
	.w7(32'hbc0eeb5f),
	.w8(32'hbaa205b5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac81213),
	.w1(32'hbc0140b9),
	.w2(32'hbbec3aa9),
	.w3(32'h3b402458),
	.w4(32'hbbdf13cf),
	.w5(32'hbc959863),
	.w6(32'h3c167c1a),
	.w7(32'h3cdcfaeb),
	.w8(32'h3c1e3bd5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb708cad),
	.w1(32'hbb0a6b2a),
	.w2(32'h3aa944f1),
	.w3(32'hbc035a38),
	.w4(32'hbb1b0d16),
	.w5(32'hbba3a4fd),
	.w6(32'h3ab99ced),
	.w7(32'h3c2d57e4),
	.w8(32'h3a5610fa),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb684419),
	.w1(32'hba82014c),
	.w2(32'hbaa2a961),
	.w3(32'hbb4b97ae),
	.w4(32'hbb106060),
	.w5(32'h3a25fede),
	.w6(32'hbb9db7e4),
	.w7(32'hbc0be4c1),
	.w8(32'hbba9a949),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195568),
	.w1(32'hbaed473b),
	.w2(32'hbbc8796b),
	.w3(32'hbb196ba8),
	.w4(32'h3b2766ff),
	.w5(32'h3bc13a07),
	.w6(32'hbbf6ca49),
	.w7(32'hbc9c20f7),
	.w8(32'hbc07afb6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa0f11),
	.w1(32'hbc5b7d54),
	.w2(32'hbc095f6e),
	.w3(32'h3a68ca15),
	.w4(32'hba857663),
	.w5(32'hbb21c339),
	.w6(32'h394b4c48),
	.w7(32'h3ab4516f),
	.w8(32'hbb46855e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9b37),
	.w1(32'h3a41b838),
	.w2(32'hbbd97b91),
	.w3(32'hbb80c205),
	.w4(32'hbb642158),
	.w5(32'hbbe3c4f7),
	.w6(32'hbb57af93),
	.w7(32'hbc35f149),
	.w8(32'hbb98ce77),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945502),
	.w1(32'h3b0cdba5),
	.w2(32'h3bc57d45),
	.w3(32'hbb51cb47),
	.w4(32'h3b079193),
	.w5(32'h3c53cfe8),
	.w6(32'hbc0abf53),
	.w7(32'hbc955ca5),
	.w8(32'hbc27a704),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09ad1c),
	.w1(32'hbc05c64f),
	.w2(32'hbbcb010f),
	.w3(32'h3b3be64b),
	.w4(32'hbaadaac0),
	.w5(32'hbb762ea5),
	.w6(32'h3b816418),
	.w7(32'h3b63387f),
	.w8(32'hba898926),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4672d0),
	.w1(32'h3a00f3b0),
	.w2(32'h3bb7d608),
	.w3(32'h3ad7df16),
	.w4(32'hba8e6cfb),
	.w5(32'hbb9e4a90),
	.w6(32'h3ba7fa4a),
	.w7(32'h3abab2a7),
	.w8(32'h38c88578),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc3fe1),
	.w1(32'hba06be7c),
	.w2(32'hba7110f2),
	.w3(32'hbc081d22),
	.w4(32'hbb804e89),
	.w5(32'hbaefabe8),
	.w6(32'hbb8ac0fa),
	.w7(32'hbc0f0e0a),
	.w8(32'hbbbc1974),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88a53e),
	.w1(32'hbc04b544),
	.w2(32'hbb7c7e9c),
	.w3(32'hbbb37969),
	.w4(32'hbbc5373f),
	.w5(32'hbb9ed602),
	.w6(32'h3aeb968c),
	.w7(32'h3c238dbb),
	.w8(32'hb94a9235),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b07c3d),
	.w1(32'h3ada624c),
	.w2(32'hbb860471),
	.w3(32'h3b1d8f91),
	.w4(32'h3bedb70b),
	.w5(32'h3afd6da2),
	.w6(32'h3af93ad6),
	.w7(32'hbbeca41b),
	.w8(32'hbb94c4b6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb22bad),
	.w1(32'h3a6a7dd6),
	.w2(32'h3ac884cd),
	.w3(32'hbaf847ce),
	.w4(32'h3b2d5426),
	.w5(32'h3bf3c20f),
	.w6(32'hbab9fc36),
	.w7(32'hba79623f),
	.w8(32'hbb91a499),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6e82e),
	.w1(32'hbac8f158),
	.w2(32'hbb362671),
	.w3(32'h3ba6b6a7),
	.w4(32'hba693064),
	.w5(32'h3b067155),
	.w6(32'hbb9de693),
	.w7(32'hbc1fc779),
	.w8(32'hbba7a7a4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6396b4),
	.w1(32'hbb91a470),
	.w2(32'hbb566e16),
	.w3(32'hbb29601a),
	.w4(32'hbbdd8d74),
	.w5(32'hbbcaf393),
	.w6(32'hbba7ba25),
	.w7(32'hbc2e2ed8),
	.w8(32'hbbe31172),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac6f9),
	.w1(32'hbb723f92),
	.w2(32'hbb1c11bb),
	.w3(32'hbc0eef3a),
	.w4(32'hbbf918bd),
	.w5(32'hbc0bddd5),
	.w6(32'hbb9d5ae5),
	.w7(32'hbbef0435),
	.w8(32'hbb9ed458),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3de6d3),
	.w1(32'h3b0c0fc7),
	.w2(32'h3ba18bad),
	.w3(32'hbb9a1e23),
	.w4(32'hbbaab306),
	.w5(32'hbbc4f254),
	.w6(32'h388f4f13),
	.w7(32'hbb58a60a),
	.w8(32'hbc1e8966),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242527),
	.w1(32'hbc374b42),
	.w2(32'hbc29d82c),
	.w3(32'hbc1c70b9),
	.w4(32'hbc2b5dda),
	.w5(32'hbca2ff19),
	.w6(32'h3c3ff0bc),
	.w7(32'h3cf9f2d1),
	.w8(32'h3c5ef60f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79830d),
	.w1(32'hbb9383ce),
	.w2(32'hbb51b910),
	.w3(32'hbc2e6bef),
	.w4(32'hbbb6936f),
	.w5(32'hbbc8f339),
	.w6(32'hbba99143),
	.w7(32'hbc11369d),
	.w8(32'hbba935fb),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05f2d8),
	.w1(32'hbb83249b),
	.w2(32'hbaa1bc79),
	.w3(32'hbc16bab1),
	.w4(32'h38b998d8),
	.w5(32'hbbed2c56),
	.w6(32'h3b559155),
	.w7(32'h3c8c8cc1),
	.w8(32'h3c00b737),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f97f0),
	.w1(32'hbbe678f1),
	.w2(32'hbb6b2d2c),
	.w3(32'hbbc4507f),
	.w4(32'hbb8b9848),
	.w5(32'hbc1b1978),
	.w6(32'h3b37caf8),
	.w7(32'h3c51adaa),
	.w8(32'h39e0b893),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8970c4),
	.w1(32'h3ad4fb52),
	.w2(32'h3bcf89e7),
	.w3(32'hbbcb869f),
	.w4(32'h39fe0672),
	.w5(32'h3c1749b2),
	.w6(32'hbb9d2453),
	.w7(32'hbc4fd09f),
	.w8(32'hbbf6debd),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db4112),
	.w1(32'hbb23e467),
	.w2(32'h3a169fee),
	.w3(32'h3a9924dc),
	.w4(32'hba9d7581),
	.w5(32'hbbd7c589),
	.w6(32'hb56b83b0),
	.w7(32'h3c2df3a6),
	.w8(32'h39fa04d9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a80b7b),
	.w1(32'h3b8cc6a3),
	.w2(32'h3af8e9f6),
	.w3(32'hbb77f7ac),
	.w4(32'h3b91aec8),
	.w5(32'h3b94d744),
	.w6(32'h3a81762a),
	.w7(32'hbb4d7f24),
	.w8(32'hbb933864),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e75f65),
	.w1(32'hbc03f807),
	.w2(32'hbb8ad7f9),
	.w3(32'h3bbf920e),
	.w4(32'hbb7adf80),
	.w5(32'hbc057186),
	.w6(32'hba247feb),
	.w7(32'h3bda417c),
	.w8(32'h3b75dc1a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb360ec4),
	.w1(32'hbb1e7789),
	.w2(32'hbaecc993),
	.w3(32'hba306051),
	.w4(32'hbba5fee9),
	.w5(32'hbb867e3c),
	.w6(32'hbbb693d7),
	.w7(32'hbc2a13eb),
	.w8(32'hbc073377),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb442001),
	.w1(32'hbc632b90),
	.w2(32'hbc0b6900),
	.w3(32'hbb99afbd),
	.w4(32'hbb89b680),
	.w5(32'hbc5dfa7a),
	.w6(32'h3ca36ef3),
	.w7(32'h3d37dd53),
	.w8(32'h3c9fce1c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8da1f),
	.w1(32'hbc056bbd),
	.w2(32'hbbb3edd2),
	.w3(32'hba05db3e),
	.w4(32'hbbb501e7),
	.w5(32'hbc2e8f0b),
	.w6(32'h3bab7b81),
	.w7(32'h3c210017),
	.w8(32'hba8fa842),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b4902),
	.w1(32'hbbd92860),
	.w2(32'hbbb0cb7f),
	.w3(32'hbb937b20),
	.w4(32'hbbfade2a),
	.w5(32'hbc03edcd),
	.w6(32'h3bbb5f47),
	.w7(32'h3c3812c2),
	.w8(32'h3bab2d4c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aaa26),
	.w1(32'hbb9cb01a),
	.w2(32'h3b2a7e63),
	.w3(32'hbbab1d2e),
	.w4(32'hb98d0d49),
	.w5(32'hbbc1cabd),
	.w6(32'hbab53e73),
	.w7(32'hbc17c5dc),
	.w8(32'hb8f3b1a5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc452e7c),
	.w1(32'hb9941e8f),
	.w2(32'hbb4b0cb5),
	.w3(32'hbab51d34),
	.w4(32'hbb32741a),
	.w5(32'hbb1aed5d),
	.w6(32'hbb587153),
	.w7(32'hbbeedbf8),
	.w8(32'hbbbe8edd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954d98),
	.w1(32'hbb02a9c3),
	.w2(32'hbb2f9b2b),
	.w3(32'hbac7be37),
	.w4(32'hbb9ab202),
	.w5(32'hbb8f488b),
	.w6(32'hbb710c7f),
	.w7(32'hbc12347a),
	.w8(32'hbbc5dcbe),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87dbc8),
	.w1(32'h3bf9f2ab),
	.w2(32'h3c03e562),
	.w3(32'hbbd8cdcf),
	.w4(32'h3be41b6a),
	.w5(32'h3c8759e6),
	.w6(32'hbb88e972),
	.w7(32'hbc8230cb),
	.w8(32'hbc0df6c9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0547ee),
	.w1(32'h3ad11fe2),
	.w2(32'h392220d4),
	.w3(32'h3b6ab9a5),
	.w4(32'h3bbe3c02),
	.w5(32'hbb4471b6),
	.w6(32'h3b65378c),
	.w7(32'h3c0a3ceb),
	.w8(32'hba3b3ab8),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81433d),
	.w1(32'hbc06bd16),
	.w2(32'hba979076),
	.w3(32'hbb22ba88),
	.w4(32'hbc4677f0),
	.w5(32'hbbde9395),
	.w6(32'h3c12e3c6),
	.w7(32'h39873990),
	.w8(32'hbc2f2e45),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52991c),
	.w1(32'h3b8bcbc9),
	.w2(32'h3b9f5023),
	.w3(32'h3b70e9f4),
	.w4(32'hbadb0052),
	.w5(32'h3a34d798),
	.w6(32'h3ba91a92),
	.w7(32'hba3753e2),
	.w8(32'hb8d5b7ad),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75bb32),
	.w1(32'h39703fd7),
	.w2(32'hbb5ff2f0),
	.w3(32'hbb2174c3),
	.w4(32'h3b562e14),
	.w5(32'hbba8afba),
	.w6(32'h3b8e3914),
	.w7(32'h3ad88c2a),
	.w8(32'h3b804213),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3056b4),
	.w1(32'hbb5c3197),
	.w2(32'hbbaa260c),
	.w3(32'hbbd22066),
	.w4(32'hbb428158),
	.w5(32'hbbcae236),
	.w6(32'hba307f08),
	.w7(32'h3b1e3967),
	.w8(32'h3acde9f7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba777f9d),
	.w1(32'hb7f3d252),
	.w2(32'hbb450d4f),
	.w3(32'hb9f2151c),
	.w4(32'h3b02cf0c),
	.w5(32'h3a8080c3),
	.w6(32'hba96097a),
	.w7(32'hbb46232c),
	.w8(32'hbb86836a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acff4e6),
	.w1(32'hbb3288cb),
	.w2(32'hbb3896c8),
	.w3(32'h3bb79fbc),
	.w4(32'hbb7654a6),
	.w5(32'hbbb8c718),
	.w6(32'hbac038a5),
	.w7(32'hbaf71fc3),
	.w8(32'hbbfc3b5a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a2226),
	.w1(32'h3b3fc8c0),
	.w2(32'h3b968866),
	.w3(32'h39057b3b),
	.w4(32'h3b44ad8d),
	.w5(32'h3c4c6ffe),
	.w6(32'h39bf4087),
	.w7(32'hbbb7cb19),
	.w8(32'hbb20b900),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39bd2b),
	.w1(32'hbc0d2cf2),
	.w2(32'hb9d8d4d6),
	.w3(32'h3bd1602a),
	.w4(32'hbbaa875c),
	.w5(32'hbbdf330e),
	.w6(32'h39cdf02d),
	.w7(32'h3c4cda5c),
	.w8(32'hbb8fefd5),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2219fb),
	.w1(32'hbace2fc3),
	.w2(32'h3bb56957),
	.w3(32'hbbba2bec),
	.w4(32'hba914f6f),
	.w5(32'h3c37754b),
	.w6(32'hbc0fdc33),
	.w7(32'hbc82513d),
	.w8(32'hbc0e5cea),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c89bf),
	.w1(32'hbbbd42b6),
	.w2(32'hbb1ba7f8),
	.w3(32'h3b5e25fa),
	.w4(32'hbb580167),
	.w5(32'hbc244a7e),
	.w6(32'h39bde96c),
	.w7(32'h3c7895e2),
	.w8(32'h3b09343c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4d33e),
	.w1(32'h3ba59046),
	.w2(32'h3c032deb),
	.w3(32'hbaeae43a),
	.w4(32'h3bfe4d6a),
	.w5(32'h3c8225a4),
	.w6(32'hbb6f393e),
	.w7(32'hbc186e81),
	.w8(32'hbb0e6d82),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c8115),
	.w1(32'h3c0d8446),
	.w2(32'h3b228590),
	.w3(32'h3b9f819b),
	.w4(32'h3c5aa21b),
	.w5(32'hbaccda2d),
	.w6(32'h3bb8869e),
	.w7(32'h3c0ca41b),
	.w8(32'h3b5e6ae8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebe628),
	.w1(32'hbc2fe519),
	.w2(32'hbbdabbe0),
	.w3(32'h3ab33b5c),
	.w4(32'hbb9a5a4f),
	.w5(32'hbc4adbfc),
	.w6(32'h3c59fd54),
	.w7(32'h3d04be68),
	.w8(32'h3c6e52dd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ed63),
	.w1(32'hbbb2f9b4),
	.w2(32'hbb5540b4),
	.w3(32'hbb06a45e),
	.w4(32'hbb1e8a1d),
	.w5(32'hbbe93029),
	.w6(32'hbb0b7cd4),
	.w7(32'h3c19c340),
	.w8(32'h3be96299),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad04bd8),
	.w1(32'h3abae740),
	.w2(32'h3b21124f),
	.w3(32'hbb52868e),
	.w4(32'h3adbac28),
	.w5(32'h3c467993),
	.w6(32'h3a9a57d8),
	.w7(32'hbb2bbdfe),
	.w8(32'h3b10a501),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe9a7),
	.w1(32'h3aa4aa34),
	.w2(32'h39138dc2),
	.w3(32'h3b5e5639),
	.w4(32'h3b05d150),
	.w5(32'h3b42082f),
	.w6(32'hb8e8aa1e),
	.w7(32'hbad1f567),
	.w8(32'hbb618dbd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60ebd3),
	.w1(32'hba8237f5),
	.w2(32'hbc0bc570),
	.w3(32'h3b908364),
	.w4(32'h3a888094),
	.w5(32'hbb69f8dc),
	.w6(32'hbb2932b6),
	.w7(32'hbc363b0c),
	.w8(32'hbbc23820),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82277a),
	.w1(32'h3b58d68b),
	.w2(32'h3bcdc601),
	.w3(32'h3a099c66),
	.w4(32'hbb97a073),
	.w5(32'h38d64afd),
	.w6(32'hb9a0720b),
	.w7(32'hbc14a816),
	.w8(32'hbbbd954a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77ae3d),
	.w1(32'hba5b5282),
	.w2(32'hbb92c1ef),
	.w3(32'hbbe01082),
	.w4(32'h3ba4cf5f),
	.w5(32'h3b9289c2),
	.w6(32'h3b302b81),
	.w7(32'h3b9eceab),
	.w8(32'hbabd1bb1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfba87e),
	.w1(32'hbbfb1ac3),
	.w2(32'hbb6cfad1),
	.w3(32'hba8bbca1),
	.w4(32'hbbd7e8f0),
	.w5(32'hbc59ae91),
	.w6(32'h3bd3703f),
	.w7(32'h3c98a88b),
	.w8(32'h3b6f2598),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb753cf5),
	.w1(32'hb98d56de),
	.w2(32'h3b3c26e4),
	.w3(32'hbbb761b5),
	.w4(32'hbaf3bb8f),
	.w5(32'h3b8623ea),
	.w6(32'hbba94416),
	.w7(32'hbc48e530),
	.w8(32'hbbcc0bbc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb395466),
	.w1(32'h3a827333),
	.w2(32'h3bb933e4),
	.w3(32'hbb9315e2),
	.w4(32'h388ee2cc),
	.w5(32'h3c014248),
	.w6(32'hbb9c68bf),
	.w7(32'hbc42f8de),
	.w8(32'hbbf25e59),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06815d),
	.w1(32'hbbe7085f),
	.w2(32'hbba2b880),
	.w3(32'h3a47d16f),
	.w4(32'hbc2798a8),
	.w5(32'hbc0fad47),
	.w6(32'hbbee55c1),
	.w7(32'hbc6bc6ea),
	.w8(32'hbc1134ea),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6bc7),
	.w1(32'hbc09ee91),
	.w2(32'hbbae7728),
	.w3(32'hbc44b6fc),
	.w4(32'hbb98a5e4),
	.w5(32'hbbf5d27c),
	.w6(32'hbb3d537b),
	.w7(32'h3be52f58),
	.w8(32'hbb06809b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42177c),
	.w1(32'h3a648e29),
	.w2(32'h3ba727d2),
	.w3(32'hba56e9d3),
	.w4(32'h3b517186),
	.w5(32'hbc34e085),
	.w6(32'h3bf6b426),
	.w7(32'h3b354b22),
	.w8(32'h3b06d3fe),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8544e),
	.w1(32'h3b365bc2),
	.w2(32'h3b2a5833),
	.w3(32'h3beaa7a9),
	.w4(32'h3bec0d04),
	.w5(32'h3ca617ac),
	.w6(32'hbbc611e0),
	.w7(32'hbca0c30c),
	.w8(32'hbc1dee50),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94ced6),
	.w1(32'hba078d12),
	.w2(32'h3b013a43),
	.w3(32'h3b9debb4),
	.w4(32'hbae5f7ca),
	.w5(32'hbc1a1c40),
	.w6(32'h3b0d60c7),
	.w7(32'h3c53d87c),
	.w8(32'h3a036b48),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4faeaf),
	.w1(32'hb9236a10),
	.w2(32'h3b8b00c1),
	.w3(32'hb9b41dad),
	.w4(32'hbba863ee),
	.w5(32'hbbc0b79f),
	.w6(32'hbb41415c),
	.w7(32'hbb404952),
	.w8(32'hbb34ce7e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cb3aa),
	.w1(32'hb75c1cb3),
	.w2(32'hbb0d2c81),
	.w3(32'hbb24f07c),
	.w4(32'h3a9fc0c4),
	.w5(32'h3bcdb1bb),
	.w6(32'hbbccdf87),
	.w7(32'hbc7b89b3),
	.w8(32'hbba74ab7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d766f),
	.w1(32'hbb38702d),
	.w2(32'hbc0c646b),
	.w3(32'hbad10e36),
	.w4(32'hba37e0a9),
	.w5(32'hbb965543),
	.w6(32'hbba2dc05),
	.w7(32'hbc4e2096),
	.w8(32'hbc09370c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9045c8),
	.w1(32'hbb1d7875),
	.w2(32'hb9b7b861),
	.w3(32'h3a32ef9e),
	.w4(32'hbb058754),
	.w5(32'hbc1202c4),
	.w6(32'hbaa04e77),
	.w7(32'h3c09703b),
	.w8(32'h3a95f2d1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336e66),
	.w1(32'hbb8b5c49),
	.w2(32'hbb576758),
	.w3(32'hbb7f90d2),
	.w4(32'hbb3cad86),
	.w5(32'hba86251f),
	.w6(32'h38f6caaa),
	.w7(32'hb96f389a),
	.w8(32'hbaa80a86),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0222ee),
	.w1(32'hbbd67e0a),
	.w2(32'hbaf19ea1),
	.w3(32'h3ae84a79),
	.w4(32'hbbbca342),
	.w5(32'hbc12af73),
	.w6(32'hbb9c3281),
	.w7(32'h3b95288d),
	.w8(32'hbbaf162d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8625c0),
	.w1(32'h3b919edb),
	.w2(32'hbb2ea95d),
	.w3(32'hbbacfd31),
	.w4(32'hbb2692bd),
	.w5(32'hbb9b9a46),
	.w6(32'hb9f04fa4),
	.w7(32'hbc1bab04),
	.w8(32'hbbb85544),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f05c0e),
	.w1(32'hbb232652),
	.w2(32'h3a716a70),
	.w3(32'hbb096689),
	.w4(32'h3a14c623),
	.w5(32'hb80e5e68),
	.w6(32'h39b50e11),
	.w7(32'h3a8d5ece),
	.w8(32'hbb911a4c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a939e6f),
	.w1(32'hba1a9add),
	.w2(32'h3a9f5a45),
	.w3(32'h3ba32e6c),
	.w4(32'hbbc8f3a8),
	.w5(32'hbc1c3660),
	.w6(32'h3797d055),
	.w7(32'h3a89c36c),
	.w8(32'hbbdf2b1b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bae10),
	.w1(32'hbacb2fb5),
	.w2(32'hbb103079),
	.w3(32'hbb11ceec),
	.w4(32'hbad1d54a),
	.w5(32'h3aade41b),
	.w6(32'hbb928897),
	.w7(32'hbc26ae3c),
	.w8(32'hbba29b3c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f490b),
	.w1(32'h3a92252a),
	.w2(32'hba222073),
	.w3(32'hbadd049f),
	.w4(32'h393b2689),
	.w5(32'hbb4b2e20),
	.w6(32'h3b3be076),
	.w7(32'h3b991046),
	.w8(32'h3ac39480),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a946d),
	.w1(32'h395b37c3),
	.w2(32'hba99046b),
	.w3(32'h3a77816b),
	.w4(32'hb700cb1a),
	.w5(32'h3b10f74c),
	.w6(32'hbbb52269),
	.w7(32'hbc772baf),
	.w8(32'hbbe0a546),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76d147),
	.w1(32'hbc1c16fa),
	.w2(32'hbc045001),
	.w3(32'hbb229fc7),
	.w4(32'hbbe6322a),
	.w5(32'hbb563b94),
	.w6(32'hbbcaf0c0),
	.w7(32'hbc44160e),
	.w8(32'hbbe16d86),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc125ad1),
	.w1(32'hbbdde6f2),
	.w2(32'hbc18c805),
	.w3(32'hbbf9eca2),
	.w4(32'hbbe041b3),
	.w5(32'hbc7f94ca),
	.w6(32'h3bb9b65a),
	.w7(32'h3c826ff5),
	.w8(32'h3bb5644c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb976),
	.w1(32'hbb38d775),
	.w2(32'h3ac3df5d),
	.w3(32'hbc0211cc),
	.w4(32'hbb5c7125),
	.w5(32'hbc0e1489),
	.w6(32'h3baf0952),
	.w7(32'h3c40204b),
	.w8(32'h3bdcf73c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c69ee),
	.w1(32'hbb4c356c),
	.w2(32'hbc202a53),
	.w3(32'hbadd2875),
	.w4(32'hb9a8fc7f),
	.w5(32'hbbd14158),
	.w6(32'hbb9386f7),
	.w7(32'hbc4347fc),
	.w8(32'hbbdc0f55),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b158c),
	.w1(32'hbbfb18e5),
	.w2(32'hbbf9253b),
	.w3(32'h3a29540b),
	.w4(32'hbaa40f8e),
	.w5(32'hbb9a700a),
	.w6(32'hbbbe037b),
	.w7(32'h3ad8bff5),
	.w8(32'hbb252228),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe85d90),
	.w1(32'h39b2aae7),
	.w2(32'h3c1d3c49),
	.w3(32'hbb0b7705),
	.w4(32'hbb95c5cc),
	.w5(32'hbb5b2137),
	.w6(32'h3bcbcdbe),
	.w7(32'h3c1bfb60),
	.w8(32'h3b1b5ed8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878a5f),
	.w1(32'h3b24b081),
	.w2(32'hbb499d34),
	.w3(32'hbb31f790),
	.w4(32'h3a91dc9c),
	.w5(32'h39c036b0),
	.w6(32'hba85c890),
	.w7(32'hbb655968),
	.w8(32'hb7110929),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6f6be),
	.w1(32'hbbdf6075),
	.w2(32'h3b91ba22),
	.w3(32'hbbcb3dcd),
	.w4(32'hbbb650df),
	.w5(32'h3ae796b0),
	.w6(32'h399005d4),
	.w7(32'h3c23b840),
	.w8(32'hbc087ca0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c0299),
	.w1(32'hbbcc4e5a),
	.w2(32'hb95d2000),
	.w3(32'h3b7e3b7e),
	.w4(32'hbb0439d5),
	.w5(32'hbc281b96),
	.w6(32'h3997a4a5),
	.w7(32'h3c5c84fe),
	.w8(32'h3abf7ba3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46825f),
	.w1(32'hbb61f95b),
	.w2(32'hbb9feed3),
	.w3(32'hbb8a6383),
	.w4(32'hbb90e337),
	.w5(32'hbbb433d3),
	.w6(32'h3afcceca),
	.w7(32'h3a991ba4),
	.w8(32'hba9bc47e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebccc3),
	.w1(32'h3a00ccd5),
	.w2(32'hba03cca6),
	.w3(32'hbace56cc),
	.w4(32'hbb5a4352),
	.w5(32'hbbd8b906),
	.w6(32'hbaab4fbf),
	.w7(32'h3bb2def7),
	.w8(32'h3ba2e21e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0240),
	.w1(32'h3b87ace2),
	.w2(32'hba90cf6e),
	.w3(32'hbbfb8f55),
	.w4(32'h3b3b7316),
	.w5(32'hbbc8689d),
	.w6(32'h3b8f7a73),
	.w7(32'hbb59e496),
	.w8(32'h3c211eab),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa06e),
	.w1(32'h3b83d4b0),
	.w2(32'h3b917e2d),
	.w3(32'hbbfaf870),
	.w4(32'h3c10fa11),
	.w5(32'h3d044838),
	.w6(32'hbc4310c6),
	.w7(32'hbd05f9ee),
	.w8(32'hbc772ffc),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb7fc4),
	.w1(32'h3adcee18),
	.w2(32'h3b9a8a54),
	.w3(32'h3be56ad5),
	.w4(32'hbac56ba5),
	.w5(32'h3bbb7309),
	.w6(32'hbb9b7448),
	.w7(32'hbc3db8a4),
	.w8(32'hbbe82e38),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf03a68),
	.w1(32'h3b00e1a5),
	.w2(32'h3b2dfb08),
	.w3(32'hbb6dcd43),
	.w4(32'h3b9c62bc),
	.w5(32'h3c7d3f51),
	.w6(32'hbb965917),
	.w7(32'hbc671753),
	.w8(32'hbbcfb97d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eb30d),
	.w1(32'h3aaa9efa),
	.w2(32'h39c90678),
	.w3(32'h3b4bd6bc),
	.w4(32'hba8fe30f),
	.w5(32'h3a9e233c),
	.w6(32'hbba6c40d),
	.w7(32'hbc055822),
	.w8(32'hbba841de),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0fdee),
	.w1(32'hbbfd0afa),
	.w2(32'hbc49ba47),
	.w3(32'hbae20e56),
	.w4(32'h3a48a821),
	.w5(32'hbbbcc189),
	.w6(32'hbb482aca),
	.w7(32'h3b8c3606),
	.w8(32'hb9f51e6b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe512fe),
	.w1(32'hbbe1e864),
	.w2(32'hbc0db70e),
	.w3(32'hba4800d6),
	.w4(32'hbb8ed3f2),
	.w5(32'h372b8f39),
	.w6(32'hbbd12047),
	.w7(32'hbc69cae0),
	.w8(32'hbc102869),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc022438),
	.w1(32'h3b2dd1af),
	.w2(32'h3b27bf8b),
	.w3(32'hbb229744),
	.w4(32'h3bb9d649),
	.w5(32'h3c8bec45),
	.w6(32'hbbb8dee8),
	.w7(32'hbc8877f9),
	.w8(32'hbbfa658f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb730dd3),
	.w1(32'hbadf4bf2),
	.w2(32'hbb3c0463),
	.w3(32'h3b748a43),
	.w4(32'h3a8b59ac),
	.w5(32'hbc183430),
	.w6(32'h3b74a6c2),
	.w7(32'h3bdaa59a),
	.w8(32'hba817553),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51324b),
	.w1(32'hba8b08d7),
	.w2(32'h3b0926e2),
	.w3(32'hbbcaafac),
	.w4(32'hbbb99504),
	.w5(32'h3b495f60),
	.w6(32'hbb0a07f6),
	.w7(32'hbc0d4c99),
	.w8(32'hbbea865f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b3ff),
	.w1(32'h3bab5014),
	.w2(32'h3b990381),
	.w3(32'hb824458c),
	.w4(32'h3c2fdb55),
	.w5(32'h3bab596e),
	.w6(32'h3bd60833),
	.w7(32'h3b032587),
	.w8(32'h3b4c31f9),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a896450),
	.w1(32'hb9cb3a8e),
	.w2(32'h3b551046),
	.w3(32'h3bf8f261),
	.w4(32'hbbbda3c9),
	.w5(32'h3ac1a726),
	.w6(32'h3807577c),
	.w7(32'hbbed8a73),
	.w8(32'hbb6a7acf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104e8d),
	.w1(32'hbc094f0e),
	.w2(32'hbc04eaaa),
	.w3(32'hbb93ff34),
	.w4(32'hb71a53d1),
	.w5(32'hbb5b7e25),
	.w6(32'hb9da6b59),
	.w7(32'h3bc283d9),
	.w8(32'hbb29054a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ef319),
	.w1(32'h3ae7e433),
	.w2(32'hbae044c8),
	.w3(32'hbb0e30c0),
	.w4(32'hb8d788e3),
	.w5(32'h3ba3053c),
	.w6(32'hbc3e4582),
	.w7(32'hbc9ded67),
	.w8(32'hbc08ffc4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02750),
	.w1(32'h3b69837d),
	.w2(32'h3b80341e),
	.w3(32'h3a15cd94),
	.w4(32'h3bfc71eb),
	.w5(32'h3cc37fcf),
	.w6(32'hbbf4d378),
	.w7(32'hbcb860d5),
	.w8(32'hbc2acbb2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa14d3),
	.w1(32'h3a59426a),
	.w2(32'h3b511f95),
	.w3(32'h3bb45218),
	.w4(32'h3af68a9e),
	.w5(32'h3c287ab0),
	.w6(32'hbbcb0962),
	.w7(32'hbc5257f5),
	.w8(32'hbbeadd3d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0130a2),
	.w1(32'h3abf2040),
	.w2(32'h3b4baf02),
	.w3(32'h3a70d5d3),
	.w4(32'h3b10d5c3),
	.w5(32'h3c469276),
	.w6(32'hbb9b0076),
	.w7(32'hbc3f3011),
	.w8(32'hbba770a3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0717b),
	.w1(32'h3a3fdf66),
	.w2(32'h3c38804a),
	.w3(32'h3af32768),
	.w4(32'h3b708cbb),
	.w5(32'h3c35471d),
	.w6(32'h3ab9be45),
	.w7(32'hba8b9033),
	.w8(32'h3a97bd7d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b784981),
	.w1(32'hbb07b007),
	.w2(32'h3ba502e4),
	.w3(32'h3c0e4954),
	.w4(32'hbb8efa5c),
	.w5(32'hb8d43841),
	.w6(32'h3bb5cc9c),
	.w7(32'h3c800f52),
	.w8(32'h3adac716),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff4f1b),
	.w1(32'hbb61841c),
	.w2(32'hbbbf1a6a),
	.w3(32'hbb512291),
	.w4(32'hbc050269),
	.w5(32'hbbe9776d),
	.w6(32'hbbd66f50),
	.w7(32'hbbf439e3),
	.w8(32'hbbc02a7f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc257),
	.w1(32'hbac68ee3),
	.w2(32'hbb192980),
	.w3(32'hbc251e5e),
	.w4(32'hbb559e23),
	.w5(32'h3a8c1352),
	.w6(32'hbb86b8bb),
	.w7(32'hbb82206b),
	.w8(32'hbb30863b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9963c1c),
	.w1(32'h3b472053),
	.w2(32'h3bdcd786),
	.w3(32'hb7ac44e9),
	.w4(32'h3b1a57b6),
	.w5(32'h3c50dd43),
	.w6(32'hbbf474ca),
	.w7(32'hbc88ebda),
	.w8(32'hbc209478),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff4382),
	.w1(32'h3b09fc7b),
	.w2(32'h3c8d58d2),
	.w3(32'h3aae9509),
	.w4(32'hbaa295d9),
	.w5(32'h3bce7538),
	.w6(32'h3c0ec694),
	.w7(32'hba704727),
	.w8(32'h394852ed),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8612dd),
	.w1(32'h3b4c4122),
	.w2(32'h3c185654),
	.w3(32'h3bca0838),
	.w4(32'h39103bce),
	.w5(32'h3b67a6ec),
	.w6(32'h3baf51fb),
	.w7(32'h3b3d6345),
	.w8(32'h3a640b49),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fe9c4),
	.w1(32'hbb9e9ff9),
	.w2(32'hbbd3b3dc),
	.w3(32'hbb81abb1),
	.w4(32'hbb502531),
	.w5(32'h3a63da35),
	.w6(32'hbc06acff),
	.w7(32'hbc6395ce),
	.w8(32'hbbc58827),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17890),
	.w1(32'hb6c69e46),
	.w2(32'h38ab21a1),
	.w3(32'hbb9fddae),
	.w4(32'h389c870c),
	.w5(32'h3937922f),
	.w6(32'h38982c21),
	.w7(32'h39222a25),
	.w8(32'h3937bf80),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fbef2),
	.w1(32'h38dd4e55),
	.w2(32'h39a45656),
	.w3(32'h3a1f0cab),
	.w4(32'h3a8e4dff),
	.w5(32'h3a710aff),
	.w6(32'hba239b7d),
	.w7(32'hba5b6736),
	.w8(32'hbac91c30),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule