module layer_10_featuremap_12(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83537),
	.w1(32'h3c6789eb),
	.w2(32'hbbb3a9c7),
	.w3(32'hbc3009d5),
	.w4(32'h3caf9135),
	.w5(32'hbc536501),
	.w6(32'hbc5aa6c4),
	.w7(32'h3c22ca49),
	.w8(32'h38c6f90a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943b3fe),
	.w1(32'h3b60e320),
	.w2(32'hbc7026d6),
	.w3(32'hbca0e121),
	.w4(32'h3be09a78),
	.w5(32'hbbfbbb46),
	.w6(32'hbc3fb542),
	.w7(32'h3a449efe),
	.w8(32'hbc7410ef),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75ca64),
	.w1(32'hbc9d17b5),
	.w2(32'hbbf42a5a),
	.w3(32'hbcbcdb22),
	.w4(32'hbcc1977d),
	.w5(32'hbbd106c9),
	.w6(32'hbca01615),
	.w7(32'hbcb7c528),
	.w8(32'hbb1e32c9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb401bd9),
	.w1(32'hba8676fe),
	.w2(32'hbc0e9559),
	.w3(32'hbbffdea7),
	.w4(32'hbbb03fb2),
	.w5(32'hbc8bc3d0),
	.w6(32'h3b18b329),
	.w7(32'h3a9c3331),
	.w8(32'hbc986129),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ad64),
	.w1(32'hbb072ee4),
	.w2(32'hbc80bf50),
	.w3(32'hbc43a777),
	.w4(32'hbbee2dcd),
	.w5(32'hbd02c2c7),
	.w6(32'hbbbebf7a),
	.w7(32'h3b155e31),
	.w8(32'hbcaa2280),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfaeac9),
	.w1(32'hbb69ab52),
	.w2(32'hbb83ba53),
	.w3(32'hbd0e262c),
	.w4(32'hbc599c52),
	.w5(32'hbbf05a9a),
	.w6(32'hbcf8ecd1),
	.w7(32'h3bc664fb),
	.w8(32'hbac5206b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7a74),
	.w1(32'hbb5028db),
	.w2(32'h3c2afa4e),
	.w3(32'hbbf8334b),
	.w4(32'h3aeeeb59),
	.w5(32'h3b00fc5d),
	.w6(32'hb9abf67c),
	.w7(32'h3b9d0612),
	.w8(32'h3bc0596c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e915d),
	.w1(32'h3c2edc2e),
	.w2(32'hba8b067f),
	.w3(32'hba87ba87),
	.w4(32'h3c688637),
	.w5(32'h3bbe878e),
	.w6(32'h3bbcc584),
	.w7(32'h3c51614a),
	.w8(32'h3c0aa8f4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39834222),
	.w1(32'h3c09ca9e),
	.w2(32'hbaeef0f1),
	.w3(32'hba34539c),
	.w4(32'hba1b8594),
	.w5(32'hba2b93ab),
	.w6(32'h3b80202f),
	.w7(32'hbba2f89e),
	.w8(32'hb7af20e7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9aca),
	.w1(32'hbb91cc88),
	.w2(32'h3b837bf2),
	.w3(32'h3bda5b7d),
	.w4(32'hbc588948),
	.w5(32'h3bdb4f55),
	.w6(32'h3b293c6f),
	.w7(32'hbcabce74),
	.w8(32'h3c0ecbef),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d2cb5),
	.w1(32'hbaa38688),
	.w2(32'hba4570da),
	.w3(32'h3b721eb9),
	.w4(32'h3b5ee04e),
	.w5(32'hbbe9e1e7),
	.w6(32'h3b0386ab),
	.w7(32'h3a48d119),
	.w8(32'hbbefaea7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3109f2),
	.w1(32'h39d2105d),
	.w2(32'h3a9a7866),
	.w3(32'hbbe88e95),
	.w4(32'h3b84dd2f),
	.w5(32'h3b1a1f95),
	.w6(32'hbb85447e),
	.w7(32'hbb5e2d5e),
	.w8(32'h3b111502),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c111010),
	.w1(32'h3bbb7db5),
	.w2(32'hb862cd88),
	.w3(32'h3b8b1b6c),
	.w4(32'h3ac427e8),
	.w5(32'h3c2a4abe),
	.w6(32'h39d74896),
	.w7(32'hbad1c003),
	.w8(32'h3b66aafa),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c2a20),
	.w1(32'hbbbb70be),
	.w2(32'hbbcde118),
	.w3(32'h3c04b770),
	.w4(32'hbabb9216),
	.w5(32'hbcb3642c),
	.w6(32'h3aca08df),
	.w7(32'hbb3d2909),
	.w8(32'hbc893e5a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2df4ac),
	.w1(32'h3ab4231f),
	.w2(32'h367815c8),
	.w3(32'hbc880e08),
	.w4(32'hbc92f966),
	.w5(32'h3ba6d335),
	.w6(32'hbbb6b29b),
	.w7(32'h39f7089c),
	.w8(32'h3bff6750),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6389d),
	.w1(32'h3b6899b1),
	.w2(32'hbabf0f8c),
	.w3(32'h3b4ff931),
	.w4(32'hb880c508),
	.w5(32'h3a635082),
	.w6(32'hbaae84cf),
	.w7(32'h3ada7c9b),
	.w8(32'h3bc844f1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac43d13),
	.w1(32'h3b0d8b9c),
	.w2(32'h3c1c0400),
	.w3(32'h3b5069cf),
	.w4(32'h3bd0662b),
	.w5(32'h3c605653),
	.w6(32'h3b183e23),
	.w7(32'h3b941f0f),
	.w8(32'h3c0bb3cc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a79aa),
	.w1(32'h3c27c9c7),
	.w2(32'hbb7e1134),
	.w3(32'h3c8013bd),
	.w4(32'h3c5ac90b),
	.w5(32'h3b995f2b),
	.w6(32'h3b07e85a),
	.w7(32'hb9aa635d),
	.w8(32'h3bb2d925),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb8310),
	.w1(32'hba350270),
	.w2(32'hbc9de279),
	.w3(32'h3beec7eb),
	.w4(32'hbb57e438),
	.w5(32'hbc818268),
	.w6(32'h3b678e2e),
	.w7(32'h3a96675c),
	.w8(32'hbb03ba08),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48d7eb),
	.w1(32'h3b0a4496),
	.w2(32'h3b1ed051),
	.w3(32'hbcae1ada),
	.w4(32'hbc6f20bb),
	.w5(32'hbb8035f0),
	.w6(32'hbc2db379),
	.w7(32'hbc44b42f),
	.w8(32'hbb0c0b4f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca10ba),
	.w1(32'h3ad0da36),
	.w2(32'hbbb624e2),
	.w3(32'hbb8dd0a2),
	.w4(32'h39ba57a1),
	.w5(32'h3bddbadf),
	.w6(32'h3aa8b770),
	.w7(32'h3baf2c93),
	.w8(32'h3c45081b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c026267),
	.w1(32'h3c2365e5),
	.w2(32'hbc2e4d47),
	.w3(32'h3c044951),
	.w4(32'h3bb7334c),
	.w5(32'hbc2369d6),
	.w6(32'h3c5f790a),
	.w7(32'h3abc9b75),
	.w8(32'hbc103df7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ae94),
	.w1(32'h3b9dc8b2),
	.w2(32'h3a2807a9),
	.w3(32'h3aa9d2a9),
	.w4(32'h3be0ed93),
	.w5(32'h3b74a821),
	.w6(32'h3c75b27e),
	.w7(32'h3c64d2f4),
	.w8(32'h3bd2bb47),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe3436),
	.w1(32'h3a64b946),
	.w2(32'h3bee252f),
	.w3(32'h3bd34415),
	.w4(32'h3abadd6a),
	.w5(32'h3c464463),
	.w6(32'h3b6fea5a),
	.w7(32'h3ab6cd68),
	.w8(32'h3bd71a90),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c435d08),
	.w1(32'h3af02dc9),
	.w2(32'hbc89712b),
	.w3(32'h3c0101d1),
	.w4(32'h3a9630a0),
	.w5(32'hbb4ccea0),
	.w6(32'h3c067227),
	.w7(32'h3b9e34fd),
	.w8(32'h3921ec57),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b43b3),
	.w1(32'h3aa71f34),
	.w2(32'h3a7ee5aa),
	.w3(32'hbb90ac03),
	.w4(32'hbc09236d),
	.w5(32'hbb2c3d6c),
	.w6(32'hba7591be),
	.w7(32'h3b29cf3e),
	.w8(32'hbb78886f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba2a79),
	.w1(32'hb96ef73d),
	.w2(32'hba1da1cb),
	.w3(32'hb8ca73af),
	.w4(32'h3b25b127),
	.w5(32'hba3a2fda),
	.w6(32'hbab9af3b),
	.w7(32'h3b64448f),
	.w8(32'h3a511a47),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4130ce),
	.w1(32'h3b3121e2),
	.w2(32'hbc946e5e),
	.w3(32'hbb3d613a),
	.w4(32'h3b252d01),
	.w5(32'hbc99762f),
	.w6(32'h3b130e40),
	.w7(32'h3c050c56),
	.w8(32'hbbd7c2d3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d4ab8),
	.w1(32'hbad2fd97),
	.w2(32'hbbd0a059),
	.w3(32'hbc49a364),
	.w4(32'h3bb37dd9),
	.w5(32'hbc0e0f71),
	.w6(32'hbba19170),
	.w7(32'h3c3848ba),
	.w8(32'hbc03c08d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30f29),
	.w1(32'h3a99c27f),
	.w2(32'hbc19c65f),
	.w3(32'hbc76725d),
	.w4(32'hba90f227),
	.w5(32'hbc2f7903),
	.w6(32'hbbd36911),
	.w7(32'h3afe95e5),
	.w8(32'hbad445d6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0325fd),
	.w1(32'h39785d7c),
	.w2(32'h3bb87641),
	.w3(32'hbc174a95),
	.w4(32'hba4ccc58),
	.w5(32'h3bb6ea6e),
	.w6(32'hbbee6527),
	.w7(32'hbb338eaa),
	.w8(32'h3b4ea741),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980f6f),
	.w1(32'hbb136d1e),
	.w2(32'hbaa805ac),
	.w3(32'h3b299c83),
	.w4(32'h3a5a97a9),
	.w5(32'h3c4fc5a3),
	.w6(32'h3c88744c),
	.w7(32'h3c35088a),
	.w8(32'h3c074f94),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034e38),
	.w1(32'h3c1ac481),
	.w2(32'h3c349200),
	.w3(32'h3b8164b8),
	.w4(32'hba925993),
	.w5(32'h3c6365bd),
	.w6(32'h3c48d98a),
	.w7(32'h3bc2c583),
	.w8(32'h3b25febf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c608894),
	.w1(32'h3a5a129b),
	.w2(32'h3a3c6917),
	.w3(32'h3c38115e),
	.w4(32'hbb364ad4),
	.w5(32'h3bf876cf),
	.w6(32'hba004e68),
	.w7(32'hbc3a6627),
	.w8(32'h3ba60a2a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab31099),
	.w1(32'h3b193ee5),
	.w2(32'h3c7dfa06),
	.w3(32'h3b8619e8),
	.w4(32'hbb0934ab),
	.w5(32'h3c9437ee),
	.w6(32'h3984df3a),
	.w7(32'hbb917141),
	.w8(32'h3ba36ebb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bbbb6),
	.w1(32'hba8b4619),
	.w2(32'hbbdb7cf7),
	.w3(32'h3c13b1ca),
	.w4(32'hbb13d12e),
	.w5(32'hbc923c7c),
	.w6(32'hb9e4abf9),
	.w7(32'hbc3ab0d0),
	.w8(32'hbc285f7c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcef816b),
	.w1(32'hbcaa6639),
	.w2(32'hbc30c5b8),
	.w3(32'hbc98f6d0),
	.w4(32'hbc4aa6ef),
	.w5(32'hbbac9b4e),
	.w6(32'h3a872a7b),
	.w7(32'hbc795750),
	.w8(32'h3c05cd69),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51140a),
	.w1(32'hbc179d30),
	.w2(32'hbc219601),
	.w3(32'hbc781bef),
	.w4(32'hbc6f412c),
	.w5(32'hbc9ff4e0),
	.w6(32'h3ae8bb10),
	.w7(32'hbb3268a4),
	.w8(32'hbbedf869),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe95dd),
	.w1(32'hbc8d4acb),
	.w2(32'hbbd36e69),
	.w3(32'hbc9307d8),
	.w4(32'hbc80660b),
	.w5(32'hbb91c346),
	.w6(32'hbb8f1228),
	.w7(32'h3b021aa7),
	.w8(32'hb9bb3b1a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f0c9b),
	.w1(32'hbc30faf2),
	.w2(32'hbb0e432e),
	.w3(32'hbc70b8bb),
	.w4(32'hbca9e1bb),
	.w5(32'h3acc62d1),
	.w6(32'hbc1f93cc),
	.w7(32'hbc6b6fc5),
	.w8(32'hbbe4efc7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0700a8),
	.w1(32'hbbe3fcd9),
	.w2(32'h3bf5b703),
	.w3(32'hbac402fb),
	.w4(32'hbc520474),
	.w5(32'h3b2cde89),
	.w6(32'hbc7c7405),
	.w7(32'hbc9bbe03),
	.w8(32'h3bd8daff),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c4c6b),
	.w1(32'hbb8de29a),
	.w2(32'h3c0f1a46),
	.w3(32'hbbfef93a),
	.w4(32'hbc209e07),
	.w5(32'h3bbe049a),
	.w6(32'hbb69f164),
	.w7(32'hbc078353),
	.w8(32'h3a0654dc),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb53639),
	.w1(32'hbb924c7e),
	.w2(32'h3a3e0238),
	.w3(32'h39819f44),
	.w4(32'hbb91431c),
	.w5(32'h3af31949),
	.w6(32'h3ad2ec8f),
	.w7(32'hba27dbaf),
	.w8(32'h3b809a40),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b47d),
	.w1(32'h3b383d8a),
	.w2(32'hbc1c929f),
	.w3(32'hb9e93278),
	.w4(32'h3a85ac58),
	.w5(32'h3c155879),
	.w6(32'h3a52692b),
	.w7(32'h3bb70212),
	.w8(32'h3c1b5481),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60761a),
	.w1(32'h3c0e3263),
	.w2(32'hbb59f16c),
	.w3(32'h3c51ef9a),
	.w4(32'h3c519402),
	.w5(32'h3b8f5af1),
	.w6(32'h3a0d33e3),
	.w7(32'h3be500f5),
	.w8(32'h3a5a0b28),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f465f),
	.w1(32'hbaf4e787),
	.w2(32'h398eb08d),
	.w3(32'hbc3ebc0b),
	.w4(32'hbc05d6e3),
	.w5(32'h3bac76ec),
	.w6(32'hbbec3a3f),
	.w7(32'hbb8a358f),
	.w8(32'h3c63c382),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b161163),
	.w1(32'h3c110cb7),
	.w2(32'h3c73d446),
	.w3(32'hba55c3ba),
	.w4(32'h3c17ef6b),
	.w5(32'h3c3cf23e),
	.w6(32'h3b986ca6),
	.w7(32'h3c4e1d70),
	.w8(32'h3bf0e64b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8deded),
	.w1(32'h3c7683f0),
	.w2(32'hb9db7bf5),
	.w3(32'h3c5d24a1),
	.w4(32'h3c5076aa),
	.w5(32'h3a4ae6a5),
	.w6(32'h3bcd287d),
	.w7(32'h3bdb7cb1),
	.w8(32'h3beec17b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c64a6),
	.w1(32'hbb6aa89e),
	.w2(32'h3ba8bc4f),
	.w3(32'hbc1a7def),
	.w4(32'hbb9b7cd9),
	.w5(32'h3c5d113d),
	.w6(32'hba3d8e22),
	.w7(32'h3af5a834),
	.w8(32'h3a31db2f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ce254),
	.w1(32'h3bb80764),
	.w2(32'h3be56dae),
	.w3(32'h3b654128),
	.w4(32'h3bd4c4cb),
	.w5(32'h3b87689f),
	.w6(32'hbb8ad1ba),
	.w7(32'hbbc66dfa),
	.w8(32'h3c1285a2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b3443),
	.w1(32'hbc2a2b6c),
	.w2(32'hbc69fd1d),
	.w3(32'h3bf48c3e),
	.w4(32'hbb6f0fe5),
	.w5(32'hbcb858ed),
	.w6(32'h3a3c03c8),
	.w7(32'hbac62181),
	.w8(32'hbc9b6991),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75ab80),
	.w1(32'hbc0d5713),
	.w2(32'h3c394b74),
	.w3(32'hbcdf8748),
	.w4(32'hbc5d6c8b),
	.w5(32'h3c5121de),
	.w6(32'hbc4732de),
	.w7(32'hbbbd09e9),
	.w8(32'h3c1dc538),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb52ec),
	.w1(32'hbb3b4261),
	.w2(32'h3bcb9d88),
	.w3(32'h3c4009a1),
	.w4(32'hbbd7b975),
	.w5(32'h3ba72efd),
	.w6(32'h3c0b8e8a),
	.w7(32'hbb647c7f),
	.w8(32'hb99f4dbc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc593f),
	.w1(32'h3c084af0),
	.w2(32'hbbffd5db),
	.w3(32'h3c20a7a4),
	.w4(32'h3c1324a3),
	.w5(32'hbcfb57b8),
	.w6(32'h3be21356),
	.w7(32'h3c12377e),
	.w8(32'hbc631f1a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7acee5),
	.w1(32'hbc030996),
	.w2(32'h3a8b124d),
	.w3(32'hbd126c4c),
	.w4(32'hbcdd5e12),
	.w5(32'h3bc37887),
	.w6(32'hbd191313),
	.w7(32'hbce60532),
	.w8(32'h3ca85563),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13d0dd),
	.w1(32'h3c52523b),
	.w2(32'hbb18a15e),
	.w3(32'h3b795dbf),
	.w4(32'h3b33001f),
	.w5(32'hbc2a3876),
	.w6(32'h3c3d7f2f),
	.w7(32'h3bc444f9),
	.w8(32'hbc1ad422),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c4f5f),
	.w1(32'hbb30ff4c),
	.w2(32'h3c108ee5),
	.w3(32'hbc9f03f9),
	.w4(32'hbc03f8e9),
	.w5(32'h3bea3d69),
	.w6(32'hbc64ad3a),
	.w7(32'hbb492e07),
	.w8(32'h3c4b34a5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b5ae),
	.w1(32'hba20dc94),
	.w2(32'h3c0ae4f6),
	.w3(32'hbb6874c0),
	.w4(32'hbbb630c6),
	.w5(32'h3c41ec3f),
	.w6(32'hbb94219e),
	.w7(32'h3ba778f2),
	.w8(32'h3b6fa90c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0500f),
	.w1(32'h3ba21fb7),
	.w2(32'h3c81c3d6),
	.w3(32'h3b054838),
	.w4(32'h3a08646a),
	.w5(32'h3ba0bbbf),
	.w6(32'hbaec62e7),
	.w7(32'hbb9f0a40),
	.w8(32'hbad55449),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b0327),
	.w1(32'h3c17091a),
	.w2(32'hbad8f5fd),
	.w3(32'hbb127244),
	.w4(32'h3b0eb94a),
	.w5(32'h3b92c883),
	.w6(32'hbb805777),
	.w7(32'h3b91e1d6),
	.w8(32'h3b2d4bb9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4386dd),
	.w1(32'h3c1e4eeb),
	.w2(32'hbc4d04f7),
	.w3(32'h3b84d713),
	.w4(32'h3c0aa7da),
	.w5(32'hbbf29573),
	.w6(32'h3b344c2b),
	.w7(32'h3ab731b5),
	.w8(32'h39803e2f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fb5e8),
	.w1(32'h3b387da6),
	.w2(32'h3c3e43ba),
	.w3(32'hbbd97b86),
	.w4(32'h3b4240d7),
	.w5(32'h3c77b4a8),
	.w6(32'h3b4a6c56),
	.w7(32'h3c07aec5),
	.w8(32'hba3ccbe9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8b2b0),
	.w1(32'h3c5eb6d5),
	.w2(32'hbb9aebba),
	.w3(32'h3c7ebd9a),
	.w4(32'h3b75de51),
	.w5(32'h39dd2616),
	.w6(32'hbb37dbac),
	.w7(32'hbbd83be8),
	.w8(32'h3b18bad9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f91ea),
	.w1(32'hb964217f),
	.w2(32'h3c72e886),
	.w3(32'hbc0afa26),
	.w4(32'h3afcf1f6),
	.w5(32'h3cb1dcb7),
	.w6(32'hbacbac20),
	.w7(32'h3ba75234),
	.w8(32'h3bc05b70),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c808862),
	.w1(32'h3b05c8d9),
	.w2(32'hbc632cd4),
	.w3(32'h3c9a5429),
	.w4(32'h3c2c6712),
	.w5(32'hbc1e5bd3),
	.w6(32'h3ab57d37),
	.w7(32'hbc2ee015),
	.w8(32'hbb27d2e8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedde6f),
	.w1(32'h3a92f46b),
	.w2(32'hbc3e5d50),
	.w3(32'hbbba218a),
	.w4(32'h39a90e39),
	.w5(32'hbbd9616a),
	.w6(32'h3b71130e),
	.w7(32'h3c1813a8),
	.w8(32'h3b0e0106),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2971ec),
	.w1(32'h39aa4898),
	.w2(32'h3bcb44a0),
	.w3(32'h3af6e055),
	.w4(32'h3c7f9668),
	.w5(32'h3c9a53d2),
	.w6(32'h3c16c712),
	.w7(32'h3c9c01b3),
	.w8(32'h3c5ea115),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c932a41),
	.w1(32'h3b31f266),
	.w2(32'h3c5af86a),
	.w3(32'h3c547a6f),
	.w4(32'h3b945487),
	.w5(32'h3c87f01d),
	.w6(32'h3b995f85),
	.w7(32'h3ba615f6),
	.w8(32'hbb535707),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf24372),
	.w1(32'h393897d6),
	.w2(32'hbca7fd35),
	.w3(32'h3ba9fc65),
	.w4(32'hbc229229),
	.w5(32'hbcca0505),
	.w6(32'hbc04ef94),
	.w7(32'hbc83568e),
	.w8(32'hbc2d7430),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc78bea),
	.w1(32'hbbac80cb),
	.w2(32'h3c122ba6),
	.w3(32'hbcf68d40),
	.w4(32'hbc27759c),
	.w5(32'h3b6de734),
	.w6(32'hbbfaf259),
	.w7(32'h3c47d833),
	.w8(32'h3bd3390f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa65f),
	.w1(32'h3b9bd87f),
	.w2(32'h3a7a4d1b),
	.w3(32'hba2afeeb),
	.w4(32'h3ba69a2c),
	.w5(32'h3b578f9c),
	.w6(32'hbbab7282),
	.w7(32'hbb586be7),
	.w8(32'h3a89da6e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe6917),
	.w1(32'hbbbe2af7),
	.w2(32'h3bf20820),
	.w3(32'h3b18837f),
	.w4(32'hbbb8af41),
	.w5(32'h3c1c0898),
	.w6(32'h3ae7a406),
	.w7(32'h3ad77364),
	.w8(32'h38d4880b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c971749),
	.w1(32'hbac3a7d9),
	.w2(32'hbb0c63f3),
	.w3(32'h3c28c490),
	.w4(32'h3b6ff210),
	.w5(32'hbac1f46d),
	.w6(32'hbc10f5ed),
	.w7(32'hbb9a68fb),
	.w8(32'h3ae31e7a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef435d),
	.w1(32'h3bc8d0de),
	.w2(32'hbb06b5c2),
	.w3(32'hbc22590e),
	.w4(32'h3b8ef688),
	.w5(32'hbb2943c6),
	.w6(32'h3abb09fe),
	.w7(32'h3c073986),
	.w8(32'h3bcac632),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01f48b),
	.w1(32'hbac4355e),
	.w2(32'h3d590639),
	.w3(32'hbc6af826),
	.w4(32'hbb94ace4),
	.w5(32'h3d5cec12),
	.w6(32'hbb51a488),
	.w7(32'h3aa7a69d),
	.w8(32'h3ad99aae),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d74d415),
	.w1(32'h3c438ab9),
	.w2(32'h3c163587),
	.w3(32'h3d2e377b),
	.w4(32'hbba2bb32),
	.w5(32'h3c239c21),
	.w6(32'hbc903643),
	.w7(32'hbd48c13d),
	.w8(32'hbbbbbc23),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a4beb),
	.w1(32'h3c1a5eda),
	.w2(32'h3bfcd626),
	.w3(32'h3c6b70f0),
	.w4(32'h3b935e3a),
	.w5(32'hbb453e6a),
	.w6(32'h3b0ad730),
	.w7(32'h3afc71bf),
	.w8(32'hbc32d4ba),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3928e7),
	.w1(32'hbb95a098),
	.w2(32'h3b1239a1),
	.w3(32'h3bac9e9f),
	.w4(32'h3bca592b),
	.w5(32'hbb056163),
	.w6(32'hbbbeaaa4),
	.w7(32'h3b6624ca),
	.w8(32'h3bac2400),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae02e7d),
	.w1(32'hbb1f6305),
	.w2(32'h3792813f),
	.w3(32'hbad3b5c0),
	.w4(32'hbb86b20a),
	.w5(32'hbb2b6920),
	.w6(32'hbbb19a68),
	.w7(32'hbb196b31),
	.w8(32'h3aa88966),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb781cb4),
	.w1(32'h3b0c987c),
	.w2(32'h3b17cf31),
	.w3(32'hbc2a4ab7),
	.w4(32'h3a917641),
	.w5(32'h3b8a1c13),
	.w6(32'hbb49ba24),
	.w7(32'h3bbf5366),
	.w8(32'h3c742d3b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f806c),
	.w1(32'hb83c4ae1),
	.w2(32'hbb10fa55),
	.w3(32'h3b7a3c09),
	.w4(32'hba1e0e7d),
	.w5(32'h3991c74e),
	.w6(32'h3a01d84f),
	.w7(32'h3a8819fc),
	.w8(32'h3a5afa86),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf3116),
	.w1(32'h3baef59d),
	.w2(32'h39807a58),
	.w3(32'hba6a32f6),
	.w4(32'h3c088513),
	.w5(32'hbc7db777),
	.w6(32'hba362988),
	.w7(32'h3bae7d93),
	.w8(32'hbc1867ad),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f4235),
	.w1(32'hba3158ce),
	.w2(32'hbbe0cfa5),
	.w3(32'hbca51fde),
	.w4(32'hb9c171f5),
	.w5(32'hbb9a481e),
	.w6(32'hbbf72be4),
	.w7(32'hbb972898),
	.w8(32'h3b12c5f2),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b3b8),
	.w1(32'hbbb7d1ee),
	.w2(32'h3b6f8b09),
	.w3(32'hbc18be45),
	.w4(32'hb9e84212),
	.w5(32'h3c62526e),
	.w6(32'hbbbc3783),
	.w7(32'hbc1fd185),
	.w8(32'h3b279eff),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a36fb),
	.w1(32'h3bf2d834),
	.w2(32'hbc21adba),
	.w3(32'h3c1e8d8a),
	.w4(32'h3b58e0e6),
	.w5(32'hbca48db8),
	.w6(32'hba8f39a4),
	.w7(32'hbbf25a9f),
	.w8(32'hbc732b6e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb03a8d),
	.w1(32'hbc10543e),
	.w2(32'hbafeb8a4),
	.w3(32'hbcf2c7d7),
	.w4(32'hbc40b19a),
	.w5(32'hbb2691bb),
	.w6(32'hbcd75494),
	.w7(32'hbbed9245),
	.w8(32'hbb633517),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5faf7a),
	.w1(32'hbb25cb0e),
	.w2(32'h3b075996),
	.w3(32'hbb822b96),
	.w4(32'hbbb1a4b0),
	.w5(32'hbb8b50cb),
	.w6(32'hba048d45),
	.w7(32'hba430440),
	.w8(32'hbbae3917),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1db5c0),
	.w1(32'hb9906630),
	.w2(32'h3bbb3813),
	.w3(32'hbbc3f21d),
	.w4(32'hbb849b89),
	.w5(32'h3c0ae44d),
	.w6(32'hbc10e8a5),
	.w7(32'hbc1029d1),
	.w8(32'h3c18b533),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d78e),
	.w1(32'hbb4c9fc2),
	.w2(32'hbb84b043),
	.w3(32'h3ba2d2b3),
	.w4(32'hbbf9c16b),
	.w5(32'h3b5e065b),
	.w6(32'h3b9c2c5e),
	.w7(32'hbb386355),
	.w8(32'h3c3a5bef),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48c5bf),
	.w1(32'h3b1b1bc8),
	.w2(32'h3c455f98),
	.w3(32'h3bddc3ff),
	.w4(32'h3c25601f),
	.w5(32'h3c00ebe4),
	.w6(32'h3cba6086),
	.w7(32'h3c59b309),
	.w8(32'h3c018f6a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bf445),
	.w1(32'h3c3dba85),
	.w2(32'hbcf90cc5),
	.w3(32'h3bd6ce6d),
	.w4(32'h3b110883),
	.w5(32'hbcd7927a),
	.w6(32'h3c0c182f),
	.w7(32'hba28fdb3),
	.w8(32'h3b384f66),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccabde3),
	.w1(32'hb92d0841),
	.w2(32'h3bb52b50),
	.w3(32'hbb9c5b78),
	.w4(32'h3c59c836),
	.w5(32'hb99e75da),
	.w6(32'h3cbdbe00),
	.w7(32'h3ceaacda),
	.w8(32'h3b72a1d5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34bb4),
	.w1(32'hba0a3ad7),
	.w2(32'hbb80d8bf),
	.w3(32'hbbea6fbd),
	.w4(32'hbbd2f913),
	.w5(32'hbb92eaf9),
	.w6(32'hbc0ae980),
	.w7(32'hbc4c7fba),
	.w8(32'hba17ff24),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb782c70),
	.w1(32'h3c01f29e),
	.w2(32'h3af879f8),
	.w3(32'hbc07f524),
	.w4(32'h3bf5b17a),
	.w5(32'h3bc5dc20),
	.w6(32'hbae9b90e),
	.w7(32'h3c1856de),
	.w8(32'h3c03f6f3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75d0b1),
	.w1(32'hbc0bf541),
	.w2(32'hbc4753ae),
	.w3(32'h3b827436),
	.w4(32'hbc3cc760),
	.w5(32'h394c0a31),
	.w6(32'hbc5cb715),
	.w7(32'hbc606cb3),
	.w8(32'h3b07eb0b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0f99d),
	.w1(32'h3bb40f76),
	.w2(32'h3c65fee7),
	.w3(32'hbab90833),
	.w4(32'hbad83ece),
	.w5(32'hbb0f5624),
	.w6(32'h3bbae32c),
	.w7(32'h3bafd1fb),
	.w8(32'hbca19135),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191aee),
	.w1(32'hbca34ffa),
	.w2(32'h3c86408c),
	.w3(32'hbc3f3228),
	.w4(32'hbd04d180),
	.w5(32'h3c4cb2d7),
	.w6(32'hbd1cb070),
	.w7(32'hbd30b27a),
	.w8(32'h3c00c733),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc462e),
	.w1(32'h3bc87002),
	.w2(32'h3afc940a),
	.w3(32'h3c5e5639),
	.w4(32'h3bd3609b),
	.w5(32'h3b9bed9a),
	.w6(32'h3b90edc5),
	.w7(32'hbb3cf12b),
	.w8(32'h3c8ee6b5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5e488),
	.w1(32'h3b05ab01),
	.w2(32'h3b8d4d68),
	.w3(32'h3c4a92f5),
	.w4(32'h3c363479),
	.w5(32'h3bd2bfd3),
	.w6(32'h3c56afe1),
	.w7(32'h3cab7b29),
	.w8(32'h3c3c1590),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471939),
	.w1(32'hbc38546d),
	.w2(32'h3c38afd3),
	.w3(32'h3b1a1fdc),
	.w4(32'hbc2d7dd6),
	.w5(32'h3c8fccad),
	.w6(32'h3c3d0b2c),
	.w7(32'hbc8928ce),
	.w8(32'hbad8fba3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c913282),
	.w1(32'hbafcbf62),
	.w2(32'h3caa0b46),
	.w3(32'h3bb8b02b),
	.w4(32'hbc7111ba),
	.w5(32'h3bf6d678),
	.w6(32'h3b00e401),
	.w7(32'hbc08e02d),
	.w8(32'h3b9c823d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb60cb9),
	.w1(32'h3b949084),
	.w2(32'h3a9581d2),
	.w3(32'h3c6cf327),
	.w4(32'h3b449c78),
	.w5(32'h3b5e59aa),
	.w6(32'h3c03cae8),
	.w7(32'hbb9d9fad),
	.w8(32'h3c04e277),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7d98),
	.w1(32'h3aad37df),
	.w2(32'h3c3bd01c),
	.w3(32'hbbf5847c),
	.w4(32'hbb945825),
	.w5(32'h3bd23227),
	.w6(32'hba935eac),
	.w7(32'hbad308cc),
	.w8(32'h3be74364),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aad72),
	.w1(32'hbb1a1a93),
	.w2(32'hbba33cad),
	.w3(32'hbbafa1e8),
	.w4(32'hba77d584),
	.w5(32'hbb4826eb),
	.w6(32'hbb9d89b0),
	.w7(32'h3b27c269),
	.w8(32'h3948e157),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb407194),
	.w1(32'h3ba65340),
	.w2(32'h3c4351b0),
	.w3(32'h3bc6b76e),
	.w4(32'h3c6742e9),
	.w5(32'h3bc2cbfc),
	.w6(32'h3c16f985),
	.w7(32'h3c216487),
	.w8(32'h3b3aad44),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b053ea7),
	.w1(32'h3a7f72a4),
	.w2(32'h3c489bed),
	.w3(32'h3b55267f),
	.w4(32'h3b713edf),
	.w5(32'h3bfdc3d1),
	.w6(32'hbaa97138),
	.w7(32'h3a86e6f1),
	.w8(32'h3b1c55bd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb84417),
	.w1(32'h3b69b68f),
	.w2(32'hba744909),
	.w3(32'h38d7010c),
	.w4(32'h3b51e102),
	.w5(32'h3ab4f896),
	.w6(32'hbafb2016),
	.w7(32'h3c0563b1),
	.w8(32'h3c072735),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c5524),
	.w1(32'hbc5b68a4),
	.w2(32'h3b84bcaf),
	.w3(32'h39fb6df5),
	.w4(32'hbb0625e7),
	.w5(32'h3b7fa0dd),
	.w6(32'h3bedccaf),
	.w7(32'h3c1aa02f),
	.w8(32'hbb40ccfb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd7a72),
	.w1(32'h3bbb4131),
	.w2(32'h3b9fd8cc),
	.w3(32'h3c237405),
	.w4(32'hba960461),
	.w5(32'h3be7531f),
	.w6(32'hbbbb148f),
	.w7(32'hbad48872),
	.w8(32'h3c0e1e1d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7973e),
	.w1(32'h3adcccf7),
	.w2(32'h3c660aa1),
	.w3(32'hbafeb4c7),
	.w4(32'h3b97ca1a),
	.w5(32'h3c7b8eca),
	.w6(32'h3c0cc1fa),
	.w7(32'h3c636b43),
	.w8(32'h3be28e17),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65d4bd),
	.w1(32'h3bd8ca67),
	.w2(32'hbbd2c55b),
	.w3(32'h3bd0d657),
	.w4(32'hbb7a8224),
	.w5(32'hbc943a77),
	.w6(32'hbaeda6b6),
	.w7(32'hba0f7d3d),
	.w8(32'hba2513ee),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4521c7),
	.w1(32'h3be8bd5e),
	.w2(32'h3c6e57e9),
	.w3(32'hbc28a4fa),
	.w4(32'h3c48bd53),
	.w5(32'h3c9af704),
	.w6(32'h3c95ec98),
	.w7(32'h3cae1f53),
	.w8(32'h3c71c236),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb940e8),
	.w1(32'h3b75b907),
	.w2(32'h3a7b4f31),
	.w3(32'h3bc1d6c5),
	.w4(32'hbba6ceaa),
	.w5(32'h3bfe147b),
	.w6(32'h3b26035d),
	.w7(32'hbc0030d2),
	.w8(32'h3c0ee65f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2566da),
	.w1(32'h3b9e4f30),
	.w2(32'h3c7a89ea),
	.w3(32'h3c143865),
	.w4(32'h3c00e381),
	.w5(32'h3d0ad374),
	.w6(32'h3cdfa0e1),
	.w7(32'h3c8efebb),
	.w8(32'h3cad6ea8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdddb83),
	.w1(32'h3cbd9ffa),
	.w2(32'hbc00699b),
	.w3(32'h3d228422),
	.w4(32'h3c9d8a2e),
	.w5(32'hbc12656c),
	.w6(32'h3c986991),
	.w7(32'h3b606852),
	.w8(32'h3af9d81f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e97e1),
	.w1(32'hbc42e152),
	.w2(32'hbc8ef1aa),
	.w3(32'hbc474794),
	.w4(32'hbc179de4),
	.w5(32'h3b79fc5b),
	.w6(32'hba4a7aea),
	.w7(32'hb94b9d50),
	.w8(32'h3b8d318d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc38d42),
	.w1(32'hbc760e98),
	.w2(32'h3a232938),
	.w3(32'hbb678615),
	.w4(32'hbbacb4eb),
	.w5(32'h3b8e77fe),
	.w6(32'hbb790c2a),
	.w7(32'hbbbc6c74),
	.w8(32'hba88fdbc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3157cf),
	.w1(32'hbb325fb8),
	.w2(32'hbb9441de),
	.w3(32'hbb227b1f),
	.w4(32'hbb999767),
	.w5(32'hbbd3a48d),
	.w6(32'hbb4225bb),
	.w7(32'hbaab3512),
	.w8(32'hbba7b800),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ad0d),
	.w1(32'h395e78d3),
	.w2(32'h3c7c3780),
	.w3(32'hbbf6c1ff),
	.w4(32'hbb136d67),
	.w5(32'h3cb02fdf),
	.w6(32'h3b75c31b),
	.w7(32'h3c4ce107),
	.w8(32'h3bc99d0f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caab87c),
	.w1(32'h3bcb5621),
	.w2(32'h3c65232c),
	.w3(32'h3c99e45b),
	.w4(32'hb9968b1a),
	.w5(32'h3cb8bd06),
	.w6(32'h3b954109),
	.w7(32'hbbdc5748),
	.w8(32'h3abf82c5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e27a2),
	.w1(32'h3b495775),
	.w2(32'hba6f89a4),
	.w3(32'h3cc0e730),
	.w4(32'h391b7608),
	.w5(32'hbb848a93),
	.w6(32'hbc07361f),
	.w7(32'hbc8e3101),
	.w8(32'hbb21a93e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04db29),
	.w1(32'h3b4dd7a0),
	.w2(32'h3c841590),
	.w3(32'hbb1f0ea0),
	.w4(32'hba8386c1),
	.w5(32'h3c8074ae),
	.w6(32'hbb3bb56a),
	.w7(32'hbb2bf495),
	.w8(32'h3bfea696),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f3393),
	.w1(32'h3c2cef82),
	.w2(32'h3cb56ba7),
	.w3(32'h3c4b107d),
	.w4(32'h3b46e989),
	.w5(32'h3d027500),
	.w6(32'h3b8ba3b0),
	.w7(32'hb9f47141),
	.w8(32'h3cd67c35),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1356a),
	.w1(32'h3c6e5433),
	.w2(32'hbc116746),
	.w3(32'h3cc6aa4d),
	.w4(32'h3c486fbc),
	.w5(32'hbc243360),
	.w6(32'h3c1fc3a4),
	.w7(32'hb95d0ad0),
	.w8(32'hbbd0faba),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe22839),
	.w1(32'hbb928791),
	.w2(32'hbb29d8ba),
	.w3(32'hbc10b76d),
	.w4(32'hbb1c4d55),
	.w5(32'hbaedaedc),
	.w6(32'hbb7abe36),
	.w7(32'h3b7f353e),
	.w8(32'hbb562dcd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba80d17),
	.w1(32'h3afd2dd8),
	.w2(32'h3b51e369),
	.w3(32'h3bb046dd),
	.w4(32'h3c5cac62),
	.w5(32'h3be53e96),
	.w6(32'h3c060a1a),
	.w7(32'h3c9d7440),
	.w8(32'h3c034440),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0668e),
	.w1(32'h3ba7c2c2),
	.w2(32'h3c33cd73),
	.w3(32'h3bd84b7e),
	.w4(32'h3c413855),
	.w5(32'h3cdcf26c),
	.w6(32'h3c19efe2),
	.w7(32'h3c237660),
	.w8(32'h3c214c46),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ecf78),
	.w1(32'hbb945f61),
	.w2(32'hba3218fc),
	.w3(32'h3c8a4f18),
	.w4(32'h3b80b9ee),
	.w5(32'h3ab27a48),
	.w6(32'h3c24d5b3),
	.w7(32'hbbc8ba23),
	.w8(32'h3bd7d9c7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b6bd),
	.w1(32'h3b074845),
	.w2(32'h3b53af53),
	.w3(32'hbbbb071d),
	.w4(32'h3a9e1252),
	.w5(32'h3c112929),
	.w6(32'h3c1d9d1d),
	.w7(32'h3b968a30),
	.w8(32'h3c00c59c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd7409),
	.w1(32'h3ab85c0f),
	.w2(32'hbd0f7c4f),
	.w3(32'hbb47070e),
	.w4(32'hbc1d824f),
	.w5(32'hbd3b1a4c),
	.w6(32'h3b116b8c),
	.w7(32'h3b5d7bb8),
	.w8(32'hbcab6117),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd65761),
	.w1(32'hbbb9389a),
	.w2(32'h3c7ae806),
	.w3(32'hbd17311b),
	.w4(32'hbb7fe981),
	.w5(32'h3c569d52),
	.w6(32'hbbf64324),
	.w7(32'hbbd1f46c),
	.w8(32'h3ba911e7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82eabc),
	.w1(32'hba75b198),
	.w2(32'hbc61274a),
	.w3(32'h3c543959),
	.w4(32'h3bae549b),
	.w5(32'hbcefe7fc),
	.w6(32'h3b41a6f2),
	.w7(32'hbbc6018f),
	.w8(32'hbc4e243a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc255622),
	.w1(32'hbc9daf78),
	.w2(32'hbc0834f2),
	.w3(32'hbcf844da),
	.w4(32'hbc9250ac),
	.w5(32'hbc932c60),
	.w6(32'hbc8622b1),
	.w7(32'hbc49664c),
	.w8(32'hbc928d62),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bed03),
	.w1(32'hbb9ce78e),
	.w2(32'h3b8c5637),
	.w3(32'hbc7d1731),
	.w4(32'hbbf8e7cd),
	.w5(32'h3a5a26ae),
	.w6(32'hbc6f5063),
	.w7(32'hbb13801d),
	.w8(32'h3b6f5089),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1905ad),
	.w1(32'h3bcb0001),
	.w2(32'hbc1ac3ad),
	.w3(32'hbbd63d50),
	.w4(32'h3b2d31d9),
	.w5(32'hbb87fbb1),
	.w6(32'hbbc32af1),
	.w7(32'h3abb36f8),
	.w8(32'h3c0a9820),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963ddf),
	.w1(32'h3b43394c),
	.w2(32'h3b96c1d6),
	.w3(32'hbbbbf68c),
	.w4(32'h3928fea0),
	.w5(32'hb97c78fb),
	.w6(32'h3b4d2d3b),
	.w7(32'h3bc8e6d0),
	.w8(32'h3b7e39b3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c2305),
	.w1(32'h3b601341),
	.w2(32'h3beb2f79),
	.w3(32'h3b5780d4),
	.w4(32'h3ab58940),
	.w5(32'h3ba95d30),
	.w6(32'h3b156f43),
	.w7(32'h3c10decf),
	.w8(32'hbb33346e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2be5e),
	.w1(32'hbb7e2034),
	.w2(32'h3ba0321c),
	.w3(32'h3c01d0a0),
	.w4(32'hbc0695d9),
	.w5(32'h3b64f213),
	.w6(32'hbb521ee8),
	.w7(32'hbc406a67),
	.w8(32'h3b49f1ea),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb52872),
	.w1(32'h3b9bb3b8),
	.w2(32'h3a9f5139),
	.w3(32'h3b68ce50),
	.w4(32'h3b68cf5a),
	.w5(32'h3c904a68),
	.w6(32'h3b801b0d),
	.w7(32'hb9f41b69),
	.w8(32'h3a2aa1ea),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c317765),
	.w1(32'h3c1da016),
	.w2(32'h3bad0fe0),
	.w3(32'h3c96fde2),
	.w4(32'h3c172221),
	.w5(32'h3bab59e5),
	.w6(32'hbb1a91da),
	.w7(32'hbb88cd15),
	.w8(32'h3c0639a4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e639b2),
	.w1(32'h3afbfe3b),
	.w2(32'h3b961506),
	.w3(32'hbb527c02),
	.w4(32'hbad57d0d),
	.w5(32'h3b51c116),
	.w6(32'hbb4902de),
	.w7(32'hbae6ca01),
	.w8(32'h3c319135),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c312849),
	.w1(32'h3c1964df),
	.w2(32'hbbb51e90),
	.w3(32'h3c35b3b3),
	.w4(32'h3c092a95),
	.w5(32'hbcbb1e83),
	.w6(32'h3cba3218),
	.w7(32'h3c7aa50f),
	.w8(32'hbc02d0a7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca58ddb),
	.w1(32'hbcad6122),
	.w2(32'h39c0c984),
	.w3(32'hbcdd6d45),
	.w4(32'hbcd25f5d),
	.w5(32'h3ab08a45),
	.w6(32'hbc9da58f),
	.w7(32'hbca70a76),
	.w8(32'h3bbfb580),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079ab6),
	.w1(32'hba647108),
	.w2(32'hbb461463),
	.w3(32'hba851235),
	.w4(32'hbacb1418),
	.w5(32'hbb94b80e),
	.w6(32'hba9b489b),
	.w7(32'h3ac56b8a),
	.w8(32'hbaffece4),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8da7d),
	.w1(32'h3b7d0d48),
	.w2(32'hbbd30126),
	.w3(32'hbb373f31),
	.w4(32'h3bc45e6e),
	.w5(32'hbc1eda56),
	.w6(32'h3a447282),
	.w7(32'h3b9919b4),
	.w8(32'h3c27a71a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe25efd),
	.w1(32'h3ba13cf9),
	.w2(32'h3b5a445f),
	.w3(32'hbc1ee139),
	.w4(32'h3bc80b44),
	.w5(32'h3ad3db65),
	.w6(32'h3c480b09),
	.w7(32'h3cd8743e),
	.w8(32'h3bc0e4cb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9de59),
	.w1(32'h3c39b641),
	.w2(32'hbbe32de1),
	.w3(32'h3c3170fd),
	.w4(32'h3c0c47ae),
	.w5(32'hbc901a07),
	.w6(32'h3c402785),
	.w7(32'h3c46aa52),
	.w8(32'hba54a255),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe97915),
	.w1(32'h39ca5bb7),
	.w2(32'h3bd7ed9d),
	.w3(32'hbc43c33b),
	.w4(32'h3a815050),
	.w5(32'h3bfd10a0),
	.w6(32'hbb33b32d),
	.w7(32'h3a544834),
	.w8(32'h3bc26156),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b09da),
	.w1(32'h3b374b1e),
	.w2(32'h3c76fb0a),
	.w3(32'hbae8d5fa),
	.w4(32'h3a48a96c),
	.w5(32'h3c87b91c),
	.w6(32'h3a758145),
	.w7(32'h3af7a1cc),
	.w8(32'h3becf83e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf1642),
	.w1(32'h3c2754fd),
	.w2(32'h3b1d1c1a),
	.w3(32'h3c4f0714),
	.w4(32'h3c2a8ca9),
	.w5(32'h3b7c1640),
	.w6(32'hbb9bb3c0),
	.w7(32'hba994672),
	.w8(32'h3b45bcf5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaf101),
	.w1(32'h3b991556),
	.w2(32'h3c387602),
	.w3(32'hbb267565),
	.w4(32'h3b90495c),
	.w5(32'h3bfd3be0),
	.w6(32'h3b7f39a9),
	.w7(32'h3bf0f1b1),
	.w8(32'h3b654b66),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61fbd6),
	.w1(32'h3bf402ea),
	.w2(32'h3b4781f7),
	.w3(32'h3bb2780f),
	.w4(32'hba8477c1),
	.w5(32'h3b07b352),
	.w6(32'hbb85036b),
	.w7(32'hbbf6a02b),
	.w8(32'h3c2516a3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fa119),
	.w1(32'h3c1a1511),
	.w2(32'h3c099398),
	.w3(32'h3c1e8f76),
	.w4(32'h3b09343c),
	.w5(32'hbb028bbe),
	.w6(32'h3c0c4655),
	.w7(32'h3c8346ca),
	.w8(32'h3b05652d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f12c),
	.w1(32'hbbfaf880),
	.w2(32'h3c03e8c0),
	.w3(32'hbba05e3b),
	.w4(32'hbc2f3b85),
	.w5(32'h3c0935ac),
	.w6(32'h3ac5b66d),
	.w7(32'hb7921220),
	.w8(32'hbbc4c0c2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00f1ce),
	.w1(32'h3b5f898c),
	.w2(32'h39c5ff0c),
	.w3(32'h3af14ef1),
	.w4(32'hbbc94af0),
	.w5(32'hbb6c16f6),
	.w6(32'hba8e35cf),
	.w7(32'hbc0b0238),
	.w8(32'h38d4f92b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b1300),
	.w1(32'h3af5aa66),
	.w2(32'hbb04f1d2),
	.w3(32'hbab96691),
	.w4(32'hbb98a168),
	.w5(32'hbb9f6443),
	.w6(32'h3b740201),
	.w7(32'h38740590),
	.w8(32'hbb6f5196),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaada087),
	.w1(32'h3acf1472),
	.w2(32'h3bfee221),
	.w3(32'hbb462838),
	.w4(32'hbbb0241b),
	.w5(32'hbb45980f),
	.w6(32'h3b1b1223),
	.w7(32'hba1d104d),
	.w8(32'h3cc26818),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d674),
	.w1(32'h3b0e8db0),
	.w2(32'h3b1c3f31),
	.w3(32'hbc826506),
	.w4(32'hbbcb657d),
	.w5(32'hbac2c68a),
	.w6(32'h3cdd2c95),
	.w7(32'h3d0da5f9),
	.w8(32'hbb3e5bd1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cca79),
	.w1(32'h3b3e7e95),
	.w2(32'hbc335b75),
	.w3(32'h3a18a25a),
	.w4(32'h3ac4a8d5),
	.w5(32'hbb871c1a),
	.w6(32'hbb342ae8),
	.w7(32'hba519d24),
	.w8(32'hbb7d228b),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9dac03),
	.w1(32'hbc7ff0c9),
	.w2(32'hbc357795),
	.w3(32'hbb888374),
	.w4(32'h3a5b8e2e),
	.w5(32'hbc1b5571),
	.w6(32'h3b2167f6),
	.w7(32'h3aff8694),
	.w8(32'hbb8e5422),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7da8),
	.w1(32'hbc67bb81),
	.w2(32'h3ac790ba),
	.w3(32'hbc3013d0),
	.w4(32'hbbfd372d),
	.w5(32'h3afcaf4b),
	.w6(32'hbbfb8ff5),
	.w7(32'hbbb376de),
	.w8(32'hbac543c2),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405f8d),
	.w1(32'hbaef638c),
	.w2(32'hbc0ab854),
	.w3(32'hbad7f23e),
	.w4(32'hbaa0aaf6),
	.w5(32'hbc1c7e45),
	.w6(32'hbbcc3ad3),
	.w7(32'hbb9fd885),
	.w8(32'hbc551ec1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11553a),
	.w1(32'h3a8d2489),
	.w2(32'hbb087f93),
	.w3(32'hbb926b13),
	.w4(32'hbba0d22c),
	.w5(32'h3a8f9900),
	.w6(32'hbc7fff7d),
	.w7(32'hbc623134),
	.w8(32'h3b3baa2f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3e22),
	.w1(32'hbb189455),
	.w2(32'hb9fed788),
	.w3(32'hba54ed94),
	.w4(32'h3a2e9532),
	.w5(32'hbce7f233),
	.w6(32'h3a2d85dc),
	.w7(32'hba45907f),
	.w8(32'h3ccbbf68),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17043c),
	.w1(32'hbc9f54a5),
	.w2(32'hba775d3d),
	.w3(32'hbce6a834),
	.w4(32'h3b298d9b),
	.w5(32'h3ab7be3c),
	.w6(32'h3c911515),
	.w7(32'h3d00d53d),
	.w8(32'hbbb8f0b1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961dfc5),
	.w1(32'hbaaee9e9),
	.w2(32'h3bc03c0e),
	.w3(32'hba7b488c),
	.w4(32'hbb982adc),
	.w5(32'h3aef101c),
	.w6(32'hbc02bfaf),
	.w7(32'hbc2a2107),
	.w8(32'hbad516e2),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34aa95),
	.w1(32'h3c355207),
	.w2(32'h3ab53366),
	.w3(32'h3a72e00c),
	.w4(32'hbb486411),
	.w5(32'hbacf20f8),
	.w6(32'hbbefce86),
	.w7(32'hbc1c3eed),
	.w8(32'h3b3cfc90),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c30dc),
	.w1(32'hbc0d3bdb),
	.w2(32'h3b373619),
	.w3(32'h3bc7fc7d),
	.w4(32'hbab6b42c),
	.w5(32'h3b96144d),
	.w6(32'hbb830c2f),
	.w7(32'hbb8b99bb),
	.w8(32'h3b74ec2d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc6ff5),
	.w1(32'h3b4777bb),
	.w2(32'h3be0046e),
	.w3(32'h3b2072c9),
	.w4(32'h3c1585af),
	.w5(32'hb7c23538),
	.w6(32'h3c2beafa),
	.w7(32'h3c126e53),
	.w8(32'h3bed3869),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8789c),
	.w1(32'h3bfff0c5),
	.w2(32'hbc3805c7),
	.w3(32'hbc28c9f4),
	.w4(32'hba860bbf),
	.w5(32'hbc1cfd61),
	.w6(32'hbb900bc3),
	.w7(32'h38e13ee4),
	.w8(32'hbc6814f5),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473c40),
	.w1(32'hbc16ab45),
	.w2(32'hbb1f44fe),
	.w3(32'hbc4bd211),
	.w4(32'hbc04804a),
	.w5(32'h3adbf02d),
	.w6(32'hbc6c3988),
	.w7(32'hbb9b0154),
	.w8(32'h3b064ffa),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea9498),
	.w1(32'hbb628391),
	.w2(32'hbba655c9),
	.w3(32'h3a813778),
	.w4(32'hba91b3af),
	.w5(32'h3c41dcf5),
	.w6(32'hb80a68de),
	.w7(32'h3985e25d),
	.w8(32'hbac123cd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76991),
	.w1(32'hbab990cc),
	.w2(32'h3c638e0a),
	.w3(32'h399f4666),
	.w4(32'hbc41bb01),
	.w5(32'h3c4049aa),
	.w6(32'h3b893e9a),
	.w7(32'h3b665b7d),
	.w8(32'h3b9908ca),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c776149),
	.w1(32'h3c545d6a),
	.w2(32'h3c01fb5b),
	.w3(32'hbb960092),
	.w4(32'hbbc8ee41),
	.w5(32'hbaef3ff4),
	.w6(32'h3c64892c),
	.w7(32'h3c925cdb),
	.w8(32'hbb191959),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80b14e),
	.w1(32'h3c5b76f3),
	.w2(32'h3b87931a),
	.w3(32'hbc107f74),
	.w4(32'hbbd947d6),
	.w5(32'hbc48b3cb),
	.w6(32'hbc6130f9),
	.w7(32'hbb955f44),
	.w8(32'h3c127e05),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c388444),
	.w1(32'h3c45a61b),
	.w2(32'hbb30172d),
	.w3(32'hbc9abef1),
	.w4(32'hbbd072a6),
	.w5(32'hb987e4d3),
	.w6(32'hbb5f4eb7),
	.w7(32'hbae5db8b),
	.w8(32'h3a8dc138),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6178b),
	.w1(32'hb9f4b371),
	.w2(32'h3b093827),
	.w3(32'h3a4d6082),
	.w4(32'hbab52232),
	.w5(32'h3c830319),
	.w6(32'h3b24e996),
	.w7(32'h3ab030cf),
	.w8(32'h3b62acc2),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b505d78),
	.w1(32'h3c8eba83),
	.w2(32'hbb111850),
	.w3(32'h3d03b38a),
	.w4(32'h3cab2e70),
	.w5(32'hbc7a4db8),
	.w6(32'h3ab8d2bd),
	.w7(32'h3ac49fab),
	.w8(32'hbba79cf0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badabe1),
	.w1(32'h3c1b4f70),
	.w2(32'h3bdf7cfe),
	.w3(32'hbc2184a3),
	.w4(32'hbc801152),
	.w5(32'hbca4dd08),
	.w6(32'hbc30f96c),
	.w7(32'h3b652d48),
	.w8(32'hbbdee8e3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba602a10),
	.w1(32'hbb945187),
	.w2(32'h3bdf2031),
	.w3(32'hbc6acc08),
	.w4(32'hbc9f92e8),
	.w5(32'hbc861470),
	.w6(32'h3b616ced),
	.w7(32'hbb146465),
	.w8(32'h3b030392),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c843312),
	.w1(32'h3c141f21),
	.w2(32'hbbb913c0),
	.w3(32'hbc65d985),
	.w4(32'hbc6cf1b1),
	.w5(32'h3b8543dc),
	.w6(32'h3b8dda41),
	.w7(32'h3c19a5e0),
	.w8(32'h3b7f05d5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc402ad1),
	.w1(32'hbb8d876d),
	.w2(32'hbb2053ea),
	.w3(32'h3bd8493b),
	.w4(32'h3be0f7af),
	.w5(32'h3c0d1f0f),
	.w6(32'hb8fef356),
	.w7(32'hba0c4852),
	.w8(32'h3c980cad),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374263),
	.w1(32'hbbe1a33f),
	.w2(32'h3b324bc7),
	.w3(32'h3c85c737),
	.w4(32'h3cf9e662),
	.w5(32'hbc1f52e5),
	.w6(32'h3cc6121e),
	.w7(32'h3cb6c78b),
	.w8(32'h3ad0b24d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3614cb),
	.w1(32'h3a1c4d85),
	.w2(32'h3b8ff392),
	.w3(32'hbc1ebd0d),
	.w4(32'hbc108197),
	.w5(32'hbbb287af),
	.w6(32'h3bff9ad4),
	.w7(32'h3c16aa94),
	.w8(32'h3adf22c7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d21ce),
	.w1(32'h3c2f9a38),
	.w2(32'hb99d077f),
	.w3(32'hbb8d47e3),
	.w4(32'hbc2e18e1),
	.w5(32'h3b577ca8),
	.w6(32'hbb1050bc),
	.w7(32'h3b922fdb),
	.w8(32'hbaa7789b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ee38),
	.w1(32'h3adb0bc4),
	.w2(32'hba4847d1),
	.w3(32'h3b5f9211),
	.w4(32'h3bc3c4d8),
	.w5(32'hba3ce6a4),
	.w6(32'hbba50036),
	.w7(32'hbb144981),
	.w8(32'hbaac2d44),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c07b),
	.w1(32'h3bc6645e),
	.w2(32'hbc030c34),
	.w3(32'hbab31b1a),
	.w4(32'h3c148acc),
	.w5(32'h38ae3edf),
	.w6(32'hbbb9a35a),
	.w7(32'h3bb6edf2),
	.w8(32'h3a72928b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ca6b1),
	.w1(32'h3c1aed95),
	.w2(32'h3b2f3928),
	.w3(32'h3c7fb0ea),
	.w4(32'h3c8df719),
	.w5(32'h3c10dafa),
	.w6(32'hbb207648),
	.w7(32'hba3075a7),
	.w8(32'h3802b016),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45f155),
	.w1(32'h3b3e10a2),
	.w2(32'h3bfa65f0),
	.w3(32'h3c0e56c5),
	.w4(32'h3b8b511a),
	.w5(32'hba88aa83),
	.w6(32'h3b7c0df1),
	.w7(32'h3c586ca5),
	.w8(32'hbb9472b2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c5cfc),
	.w1(32'h3c194ec9),
	.w2(32'h3c297548),
	.w3(32'hbbabc20a),
	.w4(32'hbb423d6e),
	.w5(32'hbbc4054f),
	.w6(32'hbb0e0acb),
	.w7(32'h3bd4235c),
	.w8(32'hbb4d829a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc871e),
	.w1(32'h3b7c02de),
	.w2(32'hbb42795b),
	.w3(32'hbc83df68),
	.w4(32'hbc63118d),
	.w5(32'hba998fd5),
	.w6(32'h3b9be4b9),
	.w7(32'h3b79d08e),
	.w8(32'hbbad4d06),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa40434),
	.w1(32'hbaf08501),
	.w2(32'h3b85d858),
	.w3(32'h3a807f4a),
	.w4(32'hbab90df1),
	.w5(32'h3c0a96b3),
	.w6(32'hbb402cca),
	.w7(32'hbbcdf62b),
	.w8(32'h3c4e5812),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68c98),
	.w1(32'hbb6a21c8),
	.w2(32'h3ae4bda7),
	.w3(32'h3ca6880f),
	.w4(32'h3c750e90),
	.w5(32'h39912014),
	.w6(32'h3c851de7),
	.w7(32'h3bd9b4d4),
	.w8(32'h3aab96d7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ec45a),
	.w1(32'h3ad311b9),
	.w2(32'h3b237952),
	.w3(32'hba27c6d7),
	.w4(32'h3a6bb6bc),
	.w5(32'h3ae45412),
	.w6(32'h3a80b413),
	.w7(32'h39c5fb5d),
	.w8(32'h3a2018d2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b331b5a),
	.w1(32'h3a85b331),
	.w2(32'hb8f5f044),
	.w3(32'hbb20f99e),
	.w4(32'hbb32cc24),
	.w5(32'hbbfe6713),
	.w6(32'h35bf16ad),
	.w7(32'h3a99642f),
	.w8(32'hbb2c7529),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c948220),
	.w1(32'h3be689c1),
	.w2(32'h3a9b4c26),
	.w3(32'hbc01d8e5),
	.w4(32'hbbe9147a),
	.w5(32'hbc1a6770),
	.w6(32'h3be4f876),
	.w7(32'hba1c7d90),
	.w8(32'h3b6399eb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be23cf0),
	.w1(32'h3c0dcd07),
	.w2(32'hbb1be0bf),
	.w3(32'hbc7f86c5),
	.w4(32'hbc27ea45),
	.w5(32'hbbe02409),
	.w6(32'hbba6eb0e),
	.w7(32'hbc12d1b8),
	.w8(32'hba95dbac),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ae14d),
	.w1(32'hb9efb187),
	.w2(32'h3b955e80),
	.w3(32'hbbb097d8),
	.w4(32'hbb7a9e61),
	.w5(32'h3baba00e),
	.w6(32'h3a093d9c),
	.w7(32'h39797fbe),
	.w8(32'h3b7783b1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c37b),
	.w1(32'h3b4e0c73),
	.w2(32'h3bb8577c),
	.w3(32'hba2daf4f),
	.w4(32'h3baafa4b),
	.w5(32'hbb182625),
	.w6(32'hbb89349e),
	.w7(32'h3b4a6a41),
	.w8(32'hbb58c1fc),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8611c5),
	.w1(32'h3c09847f),
	.w2(32'hba5ac8d3),
	.w3(32'hbbb9e5ca),
	.w4(32'hba8bbc26),
	.w5(32'hbbb2dbf2),
	.w6(32'hbbfeefa0),
	.w7(32'hbacdf1f5),
	.w8(32'hbb8f1778),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c620e3d),
	.w1(32'h3b2cd40e),
	.w2(32'hbc70b673),
	.w3(32'hbba1f043),
	.w4(32'hbc2dbe08),
	.w5(32'h3c5bf61c),
	.w6(32'h3a17e34a),
	.w7(32'hba99b17d),
	.w8(32'h3c2fa556),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc988355),
	.w1(32'hbc3d0765),
	.w2(32'hbbacba3f),
	.w3(32'h3d045851),
	.w4(32'h3d062514),
	.w5(32'hba296b45),
	.w6(32'h3c1899cd),
	.w7(32'h3c28b7b2),
	.w8(32'h3baa573e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8589e0),
	.w1(32'hbb28fcb3),
	.w2(32'hbb482dc8),
	.w3(32'h39f84c08),
	.w4(32'hb909a9b7),
	.w5(32'hbb03ed93),
	.w6(32'h3b97f64d),
	.w7(32'h3b8b3489),
	.w8(32'h3a99fe83),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b4f48),
	.w1(32'hba997b23),
	.w2(32'h3b8d9472),
	.w3(32'hbb8b7437),
	.w4(32'hbc082f72),
	.w5(32'hbc72f3b8),
	.w6(32'h3bf00d53),
	.w7(32'h3c04c094),
	.w8(32'h3c473142),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1983e4),
	.w1(32'hbb927350),
	.w2(32'hbb8bfb29),
	.w3(32'hbc259406),
	.w4(32'h3ab0c994),
	.w5(32'hbb0e272b),
	.w6(32'hbb635f55),
	.w7(32'hbc0e60e8),
	.w8(32'h3ba79516),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc290a13),
	.w1(32'hba4f3160),
	.w2(32'h3b3b0f74),
	.w3(32'hbb7da1d4),
	.w4(32'h3b38b595),
	.w5(32'hbc60a9df),
	.w6(32'hbc114417),
	.w7(32'hbb247044),
	.w8(32'h3b8c8fb0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb547d8),
	.w1(32'h3c319350),
	.w2(32'h3b529ba5),
	.w3(32'hbc5cf31a),
	.w4(32'hbc325720),
	.w5(32'hb9bccd22),
	.w6(32'h3c19cffd),
	.w7(32'h3c89b461),
	.w8(32'h3b93812f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b829),
	.w1(32'h3b4ce403),
	.w2(32'hba4f8a04),
	.w3(32'h3af1755a),
	.w4(32'h39fc80ed),
	.w5(32'hbab8caa1),
	.w6(32'h3babdcc1),
	.w7(32'h3b5cf96e),
	.w8(32'h3be2bd3f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6e3b7d),
	.w1(32'h3c4ddfbb),
	.w2(32'h3c06b64c),
	.w3(32'h3b5ddd07),
	.w4(32'h3c0aa933),
	.w5(32'h3a9f1f83),
	.w6(32'h3b8861a7),
	.w7(32'h3c48cc8a),
	.w8(32'h3a9c8a49),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa30c74),
	.w1(32'h3b5a167d),
	.w2(32'hbb3e4d5d),
	.w3(32'hbb742275),
	.w4(32'hba99d0c7),
	.w5(32'hbc622b36),
	.w6(32'hbafce57a),
	.w7(32'h3b4733dc),
	.w8(32'h3ba31a8e),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d6d4),
	.w1(32'h3baf4ce9),
	.w2(32'h3bd12ccc),
	.w3(32'hba905b92),
	.w4(32'hba87f551),
	.w5(32'hbc20f2df),
	.w6(32'h3bbe32f8),
	.w7(32'h38064635),
	.w8(32'hbba4a882),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c738fa5),
	.w1(32'h3c3a6257),
	.w2(32'h3be7dd6e),
	.w3(32'hbcc0b867),
	.w4(32'hbc950436),
	.w5(32'h3ba3e6ea),
	.w6(32'hbb896804),
	.w7(32'hbc3309ef),
	.w8(32'hbbb05499),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa242b2),
	.w1(32'h3bc742a9),
	.w2(32'h3ba0e1b2),
	.w3(32'hbc26ab4a),
	.w4(32'hbc09e36d),
	.w5(32'hbb8fe02a),
	.w6(32'hbb895b6c),
	.w7(32'h3aca8f08),
	.w8(32'h3b899b59),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14a80a),
	.w1(32'h3c1fa610),
	.w2(32'hbaac646b),
	.w3(32'hbc39e96d),
	.w4(32'hbc692b67),
	.w5(32'h3a48e9a1),
	.w6(32'hbbd4b1be),
	.w7(32'h3ba39597),
	.w8(32'h3b897f0a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72375f),
	.w1(32'h3ba28642),
	.w2(32'hba353fc7),
	.w3(32'h3b0bdca2),
	.w4(32'h3bcfef2e),
	.w5(32'hbb059256),
	.w6(32'h3a20c851),
	.w7(32'h3bd61fc3),
	.w8(32'h3b9d7cfa),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af53837),
	.w1(32'h3baff00f),
	.w2(32'h3bd9d910),
	.w3(32'h3a999b44),
	.w4(32'h3b62ecc7),
	.w5(32'hbc1fbee3),
	.w6(32'h3b35c1bd),
	.w7(32'h3bdc1205),
	.w8(32'hbb844fae),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2b6e5),
	.w1(32'h3c40bce7),
	.w2(32'h3c6942d3),
	.w3(32'hbc8c1f4e),
	.w4(32'hbc07b6d7),
	.w5(32'hbbe36c6d),
	.w6(32'hbc281269),
	.w7(32'hbad005a9),
	.w8(32'h379a0469),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7655f6),
	.w1(32'hbb04f5c7),
	.w2(32'h3bb147b3),
	.w3(32'hbc4eab23),
	.w4(32'hbc2be02f),
	.w5(32'h3b1682d6),
	.w6(32'h39d02747),
	.w7(32'h3b798e37),
	.w8(32'h3b9340c2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb8d17),
	.w1(32'h3a9c35a9),
	.w2(32'hbb1e7eba),
	.w3(32'h3ba57212),
	.w4(32'hb9a686b7),
	.w5(32'h3c256aa0),
	.w6(32'h3bcfe117),
	.w7(32'h3b146dc4),
	.w8(32'hbbc48c45),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61be20),
	.w1(32'hbc48a5b2),
	.w2(32'h3ae8cace),
	.w3(32'h3b2cf5aa),
	.w4(32'h3bca1531),
	.w5(32'h383b2646),
	.w6(32'hbc14a071),
	.w7(32'hbc9af309),
	.w8(32'h3ba9fc16),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e7a4),
	.w1(32'h3b8bd1f4),
	.w2(32'h3b343fae),
	.w3(32'h3aef9d18),
	.w4(32'h3b86ff40),
	.w5(32'h3a547bfd),
	.w6(32'h3b91ba1e),
	.w7(32'h3c1347c1),
	.w8(32'h3b3d8d5e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b624844),
	.w1(32'h3b82ee5e),
	.w2(32'h3b9bbde7),
	.w3(32'h3b26219a),
	.w4(32'h3b1860fd),
	.w5(32'hbc1aedc6),
	.w6(32'h3bac3cb6),
	.w7(32'h3bdac4fb),
	.w8(32'h3a965657),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba532fa8),
	.w1(32'hbab0cef5),
	.w2(32'hbc00e3b1),
	.w3(32'hbc79a167),
	.w4(32'hbcacc362),
	.w5(32'h3d4002a4),
	.w6(32'hbbc06820),
	.w7(32'h3904d9a4),
	.w8(32'hbc3e4ca1),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b410df9),
	.w1(32'h3c24da8e),
	.w2(32'h3ace76ae),
	.w3(32'h3d7f5244),
	.w4(32'h3ca96522),
	.w5(32'hbb750363),
	.w6(32'hbbf37945),
	.w7(32'hbc862609),
	.w8(32'h3ba01576),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e3df1),
	.w1(32'hb9584849),
	.w2(32'h3ba74d4a),
	.w3(32'hbb9fbfba),
	.w4(32'hbb01081b),
	.w5(32'hbc85bc9e),
	.w6(32'h3caac325),
	.w7(32'h3c4bd7b8),
	.w8(32'h3b013bc7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c559496),
	.w1(32'hbaf4d133),
	.w2(32'hbbeec327),
	.w3(32'hbcb676ad),
	.w4(32'hbc8768c4),
	.w5(32'hbb88f8e3),
	.w6(32'hbb92a8af),
	.w7(32'hbba744ad),
	.w8(32'hba269f7d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc403c70),
	.w1(32'hbc50e06f),
	.w2(32'h3b247526),
	.w3(32'h39a2423b),
	.w4(32'h3b2fcac2),
	.w5(32'h3bad017b),
	.w6(32'hbc20d1ab),
	.w7(32'hbac05fa9),
	.w8(32'h3bc6ee1c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c202d),
	.w1(32'h3b7e1019),
	.w2(32'hbc133b69),
	.w3(32'hbc05757b),
	.w4(32'hb9efa213),
	.w5(32'h3cc59d40),
	.w6(32'h3a20b6a0),
	.w7(32'h3b57641e),
	.w8(32'hbb9e3ad4),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0999fb),
	.w1(32'hbbc814fe),
	.w2(32'hba35bda7),
	.w3(32'h3cc2b662),
	.w4(32'h3cb55039),
	.w5(32'h3c7dc569),
	.w6(32'h3ba427f6),
	.w7(32'hbbd2edca),
	.w8(32'h3b91c18c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2bbe2),
	.w1(32'hbc25e269),
	.w2(32'h3bf1812c),
	.w3(32'h3cd3b79e),
	.w4(32'h3cef547e),
	.w5(32'h3bd47908),
	.w6(32'hbbc0338f),
	.w7(32'hbc0fb5a5),
	.w8(32'h3ad6d810),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b8c9d),
	.w1(32'h3b5d4025),
	.w2(32'h3b78d146),
	.w3(32'h3c6308a8),
	.w4(32'h3b993f42),
	.w5(32'h3c175c9a),
	.w6(32'h3c23a295),
	.w7(32'hba8edea9),
	.w8(32'hba923e66),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b9d4b),
	.w1(32'h3b079bb2),
	.w2(32'h3b72f432),
	.w3(32'h3b21c0c0),
	.w4(32'h3b8d4682),
	.w5(32'hbc301513),
	.w6(32'hbbb97cfb),
	.w7(32'h3bc52846),
	.w8(32'hbbe3c2b3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbca2f3),
	.w1(32'h3bacf085),
	.w2(32'hbb7c05e7),
	.w3(32'hbcea151b),
	.w4(32'hbca2a0e4),
	.w5(32'hba00f64f),
	.w6(32'hbc554d44),
	.w7(32'hbc0c1d2f),
	.w8(32'hba3c694a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4292ad),
	.w1(32'h3ba3b61b),
	.w2(32'hbbc2ddbf),
	.w3(32'h3a95ef55),
	.w4(32'h3b8e8a11),
	.w5(32'hbba65068),
	.w6(32'hbad6bbbd),
	.w7(32'h3b905388),
	.w8(32'hbbbb9403),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2747c),
	.w1(32'hba88e341),
	.w2(32'hbc3e9c8e),
	.w3(32'hbbb09be9),
	.w4(32'hbb39dab5),
	.w5(32'hbb23b03c),
	.w6(32'hbbbd57ed),
	.w7(32'hbb0beb2d),
	.w8(32'h3b9dfa18),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ad00),
	.w1(32'h3a2ca674),
	.w2(32'h3b761d07),
	.w3(32'hbba3c6cf),
	.w4(32'h3b829b48),
	.w5(32'hbbe6dff8),
	.w6(32'hbb393675),
	.w7(32'hbb7e76db),
	.w8(32'hbb9d6ede),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5e91a),
	.w1(32'h3a6987c0),
	.w2(32'hbbc1b375),
	.w3(32'hbc78a5a5),
	.w4(32'hbc3a00eb),
	.w5(32'h3b7d77d3),
	.w6(32'hbc162353),
	.w7(32'hbbf34284),
	.w8(32'h3bfa2476),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76c455),
	.w1(32'hbb07e930),
	.w2(32'h3bad91aa),
	.w3(32'h3c8157d7),
	.w4(32'h3c84139a),
	.w5(32'hbc92b7db),
	.w6(32'h3b32d427),
	.w7(32'h3bddab1f),
	.w8(32'hbbd9401e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2398),
	.w1(32'hba03a619),
	.w2(32'h3c5a5977),
	.w3(32'hbcb86ccc),
	.w4(32'hbc4a7852),
	.w5(32'h3af24fe9),
	.w6(32'h3bf9902f),
	.w7(32'h3b4c65cb),
	.w8(32'h3aacda9d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91c71a),
	.w1(32'h3c9c3282),
	.w2(32'h3c216ade),
	.w3(32'h3bc57776),
	.w4(32'h3c2830bc),
	.w5(32'hbb95dbe3),
	.w6(32'h3c187d7b),
	.w7(32'h3c917483),
	.w8(32'h3bb96956),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d07ee),
	.w1(32'h3c329abe),
	.w2(32'hbbca0d73),
	.w3(32'h3aba634a),
	.w4(32'hbbf9fa35),
	.w5(32'hbbc2ef40),
	.w6(32'hbb117eb6),
	.w7(32'hbb573dfa),
	.w8(32'hbbdf2436),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d964),
	.w1(32'hbbdec76b),
	.w2(32'hbb8defcd),
	.w3(32'h39bad7f9),
	.w4(32'h3bb1c2df),
	.w5(32'hbaa837a2),
	.w6(32'hbbfec36f),
	.w7(32'hbbb2c015),
	.w8(32'hbb0beb84),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ebd5),
	.w1(32'hbc196876),
	.w2(32'h3b74ecb8),
	.w3(32'hbb286e61),
	.w4(32'hbaeabf7d),
	.w5(32'h39e79575),
	.w6(32'hbc90ca87),
	.w7(32'hbcac62dc),
	.w8(32'hbaf87a17),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e56a9),
	.w1(32'h3bf7fb80),
	.w2(32'h3bde428c),
	.w3(32'h3a5e1d8d),
	.w4(32'h3af0eeae),
	.w5(32'hbbdd8bfe),
	.w6(32'hbb700da4),
	.w7(32'hbacde00a),
	.w8(32'h3c388b71),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34424a),
	.w1(32'hbb6c4c42),
	.w2(32'hbb295e23),
	.w3(32'hbbd589ef),
	.w4(32'hbb9b5bf0),
	.w5(32'hbb229247),
	.w6(32'h3c1da4a0),
	.w7(32'h3bc2896a),
	.w8(32'hbb865b12),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e074),
	.w1(32'h3b34d75f),
	.w2(32'hbc345dd8),
	.w3(32'hbaa393e3),
	.w4(32'hba0da9cb),
	.w5(32'h3b4fa0e9),
	.w6(32'hbb914623),
	.w7(32'hbb9905ac),
	.w8(32'h3bc71303),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca12668),
	.w1(32'hbc622687),
	.w2(32'h3a7be86e),
	.w3(32'h3beefa1c),
	.w4(32'h3bc6fa7f),
	.w5(32'h3ca44aeb),
	.w6(32'hbbb082b9),
	.w7(32'hbbda17b7),
	.w8(32'h3a09156c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a9443),
	.w1(32'hbbba58af),
	.w2(32'h3ba54dd6),
	.w3(32'h3cd23ff3),
	.w4(32'h3ca10ea6),
	.w5(32'h3b14e3ca),
	.w6(32'h3beab10d),
	.w7(32'h3b1c3302),
	.w8(32'hb8cd4aa6),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b273c12),
	.w1(32'hbaddaa86),
	.w2(32'h3abef679),
	.w3(32'hbc19f4d8),
	.w4(32'hbc889762),
	.w5(32'h3af0d7f8),
	.w6(32'hbb97d4c4),
	.w7(32'hba93efd7),
	.w8(32'hba213435),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d46a9),
	.w1(32'h3b6c5977),
	.w2(32'h3b945b35),
	.w3(32'h3ad01ffa),
	.w4(32'h3b67159e),
	.w5(32'h39d236d2),
	.w6(32'hbb4c4f70),
	.w7(32'hb9f71807),
	.w8(32'h3a838739),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada34c5),
	.w1(32'h3b5ba886),
	.w2(32'h3c217152),
	.w3(32'hba0c0168),
	.w4(32'hbb0e4807),
	.w5(32'hbb7554c2),
	.w6(32'hb99447ad),
	.w7(32'h3b2276d9),
	.w8(32'h3abee470),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cc35a),
	.w1(32'h3c82fb55),
	.w2(32'h3b67798d),
	.w3(32'hbc064ac7),
	.w4(32'hbc53363a),
	.w5(32'h3b1ec7dd),
	.w6(32'h3a998aa2),
	.w7(32'h3ae41207),
	.w8(32'h3a074240),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b328ff9),
	.w1(32'h3b546ae6),
	.w2(32'h3bb3282c),
	.w3(32'h3b514cfe),
	.w4(32'h3b8a90e4),
	.w5(32'hbc87ec3c),
	.w6(32'h3b2505f0),
	.w7(32'h3ba8e2a5),
	.w8(32'hbbd0476d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16b827),
	.w1(32'h3c19ee98),
	.w2(32'h3ba4a16f),
	.w3(32'hbbbb286f),
	.w4(32'hbbbcd8aa),
	.w5(32'hbc4e91b2),
	.w6(32'h3b47d8f5),
	.w7(32'h3bd84f1f),
	.w8(32'hb9fc6cc7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c910c16),
	.w1(32'h3c348a1d),
	.w2(32'hb9d18441),
	.w3(32'hbc78e3cd),
	.w4(32'hbc3f11a5),
	.w5(32'hbace6341),
	.w6(32'h3adde668),
	.w7(32'h3b313640),
	.w8(32'hbaf2cb74),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dcf97),
	.w1(32'h3c42052a),
	.w2(32'h3c001a0c),
	.w3(32'hbc2382df),
	.w4(32'hbc0be14b),
	.w5(32'h3abd1896),
	.w6(32'h3b081fa7),
	.w7(32'h3bf248d2),
	.w8(32'hbc098a48),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule