module layer_8_featuremap_147(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3339f),
	.w1(32'h3be6d73b),
	.w2(32'h3c015cb3),
	.w3(32'h3b81d9f6),
	.w4(32'h3bd0db9e),
	.w5(32'h3c143a1a),
	.w6(32'h3c1c32b5),
	.w7(32'h3c3dd203),
	.w8(32'h3c557f1a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc13436),
	.w1(32'hbbbb29be),
	.w2(32'hbb4e25ac),
	.w3(32'hbbb306dc),
	.w4(32'hbb6cf107),
	.w5(32'hba8658c4),
	.w6(32'hbb5ab7be),
	.w7(32'hbac6a6b3),
	.w8(32'h3aa12850),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd05bb4),
	.w1(32'hbbcefe04),
	.w2(32'hbbc44b21),
	.w3(32'hbbe3345a),
	.w4(32'hbbbe43b7),
	.w5(32'hbbcc97e2),
	.w6(32'hbbb832e7),
	.w7(32'hbba9a369),
	.w8(32'hbb975afc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9016a79),
	.w1(32'hb93944bc),
	.w2(32'hb8a4faab),
	.w3(32'h3931b52e),
	.w4(32'h397dfb88),
	.w5(32'h39b92980),
	.w6(32'h39225a72),
	.w7(32'h39a05085),
	.w8(32'h39eeb4b9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14b631),
	.w1(32'h3a8d44f0),
	.w2(32'hb8e1b15d),
	.w3(32'hba95d8ce),
	.w4(32'h3affe615),
	.w5(32'h3b6f9c42),
	.w6(32'hbaa59f0d),
	.w7(32'h3b0937fc),
	.w8(32'h3ba23359),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0d83),
	.w1(32'hbbd420a7),
	.w2(32'hbba06ade),
	.w3(32'hbb94bdaa),
	.w4(32'hbbc6cf0e),
	.w5(32'hbbf7557a),
	.w6(32'hbbb30015),
	.w7(32'hbbecb0ac),
	.w8(32'hbbea8d1e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36993ed1),
	.w1(32'h372f5f2d),
	.w2(32'hb85a759b),
	.w3(32'h35f6903b),
	.w4(32'hb68ddd24),
	.w5(32'hb7d4c0d1),
	.w6(32'h3814be1b),
	.w7(32'hb60b5448),
	.w8(32'hb7e564e4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc81f44),
	.w1(32'hbb10d8d6),
	.w2(32'hbb2457b7),
	.w3(32'hbb3ff9a5),
	.w4(32'h3b33c07a),
	.w5(32'h3b2ea266),
	.w6(32'hbb387666),
	.w7(32'h3b7f6ddb),
	.w8(32'h3b69241d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0a9d),
	.w1(32'hbb2f999a),
	.w2(32'h39ad2ff5),
	.w3(32'hbbd5764a),
	.w4(32'hbabc85cb),
	.w5(32'h39c300d3),
	.w6(32'h39865b20),
	.w7(32'h3b6e0819),
	.w8(32'h3bdeb05a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11b42d),
	.w1(32'hbbc5424e),
	.w2(32'hbb82c1a4),
	.w3(32'hbc021d19),
	.w4(32'hbbb8ba92),
	.w5(32'hbb90dd98),
	.w6(32'hbbb37f69),
	.w7(32'hbb53e861),
	.w8(32'hbb0bf55a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ab44f),
	.w1(32'h3bbee7b8),
	.w2(32'h3c0c8a2e),
	.w3(32'h3af5e922),
	.w4(32'h3bddf247),
	.w5(32'h3c3ae781),
	.w6(32'h3b4adb73),
	.w7(32'h3bc308de),
	.w8(32'h3c2e0d5b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f1fe),
	.w1(32'hbaa43f4f),
	.w2(32'h39229247),
	.w3(32'hbb183bd3),
	.w4(32'hbac2c45a),
	.w5(32'hb8f92edb),
	.w6(32'hba9e9255),
	.w7(32'hbab29ade),
	.w8(32'h39945b25),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4c230),
	.w1(32'hbbba54b7),
	.w2(32'hbb8eae35),
	.w3(32'hbbacce25),
	.w4(32'hbb9a5618),
	.w5(32'hbbefed84),
	.w6(32'hbb0056f3),
	.w7(32'h380de2ca),
	.w8(32'hb9c969ab),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83d98),
	.w1(32'hbab24b48),
	.w2(32'hbaa47131),
	.w3(32'hbb93f005),
	.w4(32'hbb8f13d7),
	.w5(32'hbb831460),
	.w6(32'hbaa5812c),
	.w7(32'hbb3d673d),
	.w8(32'hbb4d79b4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9c95),
	.w1(32'hb7b3c7d7),
	.w2(32'hbaf3f053),
	.w3(32'hbb2261ce),
	.w4(32'hbad302c4),
	.w5(32'hbb56032e),
	.w6(32'hba09fe4e),
	.w7(32'hbacc1bdf),
	.w8(32'hbaedccb3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91d5b0),
	.w1(32'h392861ad),
	.w2(32'h3be97d0f),
	.w3(32'hba1fb165),
	.w4(32'h3bb60e87),
	.w5(32'h3af05d6f),
	.w6(32'h3acce33e),
	.w7(32'h3ab410ca),
	.w8(32'h3928dad0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c347439),
	.w1(32'h3b607375),
	.w2(32'hba155558),
	.w3(32'hbb854093),
	.w4(32'h39c2b08e),
	.w5(32'h3c012b54),
	.w6(32'h3af7e0af),
	.w7(32'h3b666d63),
	.w8(32'h3bc9e00e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4b55),
	.w1(32'hbc27a336),
	.w2(32'hbc1b5d2e),
	.w3(32'hbb393470),
	.w4(32'hbbf9e62a),
	.w5(32'h3a2d5ada),
	.w6(32'hbbf12331),
	.w7(32'h39e0f4af),
	.w8(32'hbb4f4485),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37fab),
	.w1(32'h3c90a431),
	.w2(32'h3b823e74),
	.w3(32'h3b798358),
	.w4(32'h3c7c6ee3),
	.w5(32'h3ca95d5e),
	.w6(32'hbbdcda2b),
	.w7(32'h3b2b9f1d),
	.w8(32'h3bc8f1f7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cb620),
	.w1(32'h3b8a6927),
	.w2(32'h3c35e2f5),
	.w3(32'h3c29be55),
	.w4(32'h3ad3c7cb),
	.w5(32'h3bf34130),
	.w6(32'h384e1b58),
	.w7(32'h3c2dd1f2),
	.w8(32'h3c8f0485),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a9414),
	.w1(32'h3c0e193b),
	.w2(32'h3c1ffd09),
	.w3(32'hbc06daf8),
	.w4(32'hbb49ef1a),
	.w5(32'hb9fe42ee),
	.w6(32'hb8f142e2),
	.w7(32'h3bb2d8e0),
	.w8(32'h3ba7bd75),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1602e9),
	.w1(32'hbc7966c6),
	.w2(32'hbc1431ac),
	.w3(32'hbc48f05c),
	.w4(32'hbc59f243),
	.w5(32'hbc0de84d),
	.w6(32'hbbdf7ca5),
	.w7(32'hbb511db3),
	.w8(32'hbbd7fbd9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c2e84),
	.w1(32'h3c292e5e),
	.w2(32'h3bf9d1bf),
	.w3(32'hbbab08c0),
	.w4(32'h3b27ad9a),
	.w5(32'h3bff92bf),
	.w6(32'hba474641),
	.w7(32'h3c4dc491),
	.w8(32'h3c915c47),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81d4b6),
	.w1(32'h3c2b311e),
	.w2(32'h3aeffba6),
	.w3(32'hbc9d8890),
	.w4(32'h3c07d38c),
	.w5(32'h3bd033a7),
	.w6(32'h3a9d8a66),
	.w7(32'h3bc6d19a),
	.w8(32'h3b38cc49),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb417e4),
	.w1(32'h398f3db7),
	.w2(32'hbbcf3646),
	.w3(32'h3aa37fe9),
	.w4(32'hba5b3efa),
	.w5(32'hbb6d0ee2),
	.w6(32'h3ac1cca1),
	.w7(32'hbbf9533e),
	.w8(32'hbbafdc3c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a19f),
	.w1(32'h3c3781c6),
	.w2(32'h3babb1fb),
	.w3(32'h3bae7ef3),
	.w4(32'h3cbf50a4),
	.w5(32'h3ce2a6fa),
	.w6(32'h3bda5b32),
	.w7(32'h3c835116),
	.w8(32'h3cb33812),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab720b),
	.w1(32'hbbe81b26),
	.w2(32'h3ad1454d),
	.w3(32'h3c11c470),
	.w4(32'hbb2472f2),
	.w5(32'hb81c84f1),
	.w6(32'h3b113929),
	.w7(32'hbaf2c19d),
	.w8(32'h3983a130),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dcf221b),
	.w1(32'h3d1fd737),
	.w2(32'h3d94da58),
	.w3(32'h3ce0ea30),
	.w4(32'h3b433e8a),
	.w5(32'h3d33a765),
	.w6(32'h3d3c144a),
	.w7(32'h3d8e698e),
	.w8(32'h3da8fcd2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d10da),
	.w1(32'h3c8176d5),
	.w2(32'h3b932621),
	.w3(32'h3cb9f1f0),
	.w4(32'h3c077c3e),
	.w5(32'h3bfae333),
	.w6(32'h3d0f7600),
	.w7(32'h3c62859a),
	.w8(32'hb846ab0f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb488800),
	.w1(32'h3b033087),
	.w2(32'hbafffd31),
	.w3(32'h3b827a92),
	.w4(32'h3ba6e2c0),
	.w5(32'hbbe70a22),
	.w6(32'hbace9ecc),
	.w7(32'hbb19e118),
	.w8(32'hbc2bf85a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ea8a7),
	.w1(32'h3bd4d5d9),
	.w2(32'hbaedb1a2),
	.w3(32'h3bb2a2a4),
	.w4(32'hbb4181b6),
	.w5(32'hbbb21724),
	.w6(32'h3be7068b),
	.w7(32'hbad3912e),
	.w8(32'hbb28c14d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea02e),
	.w1(32'hba9669fc),
	.w2(32'h3bd64810),
	.w3(32'hbb82513a),
	.w4(32'hbbc1ad67),
	.w5(32'hbbe2bf91),
	.w6(32'hba312541),
	.w7(32'h3a9c235a),
	.w8(32'h39529387),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b193ce),
	.w1(32'hbae9f0ff),
	.w2(32'hbc62c708),
	.w3(32'hbc07293a),
	.w4(32'hbab156c3),
	.w5(32'hbb10edab),
	.w6(32'hbb679e9a),
	.w7(32'hbbcbf1ae),
	.w8(32'hbb56b807),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f52f3),
	.w1(32'hbbbe38f2),
	.w2(32'hb8b58097),
	.w3(32'hbc245db3),
	.w4(32'h3b8605df),
	.w5(32'h3c206807),
	.w6(32'hbc62e00f),
	.w7(32'h3b0b6b53),
	.w8(32'h3b5de1eb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4a71b),
	.w1(32'hbc7963bf),
	.w2(32'hba300986),
	.w3(32'h3c59738c),
	.w4(32'hbb5bf029),
	.w5(32'hbb471cf4),
	.w6(32'hbc43eb02),
	.w7(32'hbc0f07c8),
	.w8(32'hbb45ba1b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd88f85),
	.w1(32'h3c39c323),
	.w2(32'h3a94d953),
	.w3(32'h3c05637e),
	.w4(32'h3a068fb7),
	.w5(32'h3a21aa4e),
	.w6(32'h3c49da22),
	.w7(32'hbbb067d4),
	.w8(32'h3b7c1e42),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb358401),
	.w1(32'hba08b4d4),
	.w2(32'hbbde7aa0),
	.w3(32'hbb90ad5e),
	.w4(32'h3b378603),
	.w5(32'h3bc00ade),
	.w6(32'hbbf37c9e),
	.w7(32'hbbf34ca6),
	.w8(32'hbc308a06),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc132511),
	.w1(32'hbbf67997),
	.w2(32'hbc246562),
	.w3(32'hbbf0f174),
	.w4(32'hbb15bb4d),
	.w5(32'hb9fa265a),
	.w6(32'hbc7144ed),
	.w7(32'hbb93fe96),
	.w8(32'hbb271842),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65208d),
	.w1(32'hbb83d34f),
	.w2(32'hbb6b380d),
	.w3(32'h3b2af1b0),
	.w4(32'hbb805f17),
	.w5(32'h3bcddd82),
	.w6(32'hba72bd0f),
	.w7(32'h3bd21e89),
	.w8(32'hbb30dbef),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81f7af),
	.w1(32'hbac22ad8),
	.w2(32'h3b9dbe49),
	.w3(32'h3b1470b3),
	.w4(32'hbbaa546a),
	.w5(32'hbbfe2dd8),
	.w6(32'hbb810fa6),
	.w7(32'h3aad2ffc),
	.w8(32'h3b2a79aa),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69407c),
	.w1(32'h3baf1ffd),
	.w2(32'h3c0bcc68),
	.w3(32'hbbfe527e),
	.w4(32'h3b96adae),
	.w5(32'h3babe9d3),
	.w6(32'h3bbc1167),
	.w7(32'h3b9c2503),
	.w8(32'h3c1e8f07),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23c9dc),
	.w1(32'hbc4b4d4d),
	.w2(32'h3b8446bb),
	.w3(32'hbb368501),
	.w4(32'h3968a723),
	.w5(32'hba4d163b),
	.w6(32'hb9f3d529),
	.w7(32'hbb5ce3de),
	.w8(32'h3bf93f2d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcda243),
	.w1(32'h3bbb92f2),
	.w2(32'hbbd513f5),
	.w3(32'h3ad0f7d6),
	.w4(32'h3a06bf7b),
	.w5(32'h3b0ef528),
	.w6(32'h3c878b07),
	.w7(32'h3b3780ad),
	.w8(32'hbc5b53cb),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072c0a),
	.w1(32'h3c03b927),
	.w2(32'h3b6d6b92),
	.w3(32'h3aa36252),
	.w4(32'h3b7a0176),
	.w5(32'h3b86d8cc),
	.w6(32'hbbe1771c),
	.w7(32'h3bb78212),
	.w8(32'h3bfe9e85),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b507a85),
	.w1(32'h3b63ecc7),
	.w2(32'h3af4499e),
	.w3(32'h37c18c4a),
	.w4(32'h3b48d790),
	.w5(32'h3beb0c90),
	.w6(32'h3ac6d965),
	.w7(32'h3c18ca44),
	.w8(32'h3baaa480),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4a557),
	.w1(32'hbb03ccfa),
	.w2(32'h3b87a83b),
	.w3(32'hbaf5862b),
	.w4(32'h3b07741a),
	.w5(32'hbbaad7b8),
	.w6(32'h3aec3096),
	.w7(32'h3b23bf2e),
	.w8(32'hbbcb778a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ac2b2),
	.w1(32'h3b9ec1d9),
	.w2(32'hbb953d1a),
	.w3(32'hbc46acdc),
	.w4(32'hbb159939),
	.w5(32'hbb1e66db),
	.w6(32'h3af2024f),
	.w7(32'hbb631aa7),
	.w8(32'hbc31616e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ebd5a),
	.w1(32'hbb17927a),
	.w2(32'h3ab49531),
	.w3(32'hbbeb3178),
	.w4(32'h3a973f56),
	.w5(32'h3c23c835),
	.w6(32'hbc0f28f8),
	.w7(32'h3bd31910),
	.w8(32'h3b94eb17),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62ebfc),
	.w1(32'hbba1353d),
	.w2(32'h3bb4b85e),
	.w3(32'hbb38296e),
	.w4(32'h3b3decfe),
	.w5(32'h3bf98b74),
	.w6(32'hbc0171c0),
	.w7(32'h3c269270),
	.w8(32'h3c47e1bf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0062ed),
	.w1(32'h3bb8692b),
	.w2(32'h3c21af8f),
	.w3(32'h3b313795),
	.w4(32'h3b8072ec),
	.w5(32'h3bb1a4d2),
	.w6(32'h3ba8cffc),
	.w7(32'h3c02f1ba),
	.w8(32'h3b43c84c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9814b8),
	.w1(32'h3b60baaf),
	.w2(32'hbc66cae8),
	.w3(32'hbbcd1ccd),
	.w4(32'hb95564c3),
	.w5(32'hbac34392),
	.w6(32'hbb30b636),
	.w7(32'hbc4b11e7),
	.w8(32'h3c26785a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae177de),
	.w1(32'hbb28062c),
	.w2(32'h3c8ad295),
	.w3(32'h3b6b5e38),
	.w4(32'h3c3f97e7),
	.w5(32'h3c7a4770),
	.w6(32'hbc256e6c),
	.w7(32'h3c080827),
	.w8(32'h3c5812c1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c78f8),
	.w1(32'h3b26fd6c),
	.w2(32'h3bbca24c),
	.w3(32'h3acf4287),
	.w4(32'h3b273f80),
	.w5(32'h3beaf441),
	.w6(32'hb9d3c9b0),
	.w7(32'h3c5298ea),
	.w8(32'h3ce4d751),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb792305),
	.w1(32'hb99f9e81),
	.w2(32'h3b43735a),
	.w3(32'h3a9ea0f8),
	.w4(32'h3a96bb2c),
	.w5(32'h3a6d1c9f),
	.w6(32'h3b815ac6),
	.w7(32'h3a935d60),
	.w8(32'h3a06379a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ababd),
	.w1(32'h3adb4a48),
	.w2(32'h3a690767),
	.w3(32'hbab79211),
	.w4(32'hbb4f89b4),
	.w5(32'hbbe5d5ab),
	.w6(32'h3a924c3a),
	.w7(32'h39665f67),
	.w8(32'hbb98673a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d29b1),
	.w1(32'h3b6048a3),
	.w2(32'h3be6d944),
	.w3(32'hbc6962b3),
	.w4(32'h3b5930ef),
	.w5(32'h3c26e3f1),
	.w6(32'h3b8a263b),
	.w7(32'h3c01cd0c),
	.w8(32'h3bd20c9a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c47d7),
	.w1(32'hbc271a11),
	.w2(32'h3c3c6553),
	.w3(32'hbb6b7ae5),
	.w4(32'hbbaf6c0b),
	.w5(32'hbbcc7b41),
	.w6(32'hbc179a77),
	.w7(32'h3afc843c),
	.w8(32'h3c78e98f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e6f04),
	.w1(32'hbb065987),
	.w2(32'hba49eb58),
	.w3(32'h3bcd2a3e),
	.w4(32'h3c702d00),
	.w5(32'h3c59a029),
	.w6(32'h3c1e9ee3),
	.w7(32'h3c18edb7),
	.w8(32'h3c9d7caf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b447d42),
	.w1(32'h3c5933b7),
	.w2(32'h3b3b7d1f),
	.w3(32'h3ccee451),
	.w4(32'h3b3ee6db),
	.w5(32'h3b2cfc5a),
	.w6(32'h3caaaefb),
	.w7(32'h3b79d58e),
	.w8(32'h3baac015),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9b8f1),
	.w1(32'h3a842f3e),
	.w2(32'h3b8e7b70),
	.w3(32'hbb0f6966),
	.w4(32'h3bd7d79d),
	.w5(32'h3bfa6f5f),
	.w6(32'h399576c8),
	.w7(32'h3b55d97d),
	.w8(32'h3bcba9e2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ed707),
	.w1(32'hbb01a6d9),
	.w2(32'hbb5656a2),
	.w3(32'hb692a278),
	.w4(32'h3b55220b),
	.w5(32'hbb9d6812),
	.w6(32'hbacf44cc),
	.w7(32'hbb9ef853),
	.w8(32'h3ba29ce0),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b65e5),
	.w1(32'hbbfa0507),
	.w2(32'hbbdd1246),
	.w3(32'hbb2d59f4),
	.w4(32'hba92058a),
	.w5(32'h3ae48a30),
	.w6(32'hba8a2f0d),
	.w7(32'hbbe6c08b),
	.w8(32'hbbc0838c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10f4c8),
	.w1(32'h39b2495f),
	.w2(32'h3c366dff),
	.w3(32'h3bb473aa),
	.w4(32'h3bf8bb2d),
	.w5(32'h3c904b63),
	.w6(32'hbab2ebfc),
	.w7(32'h3c0daf47),
	.w8(32'h3c29e041),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a426290),
	.w1(32'hbb3daefb),
	.w2(32'hbb8c18ea),
	.w3(32'h3ba4d119),
	.w4(32'hbb4cb89c),
	.w5(32'hbb197478),
	.w6(32'hbb0fcfb7),
	.w7(32'h3b425960),
	.w8(32'h3b46c55d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ebbbe),
	.w1(32'hbb220c58),
	.w2(32'h3c477ba8),
	.w3(32'h3b18b903),
	.w4(32'h39a7f942),
	.w5(32'hbad8d000),
	.w6(32'h3b9d0a74),
	.w7(32'h3a9ce02e),
	.w8(32'hba16e2e9),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c377fbb),
	.w1(32'h3c8a6e4b),
	.w2(32'hbb40aeaa),
	.w3(32'hbc090287),
	.w4(32'h3a4ae610),
	.w5(32'hba3a61a0),
	.w6(32'h39cc2ef4),
	.w7(32'hbbc5dde4),
	.w8(32'hbb5f511c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376f03),
	.w1(32'h3aca181b),
	.w2(32'hba56b7ad),
	.w3(32'hbb4db2e9),
	.w4(32'h39a2f27f),
	.w5(32'h3b877d0d),
	.w6(32'hbbcddd58),
	.w7(32'h3b298507),
	.w8(32'h3bcff73e),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65fc3a),
	.w1(32'hb991cf39),
	.w2(32'hb9b09eca),
	.w3(32'h3c15baf4),
	.w4(32'h3b2409a4),
	.w5(32'h3ad78a5a),
	.w6(32'h3bc38b09),
	.w7(32'h392d91b1),
	.w8(32'h39a9f56f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12d9a7),
	.w1(32'hbc0ac2c5),
	.w2(32'h38736d7b),
	.w3(32'hba3b6479),
	.w4(32'hbb0060ba),
	.w5(32'h3a1617ff),
	.w6(32'hbbf00e1b),
	.w7(32'h3ae81875),
	.w8(32'hbb5be503),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cc30d),
	.w1(32'h3c78ecb2),
	.w2(32'h3c504ad8),
	.w3(32'hbac4fa3b),
	.w4(32'hbb110509),
	.w5(32'h3bcd8672),
	.w6(32'h3b9451d4),
	.w7(32'hbbdc1e5e),
	.w8(32'h3c552288),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a872996),
	.w1(32'hbb8b9d99),
	.w2(32'h3ae3287b),
	.w3(32'h3b998fc3),
	.w4(32'hbb152638),
	.w5(32'hbc428710),
	.w6(32'hb779032d),
	.w7(32'hbbfab9b7),
	.w8(32'hbbdbe968),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c846fae),
	.w1(32'h3c884684),
	.w2(32'hbbeb108d),
	.w3(32'hbb80789d),
	.w4(32'h3be35963),
	.w5(32'h3b5bcb2b),
	.w6(32'h3c20ccfe),
	.w7(32'h3bb97426),
	.w8(32'hbb032d10),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3ed59),
	.w1(32'hbba76c50),
	.w2(32'h3a00edf1),
	.w3(32'hbc02bb8a),
	.w4(32'h3bca9947),
	.w5(32'h3a94dc36),
	.w6(32'hbbf14e62),
	.w7(32'hbb2df6c2),
	.w8(32'h3a919f95),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f207),
	.w1(32'h3b0a47f9),
	.w2(32'h3b0318e9),
	.w3(32'hbbd0034d),
	.w4(32'hbb75d8d6),
	.w5(32'hbbd9d501),
	.w6(32'hbb12aed6),
	.w7(32'hbaecfe8b),
	.w8(32'h3c7e2c60),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7f31b),
	.w1(32'hbb51a44c),
	.w2(32'hbb8ecc39),
	.w3(32'h3b8bc397),
	.w4(32'h3b215d0d),
	.w5(32'h3c2b515b),
	.w6(32'h3c481828),
	.w7(32'h3b278774),
	.w8(32'hbbfc31cb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4c89),
	.w1(32'h3b8dcf5d),
	.w2(32'h3946a085),
	.w3(32'hb72da1dd),
	.w4(32'h3ad08391),
	.w5(32'h3b9437ec),
	.w6(32'hbb33ffa5),
	.w7(32'h3beb4998),
	.w8(32'hb95ee632),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0bbe6),
	.w1(32'h3b81a4fc),
	.w2(32'hbbf061f5),
	.w3(32'hbaf0c43f),
	.w4(32'hb9690be3),
	.w5(32'hbadf1a11),
	.w6(32'h3ab93413),
	.w7(32'hbb69f3df),
	.w8(32'hbbaa125a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb380ac),
	.w1(32'hbacecab8),
	.w2(32'h3bbcb46a),
	.w3(32'h3bb74d23),
	.w4(32'h3c085e87),
	.w5(32'h3c85490e),
	.w6(32'h3b8f38d7),
	.w7(32'h3c389b00),
	.w8(32'h3c7d6cc2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5a48),
	.w1(32'h399996ca),
	.w2(32'hba9983e9),
	.w3(32'h3b9c15a7),
	.w4(32'h39b1cb8a),
	.w5(32'h3b4114d2),
	.w6(32'h3bb65778),
	.w7(32'hb905a33e),
	.w8(32'hb9f6b982),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcc7b9),
	.w1(32'hbaae72f0),
	.w2(32'h3b62327f),
	.w3(32'hba8ce723),
	.w4(32'hb885dfd6),
	.w5(32'h3bb44791),
	.w6(32'h3a494f9b),
	.w7(32'h3c4d8710),
	.w8(32'h3c1bcd83),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b339564),
	.w1(32'hbadd11d6),
	.w2(32'hbbfd5644),
	.w3(32'h3bea669f),
	.w4(32'h3b56eea1),
	.w5(32'h3c137d62),
	.w6(32'h3c01c948),
	.w7(32'hbb9f9be7),
	.w8(32'h3c6334b3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c6d2e),
	.w1(32'h3bbaa229),
	.w2(32'hbbe3b517),
	.w3(32'hbb4902a5),
	.w4(32'h39211ae5),
	.w5(32'hbbdb28a8),
	.w6(32'hba8a3516),
	.w7(32'hbbbeb5c5),
	.w8(32'hbbaaa7f9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c5e9),
	.w1(32'h3b99505f),
	.w2(32'h3a1e9e43),
	.w3(32'hba249c24),
	.w4(32'h3b268639),
	.w5(32'h3c11eaeb),
	.w6(32'hbb31062b),
	.w7(32'h3af1a7c5),
	.w8(32'h3c05045d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4066f3),
	.w1(32'h3b5b425f),
	.w2(32'h39dde293),
	.w3(32'hbb3a128f),
	.w4(32'h39fa96b1),
	.w5(32'h3b6e0a94),
	.w6(32'hbb24e56b),
	.w7(32'h3b78454d),
	.w8(32'h3ac8f1b6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c194),
	.w1(32'hbb6c1530),
	.w2(32'h3c6bf518),
	.w3(32'h3c0d7602),
	.w4(32'h3c9fb560),
	.w5(32'h3d11e3a5),
	.w6(32'h3bdd1b40),
	.w7(32'h3cfdf9c7),
	.w8(32'h3d305093),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd53ab0),
	.w1(32'h3cbd716c),
	.w2(32'h3c2ad187),
	.w3(32'h3bc1a239),
	.w4(32'h3c853562),
	.w5(32'h3c7253ef),
	.w6(32'h3c4c783a),
	.w7(32'h3c051fab),
	.w8(32'h3c8d5579),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f9ff9),
	.w1(32'h3bc419a8),
	.w2(32'h3a1cfa91),
	.w3(32'h3bf0204f),
	.w4(32'hbba0817b),
	.w5(32'hbb7cf032),
	.w6(32'h3c1be195),
	.w7(32'hbbea6b64),
	.w8(32'hbc1c575a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bd637),
	.w1(32'hbc584f12),
	.w2(32'hbb4e4a8f),
	.w3(32'h39f06665),
	.w4(32'hbc0e2300),
	.w5(32'hbb0aef87),
	.w6(32'hbc0cecaf),
	.w7(32'hbbae507b),
	.w8(32'hbb1fee90),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06190),
	.w1(32'hbb32e3d5),
	.w2(32'h3ae751f3),
	.w3(32'h3bcb07ee),
	.w4(32'h3af675a3),
	.w5(32'h38b80e7e),
	.w6(32'h3b1a4c92),
	.w7(32'h3c832b10),
	.w8(32'h3c4189df),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b273e),
	.w1(32'hba9309db),
	.w2(32'h3c6637ba),
	.w3(32'hbb29127b),
	.w4(32'h3be0cf85),
	.w5(32'h3c0a72db),
	.w6(32'h3c38db9c),
	.w7(32'h3b5e12c4),
	.w8(32'h3c6ed72b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c199605),
	.w1(32'h3c77cd92),
	.w2(32'hbbe01f73),
	.w3(32'h3c675753),
	.w4(32'hb9bc0f93),
	.w5(32'h3c0816b7),
	.w6(32'h3c67cbdd),
	.w7(32'hbb4bd6b3),
	.w8(32'hbb8f786c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0afca8),
	.w1(32'hbb60b459),
	.w2(32'hba1ddeb5),
	.w3(32'h3bc45865),
	.w4(32'hb949414a),
	.w5(32'hbb3d0a05),
	.w6(32'h3ab0b75f),
	.w7(32'hbbd2bcb6),
	.w8(32'hbbeb9aaf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6288b),
	.w1(32'hbbb0c18f),
	.w2(32'h39ff8543),
	.w3(32'hbb6b0f43),
	.w4(32'hbb528d9c),
	.w5(32'hbc0a6a3e),
	.w6(32'hbbf53f55),
	.w7(32'hbb2f9239),
	.w8(32'h3b8dadcb),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb61dc),
	.w1(32'h3c057997),
	.w2(32'hbaeedda4),
	.w3(32'hbb950935),
	.w4(32'hbbf9f937),
	.w5(32'h39e9f783),
	.w6(32'h3c2f8fc6),
	.w7(32'hbba6d03f),
	.w8(32'h3bed6899),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1492a0),
	.w1(32'hbb381cca),
	.w2(32'h3b609759),
	.w3(32'h3c17a2ea),
	.w4(32'h3b0cc576),
	.w5(32'h3b2259cf),
	.w6(32'h3ca71e47),
	.w7(32'h3bad6e18),
	.w8(32'h3b994896),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c533b91),
	.w1(32'h3c4d78d5),
	.w2(32'h3b59b27a),
	.w3(32'h3c05375b),
	.w4(32'h3c015913),
	.w5(32'h3c0297f5),
	.w6(32'h3c1cee75),
	.w7(32'h3bab38e1),
	.w8(32'hbb1a4ca9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e3f56),
	.w1(32'hbc267f37),
	.w2(32'h3b0a9439),
	.w3(32'h3938b130),
	.w4(32'h3b4bd33c),
	.w5(32'hba63061c),
	.w6(32'hbb9fbc5c),
	.w7(32'h3c7da535),
	.w8(32'h3c93d771),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc09bd1),
	.w1(32'h3bb54319),
	.w2(32'h3adfc3e9),
	.w3(32'hbc049f51),
	.w4(32'h3c046e42),
	.w5(32'h3c8ea7c6),
	.w6(32'hbb3e032b),
	.w7(32'h3b9531d2),
	.w8(32'h3c8d4c92),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50fb25),
	.w1(32'h3c4e5e1b),
	.w2(32'h3c30ad72),
	.w3(32'h3bd87e16),
	.w4(32'h3bed8f2b),
	.w5(32'h3b7526ef),
	.w6(32'h3b9f03db),
	.w7(32'h3bf3bfa9),
	.w8(32'h3b3ff582),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9deb1),
	.w1(32'h3b6cd2d0),
	.w2(32'h3b9380f5),
	.w3(32'h3b43b7c9),
	.w4(32'hbb1b2db9),
	.w5(32'hbbb4edcd),
	.w6(32'h3ab53f77),
	.w7(32'hbba2187a),
	.w8(32'hbc22339c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85cdb7),
	.w1(32'hbc202a71),
	.w2(32'hbaa2df5f),
	.w3(32'hbb672fe8),
	.w4(32'h3b9716c3),
	.w5(32'hbac96110),
	.w6(32'hbc8ae13e),
	.w7(32'h3cae6529),
	.w8(32'h3cb85651),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8626a7),
	.w1(32'h3c33a4d5),
	.w2(32'h3b8addbe),
	.w3(32'hbb1a7e05),
	.w4(32'hbba8e0a6),
	.w5(32'hbadaecf4),
	.w6(32'h3c67919c),
	.w7(32'h3b3bc328),
	.w8(32'h3b24b929),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdeff1),
	.w1(32'hbb21b60a),
	.w2(32'h3c073c84),
	.w3(32'hbb9f3fc2),
	.w4(32'h3b51f563),
	.w5(32'hbaea60bb),
	.w6(32'hbbb2c750),
	.w7(32'h3a723ce9),
	.w8(32'h3c31d9c1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065bd5),
	.w1(32'h3af07ca1),
	.w2(32'h3bfbc422),
	.w3(32'hbabf8d62),
	.w4(32'hbc618d88),
	.w5(32'hbc479e0c),
	.w6(32'hbb8dfec3),
	.w7(32'hbc0eae6e),
	.w8(32'hbc2c492c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f426a),
	.w1(32'h3adbf34e),
	.w2(32'h3b98ae7b),
	.w3(32'hbb811518),
	.w4(32'hba7b410b),
	.w5(32'h39b158d0),
	.w6(32'hbc25bab4),
	.w7(32'h3a8bbaeb),
	.w8(32'hbb962673),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd3f06),
	.w1(32'h3c0f4e1c),
	.w2(32'h3ca20bff),
	.w3(32'h3c3aa8f2),
	.w4(32'h3bfc89fb),
	.w5(32'h3cb24a18),
	.w6(32'hbab3a619),
	.w7(32'h3c28db14),
	.w8(32'h3958ba4d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beebcca),
	.w1(32'h3b6aeb7b),
	.w2(32'h3be17e17),
	.w3(32'h3c8f953e),
	.w4(32'h3c10652c),
	.w5(32'h3c8af439),
	.w6(32'h3c35e520),
	.w7(32'h3c267f78),
	.w8(32'h3cbe375b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26b3bc),
	.w1(32'h3beb0f10),
	.w2(32'hbbfc2a54),
	.w3(32'hb95a5552),
	.w4(32'h3a0b6756),
	.w5(32'h3ade1d45),
	.w6(32'h3accaaa1),
	.w7(32'hbb3bc725),
	.w8(32'hbb4816f0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52fe16),
	.w1(32'hbc489df5),
	.w2(32'hbb112eeb),
	.w3(32'h3bae44a3),
	.w4(32'h3b4cb5e1),
	.w5(32'h3ba27bc2),
	.w6(32'hbb52c55e),
	.w7(32'hbba777cd),
	.w8(32'h3c584cce),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf011),
	.w1(32'h3bbb3599),
	.w2(32'h3c79f637),
	.w3(32'hbb4b7bc3),
	.w4(32'hbae051ac),
	.w5(32'hb9d92ebe),
	.w6(32'h3bbf879a),
	.w7(32'h3c6f2ae0),
	.w8(32'hbbe3d7c4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404e89),
	.w1(32'hbc698edc),
	.w2(32'h3b1c7306),
	.w3(32'h3c6a3652),
	.w4(32'h3ae25cbd),
	.w5(32'h3bc18f95),
	.w6(32'h3b2bf271),
	.w7(32'h3a99d565),
	.w8(32'h39c4cb97),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2dc07),
	.w1(32'hbbc5537f),
	.w2(32'h3bc51030),
	.w3(32'h3bde4f78),
	.w4(32'h3beb69b4),
	.w5(32'hbb209dde),
	.w6(32'h3b9536ad),
	.w7(32'h3b70f5d6),
	.w8(32'hbb1138b5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16651),
	.w1(32'h3be682a6),
	.w2(32'hbb98c1ab),
	.w3(32'h3bcb61cb),
	.w4(32'hbc094808),
	.w5(32'hbbf472e5),
	.w6(32'h3baae5aa),
	.w7(32'hbc0da07a),
	.w8(32'hbc6eb9df),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76ecb4),
	.w1(32'hbc159b3a),
	.w2(32'hbb7e6c44),
	.w3(32'hbb8fdd34),
	.w4(32'hbb89b251),
	.w5(32'h3b67ebcb),
	.w6(32'h3aaf5f14),
	.w7(32'hbb632815),
	.w8(32'h3a796163),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb936fd8),
	.w1(32'hbb1152b0),
	.w2(32'h3bd88a97),
	.w3(32'h3bbeafe5),
	.w4(32'hbb5d6465),
	.w5(32'h3b160147),
	.w6(32'h3c03ef04),
	.w7(32'hba2cb22f),
	.w8(32'hbc8c9bd7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc0ee0),
	.w1(32'hbaefd885),
	.w2(32'hbade1535),
	.w3(32'h3be382e7),
	.w4(32'h3c703bbc),
	.w5(32'h3be32125),
	.w6(32'hbac41492),
	.w7(32'h3c0fd66f),
	.w8(32'h3c62e4e7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca69335),
	.w1(32'h3c6d8a7d),
	.w2(32'h3af911bc),
	.w3(32'h3b83d81b),
	.w4(32'hba41c85f),
	.w5(32'h3b8d61d4),
	.w6(32'hba831269),
	.w7(32'hbb2339f4),
	.w8(32'hbb2cbc1f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ef2f),
	.w1(32'h3badaa42),
	.w2(32'hbb600b68),
	.w3(32'h3c62290c),
	.w4(32'h3a88aaf5),
	.w5(32'h3b37d8ad),
	.w6(32'h3c3d7cd3),
	.w7(32'hbb07680a),
	.w8(32'hba502530),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948173),
	.w1(32'hbad693b2),
	.w2(32'h3a8003c4),
	.w3(32'h3c07be10),
	.w4(32'h3b108cf4),
	.w5(32'hba1f5df9),
	.w6(32'h3bcb80a2),
	.w7(32'hbacdcd60),
	.w8(32'h3b89e904),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cfe33),
	.w1(32'hbb172fc7),
	.w2(32'hbba8b430),
	.w3(32'h3c09c7c3),
	.w4(32'hba23bf57),
	.w5(32'h3a98000b),
	.w6(32'hbb806796),
	.w7(32'hbbe667fa),
	.w8(32'hbbe691cf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73ef0),
	.w1(32'h38b482ef),
	.w2(32'h39e05c2b),
	.w3(32'h3b9e5a3f),
	.w4(32'hbbf5e8ed),
	.w5(32'h3ae229cd),
	.w6(32'h3983f0bf),
	.w7(32'hbb845d2b),
	.w8(32'h3a0ef474),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be05eb9),
	.w1(32'h3a9a62e2),
	.w2(32'h3ba1b34e),
	.w3(32'hbc1389d3),
	.w4(32'h3a41c043),
	.w5(32'h3b94d3e2),
	.w6(32'hbbf70ec0),
	.w7(32'hbb898bdd),
	.w8(32'h3aae431b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7c90d),
	.w1(32'h3b726a77),
	.w2(32'hbb91198d),
	.w3(32'h3c081b34),
	.w4(32'h3ab4d7da),
	.w5(32'h3af468c3),
	.w6(32'h3b0c5be4),
	.w7(32'hbae2e86d),
	.w8(32'hbb221c59),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13e62e),
	.w1(32'hbbe2f45f),
	.w2(32'h3b7c7901),
	.w3(32'h3bbd0b15),
	.w4(32'h3af4f4d8),
	.w5(32'hbba8c009),
	.w6(32'hba0acae1),
	.w7(32'hbb18b4b3),
	.w8(32'hbc0abcee),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b9a3a),
	.w1(32'hbc58bdc3),
	.w2(32'hbb570195),
	.w3(32'hb9f95a58),
	.w4(32'hbab19750),
	.w5(32'h390082e1),
	.w6(32'hbc0ee002),
	.w7(32'hbaaf17be),
	.w8(32'hbbc7412b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacf0e9),
	.w1(32'hbbfb4dcf),
	.w2(32'hbb83c5d5),
	.w3(32'h3c658ec8),
	.w4(32'h3c867dfd),
	.w5(32'h3cbff652),
	.w6(32'hbb8760a8),
	.w7(32'h3c8fda05),
	.w8(32'h3d195326),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b62d5),
	.w1(32'h3c909bb5),
	.w2(32'hbc842f28),
	.w3(32'h3c382ba4),
	.w4(32'hbc877202),
	.w5(32'hbbfcad35),
	.w6(32'h3d060995),
	.w7(32'hbc870d1a),
	.w8(32'hbc1dbeb3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37907b),
	.w1(32'hbba75047),
	.w2(32'hbb2c32de),
	.w3(32'hbb12ca0a),
	.w4(32'h39ce3d16),
	.w5(32'hbbb624b6),
	.w6(32'hbc132df1),
	.w7(32'hbbdb1275),
	.w8(32'hbc05d4a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule