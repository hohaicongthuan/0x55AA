module layer_10_featuremap_288(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4812be),
	.w1(32'hbaa78e4b),
	.w2(32'hba82bd64),
	.w3(32'hba34edf9),
	.w4(32'hba6d30e1),
	.w5(32'h394a1e6e),
	.w6(32'hb7e6c4d0),
	.w7(32'hba42415f),
	.w8(32'hba5a44c4),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9662d54),
	.w1(32'h3991e252),
	.w2(32'h3a250672),
	.w3(32'h39730a4d),
	.w4(32'hb972ec49),
	.w5(32'h3a1001f1),
	.w6(32'hb926bfa1),
	.w7(32'hb9c5dcbd),
	.w8(32'h3998642d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5197ae),
	.w1(32'h3a08f52f),
	.w2(32'h39db3549),
	.w3(32'hb986c019),
	.w4(32'h390599cd),
	.w5(32'hb97c7412),
	.w6(32'h3abcf4dd),
	.w7(32'h3a428780),
	.w8(32'h3830081a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38737876),
	.w1(32'h39812dcb),
	.w2(32'hb842dbb0),
	.w3(32'hb9a2c936),
	.w4(32'hb7d0cc48),
	.w5(32'hba88d625),
	.w6(32'hb87830dc),
	.w7(32'hb9997ad1),
	.w8(32'hbaaa4c89),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdaf12),
	.w1(32'hba47f1d3),
	.w2(32'hb9cd1f56),
	.w3(32'hbad5ce89),
	.w4(32'hbab82ac5),
	.w5(32'hba0efbea),
	.w6(32'hba84f3c9),
	.w7(32'hba933e65),
	.w8(32'h3998ec65),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dcb8c9),
	.w1(32'hb70f6263),
	.w2(32'hb8bccbef),
	.w3(32'hb9ea909b),
	.w4(32'hb9832ec1),
	.w5(32'h387a95d5),
	.w6(32'h3941ef8d),
	.w7(32'hb8eda307),
	.w8(32'h38f47bb1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399966b5),
	.w1(32'h38c9e6e9),
	.w2(32'hb8c50994),
	.w3(32'hb99ad37e),
	.w4(32'hb98f6574),
	.w5(32'hb9b46bd8),
	.w6(32'h399891d5),
	.w7(32'h39008b94),
	.w8(32'hb948853a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc6726),
	.w1(32'hba0ca501),
	.w2(32'hb9675b2f),
	.w3(32'hb9d5c073),
	.w4(32'h39f0fa08),
	.w5(32'h3a343d3a),
	.w6(32'h3a7649bc),
	.w7(32'h39a9e537),
	.w8(32'h3a110588),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f6fc),
	.w1(32'h39cfc990),
	.w2(32'h37687bc9),
	.w3(32'h39412c08),
	.w4(32'h39d0b271),
	.w5(32'hb9c0294d),
	.w6(32'hb97c7ec9),
	.w7(32'h39051d8c),
	.w8(32'h39a8d48c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c1eb5),
	.w1(32'h390222a0),
	.w2(32'hb7af0cd3),
	.w3(32'hb976316f),
	.w4(32'hb9efbebd),
	.w5(32'hb9c47fe8),
	.w6(32'hb89313b9),
	.w7(32'hb9a69011),
	.w8(32'h3a0ffce9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39955e75),
	.w1(32'h39825b2d),
	.w2(32'h3963b890),
	.w3(32'hba07a7d2),
	.w4(32'h393c4a9e),
	.w5(32'h3a94cc5f),
	.w6(32'h3a28a1c9),
	.w7(32'h3a18ae46),
	.w8(32'hba222a3a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31b8d6),
	.w1(32'hba72b191),
	.w2(32'hba2fb661),
	.w3(32'h3a1db13e),
	.w4(32'hb80fb05f),
	.w5(32'hb99b9db8),
	.w6(32'h3a39825b),
	.w7(32'hba878131),
	.w8(32'hba5c7f76),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa4de0),
	.w1(32'hb8d46a4f),
	.w2(32'hb902187d),
	.w3(32'h3a9280d5),
	.w4(32'h3a90bfb6),
	.w5(32'hba9d38c3),
	.w6(32'hb95b0a4a),
	.w7(32'hba3d552b),
	.w8(32'hbaa7b652),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f58d),
	.w1(32'hba7e839c),
	.w2(32'hb90b58e9),
	.w3(32'hba70d6ed),
	.w4(32'h38b71b96),
	.w5(32'hb924c737),
	.w6(32'hbabd7991),
	.w7(32'hb9b1f277),
	.w8(32'hb97c8b65),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2e484),
	.w1(32'hb8f33d4c),
	.w2(32'hba3c95f6),
	.w3(32'hb8df056d),
	.w4(32'h39a91257),
	.w5(32'h39d11559),
	.w6(32'hba974652),
	.w7(32'hba6674f6),
	.w8(32'hb4c5d94f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afe477),
	.w1(32'hb9399db3),
	.w2(32'h39b86a79),
	.w3(32'hb9ad8da0),
	.w4(32'hb90e8905),
	.w5(32'h39a3fd0b),
	.w6(32'hba031a04),
	.w7(32'hb90e5267),
	.w8(32'hb96bd461),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902c40d),
	.w1(32'h3a0dbee9),
	.w2(32'h39240972),
	.w3(32'hb8070fba),
	.w4(32'h39b2ed1c),
	.w5(32'h39dd3a0d),
	.w6(32'h393dee1b),
	.w7(32'hb9008d39),
	.w8(32'h396511dc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907d0fd),
	.w1(32'hba87a336),
	.w2(32'hb93baf01),
	.w3(32'hb74d8165),
	.w4(32'hba1e4e79),
	.w5(32'hba8a5ea8),
	.w6(32'hb7f99790),
	.w7(32'hb9a975fb),
	.w8(32'h397161a3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885762a),
	.w1(32'hba922518),
	.w2(32'hba727d18),
	.w3(32'hba8ba422),
	.w4(32'hba7937ad),
	.w5(32'hba47144e),
	.w6(32'h3a0b5178),
	.w7(32'hb761822b),
	.w8(32'hba40475c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bbc57),
	.w1(32'h37684689),
	.w2(32'hb93d060d),
	.w3(32'h399cd805),
	.w4(32'h39fb1b5e),
	.w5(32'h394aad84),
	.w6(32'hb9df54fe),
	.w7(32'hb9411d84),
	.w8(32'hb886dbec),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ddb25),
	.w1(32'hb9989851),
	.w2(32'h38cbb3d2),
	.w3(32'hb9bfbdeb),
	.w4(32'hb99f222a),
	.w5(32'hb9434dd5),
	.w6(32'hb98f79e2),
	.w7(32'hb8378149),
	.w8(32'hb83b4806),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d7ba1),
	.w1(32'hb867c76e),
	.w2(32'h38d14478),
	.w3(32'hb9e5b99f),
	.w4(32'h396ff0a2),
	.w5(32'h3a3e5f11),
	.w6(32'hb985c68a),
	.w7(32'h39b45f28),
	.w8(32'h39c98a1d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dd8db),
	.w1(32'hb9544f41),
	.w2(32'h3a07a331),
	.w3(32'hb8ffadd8),
	.w4(32'hba5c39a3),
	.w5(32'hba4aa8e4),
	.w6(32'h3a4e7300),
	.w7(32'hb9352c20),
	.w8(32'hbaccf9e0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba031a20),
	.w1(32'h37945bb3),
	.w2(32'hb6e66bbc),
	.w3(32'hb9e53b13),
	.w4(32'h3a291c55),
	.w5(32'h3a202d43),
	.w6(32'h39930217),
	.w7(32'h391d45bf),
	.w8(32'hba563273),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe636f),
	.w1(32'hb99f8739),
	.w2(32'h38b35c68),
	.w3(32'h391a185b),
	.w4(32'h3a2c5574),
	.w5(32'hb86f774c),
	.w6(32'h3abe63d3),
	.w7(32'h3984ae0f),
	.w8(32'hb9d25a64),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cff79c),
	.w1(32'h385041a2),
	.w2(32'hb979136d),
	.w3(32'h37c3917c),
	.w4(32'h38f001f7),
	.w5(32'hb9ad0c6e),
	.w6(32'hb94aa08d),
	.w7(32'h390b72f2),
	.w8(32'hb909325d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e65338),
	.w1(32'hb9de4bfb),
	.w2(32'hba0befb3),
	.w3(32'hba983d29),
	.w4(32'hba449b50),
	.w5(32'hb9e813da),
	.w6(32'hba0abf20),
	.w7(32'hba1a3ace),
	.w8(32'hb952e72e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d076a8),
	.w1(32'hba2a9251),
	.w2(32'hba85fb3e),
	.w3(32'hb9d9128c),
	.w4(32'hba6257d4),
	.w5(32'hba489025),
	.w6(32'hb9f1203e),
	.w7(32'hba19b3e5),
	.w8(32'hba1d82be),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b95604),
	.w1(32'hba18f50e),
	.w2(32'h3606815d),
	.w3(32'hb90c3267),
	.w4(32'h39380485),
	.w5(32'h37b29d84),
	.w6(32'hb9cd5faf),
	.w7(32'h3a0caee2),
	.w8(32'h39e4528f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f725d),
	.w1(32'h39a21bd6),
	.w2(32'h3a1d2d87),
	.w3(32'h388b88f5),
	.w4(32'h3989246d),
	.w5(32'h395685d5),
	.w6(32'hb9a47fb8),
	.w7(32'h38863f64),
	.w8(32'h3a729e1b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8a07b),
	.w1(32'h3aaeb91a),
	.w2(32'h39dd1b41),
	.w3(32'h39f47709),
	.w4(32'hba598177),
	.w5(32'h3a4e8e68),
	.w6(32'h3b3ecee1),
	.w7(32'h39949bbf),
	.w8(32'h395d888e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902d094),
	.w1(32'h39ba446b),
	.w2(32'h3887e5d7),
	.w3(32'h3ac73544),
	.w4(32'h3a9e1d3b),
	.w5(32'hb9839141),
	.w6(32'h3a5670b6),
	.w7(32'hba70550a),
	.w8(32'h3a968d03),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d52434),
	.w1(32'h38d5b43f),
	.w2(32'hbaa31acf),
	.w3(32'h3a03b8ea),
	.w4(32'hba2da2e1),
	.w5(32'hb9adfc50),
	.w6(32'h3ad97d74),
	.w7(32'hb7efe197),
	.w8(32'hb8be5fee),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a079bc),
	.w1(32'h39807b28),
	.w2(32'h3a33bf64),
	.w3(32'h39e84ec6),
	.w4(32'h39d536d6),
	.w5(32'h3a7fe1ac),
	.w6(32'h393b401b),
	.w7(32'h36868ba0),
	.w8(32'h39b9f14d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7501fc8),
	.w1(32'h351316c4),
	.w2(32'h39b38937),
	.w3(32'h3a0cc478),
	.w4(32'h3a0a07cc),
	.w5(32'hba979985),
	.w6(32'h39dadb3a),
	.w7(32'h3a1eebb4),
	.w8(32'hb9ed9797),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d989be),
	.w1(32'h393ab46e),
	.w2(32'h3909770f),
	.w3(32'hba32c9be),
	.w4(32'hb8ff92a1),
	.w5(32'hba66314b),
	.w6(32'h3a850bed),
	.w7(32'h3a972796),
	.w8(32'h3aa0ace3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954d0d8),
	.w1(32'h3a259194),
	.w2(32'hba65aca3),
	.w3(32'hb88758ca),
	.w4(32'hba8a266a),
	.w5(32'hba0d9ded),
	.w6(32'h3ad0eba9),
	.w7(32'h399fd8f3),
	.w8(32'h3904ce29),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dcf3e2),
	.w1(32'hb9e011f7),
	.w2(32'hba08e64b),
	.w3(32'hb9bac822),
	.w4(32'h39902dea),
	.w5(32'hbb0263e6),
	.w6(32'hb9b0fa7d),
	.w7(32'h3a524de2),
	.w8(32'hb838b923),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39350186),
	.w1(32'hb7e22335),
	.w2(32'hba1d8169),
	.w3(32'hbaa4e2db),
	.w4(32'hba94eb48),
	.w5(32'hb9f6225f),
	.w6(32'h3853cdb7),
	.w7(32'hb9eb7f2f),
	.w8(32'hb92efebc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a85400),
	.w1(32'hb899da6f),
	.w2(32'h39c97c2d),
	.w3(32'h3a26fc62),
	.w4(32'hb9d9951a),
	.w5(32'h39ae13a6),
	.w6(32'h388bc685),
	.w7(32'h3a7c3b6f),
	.w8(32'hb906a4c7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b7224),
	.w1(32'hba85a03b),
	.w2(32'h39bb8586),
	.w3(32'hb9a88e40),
	.w4(32'h39225e4c),
	.w5(32'hb919b957),
	.w6(32'hba852efd),
	.w7(32'hb9a00924),
	.w8(32'h390eca1c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a49ec9),
	.w1(32'hb91a979f),
	.w2(32'h3737cd5f),
	.w3(32'hba2f6ffd),
	.w4(32'hb9d1e2ed),
	.w5(32'h3a89d384),
	.w6(32'hb995efd9),
	.w7(32'h381356ff),
	.w8(32'h3a656704),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba540f),
	.w1(32'hba6bff2b),
	.w2(32'h388dd36e),
	.w3(32'hb948196a),
	.w4(32'h397d3c28),
	.w5(32'hba637968),
	.w6(32'hb9ca1e43),
	.w7(32'h3a5d941d),
	.w8(32'hbb0a2d31),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dd2c7),
	.w1(32'h389fc241),
	.w2(32'hba133f91),
	.w3(32'hbb0ae2e7),
	.w4(32'hb93f969a),
	.w5(32'h38d0b72e),
	.w6(32'hbac6157f),
	.w7(32'hb9a4a6d6),
	.w8(32'h3ab515c0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37312c89),
	.w1(32'hb87dc59f),
	.w2(32'hb9a90b58),
	.w3(32'h3a33424c),
	.w4(32'h37a065f5),
	.w5(32'hbaa391d6),
	.w6(32'h3a170fe3),
	.w7(32'h3951bbd6),
	.w8(32'hba68d221),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52f82c),
	.w1(32'hb83b382f),
	.w2(32'h38f85a09),
	.w3(32'hba799683),
	.w4(32'hba76904b),
	.w5(32'hbaab56b1),
	.w6(32'h38f6247a),
	.w7(32'h3988fe9c),
	.w8(32'hba53f274),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba071877),
	.w1(32'h39835204),
	.w2(32'hb863e76e),
	.w3(32'hba0a37f1),
	.w4(32'hba53c10d),
	.w5(32'h3a8f7dfd),
	.w6(32'hb95fc180),
	.w7(32'hba3327e9),
	.w8(32'h3a04581d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff271),
	.w1(32'hbaacf925),
	.w2(32'hba2bd5a4),
	.w3(32'h3a17e363),
	.w4(32'h39d59b9c),
	.w5(32'hb9e00cff),
	.w6(32'h39175497),
	.w7(32'h3985127e),
	.w8(32'h39ac9b31),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5826ff),
	.w1(32'hb8849644),
	.w2(32'h36a154d5),
	.w3(32'h39bcfe9a),
	.w4(32'h3a5f9cb5),
	.w5(32'h397d7849),
	.w6(32'h39e0732c),
	.w7(32'h394be0a3),
	.w8(32'h3a4235a9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0d670),
	.w1(32'h39655175),
	.w2(32'h39b2f735),
	.w3(32'hb9e5e8de),
	.w4(32'h369176be),
	.w5(32'hb98fa573),
	.w6(32'hba091879),
	.w7(32'hb925c792),
	.w8(32'hba5f5193),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28c90),
	.w1(32'h39f86566),
	.w2(32'hb8b88677),
	.w3(32'hba176f6e),
	.w4(32'h37a74d89),
	.w5(32'hb8ce68dd),
	.w6(32'h39f78e73),
	.w7(32'hb84dd5aa),
	.w8(32'hba515872),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07ae3c),
	.w1(32'hb9bbebb2),
	.w2(32'hb86ee92d),
	.w3(32'hba65750d),
	.w4(32'hba2bfcce),
	.w5(32'h3a2e6c72),
	.w6(32'hba1f4673),
	.w7(32'hb9f2c242),
	.w8(32'h3a0a5042),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab913df),
	.w1(32'hba7ffa4d),
	.w2(32'hb92ea4e9),
	.w3(32'h387f90a9),
	.w4(32'h39bd83b7),
	.w5(32'hba9e8a2a),
	.w6(32'h39ced509),
	.w7(32'hb881927b),
	.w8(32'hba0e36d0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac005f1),
	.w1(32'hbb14604a),
	.w2(32'hba1f72c5),
	.w3(32'hb931b92e),
	.w4(32'hbacf5701),
	.w5(32'hba58f391),
	.w6(32'h390c9465),
	.w7(32'hba292c06),
	.w8(32'hb9f2d5a3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98988fc),
	.w1(32'hb9cf3a25),
	.w2(32'hb97f6ebf),
	.w3(32'hb9125638),
	.w4(32'hb960cf86),
	.w5(32'hb80af81d),
	.w6(32'hb9b21c76),
	.w7(32'hb9f8441d),
	.w8(32'hb9956ef8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd2752),
	.w1(32'h38f40f4f),
	.w2(32'h3a1e92e5),
	.w3(32'hb9fb0a35),
	.w4(32'h39c154c2),
	.w5(32'h397f8b38),
	.w6(32'hb957b97a),
	.w7(32'h39edf4dd),
	.w8(32'hb9eecee2),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a74ceb),
	.w1(32'hba34c108),
	.w2(32'hb787d2e6),
	.w3(32'hb8dc9039),
	.w4(32'h3a06fab6),
	.w5(32'h39d28464),
	.w6(32'hba537887),
	.w7(32'h38b13ca0),
	.w8(32'h3a078b5d),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f7766),
	.w1(32'h34c31d4f),
	.w2(32'h3a25abbe),
	.w3(32'h3a53f7eb),
	.w4(32'h3a6c7149),
	.w5(32'h3a1b86a9),
	.w6(32'h3a12dd9f),
	.w7(32'h3abc0c1c),
	.w8(32'h3a44a8c2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1739fa),
	.w1(32'h39639eb8),
	.w2(32'h387ea306),
	.w3(32'h395fb59e),
	.w4(32'h3a037731),
	.w5(32'hb9bc96eb),
	.w6(32'h3912cf5c),
	.w7(32'h39dda499),
	.w8(32'h399c4549),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996d7d4),
	.w1(32'hb9cc502a),
	.w2(32'hba79b591),
	.w3(32'hb9896b74),
	.w4(32'hba02edc2),
	.w5(32'hba81a42d),
	.w6(32'h3a9b4bf1),
	.w7(32'h3988f89f),
	.w8(32'hb8c01a60),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea4477),
	.w1(32'hba31a851),
	.w2(32'hbab80482),
	.w3(32'hbab35e2d),
	.w4(32'hbab4304b),
	.w5(32'hba802e56),
	.w6(32'hba474d58),
	.w7(32'hba61a566),
	.w8(32'hba70022f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32159f),
	.w1(32'hb88c2544),
	.w2(32'hb996ce42),
	.w3(32'hb9f152c6),
	.w4(32'hb9ebd0f0),
	.w5(32'h39b4d07d),
	.w6(32'h38971b54),
	.w7(32'hb9a99b8b),
	.w8(32'h39e8ba7c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9765d9f),
	.w1(32'hba17018e),
	.w2(32'hb99949da),
	.w3(32'hba09ebb4),
	.w4(32'hba9213d4),
	.w5(32'h38c86f84),
	.w6(32'h39a33b44),
	.w7(32'hba0da654),
	.w8(32'hb9035de7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385be368),
	.w1(32'hb91ab91e),
	.w2(32'h3a20375a),
	.w3(32'h38280381),
	.w4(32'h398d914b),
	.w5(32'hb9b90f80),
	.w6(32'hb84739da),
	.w7(32'h39d8c418),
	.w8(32'h38b4c06c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b3e4a),
	.w1(32'hb8f80d95),
	.w2(32'hb96b94bc),
	.w3(32'hba12229b),
	.w4(32'hba19dc7e),
	.w5(32'hb8b5512b),
	.w6(32'hb99616e0),
	.w7(32'hb84dc8ac),
	.w8(32'hb98ef100),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a6348),
	.w1(32'hb920fa68),
	.w2(32'h391655ef),
	.w3(32'hb9169373),
	.w4(32'hba7b9cd4),
	.w5(32'hb9bad0c2),
	.w6(32'h3a2e4b6f),
	.w7(32'hba5a1f7e),
	.w8(32'h395f6337),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942bd26),
	.w1(32'hba4d08ec),
	.w2(32'h390e7437),
	.w3(32'hba099aed),
	.w4(32'hb999c5ec),
	.w5(32'h3991e450),
	.w6(32'h39c01704),
	.w7(32'hb99527e3),
	.w8(32'h3a2b6acd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b5ea4),
	.w1(32'h39e7a571),
	.w2(32'h392197d5),
	.w3(32'h3abc6829),
	.w4(32'h3a8d0f6d),
	.w5(32'hb9ff5e1a),
	.w6(32'h396120f3),
	.w7(32'h3998f28c),
	.w8(32'hb7a7f101),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95c0971),
	.w1(32'hba81f7cc),
	.w2(32'hbab4686d),
	.w3(32'hba3314d4),
	.w4(32'hba56658c),
	.w5(32'h38f35c0a),
	.w6(32'hb9fede95),
	.w7(32'hba273047),
	.w8(32'h389ec43e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a759),
	.w1(32'h3abe1f94),
	.w2(32'h3aa34eb8),
	.w3(32'hb9e37181),
	.w4(32'h3ae4655a),
	.w5(32'h39c7eeb6),
	.w6(32'hba3fa1f2),
	.w7(32'h3a7ee96a),
	.w8(32'h3a1c561d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7fb4),
	.w1(32'hb9bdf2ae),
	.w2(32'h3978ce3b),
	.w3(32'hb95d2156),
	.w4(32'hb56e28b8),
	.w5(32'h3990e312),
	.w6(32'h3978e6de),
	.w7(32'h39b23f7b),
	.w8(32'hba2315ed),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1cfcb),
	.w1(32'hb9f657a0),
	.w2(32'h3a04b4b9),
	.w3(32'h383947b1),
	.w4(32'hb79afdb6),
	.w5(32'h3a1b31b3),
	.w6(32'hb9617dc2),
	.w7(32'h39432eec),
	.w8(32'hba88ef0f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388db39e),
	.w1(32'h3a44f33c),
	.w2(32'h3a228b8b),
	.w3(32'h39cd79ed),
	.w4(32'hb90d5d72),
	.w5(32'hb98128c0),
	.w6(32'hb9b70d9e),
	.w7(32'hba9744b6),
	.w8(32'h38dc3ff4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396df869),
	.w1(32'hb9aec020),
	.w2(32'h3a2a6830),
	.w3(32'h3934b20e),
	.w4(32'hb9453f1f),
	.w5(32'h38ca95f3),
	.w6(32'h394d9eca),
	.w7(32'h387d464b),
	.w8(32'h39e64713),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b7453),
	.w1(32'hb9d29712),
	.w2(32'h39958d86),
	.w3(32'h399162e9),
	.w4(32'h3a18d8ba),
	.w5(32'h39ef44e6),
	.w6(32'h3a0f6b71),
	.w7(32'h38e02cc2),
	.w8(32'hb8684dc8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba340d03),
	.w1(32'hba3cfdaa),
	.w2(32'hb8129dcd),
	.w3(32'h3a29288b),
	.w4(32'h39be9af1),
	.w5(32'hb9e1799f),
	.w6(32'h39c7094d),
	.w7(32'h390f8a84),
	.w8(32'hba0ed055),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c75a3),
	.w1(32'hb88b790b),
	.w2(32'h39df01d0),
	.w3(32'hba6ad9c5),
	.w4(32'hb9004c70),
	.w5(32'hb8b7100b),
	.w6(32'h3a3e838e),
	.w7(32'h38fb2dc8),
	.w8(32'h379d02ae),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b7405),
	.w1(32'h3a397145),
	.w2(32'h39bfb668),
	.w3(32'h3a2787d6),
	.w4(32'h3a466344),
	.w5(32'hb98dce5b),
	.w6(32'h3a0b2316),
	.w7(32'h398336e3),
	.w8(32'h38f87732),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e17168),
	.w1(32'h39b2a75b),
	.w2(32'h390515c4),
	.w3(32'h3a2fccc4),
	.w4(32'h38ac7b2d),
	.w5(32'hb99c0566),
	.w6(32'h3a86c8f7),
	.w7(32'hb7a2e25a),
	.w8(32'hb97c1b07),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994ad60),
	.w1(32'h3863ca60),
	.w2(32'h38f3001f),
	.w3(32'h3898e86d),
	.w4(32'h38ebdb5a),
	.w5(32'h3a64c867),
	.w6(32'hb84bfcaa),
	.w7(32'hb9acf439),
	.w8(32'h3a2f712b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9747a),
	.w1(32'hba0ff750),
	.w2(32'h3a10e8b0),
	.w3(32'h3a81ad31),
	.w4(32'h3a902748),
	.w5(32'hb89ad6e5),
	.w6(32'hb8c96126),
	.w7(32'h3a09b10f),
	.w8(32'h39ce54bd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8e866),
	.w1(32'hb9c6c1e8),
	.w2(32'h36ac10e2),
	.w3(32'h37953091),
	.w4(32'h39337fb4),
	.w5(32'h3a43b180),
	.w6(32'h3a692392),
	.w7(32'h3a54c3d4),
	.w8(32'h38786096),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d20c24),
	.w1(32'h39f45a83),
	.w2(32'h3909ac14),
	.w3(32'h3935a8fe),
	.w4(32'h3a4d463f),
	.w5(32'hba8edc29),
	.w6(32'h3a3ccc2d),
	.w7(32'h3a49f38a),
	.w8(32'hb994fb76),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc13aa),
	.w1(32'hb9d53f28),
	.w2(32'hba9e459d),
	.w3(32'hb93cfa0a),
	.w4(32'hb9f0f5cc),
	.w5(32'h3a6b42f5),
	.w6(32'hb9db6cc3),
	.w7(32'hba2b55d4),
	.w8(32'h3a44aa66),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8b842),
	.w1(32'h3a6a9d81),
	.w2(32'h39bbe5e7),
	.w3(32'h3a21931e),
	.w4(32'h3aab0965),
	.w5(32'hbad3ba75),
	.w6(32'h3ab38082),
	.w7(32'h3a9b5a68),
	.w8(32'hba18c9bc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e8cf76),
	.w1(32'hba36c1cc),
	.w2(32'hb9d08e6a),
	.w3(32'hba7f59b5),
	.w4(32'hba4eb154),
	.w5(32'h3a01aaf2),
	.w6(32'h39d5c11e),
	.w7(32'hb9d8bdb3),
	.w8(32'h3a143f76),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c3d13),
	.w1(32'h39a86286),
	.w2(32'h3a169175),
	.w3(32'hb841d012),
	.w4(32'h39b99fab),
	.w5(32'hb9ccd939),
	.w6(32'h372ad527),
	.w7(32'h3a72f4c6),
	.w8(32'hb9e47ec9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aae073),
	.w1(32'h36dd83a4),
	.w2(32'hb9210318),
	.w3(32'h37823efc),
	.w4(32'hb9450c0e),
	.w5(32'hb99e1a07),
	.w6(32'h3992728d),
	.w7(32'hb95547cc),
	.w8(32'hb9c4fb16),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7df39),
	.w1(32'h392cfb62),
	.w2(32'hb9687f94),
	.w3(32'hb99d5e52),
	.w4(32'hb8705c81),
	.w5(32'h38d38796),
	.w6(32'hb9f34942),
	.w7(32'hb95794e0),
	.w8(32'h3a3868cf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370b83b7),
	.w1(32'h39c2406c),
	.w2(32'h39d6ad18),
	.w3(32'h39e606f6),
	.w4(32'h37bd0457),
	.w5(32'hb9e7f6ce),
	.w6(32'h3a843620),
	.w7(32'h3a5eba8a),
	.w8(32'hb810d08c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a6eb9),
	.w1(32'h39122f50),
	.w2(32'hba084e8d),
	.w3(32'hba0ee8f8),
	.w4(32'hb7852e3e),
	.w5(32'h3a1e0572),
	.w6(32'hb9670d61),
	.w7(32'hb9b7b878),
	.w8(32'h3a33ec0d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f06d05),
	.w1(32'h38de7091),
	.w2(32'hbad14890),
	.w3(32'h3a07c221),
	.w4(32'hba1e6f0a),
	.w5(32'hbab8d10a),
	.w6(32'h382891a3),
	.w7(32'hb9dcb5e9),
	.w8(32'hba9dfcb4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba3aa8),
	.w1(32'h39b1e048),
	.w2(32'hba00494f),
	.w3(32'hba85100c),
	.w4(32'h398e7726),
	.w5(32'hba6f59fa),
	.w6(32'hb93b31fc),
	.w7(32'hb99039ba),
	.w8(32'hb9b3fe76),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c9b8f),
	.w1(32'h39a5284b),
	.w2(32'hb9faab40),
	.w3(32'hba4b92a9),
	.w4(32'hbb02bcc5),
	.w5(32'h3a15a822),
	.w6(32'hba0198e8),
	.w7(32'hba415d58),
	.w8(32'h3a21ee66),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4beb1),
	.w1(32'h38aac592),
	.w2(32'h39b7684b),
	.w3(32'h3808c1cc),
	.w4(32'hba3d7ed7),
	.w5(32'h3adea2f6),
	.w6(32'hb9c08aeb),
	.w7(32'hb903ba17),
	.w8(32'h398e3de5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e67ef),
	.w1(32'h3a442b48),
	.w2(32'h3a8142fd),
	.w3(32'h3a7fc9cb),
	.w4(32'h39da6679),
	.w5(32'hba267e07),
	.w6(32'hba1d6f90),
	.w7(32'h39839408),
	.w8(32'h3989a739),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974d9db),
	.w1(32'h38d97f93),
	.w2(32'h37f34722),
	.w3(32'h384814fa),
	.w4(32'hba638dc6),
	.w5(32'h38ee16df),
	.w6(32'h3a47f9c6),
	.w7(32'h39d2cd05),
	.w8(32'hb979684f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b19f),
	.w1(32'hba16bca2),
	.w2(32'hb94ec0c6),
	.w3(32'hb83478d3),
	.w4(32'hba0d2a92),
	.w5(32'hb709e96c),
	.w6(32'hb9760fd0),
	.w7(32'hba4847ff),
	.w8(32'hb803b806),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920215d),
	.w1(32'hb9abe3ad),
	.w2(32'h3701cf6a),
	.w3(32'h38edf33c),
	.w4(32'hb9369ce0),
	.w5(32'hb8f03184),
	.w6(32'hb6a3230c),
	.w7(32'hba177cea),
	.w8(32'hb993e790),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51c706),
	.w1(32'hb8a56487),
	.w2(32'hba3651a1),
	.w3(32'hba6e59dd),
	.w4(32'hb98d09d7),
	.w5(32'hba47c2ed),
	.w6(32'hb90e19c4),
	.w7(32'h39c5382b),
	.w8(32'hb9ea86b5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93e66a7),
	.w1(32'h3a1e585d),
	.w2(32'hb94c870a),
	.w3(32'h3a069a8e),
	.w4(32'h3a8c9fe4),
	.w5(32'hb7e95239),
	.w6(32'hba8fbfc9),
	.w7(32'hb8b94328),
	.w8(32'hb908147a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16dbda),
	.w1(32'h393442ac),
	.w2(32'h3a266941),
	.w3(32'h3a1bc3fd),
	.w4(32'h394ec7d2),
	.w5(32'h3a1ad38b),
	.w6(32'hb9b0cf3d),
	.w7(32'hb88de60c),
	.w8(32'hb81604e7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a621c),
	.w1(32'hb8f4120e),
	.w2(32'hba4feddc),
	.w3(32'hb9dc7df8),
	.w4(32'hb96b8e7a),
	.w5(32'hb9f512aa),
	.w6(32'h396a2352),
	.w7(32'hb9ca789b),
	.w8(32'hb9da5898),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a323c5),
	.w1(32'h394375f7),
	.w2(32'hb952fb9e),
	.w3(32'h399d4881),
	.w4(32'h38722aba),
	.w5(32'hb818b964),
	.w6(32'h38dc715e),
	.w7(32'hb8fefca5),
	.w8(32'hb82dcad1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0eb3f),
	.w1(32'h38f2dcec),
	.w2(32'hb96c8a89),
	.w3(32'hba00b229),
	.w4(32'hba1a9bf6),
	.w5(32'hbab0007a),
	.w6(32'h3a7fb67d),
	.w7(32'hb996e54b),
	.w8(32'hbb05380e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1194f),
	.w1(32'h395dc1bf),
	.w2(32'hb83d5221),
	.w3(32'h39eb4cd5),
	.w4(32'h39a094b6),
	.w5(32'hb8834615),
	.w6(32'h381e4347),
	.w7(32'h3987f1ac),
	.w8(32'hb90b62e0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbba75),
	.w1(32'h36115c35),
	.w2(32'hb898a4be),
	.w3(32'h3852945d),
	.w4(32'hb7eac0e9),
	.w5(32'hb7686378),
	.w6(32'h38384f1e),
	.w7(32'hb7f4f706),
	.w8(32'h37e6fb9c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380b4b83),
	.w1(32'h38ad14c8),
	.w2(32'h390e4eb4),
	.w3(32'h38e5b720),
	.w4(32'h39a6003c),
	.w5(32'h39864585),
	.w6(32'hb80c3b42),
	.w7(32'h39793ddd),
	.w8(32'h3906868c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1ddf5),
	.w1(32'hb93a7033),
	.w2(32'hb9932127),
	.w3(32'h3910fe82),
	.w4(32'hb9c492ea),
	.w5(32'hb8c4b036),
	.w6(32'hb953bf0a),
	.w7(32'hb9c5fd65),
	.w8(32'hb882b12d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9b824),
	.w1(32'h3956081f),
	.w2(32'h39ca187d),
	.w3(32'hb91bfbf7),
	.w4(32'h394be910),
	.w5(32'h39b36d25),
	.w6(32'hba11b82b),
	.w7(32'hb8b14f5b),
	.w8(32'h3708c459),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901f314),
	.w1(32'h39eb31ae),
	.w2(32'h39ea14a4),
	.w3(32'hb8a3006f),
	.w4(32'hb80f65d1),
	.w5(32'h394040a7),
	.w6(32'hb9b70fd0),
	.w7(32'h39442c84),
	.w8(32'h39a21493),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95185db),
	.w1(32'h396d5862),
	.w2(32'h39cd5be5),
	.w3(32'hb998a24f),
	.w4(32'hb9ac62a7),
	.w5(32'hb72145db),
	.w6(32'hb9a4030b),
	.w7(32'hb998f55c),
	.w8(32'hb7942054),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957be27),
	.w1(32'hb8bede28),
	.w2(32'hb9b86336),
	.w3(32'hb91b97fa),
	.w4(32'hb8a11974),
	.w5(32'hb9d3482b),
	.w6(32'h39083a91),
	.w7(32'hb89556b8),
	.w8(32'hb94ed7f0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a74c5d),
	.w1(32'h3991f003),
	.w2(32'h39923957),
	.w3(32'h386f0b25),
	.w4(32'hb90d58f4),
	.w5(32'hb7eb2108),
	.w6(32'hb97aadfc),
	.w7(32'h38f2aa1a),
	.w8(32'h38ab6bd8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39169261),
	.w1(32'hb8caa40f),
	.w2(32'h38e6957b),
	.w3(32'h37a41be4),
	.w4(32'h388d7e88),
	.w5(32'h36f0576a),
	.w6(32'h381d1489),
	.w7(32'h38798c0c),
	.w8(32'h3805507e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3693365f),
	.w1(32'hb7b3bf34),
	.w2(32'h36908d85),
	.w3(32'hb65b58d6),
	.w4(32'hb58990e3),
	.w5(32'hb781b2c7),
	.w6(32'hb722792a),
	.w7(32'hb77cb20f),
	.w8(32'hb7c66073),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f10d10),
	.w1(32'hb6d41b6c),
	.w2(32'hb615317c),
	.w3(32'hb786f160),
	.w4(32'hb782e372),
	.w5(32'h378862d8),
	.w6(32'hb77b54a7),
	.w7(32'hb70055d7),
	.w8(32'hb7dacb4b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372757d6),
	.w1(32'h385e5ee6),
	.w2(32'h3679b779),
	.w3(32'h3803b611),
	.w4(32'hb63a11c0),
	.w5(32'h3929ed4f),
	.w6(32'hb6b5a5f2),
	.w7(32'hb832b672),
	.w8(32'h38b3f152),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39846066),
	.w1(32'h391e6868),
	.w2(32'h39b0f7ed),
	.w3(32'h3924efb4),
	.w4(32'h39b56675),
	.w5(32'h39ae94c5),
	.w6(32'hb6c41b2e),
	.w7(32'h38e91c31),
	.w8(32'h39405bcb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c8704),
	.w1(32'h39c6488a),
	.w2(32'h39756439),
	.w3(32'h3989d0b4),
	.w4(32'h385ae310),
	.w5(32'h3928f0dc),
	.w6(32'hb99edfc4),
	.w7(32'hb9931d20),
	.w8(32'h37d45ab8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9332106),
	.w1(32'hb7fe3ce3),
	.w2(32'hb8411668),
	.w3(32'hb8fe8fd0),
	.w4(32'hb829380d),
	.w5(32'hb860cbd5),
	.w6(32'hb893bc93),
	.w7(32'hb914d79f),
	.w8(32'hb7e7729f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a0dcd),
	.w1(32'hb9e01168),
	.w2(32'hb9a38bcd),
	.w3(32'hb7dc2f1c),
	.w4(32'hba0e554c),
	.w5(32'hb9f4fbbe),
	.w6(32'h394440b7),
	.w7(32'hb9502444),
	.w8(32'hb93ec679),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e2fc8),
	.w1(32'h391f01f7),
	.w2(32'h384c6622),
	.w3(32'hb765109f),
	.w4(32'h38ff1309),
	.w5(32'hb8da12f8),
	.w6(32'hb9599944),
	.w7(32'h37f0c62e),
	.w8(32'hb8aa5529),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb795f6a6),
	.w1(32'h373f7fe8),
	.w2(32'h372d5aff),
	.w3(32'h370a8ed4),
	.w4(32'h374090b2),
	.w5(32'h37b256bf),
	.w6(32'h364bef3a),
	.w7(32'hb6459cf8),
	.w8(32'h3731983f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86e7163),
	.w1(32'hb80309ee),
	.w2(32'hb8474d39),
	.w3(32'hb7b084d8),
	.w4(32'hb7eec256),
	.w5(32'hb788ed09),
	.w6(32'hb537e887),
	.w7(32'hb6a0e693),
	.w8(32'hb8010b47),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3651c2ad),
	.w1(32'h3743a908),
	.w2(32'hb793fbfe),
	.w3(32'h37aace7c),
	.w4(32'h37ad165d),
	.w5(32'hb6cbf52b),
	.w6(32'hb73cc5d2),
	.w7(32'hb7f715a3),
	.w8(32'hb797d427),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bc145a),
	.w1(32'hb63667f1),
	.w2(32'hb70f1ca1),
	.w3(32'h37acc341),
	.w4(32'hb8546d44),
	.w5(32'hb8563c97),
	.w6(32'hb70cd8af),
	.w7(32'hb83202cd),
	.w8(32'hb81727ac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3753c987),
	.w1(32'hb9aaa906),
	.w2(32'hb8578049),
	.w3(32'hb9b94d9e),
	.w4(32'hba3d5668),
	.w5(32'hb98dabd7),
	.w6(32'h38a42336),
	.w7(32'h381a36af),
	.w8(32'h3952b6be),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb0196),
	.w1(32'h38b6bc6d),
	.w2(32'h393eb333),
	.w3(32'h3878a92b),
	.w4(32'hb8800445),
	.w5(32'h39550df2),
	.w6(32'hb95f2b6e),
	.w7(32'h375c92d2),
	.w8(32'h39fe5ade),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4c195),
	.w1(32'hb7bf6c6e),
	.w2(32'hb745fef1),
	.w3(32'hb90720e7),
	.w4(32'hb8c289df),
	.w5(32'hb7c49e8b),
	.w6(32'hb7ce7464),
	.w7(32'hb77e181b),
	.w8(32'hb7e37ee8),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c028e8),
	.w1(32'hb8ade65c),
	.w2(32'h387ffacd),
	.w3(32'h36ab05cb),
	.w4(32'h38cd81f4),
	.w5(32'h39058873),
	.w6(32'h398da52b),
	.w7(32'h37ab412a),
	.w8(32'h37a30ebd),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373df499),
	.w1(32'h38c65bb0),
	.w2(32'h376d45f5),
	.w3(32'h3782c43c),
	.w4(32'h38732b12),
	.w5(32'h384020d2),
	.w6(32'h386753db),
	.w7(32'h38a9a9a2),
	.w8(32'hb7c2dbf1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc090b),
	.w1(32'hb80bd4db),
	.w2(32'h388d77ce),
	.w3(32'hb8b896ae),
	.w4(32'hb632c489),
	.w5(32'h38b8e8fe),
	.w6(32'hb9342444),
	.w7(32'hb88ee2d7),
	.w8(32'h38701350),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3957f6ba),
	.w1(32'hb87ac76d),
	.w2(32'h389c7da4),
	.w3(32'hb90c43b0),
	.w4(32'hb888c81b),
	.w5(32'hb913046f),
	.w6(32'hb9760dad),
	.w7(32'h37ad23c4),
	.w8(32'hb7016e52),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079af9),
	.w1(32'hba415033),
	.w2(32'h38516e81),
	.w3(32'h38536434),
	.w4(32'hba396850),
	.w5(32'hb9bb2a24),
	.w6(32'hba068d19),
	.w7(32'hba4110f0),
	.w8(32'hb7934b74),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcdd43),
	.w1(32'h388cf268),
	.w2(32'hb8da18e9),
	.w3(32'h3824ccdf),
	.w4(32'hb7a7c59f),
	.w5(32'h36eb03cc),
	.w6(32'hb9233133),
	.w7(32'hb89edff5),
	.w8(32'hb8a92043),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919cb46),
	.w1(32'h3948ff71),
	.w2(32'h3972642c),
	.w3(32'h391941bf),
	.w4(32'hb9093e23),
	.w5(32'hb8e36583),
	.w6(32'hb86e7856),
	.w7(32'hb925a722),
	.w8(32'h38145b77),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb949685d),
	.w1(32'hba89d7a5),
	.w2(32'hb9b8fee1),
	.w3(32'h37033318),
	.w4(32'hbab7eb8a),
	.w5(32'hb9acf145),
	.w6(32'h39b8628c),
	.w7(32'hba56e264),
	.w8(32'hb92a7be8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3716e642),
	.w1(32'h389fc350),
	.w2(32'h38bc6a8d),
	.w3(32'h39068bc6),
	.w4(32'h39cefa69),
	.w5(32'h38ea5f68),
	.w6(32'h38cfff6b),
	.w7(32'h3990815f),
	.w8(32'h3895386b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cadeec),
	.w1(32'h39900c80),
	.w2(32'h38a8e443),
	.w3(32'h396266f2),
	.w4(32'hb93d4cfb),
	.w5(32'hb91aa765),
	.w6(32'hb883252d),
	.w7(32'hb94a79c1),
	.w8(32'h389450f3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ae8ffe),
	.w1(32'h37867e07),
	.w2(32'h378bb302),
	.w3(32'h3727e6ac),
	.w4(32'h3807b8ef),
	.w5(32'h388b94a6),
	.w6(32'hb88141a0),
	.w7(32'h379ab62e),
	.w8(32'h38b16e25),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09e37d),
	.w1(32'h3a0dab63),
	.w2(32'h39175aa3),
	.w3(32'h38f1e16b),
	.w4(32'hb81afa68),
	.w5(32'hb904f2cc),
	.w6(32'hb9b76f94),
	.w7(32'hb831d7c1),
	.w8(32'h3895f38c),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389cc279),
	.w1(32'h39f60e6b),
	.w2(32'h39f67ef8),
	.w3(32'hb81b244c),
	.w4(32'h39a0c01f),
	.w5(32'h39ae2e35),
	.w6(32'h369737dc),
	.w7(32'h38ca4f9f),
	.w8(32'h3913eed9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368d1306),
	.w1(32'h37383622),
	.w2(32'h37c26d60),
	.w3(32'hb58c9d49),
	.w4(32'hb707debb),
	.w5(32'hb77b11c2),
	.w6(32'hb68dac16),
	.w7(32'h36b9d177),
	.w8(32'hb7a64a67),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739fd35),
	.w1(32'hb7a523fd),
	.w2(32'h3798888d),
	.w3(32'hb7aa0e01),
	.w4(32'h37a35590),
	.w5(32'h38440343),
	.w6(32'hb7afbb07),
	.w7(32'h37b252de),
	.w8(32'h37f97d5f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bae137),
	.w1(32'h378cbf8f),
	.w2(32'hb87b1251),
	.w3(32'h38c68720),
	.w4(32'h391ed699),
	.w5(32'hb78de79a),
	.w6(32'h38aa9ff3),
	.w7(32'h391d53ca),
	.w8(32'hb922e3d2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb835b75f),
	.w1(32'h392430bf),
	.w2(32'hb84d0125),
	.w3(32'hb85e7a9f),
	.w4(32'hb96e1b0f),
	.w5(32'hb8c14f7b),
	.w6(32'hb99e709a),
	.w7(32'hb9d15c7e),
	.w8(32'hb92d57d0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963dc5c),
	.w1(32'h387d514a),
	.w2(32'hb83a1622),
	.w3(32'h38c2d591),
	.w4(32'hb8326a6a),
	.w5(32'h3885395e),
	.w6(32'hb8c91e4f),
	.w7(32'h38a8b051),
	.w8(32'h397fe315),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb619f51b),
	.w1(32'h3783848b),
	.w2(32'h3791f8fc),
	.w3(32'hb71f978e),
	.w4(32'hb7b7cb25),
	.w5(32'h371832a7),
	.w6(32'hb71f84ab),
	.w7(32'hb7a39f46),
	.w8(32'hb71353f1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c20db0),
	.w1(32'h38d93417),
	.w2(32'h38278caa),
	.w3(32'h390d79f6),
	.w4(32'hb819af47),
	.w5(32'hb758986a),
	.w6(32'hb8316c20),
	.w7(32'hb95e628c),
	.w8(32'h36bb9712),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19efc5),
	.w1(32'h38be5278),
	.w2(32'hb863929e),
	.w3(32'h39904b99),
	.w4(32'hb787c43d),
	.w5(32'hb95f2d56),
	.w6(32'hb9331cb7),
	.w7(32'hb9ad1751),
	.w8(32'hb999cc49),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998aeea),
	.w1(32'hba654fa7),
	.w2(32'hb77f7dce),
	.w3(32'hb8fbf761),
	.w4(32'hba5b5516),
	.w5(32'h37e80c72),
	.w6(32'h39816468),
	.w7(32'hb9a0f0d7),
	.w8(32'h382f61bd),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399f138f),
	.w1(32'h39853df7),
	.w2(32'h39b69150),
	.w3(32'h3954192d),
	.w4(32'h37fcc80b),
	.w5(32'h39090cef),
	.w6(32'hb81d6ff4),
	.w7(32'hb92b8459),
	.w8(32'h392142cc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bdbdcd),
	.w1(32'h38665740),
	.w2(32'hb901090c),
	.w3(32'hb98bf277),
	.w4(32'hb96072dc),
	.w5(32'hb954d149),
	.w6(32'hba004fea),
	.w7(32'hb99c66cd),
	.w8(32'hb9a44308),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c697f),
	.w1(32'h3992774d),
	.w2(32'h38cfafa8),
	.w3(32'h3988b319),
	.w4(32'h3a16ab7f),
	.w5(32'h3a08fadc),
	.w6(32'h396cd203),
	.w7(32'h3954256a),
	.w8(32'h3972529a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39805884),
	.w1(32'h38e33b58),
	.w2(32'h3a11b18a),
	.w3(32'h3828782d),
	.w4(32'hb5a9f0d0),
	.w5(32'h39cdb798),
	.w6(32'hb85a2768),
	.w7(32'hb95233f8),
	.w8(32'h3939671d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384fe46d),
	.w1(32'h39efecc6),
	.w2(32'h3904a001),
	.w3(32'hb9a42a4c),
	.w4(32'hb8d8bccb),
	.w5(32'hb94a9922),
	.w6(32'hb9ab661b),
	.w7(32'hb99b6033),
	.w8(32'hb91f3d55),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e69c9d),
	.w1(32'h3918ac91),
	.w2(32'h392946ed),
	.w3(32'hb8071dc6),
	.w4(32'h3949b9f3),
	.w5(32'h393671fb),
	.w6(32'hb858f2b3),
	.w7(32'h38ebc280),
	.w8(32'h3799a4e7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92b90dc),
	.w1(32'hb880c28c),
	.w2(32'h35e051d5),
	.w3(32'hb86d898e),
	.w4(32'hb8bda53d),
	.w5(32'hb8d251bd),
	.w6(32'hb8989d49),
	.w7(32'hb7e6c2c6),
	.w8(32'h37ccf371),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8335141),
	.w1(32'hb82dfab0),
	.w2(32'h368eb416),
	.w3(32'hb8704b45),
	.w4(32'hb7537d26),
	.w5(32'h38a6a3be),
	.w6(32'h36778bb4),
	.w7(32'h3856569f),
	.w8(32'hb77a7512),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a1c28),
	.w1(32'hb930255e),
	.w2(32'h38a879cb),
	.w3(32'hb93a6a7b),
	.w4(32'hba10482f),
	.w5(32'h38a827b0),
	.w6(32'hb9850990),
	.w7(32'hb993108b),
	.w8(32'h390d0cb9),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d1636e),
	.w1(32'hb775f054),
	.w2(32'hb7b0208a),
	.w3(32'h37a599b1),
	.w4(32'h37ce68ee),
	.w5(32'hb859b726),
	.w6(32'h37bcf6be),
	.w7(32'h38097ce2),
	.w8(32'hb8293be2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b03a87),
	.w1(32'h3975348e),
	.w2(32'h39eab38f),
	.w3(32'h3843efce),
	.w4(32'h38d671be),
	.w5(32'h3959047e),
	.w6(32'hb751fa74),
	.w7(32'hb89e68af),
	.w8(32'h38ed442c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89f377b),
	.w1(32'hb83ade30),
	.w2(32'hb6e0c4e0),
	.w3(32'hb8aa529d),
	.w4(32'h378a7249),
	.w5(32'h385d99b5),
	.w6(32'hb86ef280),
	.w7(32'h38badd4d),
	.w8(32'h37e53ba4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb726321f),
	.w1(32'hb4aa1d86),
	.w2(32'hb74ab012),
	.w3(32'h37e21b04),
	.w4(32'h38807282),
	.w5(32'hb6a0e58e),
	.w6(32'hb88e2369),
	.w7(32'h38d3db38),
	.w8(32'hb8e04622),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb731e445),
	.w1(32'hb8048028),
	.w2(32'hb84b4ba0),
	.w3(32'hb84c8149),
	.w4(32'hb8bdcbc8),
	.w5(32'hb8ceb419),
	.w6(32'hb7dc427f),
	.w7(32'hb8abd90b),
	.w8(32'hb855bcd6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cfaeab),
	.w1(32'hb71dc381),
	.w2(32'h37d2c2be),
	.w3(32'hb70d6737),
	.w4(32'hb841eece),
	.w5(32'hb70f96c2),
	.w6(32'h37c4909f),
	.w7(32'hb89232f2),
	.w8(32'hb8c3de06),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb26be),
	.w1(32'h3a0a2afe),
	.w2(32'h3943e176),
	.w3(32'hb878ba54),
	.w4(32'h3819b177),
	.w5(32'h3873d59e),
	.w6(32'hb9c2c786),
	.w7(32'hb98502ea),
	.w8(32'hb9464c84),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6f2f0),
	.w1(32'h3a3dc741),
	.w2(32'h39d0df0b),
	.w3(32'hb88d991b),
	.w4(32'hb9849611),
	.w5(32'hb93043b3),
	.w6(32'hb980177b),
	.w7(32'h39412666),
	.w8(32'h387c44cb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb792caf5),
	.w1(32'hb6ad14f3),
	.w2(32'h3810290f),
	.w3(32'h36d764da),
	.w4(32'h38a14fa9),
	.w5(32'hb8abee39),
	.w6(32'h38b02cf5),
	.w7(32'h393589cd),
	.w8(32'hb911a1f3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b75964),
	.w1(32'hb9705ff8),
	.w2(32'hba214073),
	.w3(32'h39f12667),
	.w4(32'hb936a2b6),
	.w5(32'hba0575ad),
	.w6(32'h3981e9be),
	.w7(32'hb8ca5598),
	.w8(32'hb99d1b2c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ab577),
	.w1(32'hb85c71d9),
	.w2(32'h369adc42),
	.w3(32'hb8425833),
	.w4(32'h36d363dd),
	.w5(32'hb72e1f34),
	.w6(32'hb8801598),
	.w7(32'h37c23936),
	.w8(32'hb85ebf47),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8755c7d),
	.w1(32'h38a2ec43),
	.w2(32'h394899c1),
	.w3(32'h384bdd4a),
	.w4(32'h3826f1ad),
	.w5(32'h37af9671),
	.w6(32'h388a02e1),
	.w7(32'hb91aa9bd),
	.w8(32'hb8e7d73d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd125c),
	.w1(32'hb99f1c10),
	.w2(32'hb8be1daa),
	.w3(32'hb90ab22b),
	.w4(32'hb8f506fc),
	.w5(32'hb7d983a9),
	.w6(32'hb91ee12b),
	.w7(32'hb90939ba),
	.w8(32'hb82e7842),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a9683),
	.w1(32'h3997ac85),
	.w2(32'h38732590),
	.w3(32'h390c289c),
	.w4(32'hb8e73071),
	.w5(32'hb968d90d),
	.w6(32'hb8eb5c20),
	.w7(32'hb967b3d1),
	.w8(32'hb8f7295d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f704dc),
	.w1(32'h38c0f421),
	.w2(32'h394ec5cf),
	.w3(32'h37691f78),
	.w4(32'h388cc939),
	.w5(32'h3946c342),
	.w6(32'h3616b752),
	.w7(32'h38eda62f),
	.w8(32'h3929c566),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e8282),
	.w1(32'hb69dad6c),
	.w2(32'h39f9d3f7),
	.w3(32'hb9a85669),
	.w4(32'hb9aec03c),
	.w5(32'h39500859),
	.w6(32'hb9fcef62),
	.w7(32'hb9285745),
	.w8(32'h39078c66),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370929a8),
	.w1(32'h3814118d),
	.w2(32'h365753a1),
	.w3(32'h3801c3fd),
	.w4(32'h36a9e02c),
	.w5(32'h391150e8),
	.w6(32'h381632f7),
	.w7(32'h35414b14),
	.w8(32'h390a285a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36884ebc),
	.w1(32'hb8791f98),
	.w2(32'h3760a2ce),
	.w3(32'hb8e8f955),
	.w4(32'h38b4739e),
	.w5(32'h37690fea),
	.w6(32'hb83a4054),
	.w7(32'h38f1460e),
	.w8(32'h3876f74d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897ceba),
	.w1(32'hb86bbca6),
	.w2(32'h382478d8),
	.w3(32'hb88be114),
	.w4(32'hb7d446c2),
	.w5(32'h3792dcda),
	.w6(32'hb93d4c0d),
	.w7(32'hb8c0f305),
	.w8(32'hb80145a5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8865c2b),
	.w1(32'hb8fe91da),
	.w2(32'hb818d68c),
	.w3(32'h38d70860),
	.w4(32'hb873754f),
	.w5(32'hb8935095),
	.w6(32'h38549b34),
	.w7(32'hb823bb62),
	.w8(32'h37fb2176),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80d2264),
	.w1(32'h38964176),
	.w2(32'hb8e3ffc8),
	.w3(32'h3841f28d),
	.w4(32'hb8dd6306),
	.w5(32'hb70b8ea0),
	.w6(32'h388e9fea),
	.w7(32'hb9139eb0),
	.w8(32'hb7855eca),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ab1db9),
	.w1(32'hb82b48c2),
	.w2(32'hb7ec8294),
	.w3(32'hb7dc2fb6),
	.w4(32'h376bda1e),
	.w5(32'h38423737),
	.w6(32'hb7b39033),
	.w7(32'h3533f0f8),
	.w8(32'h38373fef),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9291f27),
	.w1(32'hb9cbd7da),
	.w2(32'h3963567d),
	.w3(32'hb895b3ae),
	.w4(32'hb839f0eb),
	.w5(32'h37c66fbb),
	.w6(32'h39f50166),
	.w7(32'h38504a9c),
	.w8(32'h38b2d092),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce4757),
	.w1(32'hba2a348b),
	.w2(32'hb9813e90),
	.w3(32'hb9ba49b8),
	.w4(32'hb9bc77e0),
	.w5(32'hb98f8884),
	.w6(32'h398c9726),
	.w7(32'h38581565),
	.w8(32'hb7b9f428),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386bb41a),
	.w1(32'h39928b09),
	.w2(32'hb9b897f0),
	.w3(32'hb7e5dce0),
	.w4(32'h3941dda7),
	.w5(32'hb9bf5e94),
	.w6(32'h391780b3),
	.w7(32'h38180809),
	.w8(32'hb9bdacc6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a23ff),
	.w1(32'h3920b061),
	.w2(32'hb7bec1c2),
	.w3(32'hb7869fe1),
	.w4(32'h386bd2d4),
	.w5(32'h384377b7),
	.w6(32'h38d784a6),
	.w7(32'h390ccd64),
	.w8(32'h388b3339),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a0d2b),
	.w1(32'hb9d95a39),
	.w2(32'hba0fcc8c),
	.w3(32'hb9305277),
	.w4(32'hba4d4f56),
	.w5(32'hb9b35f9a),
	.w6(32'h39392d8a),
	.w7(32'hb92858f6),
	.w8(32'h399ec2f5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396365e0),
	.w1(32'h39b87a52),
	.w2(32'h39be23e6),
	.w3(32'h39869ef6),
	.w4(32'h399296bf),
	.w5(32'h3967d119),
	.w6(32'h38e77c7f),
	.w7(32'h38e37a31),
	.w8(32'h38900b1f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dde591),
	.w1(32'hb89cdd18),
	.w2(32'hb8aa3744),
	.w3(32'hb83e8cb6),
	.w4(32'hb88893e7),
	.w5(32'hb8d927e4),
	.w6(32'hb79bb967),
	.w7(32'hb79bc136),
	.w8(32'hb90f3aa0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7847178),
	.w1(32'hb5e4e2fa),
	.w2(32'h3816199c),
	.w3(32'h37be2a1b),
	.w4(32'h38800b96),
	.w5(32'h37a1bcf4),
	.w6(32'hb80d335d),
	.w7(32'hb719a209),
	.w8(32'h378c90ba),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7e6c1),
	.w1(32'h38528bb6),
	.w2(32'h38557d97),
	.w3(32'hb6acffa7),
	.w4(32'h39185ff2),
	.w5(32'h37e9d348),
	.w6(32'h3880ac3c),
	.w7(32'h389673fa),
	.w8(32'hb7a63e07),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38323ca0),
	.w1(32'hb8810ebb),
	.w2(32'hb80461ef),
	.w3(32'hb862ab42),
	.w4(32'h37f7f2b4),
	.w5(32'h36591496),
	.w6(32'hb8853a0c),
	.w7(32'h3765645f),
	.w8(32'hb7f96965),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853c705),
	.w1(32'hb79e0897),
	.w2(32'hb957c8c3),
	.w3(32'hb87f9dd4),
	.w4(32'hb927eb94),
	.w5(32'hb88e6b6f),
	.w6(32'h38e3a29d),
	.w7(32'hb83b2cb4),
	.w8(32'h38d436e7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f002a),
	.w1(32'hb9827eab),
	.w2(32'hb98c136a),
	.w3(32'hb87e3bec),
	.w4(32'hb987b632),
	.w5(32'hb9965407),
	.w6(32'hb8cefd67),
	.w7(32'h36f57f22),
	.w8(32'h388f7477),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39393731),
	.w1(32'h39abe451),
	.w2(32'h384de532),
	.w3(32'hb83469b3),
	.w4(32'h395d49fb),
	.w5(32'h394d6cb1),
	.w6(32'hb968376d),
	.w7(32'h38a257d9),
	.w8(32'h392a1c31),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca15fe),
	.w1(32'hb889ba63),
	.w2(32'h39091364),
	.w3(32'hb9579877),
	.w4(32'hb83508b3),
	.w5(32'hb797483a),
	.w6(32'hb8f34df9),
	.w7(32'h38385060),
	.w8(32'h3743e05c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e93574),
	.w1(32'hb9b22020),
	.w2(32'hb9f9a5b6),
	.w3(32'h38b252e1),
	.w4(32'hb96a3b78),
	.w5(32'hb9a9ef0e),
	.w6(32'h388e6dd0),
	.w7(32'hb88cd7b5),
	.w8(32'hb8f32e52),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f517b),
	.w1(32'hb899cfaa),
	.w2(32'hb97fe84a),
	.w3(32'h38ef720c),
	.w4(32'h373fa291),
	.w5(32'hb9aa0aea),
	.w6(32'h3960f8e9),
	.w7(32'h39024436),
	.w8(32'hb91859ec),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78df8d5),
	.w1(32'hb6acbf79),
	.w2(32'h36d32926),
	.w3(32'hb7b23d72),
	.w4(32'hb70dd213),
	.w5(32'hb6d5735b),
	.w6(32'hb67ce6ca),
	.w7(32'h373c60c8),
	.w8(32'h35a22497),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8175ec8),
	.w1(32'h3628b105),
	.w2(32'hb8483fb0),
	.w3(32'h38cab08c),
	.w4(32'hb958d13b),
	.w5(32'hb8592adf),
	.w6(32'h39944579),
	.w7(32'h388c843c),
	.w8(32'hb997262f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c438e0),
	.w1(32'h3820bd18),
	.w2(32'h3740fa46),
	.w3(32'h3863a030),
	.w4(32'h3834d71b),
	.w5(32'h365eb6bc),
	.w6(32'h38425621),
	.w7(32'h375fd214),
	.w8(32'h372b21bc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b2163),
	.w1(32'hb8ee3f6f),
	.w2(32'hb949b10f),
	.w3(32'hb7c3927f),
	.w4(32'hb8978a86),
	.w5(32'hb7d16070),
	.w6(32'h37c8c127),
	.w7(32'h3883b509),
	.w8(32'h38486d24),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5555b),
	.w1(32'h371991fd),
	.w2(32'hb812047b),
	.w3(32'hb9d6fb7c),
	.w4(32'hb892578b),
	.w5(32'hb840e328),
	.w6(32'hba0e0b29),
	.w7(32'hb90257e4),
	.w8(32'hb9abbd06),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c3860),
	.w1(32'h38e8324c),
	.w2(32'hb7e7b5ae),
	.w3(32'h381c176b),
	.w4(32'h38841c0a),
	.w5(32'hb72a6a61),
	.w6(32'hb93f6c10),
	.w7(32'hb8f51df9),
	.w8(32'hb91dbdd5),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c3dc4d),
	.w1(32'hb78a41d9),
	.w2(32'h384283bd),
	.w3(32'hb84245cd),
	.w4(32'h388a5f43),
	.w5(32'hb72202a3),
	.w6(32'hb79a7637),
	.w7(32'h38379fc1),
	.w8(32'h382afb9f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39940a60),
	.w1(32'h3567a510),
	.w2(32'hb98853f4),
	.w3(32'h38990299),
	.w4(32'hb841bf03),
	.w5(32'hb8b66698),
	.w6(32'hb85d96bd),
	.w7(32'h378ab5b8),
	.w8(32'hb890a83c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd43e8),
	.w1(32'h398db97a),
	.w2(32'h39a25c86),
	.w3(32'h38ddfcc3),
	.w4(32'h38e6da52),
	.w5(32'h394449cb),
	.w6(32'hb8c6f9ee),
	.w7(32'hb8c63568),
	.w8(32'h390f8b55),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3898776d),
	.w1(32'h3888da5a),
	.w2(32'hb9658165),
	.w3(32'hb9111e55),
	.w4(32'hb931741d),
	.w5(32'hb978e549),
	.w6(32'hb945c618),
	.w7(32'h37892e2b),
	.w8(32'hb82d439d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378369ea),
	.w1(32'hb79914cf),
	.w2(32'h37a2aea2),
	.w3(32'h383ffe79),
	.w4(32'h38429a91),
	.w5(32'h3882c186),
	.w6(32'hb794512e),
	.w7(32'hb71fdfe9),
	.w8(32'h3830c29c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861bd4e),
	.w1(32'hb8746d53),
	.w2(32'h381aa80f),
	.w3(32'hb7e3f31d),
	.w4(32'h37813d91),
	.w5(32'h3739743a),
	.w6(32'hb80b27e0),
	.w7(32'h374d4b1d),
	.w8(32'h38185a59),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ae711),
	.w1(32'hb907ea89),
	.w2(32'hb960c7b3),
	.w3(32'hb99ef44e),
	.w4(32'hb92a50c1),
	.w5(32'hb989da4d),
	.w6(32'hb993e88f),
	.w7(32'hb9262b96),
	.w8(32'hb904f6ee),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e09e9),
	.w1(32'hb9f1027a),
	.w2(32'hb9805b8d),
	.w3(32'hb9ec4a5f),
	.w4(32'hba740dd6),
	.w5(32'hba1300e1),
	.w6(32'hb8aff284),
	.w7(32'hb9984d43),
	.w8(32'hb989c04c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdef7d),
	.w1(32'h38b05ecf),
	.w2(32'h39df4b5a),
	.w3(32'h3904a96a),
	.w4(32'h39cd67b4),
	.w5(32'h394ab44e),
	.w6(32'h39063924),
	.w7(32'h390bf761),
	.w8(32'h3916fcf9),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cceea4),
	.w1(32'hb9da71b6),
	.w2(32'hb973a604),
	.w3(32'h38f1ee20),
	.w4(32'hba01a9e2),
	.w5(32'hb94a8485),
	.w6(32'h39618478),
	.w7(32'hb98f006a),
	.w8(32'hb8c1d3e6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37452a3e),
	.w1(32'h372790f0),
	.w2(32'hb71b1b16),
	.w3(32'h3845b21e),
	.w4(32'h37e07f4f),
	.w5(32'hb778bb37),
	.w6(32'hb7e69327),
	.w7(32'hb81f6275),
	.w8(32'hb7a8407f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6b88f),
	.w1(32'hb80e993d),
	.w2(32'hb81185d4),
	.w3(32'hb971b39d),
	.w4(32'hb9420bf3),
	.w5(32'hb89178c0),
	.w6(32'hb98497ed),
	.w7(32'hb8fee57b),
	.w8(32'hb85c87b5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a57387),
	.w1(32'h39732d4e),
	.w2(32'hba9d25c6),
	.w3(32'hb8e88c15),
	.w4(32'hb89bf9e5),
	.w5(32'hba831895),
	.w6(32'h3908fb34),
	.w7(32'h392fe3ac),
	.w8(32'hba0a740c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98db0c9),
	.w1(32'hba922a97),
	.w2(32'hba4a57e2),
	.w3(32'hb9b99b22),
	.w4(32'hba8a2f82),
	.w5(32'hba302d5a),
	.w6(32'h399da737),
	.w7(32'hb9471a44),
	.w8(32'hb8953a25),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba422231),
	.w1(32'hb9cdfd7e),
	.w2(32'hba07d89b),
	.w3(32'hba0d66d6),
	.w4(32'hb9786716),
	.w5(32'hba22c9dd),
	.w6(32'hb92cf481),
	.w7(32'hb8acb9b0),
	.w8(32'hb9c0b9ce),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798a133),
	.w1(32'h38dd1448),
	.w2(32'h3841b0fb),
	.w3(32'hb7e7cdbf),
	.w4(32'h3939eded),
	.w5(32'h3905e142),
	.w6(32'hb92c7d03),
	.w7(32'h389a8671),
	.w8(32'hb7c41ae5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9b803),
	.w1(32'h3975abb1),
	.w2(32'h389775eb),
	.w3(32'hb8b32136),
	.w4(32'h3742ceb8),
	.w5(32'h3775f811),
	.w6(32'hb9b0f179),
	.w7(32'hb9017686),
	.w8(32'hb84cb65b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a9ccef),
	.w1(32'h371dcdb7),
	.w2(32'h36a6275f),
	.w3(32'h3793c10b),
	.w4(32'h370f486f),
	.w5(32'hb807d07d),
	.w6(32'h3763878c),
	.w7(32'h36e02e70),
	.w8(32'hb6b92ff0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cb798e),
	.w1(32'hb72831f1),
	.w2(32'hb7ec6ca6),
	.w3(32'hb6b7b421),
	.w4(32'hb787ad9a),
	.w5(32'h37930421),
	.w6(32'h37636737),
	.w7(32'hb77ac8a6),
	.w8(32'h3831d805),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e0bbdf),
	.w1(32'hb8183936),
	.w2(32'hb89cfb0d),
	.w3(32'hb6b5c335),
	.w4(32'hb8549992),
	.w5(32'h38611daf),
	.w6(32'h37ec1051),
	.w7(32'hb7cd090e),
	.w8(32'h381020b1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891c31d),
	.w1(32'hb8069fdf),
	.w2(32'h38f0a8a6),
	.w3(32'hb80f7454),
	.w4(32'h3891b7be),
	.w5(32'hba96a0be),
	.w6(32'hb8c4c465),
	.w7(32'h3888cda9),
	.w8(32'hb7ece010),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3e946),
	.w1(32'h3a9ed8df),
	.w2(32'h3aacd5ca),
	.w3(32'hba0cc1f1),
	.w4(32'h3a4abb5d),
	.w5(32'h390c4d81),
	.w6(32'h3b113abe),
	.w7(32'h3b2692b6),
	.w8(32'hb99e54b6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0003b3),
	.w1(32'hbb8b9c67),
	.w2(32'h3a702f5a),
	.w3(32'hbb978584),
	.w4(32'hb9fcdae1),
	.w5(32'hb9fba1e6),
	.w6(32'h3a422ee0),
	.w7(32'hbb357335),
	.w8(32'hb906ce37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2dc00),
	.w1(32'hbb5b6c9b),
	.w2(32'hbb94b80c),
	.w3(32'hbaeba1a1),
	.w4(32'h3af3e94c),
	.w5(32'hba3c204d),
	.w6(32'hba85ed1c),
	.w7(32'hbaee1416),
	.w8(32'hbb16ca23),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2392f8),
	.w1(32'hb905b460),
	.w2(32'hbc021d41),
	.w3(32'hbb06d7ef),
	.w4(32'h3b24946f),
	.w5(32'h3af6559f),
	.w6(32'hbbdfc129),
	.w7(32'hbb846670),
	.w8(32'hb989f98d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb705dc2),
	.w1(32'hbb37ce70),
	.w2(32'hbb03235d),
	.w3(32'hba2dc906),
	.w4(32'h3b32a240),
	.w5(32'hbc0ee2d7),
	.w6(32'hbb3c80b2),
	.w7(32'hba6d4144),
	.w8(32'hbc16675f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7b4d2),
	.w1(32'hbba003f5),
	.w2(32'hbc083b61),
	.w3(32'hbbec7175),
	.w4(32'hbc2c938c),
	.w5(32'hba968a13),
	.w6(32'hbbb4bff1),
	.w7(32'hbc05cba7),
	.w8(32'h3ad03098),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb72909),
	.w1(32'hbb885e55),
	.w2(32'hbb565aa1),
	.w3(32'hbb0cbb58),
	.w4(32'h3b86615b),
	.w5(32'hbb3202f5),
	.w6(32'hbaf6c7ee),
	.w7(32'hbb4ead67),
	.w8(32'hbaa8b3f2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac005),
	.w1(32'hbb6dd6ee),
	.w2(32'h3add93da),
	.w3(32'hbaea936c),
	.w4(32'h3ba06266),
	.w5(32'hbb2d44a2),
	.w6(32'h3ac1d96b),
	.w7(32'h3b8af8b2),
	.w8(32'h3b24b6c4),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8662d),
	.w1(32'h3a841812),
	.w2(32'hba65ce3c),
	.w3(32'hbb952fd9),
	.w4(32'h3a9b306c),
	.w5(32'h39a35458),
	.w6(32'hbac7732a),
	.w7(32'h3bafa0ae),
	.w8(32'hbbac4c02),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acc46),
	.w1(32'hbada4f24),
	.w2(32'hbb1b7d8f),
	.w3(32'hbb98dc26),
	.w4(32'hbb338c55),
	.w5(32'h3a2b37f1),
	.w6(32'hbbb09518),
	.w7(32'hbb9df114),
	.w8(32'h3b0c8f85),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc5ae),
	.w1(32'h3ba30727),
	.w2(32'h3b547fb2),
	.w3(32'h3b52463f),
	.w4(32'h3b12936b),
	.w5(32'h3b9828fd),
	.w6(32'h3bb59e1b),
	.w7(32'h3b914243),
	.w8(32'hbaa5b9e5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba504bd8),
	.w1(32'h3a093829),
	.w2(32'h3b8950dc),
	.w3(32'h3b690837),
	.w4(32'h3b8df9a2),
	.w5(32'hb996c349),
	.w6(32'hba2dc313),
	.w7(32'h3af80699),
	.w8(32'hb9d90d94),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b8844),
	.w1(32'h3b053826),
	.w2(32'h39d1c469),
	.w3(32'hba42684d),
	.w4(32'h3a54ad37),
	.w5(32'h3b6f271e),
	.w6(32'h3bd8a282),
	.w7(32'h3b8d333e),
	.w8(32'h3b1de024),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842790),
	.w1(32'hb994b385),
	.w2(32'h3ad42a28),
	.w3(32'hbabad42e),
	.w4(32'hbb313f7f),
	.w5(32'h3b98242e),
	.w6(32'hbac6713b),
	.w7(32'hba9d7a72),
	.w8(32'h3bf283ea),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2cf0a),
	.w1(32'h3bb8766d),
	.w2(32'h3be6be86),
	.w3(32'h3b90ffa8),
	.w4(32'h3ba2d7d2),
	.w5(32'h3ae18fb3),
	.w6(32'h3c011eef),
	.w7(32'h3bdf7338),
	.w8(32'h3bee3a4f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b667f65),
	.w1(32'hba5069bf),
	.w2(32'hba4be64c),
	.w3(32'h3b307027),
	.w4(32'h3a7aad1f),
	.w5(32'hbb6da275),
	.w6(32'hbb02bae2),
	.w7(32'h3b399fc3),
	.w8(32'hbbe8434b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cc9b8),
	.w1(32'hbb7d4df6),
	.w2(32'h3aeb08d8),
	.w3(32'hbaa1a7a4),
	.w4(32'h3b471e1a),
	.w5(32'h3b476e5e),
	.w6(32'hbb30880f),
	.w7(32'hb927e879),
	.w8(32'hb962609a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15fae3),
	.w1(32'hb9aee544),
	.w2(32'hbb779749),
	.w3(32'hbaf96af1),
	.w4(32'h3a2b1f0d),
	.w5(32'h3bbaaf36),
	.w6(32'hbba0d21e),
	.w7(32'hba111551),
	.w8(32'h3b538272),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0852ad),
	.w1(32'h3b519b73),
	.w2(32'h3ac145f9),
	.w3(32'h3bc61104),
	.w4(32'h3aa5d7ad),
	.w5(32'hba441c41),
	.w6(32'h3bc5391d),
	.w7(32'h3aac642b),
	.w8(32'h3b90d116),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c103bf4),
	.w1(32'hba58aaf1),
	.w2(32'h34eed22a),
	.w3(32'hbb85e338),
	.w4(32'hbac552c7),
	.w5(32'h3ac8918d),
	.w6(32'hb99d18d1),
	.w7(32'hbb1b4814),
	.w8(32'h3a8844b9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00e4d3),
	.w1(32'hbab9459b),
	.w2(32'hb9e9608f),
	.w3(32'hb9f9256d),
	.w4(32'hba8e66f1),
	.w5(32'hbab6615b),
	.w6(32'h39d8315d),
	.w7(32'hba92558d),
	.w8(32'hbaf433ea),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb005d),
	.w1(32'h3b0825e8),
	.w2(32'hbb453234),
	.w3(32'hbb10d01c),
	.w4(32'hbb8c2c18),
	.w5(32'hb986e9b2),
	.w6(32'hbb02329a),
	.w7(32'hbb56c901),
	.w8(32'hbb21beea),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa81ce5),
	.w1(32'h3b797e76),
	.w2(32'h3b69c243),
	.w3(32'h3b31cf09),
	.w4(32'hba5bf0ce),
	.w5(32'h3b538f95),
	.w6(32'hbb12d775),
	.w7(32'h39e56191),
	.w8(32'hbae35e4d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03a0b6),
	.w1(32'h3c13da20),
	.w2(32'h3b36abfb),
	.w3(32'h3c49d351),
	.w4(32'hbb379afa),
	.w5(32'hbbb11ede),
	.w6(32'h3c4b820c),
	.w7(32'h3a47c7ae),
	.w8(32'hbbfaac7d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a32f),
	.w1(32'hbb83c4ed),
	.w2(32'h3b5c179d),
	.w3(32'hbc29c8fc),
	.w4(32'hba3b6b98),
	.w5(32'h3c113111),
	.w6(32'hbc7b67c8),
	.w7(32'hbb5e92f5),
	.w8(32'hba6c5849),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55cbd4),
	.w1(32'h3c3001b2),
	.w2(32'h3b4cf897),
	.w3(32'h3c0d0463),
	.w4(32'h3a1da168),
	.w5(32'hbbce5761),
	.w6(32'h3c42b606),
	.w7(32'h3ad27f27),
	.w8(32'hbbfbb4ef),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa79b),
	.w1(32'hbb9b1dc5),
	.w2(32'hbb1cbc40),
	.w3(32'hbc11019c),
	.w4(32'hb9ce1b60),
	.w5(32'h3be5309b),
	.w6(32'hbc44e180),
	.w7(32'hbba2ccb0),
	.w8(32'h3bfe4463),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ee42),
	.w1(32'h3bc11ce4),
	.w2(32'h39cc62c4),
	.w3(32'h3acfb677),
	.w4(32'hba112c35),
	.w5(32'h39661ec4),
	.w6(32'h3bcfb247),
	.w7(32'hbaa03b06),
	.w8(32'hbbf675b2),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6b7ef),
	.w1(32'hbaed0b80),
	.w2(32'hba9cd12f),
	.w3(32'hbb7a6480),
	.w4(32'h3a828be1),
	.w5(32'h3a012893),
	.w6(32'hbc11752e),
	.w7(32'hbbcf9213),
	.w8(32'hb8aeb6c7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf259),
	.w1(32'h3b7ef6c4),
	.w2(32'h3bbb25f7),
	.w3(32'h3b7f79f0),
	.w4(32'h3b77b14f),
	.w5(32'hbba5faa5),
	.w6(32'h3b92219c),
	.w7(32'h3ba17571),
	.w8(32'hbbd9e969),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule