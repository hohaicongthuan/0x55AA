module layer_10_featuremap_239(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f646),
	.w1(32'hbbe09ac0),
	.w2(32'hbbf9146e),
	.w3(32'hb95f5737),
	.w4(32'hba4358fe),
	.w5(32'h3a89dc7e),
	.w6(32'h3770e37b),
	.w7(32'h39e089d8),
	.w8(32'h3c1bbcd7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae155a),
	.w1(32'hbb890483),
	.w2(32'hbc483b9f),
	.w3(32'h3b813fe6),
	.w4(32'hbbad458f),
	.w5(32'hbb9dbc1e),
	.w6(32'h3c43f730),
	.w7(32'hbbde7de3),
	.w8(32'hbb21c951),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06fca2),
	.w1(32'hbbec8525),
	.w2(32'hbb20e5d0),
	.w3(32'hbbf615d1),
	.w4(32'hbba525de),
	.w5(32'hbc3ce52b),
	.w6(32'h3bf954a2),
	.w7(32'h39a6d6c2),
	.w8(32'hb8df5dbb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacd908),
	.w1(32'h3b83b232),
	.w2(32'h3c0888e1),
	.w3(32'hbbcd818d),
	.w4(32'h3b5ab98f),
	.w5(32'h3b2c19ae),
	.w6(32'hbc066482),
	.w7(32'h3c24f979),
	.w8(32'hbc7fe715),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c426d),
	.w1(32'hbaf9d477),
	.w2(32'h3c4305f7),
	.w3(32'hbc1d79ff),
	.w4(32'hb9680fb0),
	.w5(32'hbc47b9d8),
	.w6(32'hbcd8affe),
	.w7(32'h3beedeaa),
	.w8(32'hbc01fd2d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd97d45),
	.w1(32'hbbc6cfce),
	.w2(32'hbb5ed08e),
	.w3(32'hbbb7233c),
	.w4(32'hba3dd526),
	.w5(32'h3b30ce6d),
	.w6(32'hbc05a312),
	.w7(32'hbb0325cf),
	.w8(32'h3b8d8dc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef8487),
	.w1(32'hbbe879ef),
	.w2(32'hbc32cd80),
	.w3(32'h3ac209fb),
	.w4(32'hbbf471ff),
	.w5(32'hbc5601b9),
	.w6(32'h3b61e744),
	.w7(32'hbb569908),
	.w8(32'hbbea5285),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeac820),
	.w1(32'hb8e083c3),
	.w2(32'h3b1960cb),
	.w3(32'hbbc6ebc0),
	.w4(32'hbb5b7973),
	.w5(32'h3c07daa1),
	.w6(32'h3a8ceb14),
	.w7(32'hbab48918),
	.w8(32'h3c3aba0f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc2ab0),
	.w1(32'hbc1f5fff),
	.w2(32'hbc8bc43e),
	.w3(32'h3ba5e684),
	.w4(32'hbb74c35c),
	.w5(32'hbc49d2bc),
	.w6(32'hb9b81265),
	.w7(32'hbc4c7299),
	.w8(32'hbbf8cda3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b97e8),
	.w1(32'hbbc14a11),
	.w2(32'hba75d871),
	.w3(32'hbbcb0737),
	.w4(32'h3ab187f4),
	.w5(32'hbc2a0fa5),
	.w6(32'hbb599c78),
	.w7(32'h3bb24f3d),
	.w8(32'hbbd1023a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2754a),
	.w1(32'hbb7e0e96),
	.w2(32'h3ba0bbdf),
	.w3(32'hbbb4408b),
	.w4(32'hbb356f4c),
	.w5(32'h3bce9299),
	.w6(32'hbc70e3dd),
	.w7(32'h3b89bc26),
	.w8(32'hbb0c4877),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5c93a),
	.w1(32'hbc266972),
	.w2(32'hbc47cc70),
	.w3(32'h3ae8231f),
	.w4(32'hbc417d0b),
	.w5(32'h3bdab7b9),
	.w6(32'h3c87ae8d),
	.w7(32'hbbd4a816),
	.w8(32'h3c1fd484),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3aed01),
	.w1(32'hbc602511),
	.w2(32'hbc9c2542),
	.w3(32'h3c130b8e),
	.w4(32'hbbea407e),
	.w5(32'h3c0e0cd7),
	.w6(32'hbc1064fd),
	.w7(32'hbc132e3c),
	.w8(32'h3adc9e03),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb073cb6),
	.w1(32'hbbea7181),
	.w2(32'h3b5a10ce),
	.w3(32'hbb830ec8),
	.w4(32'hbb6d3c03),
	.w5(32'hbc313d41),
	.w6(32'h3b64f187),
	.w7(32'hbb7a2326),
	.w8(32'h3b6c1a0e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24cea7),
	.w1(32'hbc113e7b),
	.w2(32'hbb49a4c7),
	.w3(32'h3ac1ae8c),
	.w4(32'hba90eec2),
	.w5(32'h3c2b522e),
	.w6(32'hbc269eb9),
	.w7(32'hbbd36ce2),
	.w8(32'h3babb930),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb6c7f),
	.w1(32'hbc90053a),
	.w2(32'hbbc9b665),
	.w3(32'h3b523f61),
	.w4(32'h3a88cbc3),
	.w5(32'h3a146cb1),
	.w6(32'hbbaf40c2),
	.w7(32'hbae75529),
	.w8(32'hba177b4d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a24b8),
	.w1(32'hbc61efc6),
	.w2(32'hbc8790fe),
	.w3(32'h3c675d7b),
	.w4(32'hbb9c778f),
	.w5(32'hbbbb8fcb),
	.w6(32'hbaad0fb5),
	.w7(32'hbc5b601f),
	.w8(32'h3a744136),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb075688),
	.w1(32'h3824c73f),
	.w2(32'h3bcdace9),
	.w3(32'hbaad6cf6),
	.w4(32'h3b8a5ace),
	.w5(32'hbb44e1a2),
	.w6(32'h3a310db0),
	.w7(32'h3c538353),
	.w8(32'hbb57c1e6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fbb01),
	.w1(32'h3c17ab38),
	.w2(32'h3c4f2bb0),
	.w3(32'hbc7b7da7),
	.w4(32'hbb497b48),
	.w5(32'hbb848c74),
	.w6(32'hbc4714f0),
	.w7(32'h3c971e9e),
	.w8(32'h3a6deb85),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fba92),
	.w1(32'hbb3eef0d),
	.w2(32'h3b85a522),
	.w3(32'hbbe89844),
	.w4(32'h3adad7c6),
	.w5(32'h3b538697),
	.w6(32'hbbb00ddf),
	.w7(32'h3b9839c0),
	.w8(32'h3a712568),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390936af),
	.w1(32'hbb1dda02),
	.w2(32'h3a95a65d),
	.w3(32'h3bb7f635),
	.w4(32'h3bb74186),
	.w5(32'hbb95d947),
	.w6(32'h3c34b864),
	.w7(32'h3be6cd1d),
	.w8(32'hbb81ddd4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96b06d),
	.w1(32'h3b1dc39f),
	.w2(32'hb9a06896),
	.w3(32'hbb87ebc3),
	.w4(32'h3ad7a650),
	.w5(32'hbaea1e7f),
	.w6(32'hbb108903),
	.w7(32'h3b2c5d3d),
	.w8(32'h3a70afc8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be380a3),
	.w1(32'hbbd2efc4),
	.w2(32'hbc60b093),
	.w3(32'hba2de918),
	.w4(32'h39581f3e),
	.w5(32'h3c52d9c9),
	.w6(32'h3cdb59e9),
	.w7(32'hbb156832),
	.w8(32'h3b7b5272),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b887ec7),
	.w1(32'h398d595e),
	.w2(32'hb953411d),
	.w3(32'h395dfd10),
	.w4(32'h3bb18f29),
	.w5(32'h3b8753b5),
	.w6(32'hbb24f219),
	.w7(32'h3b9efb28),
	.w8(32'hbbc64e7a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c820c8),
	.w1(32'hbc0be33d),
	.w2(32'h3a9f5a61),
	.w3(32'h3a9c0aad),
	.w4(32'hbb13c13d),
	.w5(32'hbc486617),
	.w6(32'hbbfda031),
	.w7(32'h3baa8b62),
	.w8(32'hbb126196),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d17b5),
	.w1(32'hbb91bf77),
	.w2(32'hbacb869b),
	.w3(32'h3b87e867),
	.w4(32'h3abb028c),
	.w5(32'h3c63fe12),
	.w6(32'h3a06b73c),
	.w7(32'hba92d39a),
	.w8(32'h3b9b1672),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab748f1),
	.w1(32'h3aa67d34),
	.w2(32'h38489ccc),
	.w3(32'h3b8ffa09),
	.w4(32'hb98d59b6),
	.w5(32'hbafad8c3),
	.w6(32'h3b38fd97),
	.w7(32'hbb7e4e52),
	.w8(32'hbb17355a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4489af),
	.w1(32'hbc4521a5),
	.w2(32'hbc32079e),
	.w3(32'hbbea767d),
	.w4(32'hbc0e38c9),
	.w5(32'h3a9d1223),
	.w6(32'hbc0fc024),
	.w7(32'hbbfa3e16),
	.w8(32'h3b32f03f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff0e21),
	.w1(32'hbb9ad4c5),
	.w2(32'h3ba050b2),
	.w3(32'hbbe4e685),
	.w4(32'hba9883cd),
	.w5(32'h3a6605a3),
	.w6(32'hbbc3b20e),
	.w7(32'h3bf8161a),
	.w8(32'h3b5e5484),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d23a6),
	.w1(32'h3ab46876),
	.w2(32'hbae327a9),
	.w3(32'hbb6f4dbf),
	.w4(32'hbb9a1b49),
	.w5(32'hba96424d),
	.w6(32'h391b51eb),
	.w7(32'hbb07d463),
	.w8(32'h3c1ae20b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7d20),
	.w1(32'hbbe40296),
	.w2(32'hbbb199e7),
	.w3(32'h3b101770),
	.w4(32'hbbb34a6e),
	.w5(32'h3b47a29d),
	.w6(32'h3b452812),
	.w7(32'hbc3f13be),
	.w8(32'h3b2cff1c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e109d),
	.w1(32'hbc73252a),
	.w2(32'h3a2e5d23),
	.w3(32'hbb130e3b),
	.w4(32'hbb33d8c1),
	.w5(32'h3c03cc49),
	.w6(32'hbc48a332),
	.w7(32'hbb29b0bd),
	.w8(32'h38a316d1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca5f24),
	.w1(32'hbba44eee),
	.w2(32'h3b44428a),
	.w3(32'hbbcac225),
	.w4(32'hb96f13ab),
	.w5(32'hbb533176),
	.w6(32'h3b1e9550),
	.w7(32'h3a29a9e9),
	.w8(32'h3aa717fb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c8012),
	.w1(32'h3a8491ee),
	.w2(32'hbae15a16),
	.w3(32'hbb86481d),
	.w4(32'h38b0cb82),
	.w5(32'h383e2501),
	.w6(32'hbb92ff48),
	.w7(32'h3c3cf893),
	.w8(32'hbb88ce4e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86146a),
	.w1(32'hbbaac793),
	.w2(32'hbb23db08),
	.w3(32'h3ae09aa4),
	.w4(32'h3b8ac53f),
	.w5(32'hbb07bf5b),
	.w6(32'hbc5d653b),
	.w7(32'hbb56d96e),
	.w8(32'hba8f07cd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6094a6),
	.w1(32'hbbd4814b),
	.w2(32'hbb9efc47),
	.w3(32'hbac700f1),
	.w4(32'h3a95eee7),
	.w5(32'hbb5c15f6),
	.w6(32'h3bea81fb),
	.w7(32'h3b8179d8),
	.w8(32'hbc074232),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4280d),
	.w1(32'hbb4737d2),
	.w2(32'hbc76d60e),
	.w3(32'h3b268b93),
	.w4(32'hbc2395ae),
	.w5(32'hbc15fc8e),
	.w6(32'hbc3e6849),
	.w7(32'hbbe000d2),
	.w8(32'hba608766),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99d54f),
	.w1(32'h3c658278),
	.w2(32'h3b9a02bc),
	.w3(32'hba86f3b8),
	.w4(32'hbb70b3b0),
	.w5(32'h3be1305d),
	.w6(32'hbb26523a),
	.w7(32'h3b69c454),
	.w8(32'h3c50ab60),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0b657),
	.w1(32'h3b521281),
	.w2(32'hbb400066),
	.w3(32'h3b464737),
	.w4(32'h3ba208b7),
	.w5(32'hbd1d715e),
	.w6(32'hbc1472a6),
	.w7(32'hb7e9b937),
	.w8(32'hbd391de8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6e4cd),
	.w1(32'h3cf6ec9b),
	.w2(32'h3c998855),
	.w3(32'hbc8aed54),
	.w4(32'h3ae297ae),
	.w5(32'h3c035f50),
	.w6(32'h3c3aa594),
	.w7(32'h3cec14f1),
	.w8(32'h3ba045e3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98327d7),
	.w1(32'hbaf12890),
	.w2(32'hbb966d01),
	.w3(32'h3acd3a71),
	.w4(32'hb997c400),
	.w5(32'hbaccb926),
	.w6(32'h3cc4a68b),
	.w7(32'hbad5b305),
	.w8(32'h39c158ac),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e64c1),
	.w1(32'hb961d53a),
	.w2(32'h3b591ad3),
	.w3(32'h3b2526b7),
	.w4(32'h3b4d6ceb),
	.w5(32'h3b61851b),
	.w6(32'hbb1acd76),
	.w7(32'h3b56bc98),
	.w8(32'h3b6c4d4e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6d18a),
	.w1(32'h3b40fa12),
	.w2(32'hba807a2b),
	.w3(32'h3b55ab4d),
	.w4(32'h39e732e9),
	.w5(32'h3c3b40fc),
	.w6(32'hba1c7e5c),
	.w7(32'hb8bde0fd),
	.w8(32'h3c98b532),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b579e9e),
	.w1(32'hbc54c2db),
	.w2(32'hbca1de83),
	.w3(32'h3c87ce5f),
	.w4(32'h3a5ee427),
	.w5(32'hbca5d0df),
	.w6(32'h3c04a5d5),
	.w7(32'hbc40f98e),
	.w8(32'hbcd755f7),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28a9a3),
	.w1(32'h3c459174),
	.w2(32'h3cd0f226),
	.w3(32'hbccdad86),
	.w4(32'hbbd48c0b),
	.w5(32'hbb17405c),
	.w6(32'hbcd97b98),
	.w7(32'h3cbf7bcc),
	.w8(32'hbaed4746),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7b412),
	.w1(32'h3a233c1c),
	.w2(32'h3b5230fd),
	.w3(32'hbaba6538),
	.w4(32'h3b8d817c),
	.w5(32'hbb658d70),
	.w6(32'hbb5a48d5),
	.w7(32'h3c0af3bf),
	.w8(32'hbbf1c222),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c23d),
	.w1(32'h3c3a1b35),
	.w2(32'h3c38d347),
	.w3(32'hbb55544e),
	.w4(32'h3b4d6d0f),
	.w5(32'h3c37ec04),
	.w6(32'h3aad3a41),
	.w7(32'h3c0d983a),
	.w8(32'h3c63d31b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839d0e),
	.w1(32'hbc878c78),
	.w2(32'hbc946bbe),
	.w3(32'h3c83611d),
	.w4(32'hbabe9fa6),
	.w5(32'h3c3b942b),
	.w6(32'h3bf7cc20),
	.w7(32'hbc8b72bf),
	.w8(32'h3cb77d53),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf004e4),
	.w1(32'hbbd2e5da),
	.w2(32'hbc1138ab),
	.w3(32'h3c031775),
	.w4(32'hba210694),
	.w5(32'h3b2a47bc),
	.w6(32'hbb03bfb4),
	.w7(32'hbc04682d),
	.w8(32'h3b46f852),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98f5b5),
	.w1(32'h3ae58fea),
	.w2(32'h3a864208),
	.w3(32'h39bbcf1c),
	.w4(32'h3b8cbca8),
	.w5(32'h3c1f1732),
	.w6(32'h3ae3d852),
	.w7(32'h3a56feaa),
	.w8(32'hbc3f863c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1abb6a),
	.w1(32'h399e49a1),
	.w2(32'hbb67793f),
	.w3(32'hbcbb7bd9),
	.w4(32'hbb45ea90),
	.w5(32'hbb082992),
	.w6(32'hbc115f88),
	.w7(32'hbbdc9f5c),
	.w8(32'h3bcd2f60),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4988),
	.w1(32'h3c14a29f),
	.w2(32'h3ba9e42c),
	.w3(32'hbb96fd96),
	.w4(32'h3b99d1c0),
	.w5(32'h3b0eb153),
	.w6(32'hbadee6d9),
	.w7(32'h3c029d35),
	.w8(32'h3ad41920),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0255b6),
	.w1(32'hba10be58),
	.w2(32'h3a26763e),
	.w3(32'hbb9f386d),
	.w4(32'hba78dab7),
	.w5(32'hbb1e26db),
	.w6(32'h3bc584a8),
	.w7(32'hb94fc658),
	.w8(32'hbc0127fe),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08c87e),
	.w1(32'hbc05b86e),
	.w2(32'hbc0b3020),
	.w3(32'h3b2b9e58),
	.w4(32'hbba0aeba),
	.w5(32'h3b03382b),
	.w6(32'h3c214918),
	.w7(32'hbc69b329),
	.w8(32'h3bd89288),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc251ea),
	.w1(32'hbad817be),
	.w2(32'h3bf3bdf2),
	.w3(32'hbaba5ce7),
	.w4(32'h3c046b0d),
	.w5(32'hbb1024fe),
	.w6(32'hbba40d28),
	.w7(32'h3aebd9a9),
	.w8(32'hbb99b075),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a11f3),
	.w1(32'hbaf97b5f),
	.w2(32'h3b8faebf),
	.w3(32'hbb040ae5),
	.w4(32'h3a1400ec),
	.w5(32'h3bf0061e),
	.w6(32'hbaf8e019),
	.w7(32'h3bb88b2e),
	.w8(32'h3ad0d147),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6287fc),
	.w1(32'hbc52b497),
	.w2(32'hbc08f8fe),
	.w3(32'h3b6c525f),
	.w4(32'hb86f7032),
	.w5(32'h3a1ee7e3),
	.w6(32'h3b3f4ce0),
	.w7(32'hbc06585d),
	.w8(32'h3a63a7d2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3634ae),
	.w1(32'hbc2e529c),
	.w2(32'h3bd3ad6f),
	.w3(32'hbbeede8f),
	.w4(32'hbabbaceb),
	.w5(32'h3bb7b172),
	.w6(32'hbc50a868),
	.w7(32'h3a12a5d1),
	.w8(32'h3ba9779a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a020b30),
	.w1(32'hba52ec8f),
	.w2(32'hbbc53a00),
	.w3(32'h3b14aad1),
	.w4(32'h3b5feb52),
	.w5(32'hbb9101cf),
	.w6(32'h3afe7e2a),
	.w7(32'hbb84d901),
	.w8(32'h3aecab0c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c852466),
	.w1(32'h3c4eebeb),
	.w2(32'h3b874bbf),
	.w3(32'hbc79b437),
	.w4(32'hbbe2f562),
	.w5(32'h3bd9054e),
	.w6(32'hbc6f6d8d),
	.w7(32'h3c43e339),
	.w8(32'h3c08400d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9e798),
	.w1(32'hbb5b5f3e),
	.w2(32'hbb2f6a9f),
	.w3(32'h3bd92e00),
	.w4(32'h3b859078),
	.w5(32'hbb447933),
	.w6(32'h3b780932),
	.w7(32'hbb3728f2),
	.w8(32'h3c2d998e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a167656),
	.w1(32'hbb8d6d42),
	.w2(32'hba34fef6),
	.w3(32'h3b0c1994),
	.w4(32'h3b8f096b),
	.w5(32'h3c88feba),
	.w6(32'h392e2cb8),
	.w7(32'h3b471618),
	.w8(32'hbbb85605),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2432f2),
	.w1(32'hbb489800),
	.w2(32'hbaef137c),
	.w3(32'h3c0213e5),
	.w4(32'h3b83aff3),
	.w5(32'h3b04cff8),
	.w6(32'hbbfdf2dc),
	.w7(32'hba9fccdb),
	.w8(32'hb995927d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36762c),
	.w1(32'hbb1df095),
	.w2(32'hbbddaac5),
	.w3(32'h3a842d28),
	.w4(32'h3a0aeff8),
	.w5(32'hba8ad0bb),
	.w6(32'h3b9b4a43),
	.w7(32'hbc0f4b20),
	.w8(32'hbac200f4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd07bf7),
	.w1(32'h3b5f23fa),
	.w2(32'h3a954447),
	.w3(32'hbad79a74),
	.w4(32'h3be2e5c6),
	.w5(32'h3b206cd5),
	.w6(32'hbbb0744c),
	.w7(32'hbaf19a0f),
	.w8(32'hbb3d2205),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96adfc),
	.w1(32'h3bbce3c0),
	.w2(32'h3b788fb3),
	.w3(32'hb9b64daa),
	.w4(32'h3a991659),
	.w5(32'hbb5e5f21),
	.w6(32'h3b298c12),
	.w7(32'hbb728429),
	.w8(32'h3aedd5e3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5550),
	.w1(32'hbc4fd2e0),
	.w2(32'h3aec20c9),
	.w3(32'hbb225136),
	.w4(32'hbbe6937f),
	.w5(32'h3c49e407),
	.w6(32'hbc116ecf),
	.w7(32'hbbb01851),
	.w8(32'h3c6a0219),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be87f24),
	.w1(32'hbca05bca),
	.w2(32'hbca126da),
	.w3(32'h3c920431),
	.w4(32'hbb37294d),
	.w5(32'h3b4ac406),
	.w6(32'h3c226533),
	.w7(32'hbc9b55c6),
	.w8(32'hbbc8e33f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fb144),
	.w1(32'hbb48dada),
	.w2(32'hbb933e91),
	.w3(32'hbc6f26e3),
	.w4(32'hba8c5413),
	.w5(32'h3c088b2f),
	.w6(32'hbc0277fa),
	.w7(32'h3b504a37),
	.w8(32'h3c8a3b7a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e4cf0),
	.w1(32'hbb56c15a),
	.w2(32'hbbe67f7f),
	.w3(32'h3b42de67),
	.w4(32'hbb8891a2),
	.w5(32'h3b030507),
	.w6(32'hbc824edc),
	.w7(32'hbc12b26f),
	.w8(32'hbb3a8b40),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2b9c3),
	.w1(32'h3b6e1bb4),
	.w2(32'hbb75911f),
	.w3(32'h3a76da62),
	.w4(32'h38f52235),
	.w5(32'h3b9322f6),
	.w6(32'hbac4b269),
	.w7(32'hbbdc9d86),
	.w8(32'hbc1e1025),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf3e29),
	.w1(32'hbb2b7a75),
	.w2(32'h3b9e97c9),
	.w3(32'h3c068bbf),
	.w4(32'h3bcdc6c5),
	.w5(32'hbb397adf),
	.w6(32'h3c365cd2),
	.w7(32'hbb019114),
	.w8(32'h3c398c88),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4229e3),
	.w1(32'hbb96d607),
	.w2(32'hbba02738),
	.w3(32'h3b04915f),
	.w4(32'h3b957cbc),
	.w5(32'hbb2398c1),
	.w6(32'hbadecd45),
	.w7(32'hbc47c46c),
	.w8(32'hbb11d94e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad04bf),
	.w1(32'h3b844d8f),
	.w2(32'h3b82d819),
	.w3(32'h3c058d4a),
	.w4(32'hbabac915),
	.w5(32'h3c0d5af4),
	.w6(32'h3b86eaf7),
	.w7(32'h3bb04611),
	.w8(32'h3c10f656),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13dd03),
	.w1(32'hbc87fe33),
	.w2(32'hbbfd0d44),
	.w3(32'hbb670257),
	.w4(32'hbc4d5045),
	.w5(32'h3be78967),
	.w6(32'hbc90b6c0),
	.w7(32'hbc293fda),
	.w8(32'h3bb890f6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d42a6),
	.w1(32'h39cc31cd),
	.w2(32'hbbe268c6),
	.w3(32'hb991d6db),
	.w4(32'hba93739b),
	.w5(32'h3b519137),
	.w6(32'h3b9e1e33),
	.w7(32'h3b45078e),
	.w8(32'h398ae562),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7475c9),
	.w1(32'hbba338ae),
	.w2(32'hbc0ca2fc),
	.w3(32'h378ebb11),
	.w4(32'h3a0acaee),
	.w5(32'hbbff7f07),
	.w6(32'h3cbb50ba),
	.w7(32'hbaa4df5d),
	.w8(32'hbac51875),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e303b),
	.w1(32'h3b4e2152),
	.w2(32'h3c8613e6),
	.w3(32'hbc71e3a4),
	.w4(32'h3b5ba4fe),
	.w5(32'hbce3b31e),
	.w6(32'hbc30daef),
	.w7(32'h3cce1d4f),
	.w8(32'hbcc7d62b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40751),
	.w1(32'h3c89b1d3),
	.w2(32'h3c35fc00),
	.w3(32'hbcaabcfb),
	.w4(32'h3abacdab),
	.w5(32'hba2ec175),
	.w6(32'h3c26fc28),
	.w7(32'h3ccf51ff),
	.w8(32'h3bd9817d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02580e),
	.w1(32'hbcbc6053),
	.w2(32'hbcb53196),
	.w3(32'h3bc03197),
	.w4(32'hbba024b6),
	.w5(32'h3aef277a),
	.w6(32'hbbf0d108),
	.w7(32'hbc8c11f2),
	.w8(32'hbc52926c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7325a),
	.w1(32'h3c77e0fc),
	.w2(32'hbb2c89a9),
	.w3(32'h3b4702c1),
	.w4(32'hba251b9b),
	.w5(32'hbb8b045d),
	.w6(32'h3c9cb99e),
	.w7(32'h3ba18511),
	.w8(32'hbb1eb8ea),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9f8ff),
	.w1(32'h3b2ebde7),
	.w2(32'h3938f9e1),
	.w3(32'h3bcee7be),
	.w4(32'hb9fe7ffc),
	.w5(32'hbb538d56),
	.w6(32'h3ab9597a),
	.w7(32'h3b5ac335),
	.w8(32'hbc17bed9),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb752e84),
	.w1(32'h3b41f5d1),
	.w2(32'hbbfd0f43),
	.w3(32'hbc2268a8),
	.w4(32'hbbf92a2d),
	.w5(32'hbb4c4642),
	.w6(32'h3c9b430c),
	.w7(32'hba91f806),
	.w8(32'hbb951d43),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6266d),
	.w1(32'hbb74e15d),
	.w2(32'h3c3703e5),
	.w3(32'hbba21242),
	.w4(32'hbba40868),
	.w5(32'h3ad414bb),
	.w6(32'hbc0808a6),
	.w7(32'h3b215e88),
	.w8(32'h3aedaefa),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065ca3),
	.w1(32'h3b9a1b41),
	.w2(32'hbc01bf97),
	.w3(32'h3b2deeed),
	.w4(32'hb90100fa),
	.w5(32'h3b76f5d4),
	.w6(32'h3d0ddcc6),
	.w7(32'h3ba5e940),
	.w8(32'h3a21ee5e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39757851),
	.w1(32'h3b8050a3),
	.w2(32'h3bcf7109),
	.w3(32'h3b869c8b),
	.w4(32'h39cdd0e2),
	.w5(32'h3bf0ff50),
	.w6(32'hbb9d67d8),
	.w7(32'h3b867e6f),
	.w8(32'hbb5eebac),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b61c6d),
	.w1(32'hbb670091),
	.w2(32'h3a77673b),
	.w3(32'h3ba31779),
	.w4(32'hbbb157da),
	.w5(32'hbb40fb94),
	.w6(32'hbaa865b9),
	.w7(32'h3a84fa54),
	.w8(32'h3a71e18b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89da7),
	.w1(32'hbc0fb3f9),
	.w2(32'hbb9b20ca),
	.w3(32'h3b658916),
	.w4(32'hba9d2197),
	.w5(32'hbb216e8c),
	.w6(32'hbaa86c34),
	.w7(32'hbc08bf6e),
	.w8(32'h3b09de2e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49e6ff),
	.w1(32'hbbca4cba),
	.w2(32'hbc1ab7af),
	.w3(32'h3c16ebe5),
	.w4(32'hba00beab),
	.w5(32'hbae34712),
	.w6(32'h3bd1e5bb),
	.w7(32'hbbe02b46),
	.w8(32'hbb0c4639),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58cc52),
	.w1(32'h396e7ce2),
	.w2(32'h3be1760e),
	.w3(32'hbb1340ea),
	.w4(32'hbae9b463),
	.w5(32'hb7e33fe5),
	.w6(32'h3b8cedd9),
	.w7(32'h3c1c7683),
	.w8(32'hb8a68780),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ddc9),
	.w1(32'h3c26df8b),
	.w2(32'h3aab0d03),
	.w3(32'hb9b70c23),
	.w4(32'h3befa75c),
	.w5(32'hbc1fcfe6),
	.w6(32'h3a878772),
	.w7(32'h3af54529),
	.w8(32'hbc147e29),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3bbf7),
	.w1(32'hbb188a37),
	.w2(32'hbb475468),
	.w3(32'h3af3c236),
	.w4(32'hbb84a5eb),
	.w5(32'h3b7dfb44),
	.w6(32'h3c3a90dc),
	.w7(32'hb9b7d94d),
	.w8(32'hba613126),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57d3c),
	.w1(32'hbb9bbb4d),
	.w2(32'hbb93ade9),
	.w3(32'h3b2b1b9a),
	.w4(32'hbb9a83aa),
	.w5(32'hbc16d8de),
	.w6(32'hbc31aaef),
	.w7(32'hbc19342f),
	.w8(32'hbba73416),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba25395),
	.w1(32'hbbaf0d14),
	.w2(32'h3b5e27d6),
	.w3(32'h3b2a65d8),
	.w4(32'h3afe7899),
	.w5(32'h3b0536b1),
	.w6(32'h3b197518),
	.w7(32'h3b02e1ed),
	.w8(32'h39975779),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb988dab),
	.w1(32'h3965c2ed),
	.w2(32'h3bb17188),
	.w3(32'hba9a8519),
	.w4(32'hb92f419d),
	.w5(32'h3baa6108),
	.w6(32'hbb58ac61),
	.w7(32'h3bc249f9),
	.w8(32'hbbb92b17),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b804c6b),
	.w1(32'h3c611da9),
	.w2(32'h3c248fad),
	.w3(32'hbc5d9b33),
	.w4(32'hbba8a9af),
	.w5(32'hbd1c0258),
	.w6(32'hbc88a322),
	.w7(32'h3bc56745),
	.w8(32'hbd08e250),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944ff51),
	.w1(32'h3d214fd3),
	.w2(32'h3cdcb94b),
	.w3(32'hbd0ebb9e),
	.w4(32'h3b4beff2),
	.w5(32'h3bbf67b9),
	.w6(32'h3c037c00),
	.w7(32'h3d33e81f),
	.w8(32'hbc2599e2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08380),
	.w1(32'hbab16322),
	.w2(32'hbc141859),
	.w3(32'hbb5520f2),
	.w4(32'hbba4d25d),
	.w5(32'h3ace2319),
	.w6(32'h3c50778d),
	.w7(32'hbb3ea8e1),
	.w8(32'h3aea9e17),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952bd61),
	.w1(32'hbb3782cd),
	.w2(32'hbb9d5cbb),
	.w3(32'h3aff0574),
	.w4(32'hba2939da),
	.w5(32'hbadae818),
	.w6(32'h3b29d9a5),
	.w7(32'h3aa534ca),
	.w8(32'hbb11e9c4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f732a),
	.w1(32'hbbab9f52),
	.w2(32'hbc32e4b5),
	.w3(32'h3b7a07d3),
	.w4(32'hbb56b60c),
	.w5(32'hbbcccdad),
	.w6(32'h3b4fc249),
	.w7(32'hb993c20c),
	.w8(32'hbbdda4e8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a035151),
	.w1(32'h3b829eed),
	.w2(32'hb8b0ace4),
	.w3(32'hbae934c7),
	.w4(32'h3ad1cf4a),
	.w5(32'hbb2be7bb),
	.w6(32'hb9b7b393),
	.w7(32'h3bb1962e),
	.w8(32'h3ab6700c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996505d),
	.w1(32'h3aa5c48a),
	.w2(32'h3a2697b7),
	.w3(32'hba928589),
	.w4(32'h3a215772),
	.w5(32'hba805bcf),
	.w6(32'hbb1999a5),
	.w7(32'h372a9d0e),
	.w8(32'hbb40991a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf31e1),
	.w1(32'hbb8ff835),
	.w2(32'hbc09be99),
	.w3(32'h3b8a7cee),
	.w4(32'hbb4d5c0f),
	.w5(32'hbbc55e65),
	.w6(32'h3b74bd2f),
	.w7(32'hbafadb56),
	.w8(32'hbb9772de),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a473e),
	.w1(32'h38a06f65),
	.w2(32'h3768c226),
	.w3(32'h37743755),
	.w4(32'hb89d9e4e),
	.w5(32'h37d05137),
	.w6(32'hb859d702),
	.w7(32'hb86719fb),
	.w8(32'h36bf2963),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8260cb),
	.w1(32'hbb4d060e),
	.w2(32'hbc06004e),
	.w3(32'h3b2de965),
	.w4(32'hbb93afc6),
	.w5(32'hbbd7563a),
	.w6(32'h3b1a6f16),
	.w7(32'hba0f046e),
	.w8(32'hbb9ecf92),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5f3c1),
	.w1(32'hb9834762),
	.w2(32'hbba1c448),
	.w3(32'h3a34f00c),
	.w4(32'hbaf499f3),
	.w5(32'hbb51e2c2),
	.w6(32'h3b475edb),
	.w7(32'h3a7c9424),
	.w8(32'hbb23cc9a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f836e2),
	.w1(32'h38a152a1),
	.w2(32'h3910691e),
	.w3(32'hb974da78),
	.w4(32'h38414cd2),
	.w5(32'h38b2c1f7),
	.w6(32'hb943dea3),
	.w7(32'h391772b9),
	.w8(32'h3930151d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73cf02),
	.w1(32'hbafc6637),
	.w2(32'hba4b9f5c),
	.w3(32'hbac86e51),
	.w4(32'hbaec196c),
	.w5(32'hbaa7f897),
	.w6(32'hba4c172e),
	.w7(32'h39d02dcf),
	.w8(32'hba0ae46d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7db4f),
	.w1(32'hbb1ee9a8),
	.w2(32'hba3b9a93),
	.w3(32'h39b906c6),
	.w4(32'hba20b3c6),
	.w5(32'h3a6044eb),
	.w6(32'h3afd4b27),
	.w7(32'h3a7071b9),
	.w8(32'h3a8b3df5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38941844),
	.w1(32'h3a950946),
	.w2(32'h398eecf9),
	.w3(32'hba0b69b0),
	.w4(32'h3a4da972),
	.w5(32'hba609068),
	.w6(32'hbab105cd),
	.w7(32'h3a47b8d3),
	.w8(32'hbab5086d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8236c0d),
	.w1(32'h3ad2ac2d),
	.w2(32'h3af4ea54),
	.w3(32'hbaef9f6d),
	.w4(32'h38adb5af),
	.w5(32'h370cea7e),
	.w6(32'hbab6f5a9),
	.w7(32'h3aa8a3da),
	.w8(32'h3a5412c2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2b5c9),
	.w1(32'h3a84aed5),
	.w2(32'h39e76251),
	.w3(32'h39d6862c),
	.w4(32'h399585d8),
	.w5(32'hba8a0b01),
	.w6(32'hbad32eaa),
	.w7(32'hba74ad99),
	.w8(32'hbad1ff77),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b805ebb),
	.w1(32'h3a8f02a1),
	.w2(32'hb9869e24),
	.w3(32'h3b903701),
	.w4(32'h3b033a07),
	.w5(32'h39cda3ab),
	.w6(32'h3b91a5bc),
	.w7(32'h3b6cde36),
	.w8(32'h3b14e9c7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c5d7),
	.w1(32'hbbc59af3),
	.w2(32'hbb371158),
	.w3(32'hbb590083),
	.w4(32'hbb0e8f3e),
	.w5(32'h39c576c5),
	.w6(32'hbb528f87),
	.w7(32'hbabfe086),
	.w8(32'hb93268dd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5423f8),
	.w1(32'h3a067b05),
	.w2(32'h39b97a78),
	.w3(32'h39d88d91),
	.w4(32'h3a05b4a5),
	.w5(32'hb8f97fb4),
	.w6(32'h38005c8e),
	.w7(32'h39b84ad7),
	.w8(32'hba199ea4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e67b2),
	.w1(32'hb769a79c),
	.w2(32'hb87c044b),
	.w3(32'hb7d2688c),
	.w4(32'h36f45915),
	.w5(32'hb862eb4e),
	.w6(32'hb8b4a416),
	.w7(32'hb81bfeb4),
	.w8(32'hb832c73f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e9d5e),
	.w1(32'hba44b04b),
	.w2(32'hb90fa92e),
	.w3(32'hb9ed6cf1),
	.w4(32'hba27dc72),
	.w5(32'hb9e581c4),
	.w6(32'hba6e3772),
	.w7(32'hba753270),
	.w8(32'hba08df8e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dac46e),
	.w1(32'h3883828a),
	.w2(32'hb708b6d2),
	.w3(32'h369f953f),
	.w4(32'h37ead056),
	.w5(32'h3673ae69),
	.w6(32'h374505b9),
	.w7(32'h370523ee),
	.w8(32'hb715bc8f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361e596d),
	.w1(32'hb8d46a7d),
	.w2(32'hb850fc42),
	.w3(32'hb88c2bb0),
	.w4(32'hb8612936),
	.w5(32'h37db5c90),
	.w6(32'hb8ca5874),
	.w7(32'hb8b17a52),
	.w8(32'h38412ab2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e24fb),
	.w1(32'h3a026bad),
	.w2(32'h37ba372d),
	.w3(32'h3a011876),
	.w4(32'h3a837671),
	.w5(32'h383ada53),
	.w6(32'h38fabbb1),
	.w7(32'h3a625522),
	.w8(32'hba4fdab2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bde49),
	.w1(32'h391eb570),
	.w2(32'h3919239c),
	.w3(32'h387e57fa),
	.w4(32'hb7312538),
	.w5(32'h3913da31),
	.w6(32'h3898a5bc),
	.w7(32'h38cee8bd),
	.w8(32'h39385655),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a524c46),
	.w1(32'hba706b55),
	.w2(32'hbafac527),
	.w3(32'h3a340c24),
	.w4(32'hb9e5f950),
	.w5(32'hb9ab8317),
	.w6(32'h3ac9e69b),
	.w7(32'h3925ebd7),
	.w8(32'h39f53bfd),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a1b6),
	.w1(32'h3a82744b),
	.w2(32'h3b0cb16d),
	.w3(32'hbb5c33d3),
	.w4(32'hba601b0f),
	.w5(32'hbb07f34d),
	.w6(32'hbb87cf74),
	.w7(32'hba573435),
	.w8(32'hbae3127d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813ffc1),
	.w1(32'hb6378e44),
	.w2(32'h383e99cc),
	.w3(32'h37c6c484),
	.w4(32'hb72c20aa),
	.w5(32'hb8200f1a),
	.w6(32'hb7105e14),
	.w7(32'hb7f0fce6),
	.w8(32'hb86c0db9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728b3a1),
	.w1(32'h3798fc8b),
	.w2(32'hb78d7361),
	.w3(32'hb82dbc33),
	.w4(32'hb7cb4f9a),
	.w5(32'hb898a627),
	.w6(32'hb83129c7),
	.w7(32'hb5d743ff),
	.w8(32'hb6a3f8bc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35bc1980),
	.w1(32'h36aad795),
	.w2(32'h37479256),
	.w3(32'h3673bb12),
	.w4(32'h37a639b1),
	.w5(32'h37139f13),
	.w6(32'h35e22aa3),
	.w7(32'h3694e50a),
	.w8(32'h36accf5f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913095f),
	.w1(32'hb92586c5),
	.w2(32'hb7cd89ef),
	.w3(32'h39791088),
	.w4(32'hb96bbfb9),
	.w5(32'hb9005b48),
	.w6(32'h38dfc324),
	.w7(32'hb99b5b05),
	.w8(32'hb9bd4c32),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84ea6c),
	.w1(32'hbbfc13b9),
	.w2(32'hbb664bb3),
	.w3(32'h3b355f59),
	.w4(32'hb930e766),
	.w5(32'h3aa310fb),
	.w6(32'h3c14c709),
	.w7(32'h3b6a971a),
	.w8(32'h3b693a87),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb345e65),
	.w1(32'hbb81695e),
	.w2(32'hbadaf53f),
	.w3(32'h3a933309),
	.w4(32'h3a3c0675),
	.w5(32'h3aecc9e8),
	.w6(32'h3b2d525b),
	.w7(32'h3a12fc8b),
	.w8(32'h3af500a6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b7a715),
	.w1(32'hba1a48c1),
	.w2(32'hb9c04690),
	.w3(32'h391fd105),
	.w4(32'hb9de8168),
	.w5(32'hb9f62713),
	.w6(32'h390c67c1),
	.w7(32'hb948816e),
	.w8(32'h37c9e75e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba084eab),
	.w1(32'hba1064b2),
	.w2(32'h399d042b),
	.w3(32'h383bdd3a),
	.w4(32'hb92d996f),
	.w5(32'h3a1c25fb),
	.w6(32'hb880baf4),
	.w7(32'hba2d87f6),
	.w8(32'hb910ccf1),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397108d3),
	.w1(32'h39ba42b6),
	.w2(32'h3794fa97),
	.w3(32'hb7f17478),
	.w4(32'h3959b285),
	.w5(32'hba221635),
	.w6(32'hba21f3b0),
	.w7(32'h38697c6a),
	.w8(32'hba1d7e93),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d520e),
	.w1(32'hba7f3a1f),
	.w2(32'hb9e11251),
	.w3(32'hb9aaf7b4),
	.w4(32'h3a5fa0ee),
	.w5(32'h3a3f9cde),
	.w6(32'hb9fe3411),
	.w7(32'hb9871e9b),
	.w8(32'h39b9c6c6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c6122),
	.w1(32'hbb1d5aec),
	.w2(32'hba31a468),
	.w3(32'hbb33f93d),
	.w4(32'hbada6fc1),
	.w5(32'hbb1a48fa),
	.w6(32'hbb4d0183),
	.w7(32'hba842206),
	.w8(32'hbb12c527),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb110eb1),
	.w1(32'hbbbd3c61),
	.w2(32'hbb9d2579),
	.w3(32'h3b1562cf),
	.w4(32'hb8b9e604),
	.w5(32'h393491db),
	.w6(32'h3af39f6f),
	.w7(32'h3994da6c),
	.w8(32'h3ad056b4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0589e4),
	.w1(32'h3ab80df5),
	.w2(32'h3a6aec85),
	.w3(32'hb9ed99f5),
	.w4(32'h392334c1),
	.w5(32'hba783685),
	.w6(32'hba7b7a88),
	.w7(32'h3a1fd04e),
	.w8(32'hba003aa2),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e065b9),
	.w1(32'hbb04e0a3),
	.w2(32'hbb206d57),
	.w3(32'h3a7d9e8a),
	.w4(32'hba1900eb),
	.w5(32'hba972599),
	.w6(32'h3a324d47),
	.w7(32'hb9730092),
	.w8(32'hba8d8548),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c39c),
	.w1(32'hbb46a15d),
	.w2(32'hbb8ceb97),
	.w3(32'h3b287e3f),
	.w4(32'hba3c0ae0),
	.w5(32'hb8ed4e97),
	.w6(32'h3b2b2ac1),
	.w7(32'hba05b1e1),
	.w8(32'h3ac7a7df),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16cfad),
	.w1(32'h3aaee812),
	.w2(32'h3ac69e67),
	.w3(32'h3ae0a4b5),
	.w4(32'h3a1b7153),
	.w5(32'h3a5aece7),
	.w6(32'h3a4955aa),
	.w7(32'h33ffa820),
	.w8(32'hba9f06db),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8701f75),
	.w1(32'hbb18b0c0),
	.w2(32'hbb22cae0),
	.w3(32'h3a34b11c),
	.w4(32'hba01c401),
	.w5(32'hb7c4a885),
	.w6(32'h3a9a4d53),
	.w7(32'h3894e6b7),
	.w8(32'hb9361c6c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9053368),
	.w1(32'hb732d90c),
	.w2(32'hb8337089),
	.w3(32'h38ac8f74),
	.w4(32'h39171533),
	.w5(32'hb83ee633),
	.w6(32'hb7186233),
	.w7(32'h395ed224),
	.w8(32'hb90c494a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d8a12),
	.w1(32'h3b8af40c),
	.w2(32'h3bc69222),
	.w3(32'hbba606c6),
	.w4(32'hbaa3f0b6),
	.w5(32'hbacc37c5),
	.w6(32'hbbb8aff1),
	.w7(32'h3a90bcbe),
	.w8(32'h3aa76cd4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84e3a7),
	.w1(32'h3a9cd5c5),
	.w2(32'h3a2046eb),
	.w3(32'h39c7d5af),
	.w4(32'h3a1c0264),
	.w5(32'h3992033a),
	.w6(32'h39a8771f),
	.w7(32'h397aef91),
	.w8(32'h39dee6c8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900fdeb),
	.w1(32'hb8ae63c7),
	.w2(32'hb7eba0af),
	.w3(32'hb8b960be),
	.w4(32'hb93eb5d9),
	.w5(32'hb91fbb29),
	.w6(32'hb906ed97),
	.w7(32'hb91ad62b),
	.w8(32'hb8976105),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8369336),
	.w1(32'h37d19462),
	.w2(32'h388a35de),
	.w3(32'hb703843f),
	.w4(32'h384c0947),
	.w5(32'h389e2ceb),
	.w6(32'hb7c2ec2b),
	.w7(32'hb7a58d88),
	.w8(32'hb70f623d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370af066),
	.w1(32'h382af567),
	.w2(32'h38dd2659),
	.w3(32'hb9ef5667),
	.w4(32'hb93edc80),
	.w5(32'h35a7c794),
	.w6(32'hb8ccfa7f),
	.w7(32'h391966d2),
	.w8(32'hb9f90dd1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b376465),
	.w1(32'h3b13ca8c),
	.w2(32'h3ab80452),
	.w3(32'h3ac3277a),
	.w4(32'h3a9b48b6),
	.w5(32'hb9535d6c),
	.w6(32'h3a777aaf),
	.w7(32'h3a907e06),
	.w8(32'hba27d7e2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad102a3),
	.w1(32'hbade4cba),
	.w2(32'hba11542f),
	.w3(32'h37caa984),
	.w4(32'h3a21d106),
	.w5(32'h3a52c77c),
	.w6(32'h3a1dd585),
	.w7(32'h3ac9b7e3),
	.w8(32'h3a8de6dc),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83470bd),
	.w1(32'h37430da9),
	.w2(32'h386456f0),
	.w3(32'hb7e711c7),
	.w4(32'h386bdde0),
	.w5(32'h38321245),
	.w6(32'hb7fa6312),
	.w7(32'h386cd988),
	.w8(32'h3849d849),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bbdb8),
	.w1(32'hbb27545b),
	.w2(32'hbae75c1b),
	.w3(32'hba07d8a6),
	.w4(32'hba1e4f3c),
	.w5(32'h39360abb),
	.w6(32'h3a91f4ea),
	.w7(32'h3994cbac),
	.w8(32'h3a27bbfd),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a5241),
	.w1(32'hb80dc1b4),
	.w2(32'hb707f508),
	.w3(32'h3a35f117),
	.w4(32'h39cc79fd),
	.w5(32'h38bd137d),
	.w6(32'h3a5f0f66),
	.w7(32'h3a41787c),
	.w8(32'hb9ae2787),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05d1f5),
	.w1(32'hbb82506a),
	.w2(32'hbb410a1a),
	.w3(32'h3b13403f),
	.w4(32'hbaeaf023),
	.w5(32'hbabdee27),
	.w6(32'h3b08cfca),
	.w7(32'h393fdd1c),
	.w8(32'h3a493cb5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e02f),
	.w1(32'h3af640cf),
	.w2(32'h3b9799e2),
	.w3(32'hbb67e19b),
	.w4(32'h3abc234d),
	.w5(32'h3afece86),
	.w6(32'hbb82f2f7),
	.w7(32'h3af46abf),
	.w8(32'h3a56e427),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dba7ea),
	.w1(32'hba96570c),
	.w2(32'hba68d13c),
	.w3(32'hba8c7529),
	.w4(32'hbad6b098),
	.w5(32'hbaef7d4a),
	.w6(32'hba467073),
	.w7(32'hba80631c),
	.w8(32'hbaaef380),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a410a),
	.w1(32'h3907d374),
	.w2(32'hb816187f),
	.w3(32'hb8077e4c),
	.w4(32'h3886bf59),
	.w5(32'hb8a2c7ed),
	.w6(32'hb9496bdc),
	.w7(32'hb8906421),
	.w8(32'hb90669a5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac36478),
	.w1(32'h3b157f26),
	.w2(32'h3ab3a6ba),
	.w3(32'h398a319a),
	.w4(32'h3aacf16a),
	.w5(32'hb984504d),
	.w6(32'hb9374d90),
	.w7(32'h3a547ec4),
	.w8(32'hba6358ca),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add1646),
	.w1(32'h3ad5ca73),
	.w2(32'h3a364e4e),
	.w3(32'h37cbd805),
	.w4(32'h39da2ad1),
	.w5(32'hbaad597e),
	.w6(32'hba2c3350),
	.w7(32'h3a75aac7),
	.w8(32'hbaa9ad0e),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba250f0c),
	.w1(32'h3aa143a2),
	.w2(32'h3a022190),
	.w3(32'hbac8991c),
	.w4(32'h39a747a8),
	.w5(32'hba1ba66a),
	.w6(32'hbaea2cff),
	.w7(32'h39a4c9c7),
	.w8(32'h38e79df0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a4cd6),
	.w1(32'hba400449),
	.w2(32'hbaa26c92),
	.w3(32'h398d61e8),
	.w4(32'hba412a79),
	.w5(32'hba5a6c33),
	.w6(32'h396c73f2),
	.w7(32'hb9093195),
	.w8(32'h39717dbc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3817acd9),
	.w1(32'hb97f7323),
	.w2(32'hb944e466),
	.w3(32'hb8bfc4fd),
	.w4(32'hba0e354b),
	.w5(32'hb9a60fb4),
	.w6(32'hb9c26563),
	.w7(32'hb9c7dece),
	.w8(32'hb9091acb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53f2b1),
	.w1(32'hbb22f0b0),
	.w2(32'hbadad1ec),
	.w3(32'h3aeae115),
	.w4(32'h38e21fae),
	.w5(32'h39844524),
	.w6(32'h3b1fbad1),
	.w7(32'h3aa0949a),
	.w8(32'h3a262f64),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38833d74),
	.w1(32'hba190b31),
	.w2(32'hba3600bd),
	.w3(32'h3a0fe202),
	.w4(32'hb9373096),
	.w5(32'hb907e856),
	.w6(32'h3acd0e77),
	.w7(32'h3a64366d),
	.w8(32'h3a301168),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cef4e),
	.w1(32'h3ab2e8bb),
	.w2(32'h3ac8046a),
	.w3(32'hba7ecc47),
	.w4(32'h3a8d6ab4),
	.w5(32'h3a41dd0b),
	.w6(32'hba7f3605),
	.w7(32'h3ab094bd),
	.w8(32'h37a3cd6f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d87c6),
	.w1(32'hb6e7cd76),
	.w2(32'h386d34f7),
	.w3(32'h38993ce2),
	.w4(32'h38bdb6a0),
	.w5(32'h378abda7),
	.w6(32'h37e9f2a9),
	.w7(32'h37ef13ab),
	.w8(32'hb7fbe4ff),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c0750),
	.w1(32'hbb12244b),
	.w2(32'hbab6c1c6),
	.w3(32'h38c3fbbe),
	.w4(32'h390db100),
	.w5(32'h39c104a6),
	.w6(32'h3abb9582),
	.w7(32'h3aa2820c),
	.w8(32'h3a461466),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ae689),
	.w1(32'h35a65453),
	.w2(32'h37e4fe79),
	.w3(32'h37c73cb2),
	.w4(32'h37ae4050),
	.w5(32'h382d03b4),
	.w6(32'h37088598),
	.w7(32'h36f1baa2),
	.w8(32'h362d8299),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880c6cf),
	.w1(32'h37759b97),
	.w2(32'h38b72aad),
	.w3(32'hb86fd268),
	.w4(32'h3794308f),
	.w5(32'h38bccef5),
	.w6(32'hb92739dc),
	.w7(32'hb8f06cff),
	.w8(32'h391ee6d9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91e101),
	.w1(32'h3abeb1f7),
	.w2(32'h3aa3e932),
	.w3(32'hb94f6151),
	.w4(32'h39fff759),
	.w5(32'hb959dd9e),
	.w6(32'hb990a545),
	.w7(32'h3a01a300),
	.w8(32'hb91fc069),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f9246),
	.w1(32'hb90eeac0),
	.w2(32'hbb445826),
	.w3(32'h3b8e218a),
	.w4(32'h3ae3c3b3),
	.w5(32'hb961ff20),
	.w6(32'h3be95494),
	.w7(32'h3b6078ba),
	.w8(32'h3a8f5955),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c659a),
	.w1(32'hb8c536ce),
	.w2(32'hb9d2410c),
	.w3(32'hba2c4220),
	.w4(32'hb9d1bfcf),
	.w5(32'hba43e0ea),
	.w6(32'hba1d9b90),
	.w7(32'hb9281be7),
	.w8(32'hba132d4e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06808e),
	.w1(32'h3a2917f8),
	.w2(32'h3a0899a7),
	.w3(32'hbabf13e5),
	.w4(32'hb8854e7b),
	.w5(32'hba87ce6d),
	.w6(32'hbacc35bc),
	.w7(32'hb8aff72d),
	.w8(32'hbaafd8e8),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0624),
	.w1(32'hba691852),
	.w2(32'hba4c3338),
	.w3(32'hbaf1f70c),
	.w4(32'hb9ad1a5c),
	.w5(32'h38270d84),
	.w6(32'hba64bf67),
	.w7(32'hb7d3afc4),
	.w8(32'h39ddbdcd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1815),
	.w1(32'hbadd86c3),
	.w2(32'hba415a03),
	.w3(32'hba4e20c1),
	.w4(32'h39c74829),
	.w5(32'h3ae30a22),
	.w6(32'h3afcf92b),
	.w7(32'h3b074043),
	.w8(32'h3b292111),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bb8fc),
	.w1(32'hbae2bb06),
	.w2(32'hbaa8d467),
	.w3(32'hb9583c6f),
	.w4(32'hb9a9e9e4),
	.w5(32'hb8b8e441),
	.w6(32'h3aa3bbee),
	.w7(32'h39c243f7),
	.w8(32'hb840b4e3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac20cb0),
	.w1(32'hbb4179eb),
	.w2(32'hbae51c92),
	.w3(32'h3a2cb876),
	.w4(32'h391b960f),
	.w5(32'h3a9607d8),
	.w6(32'h3ac7cd6a),
	.w7(32'h39b1e0a7),
	.w8(32'h3ac71b22),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b9fea),
	.w1(32'hb70f018d),
	.w2(32'h38621a09),
	.w3(32'h366f7828),
	.w4(32'h36724fe4),
	.w5(32'h37bf2122),
	.w6(32'hb61b30f5),
	.w7(32'h36c3e19a),
	.w8(32'hb75fdc37),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e5551),
	.w1(32'hbb04b513),
	.w2(32'hb9f91964),
	.w3(32'hba10ea65),
	.w4(32'hb80116dc),
	.w5(32'h39b76ed7),
	.w6(32'hba16872b),
	.w7(32'hba192dfd),
	.w8(32'hb8d85611),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cefac0),
	.w1(32'hb706c499),
	.w2(32'h375805f2),
	.w3(32'hb6d5dc3d),
	.w4(32'hb70c2a13),
	.w5(32'h384e740f),
	.w6(32'hb6d7b028),
	.w7(32'hb6519800),
	.w8(32'h37b3fac2),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e68ce1),
	.w1(32'hb826522c),
	.w2(32'hb8d14100),
	.w3(32'hb8be2497),
	.w4(32'hb9a67f75),
	.w5(32'hb9860c25),
	.w6(32'hb976e539),
	.w7(32'hba3464c3),
	.w8(32'hba39a961),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930f765),
	.w1(32'h3a0b1318),
	.w2(32'h3a1c21ca),
	.w3(32'hb9ff6b66),
	.w4(32'h39b836fc),
	.w5(32'hb90d8ced),
	.w6(32'hba4c1b5d),
	.w7(32'hb92dc59f),
	.w8(32'hb89934c0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55cd15),
	.w1(32'hbb805d93),
	.w2(32'hbaa4c3d3),
	.w3(32'hbb1553df),
	.w4(32'hba992165),
	.w5(32'h3819a4a3),
	.w6(32'hbaf45099),
	.w7(32'hb9a64f4d),
	.w8(32'h39c46b9b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7424007),
	.w1(32'h3820b2ca),
	.w2(32'hb798652e),
	.w3(32'h37d2cba2),
	.w4(32'hb77c024e),
	.w5(32'h36e99b85),
	.w6(32'h377e8e9e),
	.w7(32'hb74b60a0),
	.w8(32'h377c78d5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7593e47),
	.w1(32'h37621968),
	.w2(32'h37c402de),
	.w3(32'h36b5038c),
	.w4(32'h37de0f65),
	.w5(32'h383d1e4a),
	.w6(32'hb5e4f083),
	.w7(32'h3687645a),
	.w8(32'hb7fa08d3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2331ab),
	.w1(32'h3836f039),
	.w2(32'h3a4438ae),
	.w3(32'hba788184),
	.w4(32'hb910314d),
	.w5(32'hb9f0da81),
	.w6(32'hba46c0fd),
	.w7(32'h38f4037f),
	.w8(32'hba5a3a44),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079ce1),
	.w1(32'hbb98f18b),
	.w2(32'hbb8db96e),
	.w3(32'h3a3ba42c),
	.w4(32'hbb7ec321),
	.w5(32'hbb9a3a1a),
	.w6(32'h366fcfc7),
	.w7(32'hbb4e18c3),
	.w8(32'hbba88d94),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba471c7e),
	.w1(32'hbafb50c8),
	.w2(32'hbb9c431c),
	.w3(32'h3a9296ef),
	.w4(32'hbb78d365),
	.w5(32'hbb8fce4b),
	.w6(32'h3a8640df),
	.w7(32'h39735da1),
	.w8(32'hbb314c36),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccbfda),
	.w1(32'h389bf93e),
	.w2(32'hb661196e),
	.w3(32'h37eb1d02),
	.w4(32'h385266eb),
	.w5(32'h39334ee2),
	.w6(32'hb8551a88),
	.w7(32'h3975d50e),
	.w8(32'h3989a2ed),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8d0d8),
	.w1(32'hbb9a5719),
	.w2(32'hba9260d4),
	.w3(32'h3aedb587),
	.w4(32'h3a8e2ea5),
	.w5(32'h3bc95ed9),
	.w6(32'h3ba8a541),
	.w7(32'h3b8bd7c7),
	.w8(32'h3bbfb1d4),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf2335),
	.w1(32'h3abe366f),
	.w2(32'h3b19b878),
	.w3(32'hbb87aec2),
	.w4(32'hba1b66d0),
	.w5(32'hbad72000),
	.w6(32'hbb99a71d),
	.w7(32'h3a73d392),
	.w8(32'h37a8ad83),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81bf0ad),
	.w1(32'hbac59ed6),
	.w2(32'hbb202f1c),
	.w3(32'h3a7b1d8d),
	.w4(32'hba602e2b),
	.w5(32'hbac545f9),
	.w6(32'h3ac412d4),
	.w7(32'h3980c4c3),
	.w8(32'hba42aca6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8336cb3),
	.w1(32'hb7432cbd),
	.w2(32'hb6990a21),
	.w3(32'hb6aded73),
	.w4(32'hb5752cd6),
	.w5(32'h379ab53f),
	.w6(32'hb87c3041),
	.w7(32'hb80b0a52),
	.w8(32'h37ef9770),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374b4828),
	.w1(32'h37f1af51),
	.w2(32'hb7eebec5),
	.w3(32'h3812c9b0),
	.w4(32'h36cf9665),
	.w5(32'h37cd4963),
	.w6(32'h3748fc77),
	.w7(32'hb849a420),
	.w8(32'hb784e30b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5429f9c),
	.w1(32'hb7a8e5b4),
	.w2(32'hb74627e5),
	.w3(32'h370bb5c2),
	.w4(32'h376edd7b),
	.w5(32'h37f6148f),
	.w6(32'h37100e3f),
	.w7(32'hb7632139),
	.w8(32'hb79118b3),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab0590),
	.w1(32'hbad71456),
	.w2(32'hbb7e4146),
	.w3(32'h3aa5c8fc),
	.w4(32'hba913e5c),
	.w5(32'hbb340968),
	.w6(32'h3b244631),
	.w7(32'h3a0f6d5f),
	.w8(32'hba4fdbb3),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9bf78),
	.w1(32'h39ba0e56),
	.w2(32'hba432c95),
	.w3(32'h3af5e93e),
	.w4(32'h3aa7a979),
	.w5(32'h3839f94a),
	.w6(32'h3b013623),
	.w7(32'h3a63e48b),
	.w8(32'hb96cda6a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5004),
	.w1(32'h39fdf2af),
	.w2(32'h3a19ecbf),
	.w3(32'hba886bf6),
	.w4(32'hb9d36b8d),
	.w5(32'hbabd50e8),
	.w6(32'hbaf8c83c),
	.w7(32'hb939802a),
	.w8(32'hbb189429),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923f50e),
	.w1(32'h39c5322b),
	.w2(32'h3a162baf),
	.w3(32'hb9966cdb),
	.w4(32'h3915d543),
	.w5(32'hb6342b39),
	.w6(32'hb9b33dc2),
	.w7(32'h3810ce70),
	.w8(32'hb9331084),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a9f94),
	.w1(32'hbb28497f),
	.w2(32'hbafc5132),
	.w3(32'h3b1d2e81),
	.w4(32'h398bf784),
	.w5(32'h3a4f647f),
	.w6(32'h3b42cdff),
	.w7(32'h3ab08f23),
	.w8(32'h3a44e4a7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9120117),
	.w1(32'hba00ff83),
	.w2(32'hbb01cf8e),
	.w3(32'h3a45417c),
	.w4(32'hba27c493),
	.w5(32'hbac1a041),
	.w6(32'h3a623ab1),
	.w7(32'hba0516e3),
	.w8(32'hbb096110),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8030a54),
	.w1(32'hb6db6846),
	.w2(32'hb694ca95),
	.w3(32'hb6d90eb4),
	.w4(32'h3698d124),
	.w5(32'hb6a4aca9),
	.w6(32'hb6583f52),
	.w7(32'hb6380d95),
	.w8(32'hb503d813),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb157e76),
	.w1(32'hbb5702a6),
	.w2(32'hbaab0273),
	.w3(32'hbb144bd4),
	.w4(32'hbb25d681),
	.w5(32'h3803809c),
	.w6(32'hbb06ebd4),
	.w7(32'hbaf9782c),
	.w8(32'hba9ab123),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7819fdf),
	.w1(32'hb754fd75),
	.w2(32'h375f5bf2),
	.w3(32'hb7c4f0ce),
	.w4(32'h37b1aafb),
	.w5(32'h380d3130),
	.w6(32'hb882f887),
	.w7(32'hb752c8d2),
	.w8(32'h379a5287),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef29a0),
	.w1(32'hbab86452),
	.w2(32'hb961ec9a),
	.w3(32'h3a8ff3f6),
	.w4(32'h3a187e3c),
	.w5(32'h3a3d24ec),
	.w6(32'h3aaba067),
	.w7(32'h39862ab5),
	.w8(32'h3a1af11a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa323c0),
	.w1(32'h3b0815e3),
	.w2(32'h3a59be8b),
	.w3(32'hba755371),
	.w4(32'h37e301f7),
	.w5(32'hbb0f3a45),
	.w6(32'hbafa596b),
	.w7(32'h3a1d8cb7),
	.w8(32'hbadfe1eb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a977398),
	.w1(32'h3a6b880a),
	.w2(32'h39faf26e),
	.w3(32'h399cd5ab),
	.w4(32'h38dff51d),
	.w5(32'hba439ac0),
	.w6(32'hb941a57d),
	.w7(32'h39890b7f),
	.w8(32'hba989bc3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97d085d),
	.w1(32'hb8e3fec0),
	.w2(32'hb981de6b),
	.w3(32'hb93236f7),
	.w4(32'hb95c8794),
	.w5(32'hba18d886),
	.w6(32'hb95d7e4c),
	.w7(32'hb938b829),
	.w8(32'hb9db1248),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4c619),
	.w1(32'h3a8b2a4f),
	.w2(32'h3ac91bbf),
	.w3(32'hba9648ad),
	.w4(32'h39822e76),
	.w5(32'hbac6bc41),
	.w6(32'hbb299953),
	.w7(32'hb933edd6),
	.w8(32'hbb1abae2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b7c46),
	.w1(32'hbadef85f),
	.w2(32'hba96df3c),
	.w3(32'h375c5d82),
	.w4(32'h39dd96f7),
	.w5(32'h3a3860c8),
	.w6(32'h39500d55),
	.w7(32'h39f26ac5),
	.w8(32'h3a036e76),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7013),
	.w1(32'hba9df476),
	.w2(32'hbab93cef),
	.w3(32'h3a2e5c4a),
	.w4(32'h3a407969),
	.w5(32'h3a858dda),
	.w6(32'h3b059e3d),
	.w7(32'h3b0c7b61),
	.w8(32'h3a2952f5),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb657cad4),
	.w1(32'hb7ff878a),
	.w2(32'hb86f6e76),
	.w3(32'hb7f25430),
	.w4(32'hb859cab2),
	.w5(32'hb89eb19d),
	.w6(32'hb81aae11),
	.w7(32'hb87c9260),
	.w8(32'h377661af),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9802d8b),
	.w1(32'hb8179a27),
	.w2(32'hb8cd7d87),
	.w3(32'hb99e573f),
	.w4(32'h392d7e80),
	.w5(32'h38ff0f0f),
	.w6(32'hb984c5f3),
	.w7(32'h38cf3259),
	.w8(32'h391ee94e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10db11),
	.w1(32'hb912ba83),
	.w2(32'hbb16009b),
	.w3(32'h3ba5f18c),
	.w4(32'h3b2d0656),
	.w5(32'hba98a3f8),
	.w6(32'h3bfad0c1),
	.w7(32'h3b346a8c),
	.w8(32'hbaaa358f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a581),
	.w1(32'hba07fcbb),
	.w2(32'hba25c966),
	.w3(32'h3b4e2b1f),
	.w4(32'h3ab0f102),
	.w5(32'h3acf9bc9),
	.w6(32'h3b7dfe35),
	.w7(32'h3aa92bc3),
	.w8(32'h3a58059b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a719c4c),
	.w1(32'h3a6ee1a1),
	.w2(32'h3a1490d5),
	.w3(32'h3a91eaeb),
	.w4(32'h3a85d0fd),
	.w5(32'h393e5d59),
	.w6(32'h39ff39d2),
	.w7(32'h39ecd331),
	.w8(32'hbace28fc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aa128),
	.w1(32'hbbd6b304),
	.w2(32'hbb70d618),
	.w3(32'hb9dea9ff),
	.w4(32'hbaecbeda),
	.w5(32'hbae26bb7),
	.w6(32'h37f0b441),
	.w7(32'hbad69a5a),
	.w8(32'hbb425544),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7a966),
	.w1(32'hba4934bf),
	.w2(32'hb91090ea),
	.w3(32'hb9dbe32d),
	.w4(32'hba0b5eb8),
	.w5(32'h398f7fb9),
	.w6(32'hb967ec6e),
	.w7(32'hb9334ad3),
	.w8(32'h3993a3a0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e4202),
	.w1(32'hba91ec80),
	.w2(32'hba0143f2),
	.w3(32'h37c3137d),
	.w4(32'hb9b7ae6b),
	.w5(32'h39ae8a51),
	.w6(32'h3a027be1),
	.w7(32'hb9264b9e),
	.w8(32'h397c89e0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b481d7c),
	.w1(32'hbadc5954),
	.w2(32'hbc30cacc),
	.w3(32'h3b4f54b8),
	.w4(32'hbb176af2),
	.w5(32'hbbec276b),
	.w6(32'h3c20d3bc),
	.w7(32'h3b570d68),
	.w8(32'hbb17efee),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95a578),
	.w1(32'hbb4ffac0),
	.w2(32'hbae29680),
	.w3(32'h3ad5cbf6),
	.w4(32'h3a9f042e),
	.w5(32'h3b863c81),
	.w6(32'h3b47dcf5),
	.w7(32'h3b35944a),
	.w8(32'h3b89cd41),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bd6b0),
	.w1(32'hbaf82e54),
	.w2(32'hbb6743f4),
	.w3(32'h3b9b28c7),
	.w4(32'hba6294a2),
	.w5(32'hbb295269),
	.w6(32'h3b693ab6),
	.w7(32'h39a0106b),
	.w8(32'hb89d1192),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00dc0d),
	.w1(32'h3b36dde1),
	.w2(32'h3aac81ad),
	.w3(32'hbae72a3a),
	.w4(32'h39e0fd43),
	.w5(32'hba2b7965),
	.w6(32'hbb09a048),
	.w7(32'h3a44a2d2),
	.w8(32'hb70e5ed3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a898),
	.w1(32'h39721c25),
	.w2(32'h39c5331d),
	.w3(32'hbb247732),
	.w4(32'hba478a2e),
	.w5(32'hbb0be9bc),
	.w6(32'hbb75e00b),
	.w7(32'hba2588f7),
	.w8(32'hbaeb65e0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c04e5b),
	.w1(32'hb6b1067b),
	.w2(32'h37b0437b),
	.w3(32'hb5287b9d),
	.w4(32'hb5d8af33),
	.w5(32'hb752ddfb),
	.w6(32'hb7215137),
	.w7(32'h37032141),
	.w8(32'hb730e579),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33ce4f58),
	.w1(32'hb805fcbb),
	.w2(32'hb7f9186c),
	.w3(32'h360e0c0c),
	.w4(32'h379c3408),
	.w5(32'hb6656ad9),
	.w6(32'hb6f9fcf0),
	.w7(32'h36f2e424),
	.w8(32'h3688f356),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a856c),
	.w1(32'hb9b26537),
	.w2(32'h391ae189),
	.w3(32'h3a8e7e3c),
	.w4(32'h3a147e62),
	.w5(32'h3a163232),
	.w6(32'h3ad835d7),
	.w7(32'h3aaf828b),
	.w8(32'h3a5420d1),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37394bfb),
	.w1(32'hb832a445),
	.w2(32'h37acba34),
	.w3(32'hb7c4017f),
	.w4(32'hb86e3b01),
	.w5(32'h37acb292),
	.w6(32'hb77fb4f4),
	.w7(32'hb7e34a08),
	.w8(32'h3701cfde),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ded926),
	.w1(32'hbb12d943),
	.w2(32'hbb1e5545),
	.w3(32'hb8f8ac48),
	.w4(32'hbad630e8),
	.w5(32'hbafa6ac0),
	.w6(32'h3ae33bc4),
	.w7(32'hb7a56f89),
	.w8(32'hb9f4645a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824546),
	.w1(32'hbb4d6154),
	.w2(32'hba9a4926),
	.w3(32'h3a906152),
	.w4(32'hba8ece75),
	.w5(32'h3a4b9b9a),
	.w6(32'h3ab57c51),
	.w7(32'hb9c54b1a),
	.w8(32'hb9d5187d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a42b),
	.w1(32'h39de0d25),
	.w2(32'h39d00d96),
	.w3(32'h3a20b3eb),
	.w4(32'h394925bb),
	.w5(32'hb9221898),
	.w6(32'h3a279449),
	.w7(32'h38e07812),
	.w8(32'hba53fa43),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c548fb),
	.w1(32'h3801cd5a),
	.w2(32'h37f2023e),
	.w3(32'h388e52aa),
	.w4(32'h389d8b9c),
	.w5(32'hb790fd81),
	.w6(32'hb8a38cb2),
	.w7(32'hb818e61e),
	.w8(32'hb79420b2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801f70),
	.w1(32'hbbce66b4),
	.w2(32'hbc191d61),
	.w3(32'h3b8bd268),
	.w4(32'hbb0d706f),
	.w5(32'hbb91f0ca),
	.w6(32'h3bac1770),
	.w7(32'hbaae8d91),
	.w8(32'hb8237ba6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beb8d9),
	.w1(32'hbac0e9c5),
	.w2(32'hbaa03b3c),
	.w3(32'h3a50089c),
	.w4(32'hb8523012),
	.w5(32'h3a17efaa),
	.w6(32'h3a7e51ca),
	.w7(32'h39ba886e),
	.w8(32'h3a5254cd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f5b2fc),
	.w1(32'hb75bb362),
	.w2(32'h38967ee8),
	.w3(32'hb8bb9088),
	.w4(32'h3670eac9),
	.w5(32'h37d59173),
	.w6(32'hb9137c99),
	.w7(32'hb8e407aa),
	.w8(32'hb798e3ab),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898ca59),
	.w1(32'hbacb6991),
	.w2(32'hbaf3c653),
	.w3(32'h3b010d24),
	.w4(32'h3a266279),
	.w5(32'h3979af0b),
	.w6(32'h3b403f2e),
	.w7(32'h3b151409),
	.w8(32'h3ac42401),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb686d5db),
	.w1(32'hb7ab2a9e),
	.w2(32'hb78810dc),
	.w3(32'hb7d3c5e8),
	.w4(32'hb7b1f4b3),
	.w5(32'hb6e7cf5d),
	.w6(32'hb7bdc1f5),
	.w7(32'hb78f5053),
	.w8(32'hb75c0749),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f493fc),
	.w1(32'hb9142a8c),
	.w2(32'hb8c05848),
	.w3(32'h37c1d87a),
	.w4(32'hb8b52133),
	.w5(32'h38cd0e64),
	.w6(32'hb7ccf9f2),
	.w7(32'hb981670b),
	.w8(32'hb6fe5728),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f69b24),
	.w1(32'h38021cf8),
	.w2(32'h37359021),
	.w3(32'h384640d6),
	.w4(32'h37e21da4),
	.w5(32'hb70c4307),
	.w6(32'h37e4ec51),
	.w7(32'hb6018220),
	.w8(32'hb8304d3c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38396247),
	.w1(32'h3556fb1d),
	.w2(32'hb79c5b8c),
	.w3(32'h38a707dc),
	.w4(32'h383f5532),
	.w5(32'hb6c7f39a),
	.w6(32'h382f7bf7),
	.w7(32'h36057e6d),
	.w8(32'h3745d2bb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f4b01),
	.w1(32'h3a858ebc),
	.w2(32'h39118b8d),
	.w3(32'hb9fc44fb),
	.w4(32'h3833a84b),
	.w5(32'hba3a851b),
	.w6(32'hb9ca5c61),
	.w7(32'h3964095f),
	.w8(32'hb9e7c3e6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7699f8),
	.w1(32'hbba8d7f9),
	.w2(32'hbb7d9e95),
	.w3(32'hbadcb14a),
	.w4(32'hbaec2d6e),
	.w5(32'hba9e0957),
	.w6(32'hb844311e),
	.w7(32'hb94fc36f),
	.w8(32'hb8536996),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba196aea),
	.w1(32'hbaf8bee3),
	.w2(32'hbab6ca9b),
	.w3(32'h3af95a02),
	.w4(32'h3a8d0327),
	.w5(32'h3aa2f760),
	.w6(32'h3b2941ff),
	.w7(32'h3abb98eb),
	.w8(32'h3b0b1254),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb484d61),
	.w1(32'hbb5a3601),
	.w2(32'hbb0e2160),
	.w3(32'h3a35ce07),
	.w4(32'h398a6a72),
	.w5(32'h3abd9c11),
	.w6(32'h3ae40a4a),
	.w7(32'h3ace4927),
	.w8(32'h3b13e28b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb737e1bd),
	.w1(32'h37dd95ff),
	.w2(32'hb74ef4c5),
	.w3(32'hb7d6071e),
	.w4(32'hb78638b6),
	.w5(32'h363d270e),
	.w6(32'hb7d235fd),
	.w7(32'hb76d3c3d),
	.w8(32'hb84e06eb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba112de2),
	.w1(32'hba165c6b),
	.w2(32'hb9d14e6f),
	.w3(32'hb9221f8c),
	.w4(32'hb9901dc4),
	.w5(32'hb88db29f),
	.w6(32'hb84f3294),
	.w7(32'hb9514b7a),
	.w8(32'hb8bb00f5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370dd0fe),
	.w1(32'h3720263c),
	.w2(32'h372cce8a),
	.w3(32'hb72ca512),
	.w4(32'h36c9c67f),
	.w5(32'h3810e3ba),
	.w6(32'h370fed30),
	.w7(32'h370317ba),
	.w8(32'hb847f4d9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38108450),
	.w1(32'h37a152f7),
	.w2(32'h364f51ea),
	.w3(32'h381db799),
	.w4(32'h38271647),
	.w5(32'h379a5c78),
	.w6(32'hb87b7350),
	.w7(32'hb8510ca5),
	.w8(32'hb83eca26),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60d23e),
	.w1(32'hbb2118a9),
	.w2(32'hb9db914c),
	.w3(32'h38081e6d),
	.w4(32'h3a73b086),
	.w5(32'h3b0d43b4),
	.w6(32'h3a752864),
	.w7(32'hb9ab80b4),
	.w8(32'h3b076956),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d32e11),
	.w1(32'h37fb7480),
	.w2(32'hb7c4c573),
	.w3(32'h372c4bd2),
	.w4(32'h36485779),
	.w5(32'hb724889b),
	.w6(32'h36b66eb2),
	.w7(32'hb8182467),
	.w8(32'hb656b1c5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4a7b2),
	.w1(32'hb92026fd),
	.w2(32'hb9a85df4),
	.w3(32'hb9e42f14),
	.w4(32'hb98f3c3c),
	.w5(32'hba080c17),
	.w6(32'hb9d7f8c6),
	.w7(32'hb94719b6),
	.w8(32'hb9b99cc7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf8a7e),
	.w1(32'hbaa715f2),
	.w2(32'hba1169c6),
	.w3(32'hba998c8b),
	.w4(32'hba769d63),
	.w5(32'hba05ba33),
	.w6(32'hb5b2a620),
	.w7(32'h396ca498),
	.w8(32'h3963c04d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5af2f),
	.w1(32'hb3e8b5bf),
	.w2(32'h36a8ac41),
	.w3(32'h375fd741),
	.w4(32'hb7470afd),
	.w5(32'h377333a1),
	.w6(32'hb4d0363f),
	.w7(32'hb787757e),
	.w8(32'hb7b8a339),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb827ac08),
	.w1(32'hba58ac4e),
	.w2(32'hb9a57697),
	.w3(32'h3a36b266),
	.w4(32'hb8aa6e32),
	.w5(32'h39d525ef),
	.w6(32'h3a7fd9fe),
	.w7(32'h3a061e37),
	.w8(32'h3a03d56e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f756d),
	.w1(32'hba007139),
	.w2(32'hb93f1841),
	.w3(32'hba24d25b),
	.w4(32'hb9a5390b),
	.w5(32'h393c5248),
	.w6(32'hba10348e),
	.w7(32'hb998dfb9),
	.w8(32'h39283657),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8054),
	.w1(32'hbbb90f59),
	.w2(32'hbae5febf),
	.w3(32'hbb87bfc7),
	.w4(32'h39bb0e41),
	.w5(32'h3b0490b1),
	.w6(32'hbadcdaa0),
	.w7(32'h3b572a53),
	.w8(32'h3bb5aa7c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ec5939),
	.w1(32'hb8415c93),
	.w2(32'hb8e9ed41),
	.w3(32'h383719e7),
	.w4(32'hb6efd959),
	.w5(32'hb872566a),
	.w6(32'h3939f50e),
	.w7(32'h38fae480),
	.w8(32'h380d083c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6551da),
	.w1(32'h3b1f8548),
	.w2(32'h3abdb2c7),
	.w3(32'h3b0153b7),
	.w4(32'h3b2863c9),
	.w5(32'hb9f97e7d),
	.w6(32'h3b035ae8),
	.w7(32'h3aeed711),
	.w8(32'hba0f6696),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule