module layer_8_featuremap_78(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2316a),
	.w1(32'hba7bf82e),
	.w2(32'h3b7fd9b8),
	.w3(32'hbaade0e6),
	.w4(32'hba2afad6),
	.w5(32'h3b9a9fc8),
	.w6(32'hbb197367),
	.w7(32'hbad1ca5e),
	.w8(32'hba1b29a2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fbb80),
	.w1(32'h3b8f86e2),
	.w2(32'h3bc86804),
	.w3(32'h3bd27510),
	.w4(32'h3bc036f4),
	.w5(32'h3bda9cb6),
	.w6(32'h3bb54897),
	.w7(32'h3bcccb80),
	.w8(32'h3bea32d0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59dad),
	.w1(32'h3b809165),
	.w2(32'h3b22b266),
	.w3(32'h3b8a1ac6),
	.w4(32'h3b6ab160),
	.w5(32'h3b4263b4),
	.w6(32'h3bb8fd69),
	.w7(32'h3ba6d421),
	.w8(32'h3b8a4b53),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3f392),
	.w1(32'h3bef8d87),
	.w2(32'h3bc8d9e1),
	.w3(32'h3b8fee1a),
	.w4(32'h3bde345e),
	.w5(32'h3bc3e429),
	.w6(32'hbae0d571),
	.w7(32'hb8cc6a1a),
	.w8(32'h3b4d2389),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22c64),
	.w1(32'h3bf9009c),
	.w2(32'h3bb9748a),
	.w3(32'h3b7b7c02),
	.w4(32'h3b8c4a54),
	.w5(32'h3b9d4d80),
	.w6(32'h3b72b8c3),
	.w7(32'h3b1e6864),
	.w8(32'h3b38a1a0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48bb6f),
	.w1(32'h3bc88335),
	.w2(32'h3bb67a69),
	.w3(32'hbb0f8632),
	.w4(32'hbb5e54f6),
	.w5(32'hbb284973),
	.w6(32'h3b50d2d8),
	.w7(32'h3a78365c),
	.w8(32'h3b49e419),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c0418),
	.w1(32'h3b90afc3),
	.w2(32'h3b865b35),
	.w3(32'h3b749776),
	.w4(32'h3b5ea19d),
	.w5(32'h3b33212e),
	.w6(32'h3b3c2075),
	.w7(32'h3b389121),
	.w8(32'h3984581a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda3baf),
	.w1(32'h3c8a00af),
	.w2(32'h3c635ad5),
	.w3(32'h3b86e3f4),
	.w4(32'h3c21e4ec),
	.w5(32'h3c2a0a4e),
	.w6(32'h3b9b9a6a),
	.w7(32'h3be13b9e),
	.w8(32'h3c165414),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfbcd7),
	.w1(32'h3b134b35),
	.w2(32'h3ba462db),
	.w3(32'h3bf27d6e),
	.w4(32'h3bc4c96b),
	.w5(32'h3befdb42),
	.w6(32'h3b88b870),
	.w7(32'h3b61af20),
	.w8(32'h3aef24eb),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0db949),
	.w1(32'h3c449af6),
	.w2(32'h3b8f7aa2),
	.w3(32'h3c035c4f),
	.w4(32'h3c69b3d6),
	.w5(32'h3c3887b8),
	.w6(32'hbbb2c33b),
	.w7(32'hbba40d01),
	.w8(32'h3a6d8330),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80968f),
	.w1(32'h3b45c466),
	.w2(32'h3b84bed5),
	.w3(32'hbb95d357),
	.w4(32'h39a94a14),
	.w5(32'h3b858c59),
	.w6(32'hbb5233f0),
	.w7(32'hbb48ccf2),
	.w8(32'h3bcfd44a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae04793),
	.w1(32'h3b5b73a7),
	.w2(32'h3bc74c11),
	.w3(32'h3b505191),
	.w4(32'h3b97db74),
	.w5(32'h3bec96c9),
	.w6(32'h3a624df7),
	.w7(32'hb9f9db64),
	.w8(32'h3a4b6cf7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be14371),
	.w1(32'h3c0eb605),
	.w2(32'h3bd6adb2),
	.w3(32'h3b910a8d),
	.w4(32'h3b923acb),
	.w5(32'h3b1df4d5),
	.w6(32'h3b5fc5cd),
	.w7(32'h38361901),
	.w8(32'hbace730c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa24be8),
	.w1(32'h3b96329d),
	.w2(32'h3bd3a357),
	.w3(32'hbbd91f48),
	.w4(32'hbb4264e6),
	.w5(32'h3a2eadcd),
	.w6(32'h3ad1afd9),
	.w7(32'h3b3fda95),
	.w8(32'hbad31790),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5fbcc),
	.w1(32'h3bbf7dad),
	.w2(32'h3baf1586),
	.w3(32'hbb02f91e),
	.w4(32'h3a8ee862),
	.w5(32'h3b02da0f),
	.w6(32'h3b2a4e9c),
	.w7(32'h3b063203),
	.w8(32'h3b132e26),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63eb3c),
	.w1(32'h3b84e711),
	.w2(32'h3b0c152b),
	.w3(32'h3b19c1e0),
	.w4(32'h3addb1a1),
	.w5(32'h3af94a2e),
	.w6(32'h3b1293d9),
	.w7(32'h3a86e556),
	.w8(32'hbac51afb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0624be),
	.w1(32'hbc24f4ba),
	.w2(32'hbc1a82c8),
	.w3(32'hbb5a83ab),
	.w4(32'hba44acc4),
	.w5(32'hbaff2022),
	.w6(32'hbbc75206),
	.w7(32'hbb9bbf36),
	.w8(32'h3b3e6a8e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19abc6),
	.w1(32'h3c0380d8),
	.w2(32'h3bbb295b),
	.w3(32'h3a93e923),
	.w4(32'h3b6bc0d9),
	.w5(32'h3ba5e044),
	.w6(32'h3ba5687f),
	.w7(32'h3b153fe8),
	.w8(32'h3bae4a0f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea0161),
	.w1(32'h3c9cc645),
	.w2(32'h3c3c4aec),
	.w3(32'hbc030973),
	.w4(32'h3c64866f),
	.w5(32'h3cac3139),
	.w6(32'hbb547dfd),
	.w7(32'hbb2242fd),
	.w8(32'h3afd3872),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43d563),
	.w1(32'hbc738c23),
	.w2(32'hbbfff1cb),
	.w3(32'hbc84be7c),
	.w4(32'hbcaf1425),
	.w5(32'hbc169da9),
	.w6(32'hbb0d23b2),
	.w7(32'hbbb00611),
	.w8(32'h3adf2721),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a22e9),
	.w1(32'h3ae39c7d),
	.w2(32'hbb119d0c),
	.w3(32'hbb116817),
	.w4(32'hbb3b4bc5),
	.w5(32'hbb351773),
	.w6(32'hbb632294),
	.w7(32'hbc0b4f27),
	.w8(32'hbbd53cd1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99d897),
	.w1(32'h3b1caf9c),
	.w2(32'h3a9364bb),
	.w3(32'hbba28bc4),
	.w4(32'hbba8b271),
	.w5(32'hbb2adcfc),
	.w6(32'hb8991e00),
	.w7(32'hbb0bc8a8),
	.w8(32'h3b89e869),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf37122),
	.w1(32'hbc650cd9),
	.w2(32'h3b55709d),
	.w3(32'hbc878a58),
	.w4(32'hbc1e54ca),
	.w5(32'h3c626aea),
	.w6(32'hbcb33890),
	.w7(32'hbbfc32dd),
	.w8(32'h3c25b7d0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4580c8),
	.w1(32'h3c111b9e),
	.w2(32'h3c066b84),
	.w3(32'h3b56af40),
	.w4(32'h3bcf993a),
	.w5(32'h3b84a661),
	.w6(32'h3b9b77d1),
	.w7(32'h3b989905),
	.w8(32'h3b6ccdfd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9544c0),
	.w1(32'h3bf325a4),
	.w2(32'h3b49ee72),
	.w3(32'h3b94546e),
	.w4(32'h3bd28201),
	.w5(32'h3b9af85b),
	.w6(32'h3bc7b5c0),
	.w7(32'h3b25c7a3),
	.w8(32'h3a8ab832),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e0555),
	.w1(32'hbc0014ef),
	.w2(32'hbaf305a7),
	.w3(32'hb949604c),
	.w4(32'h3a8f7664),
	.w5(32'h3bcad5ce),
	.w6(32'hbc020ed9),
	.w7(32'h39d335a9),
	.w8(32'h3c18ace3),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e9c13),
	.w1(32'hbbbd5ad1),
	.w2(32'hbb6fd06b),
	.w3(32'h3aef3b37),
	.w4(32'hbac223b3),
	.w5(32'hbaeb9f2c),
	.w6(32'hbb7622a6),
	.w7(32'hbb294e9d),
	.w8(32'hba60d6ef),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c734a33),
	.w1(32'h3cbb921d),
	.w2(32'h3b7e73a6),
	.w3(32'hbcd39bbe),
	.w4(32'hbc529cff),
	.w5(32'h3d1742a9),
	.w6(32'hbc59a327),
	.w7(32'hbc31476e),
	.w8(32'h3c6d81ae),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6381e),
	.w1(32'h3be723ac),
	.w2(32'h3b96ca7c),
	.w3(32'hbab0bf09),
	.w4(32'h3b8d19e6),
	.w5(32'h3c03bcf8),
	.w6(32'hb9838e4f),
	.w7(32'hba8d453b),
	.w8(32'h3b9ab590),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4af7d),
	.w1(32'h3ae1ddcf),
	.w2(32'h3ad13763),
	.w3(32'h3ad2feb6),
	.w4(32'h3ab20232),
	.w5(32'h3ac7e18f),
	.w6(32'h3aed30d3),
	.w7(32'h3a868f31),
	.w8(32'h3b2839c1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a59bb),
	.w1(32'h3be86926),
	.w2(32'h3b973e11),
	.w3(32'h3b54ebd7),
	.w4(32'h3bad74c1),
	.w5(32'h3b9ec264),
	.w6(32'h3bd308f8),
	.w7(32'h3b306842),
	.w8(32'hbb8dbfe6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d4327),
	.w1(32'h3bace8cf),
	.w2(32'hb9039d8e),
	.w3(32'hba707ca5),
	.w4(32'h3b61798e),
	.w5(32'hb9249815),
	.w6(32'h3afaf478),
	.w7(32'hbb0d18e9),
	.w8(32'hba8297bd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a293a13),
	.w1(32'h3b9e66f0),
	.w2(32'h3bbcf1dd),
	.w3(32'h3b2fc7f0),
	.w4(32'h3b405118),
	.w5(32'h3aa637e8),
	.w6(32'hba513719),
	.w7(32'hba9f5c1c),
	.w8(32'hbacc2d69),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1c84),
	.w1(32'hbb0f7af6),
	.w2(32'hbb5b5d8b),
	.w3(32'hbb7acc6a),
	.w4(32'hbb95b210),
	.w5(32'hbb09f663),
	.w6(32'h3b6b1e53),
	.w7(32'hbb91a074),
	.w8(32'hbac4c127),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cb9b5),
	.w1(32'h3b21b46b),
	.w2(32'h3bc342b5),
	.w3(32'hbc05340c),
	.w4(32'hbbddaf7c),
	.w5(32'hbb0a076c),
	.w6(32'h3a94a7bf),
	.w7(32'h3a634c63),
	.w8(32'h3af4d4c7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00c7ac),
	.w1(32'h3c2d4295),
	.w2(32'h3c2db496),
	.w3(32'h3b9f5e8f),
	.w4(32'h3bd2739b),
	.w5(32'h3c3ce574),
	.w6(32'h3bb1602f),
	.w7(32'h3baa1429),
	.w8(32'h3ba16089),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a455ac8),
	.w1(32'h3a36078a),
	.w2(32'h397f1e0f),
	.w3(32'hb9d30ff2),
	.w4(32'h3a8c4835),
	.w5(32'h3a256d2a),
	.w6(32'h3a89f707),
	.w7(32'h38c789a1),
	.w8(32'h3a8ec5de),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48c38b),
	.w1(32'h3b4ae3e3),
	.w2(32'h3b6e7089),
	.w3(32'h3b005d8e),
	.w4(32'h3b2c19e6),
	.w5(32'h3b7f1690),
	.w6(32'h3ab68a57),
	.w7(32'h3b05af68),
	.w8(32'h3a90b10f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0f84b),
	.w1(32'h3c43605e),
	.w2(32'h3c2d14d8),
	.w3(32'hbb5955d2),
	.w4(32'h3b2d0468),
	.w5(32'h3b8c6be6),
	.w6(32'h3bb3c23e),
	.w7(32'h3b649cc3),
	.w8(32'h3a304cf0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7b13d),
	.w1(32'h3aa74fec),
	.w2(32'hb9ff4f8f),
	.w3(32'hba5bc8c9),
	.w4(32'h39fa0a68),
	.w5(32'hba77d2a7),
	.w6(32'h39388a5f),
	.w7(32'hbac4ab7f),
	.w8(32'hba2a7dd6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2d115),
	.w1(32'h3bb6d204),
	.w2(32'h3c51a7ec),
	.w3(32'h3c66ebc7),
	.w4(32'h3c802fd1),
	.w5(32'h3cb8b905),
	.w6(32'h3bf7fa70),
	.w7(32'h3c1f224f),
	.w8(32'h3c985d7b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eeed6),
	.w1(32'h3b4e7d14),
	.w2(32'h3b2c42bc),
	.w3(32'h3b5223b9),
	.w4(32'h3b8cca79),
	.w5(32'h3b90d2a1),
	.w6(32'h3b331617),
	.w7(32'h3b2278c9),
	.w8(32'h3b35863b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f75220),
	.w1(32'h3910fcdf),
	.w2(32'hb96c0bfe),
	.w3(32'h39cec193),
	.w4(32'hb8c8e84f),
	.w5(32'hb996fbb5),
	.w6(32'h39d1f834),
	.w7(32'hb8ed928c),
	.w8(32'hb9ecee31),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a141034),
	.w1(32'hbad459a0),
	.w2(32'hb980763a),
	.w3(32'hba346da7),
	.w4(32'hba030e0b),
	.w5(32'h3b371ba1),
	.w6(32'hbad8ee14),
	.w7(32'hbab291d9),
	.w8(32'h3a699b6c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e2d07),
	.w1(32'h3a2c103e),
	.w2(32'h3b6b1c5b),
	.w3(32'hbafadbce),
	.w4(32'h3a91aced),
	.w5(32'h3c0cd584),
	.w6(32'hbb11a7da),
	.w7(32'hb9bcf1c3),
	.w8(32'h3b21a30d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3702a060),
	.w1(32'h3ac719c1),
	.w2(32'h3af1774c),
	.w3(32'h3a82d3e7),
	.w4(32'h3b4984af),
	.w5(32'h3b53be4d),
	.w6(32'h3acd5c20),
	.w7(32'h3a678575),
	.w8(32'h39d4440d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80e688c),
	.w1(32'hb6ff20d4),
	.w2(32'h37f20fc1),
	.w3(32'hb7b8f6a9),
	.w4(32'h378a5c4c),
	.w5(32'h37d7ac66),
	.w6(32'hb7fcbdbc),
	.w7(32'h380d351d),
	.w8(32'hb694c9dd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaea581),
	.w1(32'hbbde83b3),
	.w2(32'h3a8bb9cf),
	.w3(32'hbc367a14),
	.w4(32'hbbd9ebd1),
	.w5(32'h3bbfae9d),
	.w6(32'hbc197c4e),
	.w7(32'hbb857175),
	.w8(32'h398769f6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8aaf9c),
	.w1(32'h3ab65cb2),
	.w2(32'h3a644a6d),
	.w3(32'h3b176128),
	.w4(32'h3b0c95b6),
	.w5(32'h3add6939),
	.w6(32'h3b4e2f52),
	.w7(32'h3aecc573),
	.w8(32'h3af25bc0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba606fa8),
	.w1(32'hbae8c058),
	.w2(32'h3b0e0e55),
	.w3(32'h3a15b0b4),
	.w4(32'h3af505f5),
	.w5(32'h3bb8d981),
	.w6(32'hb968e939),
	.w7(32'hba8a4947),
	.w8(32'h3b67372c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77d966),
	.w1(32'h3b859a5a),
	.w2(32'h3ba944cf),
	.w3(32'h3ba6d4ed),
	.w4(32'h3b6f47b2),
	.w5(32'h3b3cf72f),
	.w6(32'h3b382a0a),
	.w7(32'h399074f7),
	.w8(32'hb9249c7a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cf310),
	.w1(32'h3986b5b4),
	.w2(32'h3bd3f3c7),
	.w3(32'hbb2fbb95),
	.w4(32'h39e4468a),
	.w5(32'h3c60d44f),
	.w6(32'hbbc306a0),
	.w7(32'h3bca2de2),
	.w8(32'h3c8e49bb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba83bc3),
	.w1(32'hbb84884a),
	.w2(32'hbadee5d9),
	.w3(32'hbb965646),
	.w4(32'hbb8d1da6),
	.w5(32'hbad3f4ec),
	.w6(32'hbb158788),
	.w7(32'h3a11b87e),
	.w8(32'h3b0293ad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874741),
	.w1(32'h384be0f5),
	.w2(32'h3bd7bb04),
	.w3(32'h3ad7cf04),
	.w4(32'h3b463714),
	.w5(32'h3c012422),
	.w6(32'h3a766655),
	.w7(32'h3a836915),
	.w8(32'h3ac810c9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d166b),
	.w1(32'h37a19f62),
	.w2(32'h38dcf3ff),
	.w3(32'hb817744e),
	.w4(32'h380cf75d),
	.w5(32'h390a7ccc),
	.w6(32'hb8791bf5),
	.w7(32'h38ef5f28),
	.w8(32'h3881b2ff),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadde29e),
	.w1(32'hbabeee76),
	.w2(32'h3c0ac3ff),
	.w3(32'hbbbb7c78),
	.w4(32'h3a49cca0),
	.w5(32'h3c53a63b),
	.w6(32'hbbda4ea8),
	.w7(32'hbb9f0c1e),
	.w8(32'hbaa78e2f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7263e),
	.w1(32'hbac0f23c),
	.w2(32'hba87ef86),
	.w3(32'hba93ee43),
	.w4(32'hbb4cbd41),
	.w5(32'hbb467639),
	.w6(32'hbb6ecf33),
	.w7(32'hbb8ee5b9),
	.w8(32'hbb72ab4b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba35e7c),
	.w1(32'h3b1ba5f1),
	.w2(32'h3afa3207),
	.w3(32'h3b94e0a7),
	.w4(32'h3ba263b9),
	.w5(32'h3bf4510f),
	.w6(32'h3b13ca76),
	.w7(32'h3b3d0c8f),
	.w8(32'h3bb387cd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6ed1e),
	.w1(32'hba110910),
	.w2(32'h384c045b),
	.w3(32'hbb0fd3a8),
	.w4(32'hbb17fe1c),
	.w5(32'h3b14bec4),
	.w6(32'hbb0cc044),
	.w7(32'hbad0b247),
	.w8(32'h3a21af45),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6551d),
	.w1(32'h38fd4053),
	.w2(32'h3a6712d0),
	.w3(32'h3a58b334),
	.w4(32'h3a03ecf7),
	.w5(32'h3ac5c11b),
	.w6(32'h3a6100ed),
	.w7(32'h3ae8d4b3),
	.w8(32'h3b27f7d5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb843519c),
	.w1(32'h391f010d),
	.w2(32'h391164f7),
	.w3(32'h38949c5e),
	.w4(32'h3963b4bd),
	.w5(32'h39909405),
	.w6(32'hb98e5641),
	.w7(32'hb914b4b2),
	.w8(32'hb8e1d690),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0853fe),
	.w1(32'hb9fb70f2),
	.w2(32'h38b07235),
	.w3(32'hba2eaa43),
	.w4(32'hb9df0546),
	.w5(32'hb7b5426c),
	.w6(32'hba3b327a),
	.w7(32'hba0818a3),
	.w8(32'hb9ba3773),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f32469),
	.w1(32'h3b77a28c),
	.w2(32'h3c24a280),
	.w3(32'h3b8d2e33),
	.w4(32'h3c0220a9),
	.w5(32'h3c63d6a7),
	.w6(32'h3a4b72a9),
	.w7(32'h3b0f7aff),
	.w8(32'h3be1464e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918f7c7),
	.w1(32'h3a592467),
	.w2(32'h3abee474),
	.w3(32'h3a189094),
	.w4(32'h3a688c28),
	.w5(32'h3b0223e8),
	.w6(32'h3ad865a1),
	.w7(32'h3b3cd17c),
	.w8(32'h3b344ef0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a6073),
	.w1(32'hbacf57cc),
	.w2(32'hbb16d881),
	.w3(32'hba98c605),
	.w4(32'hbaf68cf3),
	.w5(32'hbb10ac6e),
	.w6(32'hbac86897),
	.w7(32'hbb2d4388),
	.w8(32'hbb0ca3d1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761635),
	.w1(32'h3b1df3f0),
	.w2(32'h3b404ea7),
	.w3(32'h3b13718c),
	.w4(32'h3b143f77),
	.w5(32'h3b8de8c9),
	.w6(32'h3ab908da),
	.w7(32'h3b27903d),
	.w8(32'h3b6a7fd3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fad04),
	.w1(32'h3b180aa9),
	.w2(32'h3b5c900f),
	.w3(32'h3b284d7d),
	.w4(32'h3a8918ca),
	.w5(32'h3b65b43b),
	.w6(32'h3b0894e4),
	.w7(32'h3b1c7d76),
	.w8(32'h3b9ce870),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2943cf),
	.w1(32'hbac1dfad),
	.w2(32'h3a71a8e4),
	.w3(32'hbaab7c10),
	.w4(32'hb9d907d1),
	.w5(32'h3b07dd21),
	.w6(32'hbae32c11),
	.w7(32'hbb5f72e3),
	.w8(32'hbb484236),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1c310),
	.w1(32'hb9667c71),
	.w2(32'hb971862d),
	.w3(32'hb985427b),
	.w4(32'hb8d5fd54),
	.w5(32'hb938672a),
	.w6(32'hb9408b95),
	.w7(32'hb8e660d8),
	.w8(32'hb8b03ac7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4167c),
	.w1(32'hbbca5e8b),
	.w2(32'hbb90798b),
	.w3(32'hbbe8135e),
	.w4(32'hbc4f0a3d),
	.w5(32'h3b948597),
	.w6(32'hbc10d738),
	.w7(32'hbbdcfd4a),
	.w8(32'h3b1dd452),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4b10f),
	.w1(32'h38a68fb1),
	.w2(32'hb8ad2d91),
	.w3(32'h3897abd2),
	.w4(32'h38e88dbd),
	.w5(32'hb8016991),
	.w6(32'h38a21289),
	.w7(32'h36c8966d),
	.w8(32'hb8c4a784),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaefb69a),
	.w1(32'hbaaeaebd),
	.w2(32'hba370d10),
	.w3(32'h3a418314),
	.w4(32'h3a97896c),
	.w5(32'h3b1ffa96),
	.w6(32'h3a874f02),
	.w7(32'h3b8f9d5b),
	.w8(32'h3bae9418),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b300bc),
	.w1(32'h3a197a3f),
	.w2(32'h38f370f5),
	.w3(32'h3a17ddc7),
	.w4(32'h3a4914bf),
	.w5(32'h39f4f9cc),
	.w6(32'h3a267c78),
	.w7(32'h3a63cb7e),
	.w8(32'h39af9642),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba839ee),
	.w1(32'h3bd80d1e),
	.w2(32'h3be77c1f),
	.w3(32'h3c07d162),
	.w4(32'h3c10736e),
	.w5(32'h3c11d1b0),
	.w6(32'h3b6025d3),
	.w7(32'h3b57f520),
	.w8(32'h3b16abee),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eb396b),
	.w1(32'h3755e770),
	.w2(32'h37f9f2d7),
	.w3(32'hb83d17ab),
	.w4(32'h36f3bf07),
	.w5(32'h37de4649),
	.w6(32'hb886fb8b),
	.w7(32'hb7cbc8b9),
	.w8(32'h375c9a4b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ed23a),
	.w1(32'hbb87e571),
	.w2(32'hbade6c32),
	.w3(32'hbb467eb2),
	.w4(32'hbba3d5a4),
	.w5(32'hbaf201d2),
	.w6(32'hbbb63a79),
	.w7(32'hbb9e1792),
	.w8(32'hb9d8e250),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883716e),
	.w1(32'h38553b62),
	.w2(32'h3873630d),
	.w3(32'h389c7be8),
	.w4(32'h389a9823),
	.w5(32'h387bd51a),
	.w6(32'h387c5de2),
	.w7(32'h384a782f),
	.w8(32'h37898263),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943e7de),
	.w1(32'hbad72087),
	.w2(32'h3a9f69e1),
	.w3(32'hbb841809),
	.w4(32'hb9663dc9),
	.w5(32'h3be3ee71),
	.w6(32'hbba64261),
	.w7(32'hba26f78f),
	.w8(32'h3b45a461),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39623cdd),
	.w1(32'h3b287ae5),
	.w2(32'h3b9672fc),
	.w3(32'h3b0bc962),
	.w4(32'h3b8f011a),
	.w5(32'h3bea85dc),
	.w6(32'h3a590aa2),
	.w7(32'h3b33c695),
	.w8(32'h3b23ab08),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a123ee6),
	.w1(32'h3a188f77),
	.w2(32'h39c2908c),
	.w3(32'h38811f0b),
	.w4(32'h3949704b),
	.w5(32'h397f6614),
	.w6(32'hb8e372ec),
	.w7(32'hb8dfc227),
	.w8(32'h3940968a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c63252),
	.w1(32'hb8b17f80),
	.w2(32'hb937c2eb),
	.w3(32'hb8d86088),
	.w4(32'hb82b14eb),
	.w5(32'hb929e1b3),
	.w6(32'hb8bfaf12),
	.w7(32'hb895b865),
	.w8(32'hb918c547),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38ad91),
	.w1(32'h3a52e692),
	.w2(32'h39da5bd8),
	.w3(32'h3aa85da4),
	.w4(32'h39a67e98),
	.w5(32'h3a87f831),
	.w6(32'h3acee5c8),
	.w7(32'h3b61fea7),
	.w8(32'h3bd52847),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaaed5),
	.w1(32'hbb100bac),
	.w2(32'h3a8dc8bd),
	.w3(32'h398a0ffc),
	.w4(32'h3ac45ed7),
	.w5(32'h3bd8c130),
	.w6(32'h388708d2),
	.w7(32'h3acca4fe),
	.w8(32'h3bb77c35),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c014bfd),
	.w1(32'h3c0fa08f),
	.w2(32'h3c87063b),
	.w3(32'h3c906c2a),
	.w4(32'h3c925ca5),
	.w5(32'h3c9646dd),
	.w6(32'h3c6a91e8),
	.w7(32'h3c341da7),
	.w8(32'h3c3b45bf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700624),
	.w1(32'hbbcf0b24),
	.w2(32'h3ac90247),
	.w3(32'hbb55ce4c),
	.w4(32'h3ab07d5f),
	.w5(32'h3c7511aa),
	.w6(32'hbbcb92e0),
	.w7(32'hba4be9aa),
	.w8(32'h3c01038d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85ac6d),
	.w1(32'hbb68890b),
	.w2(32'h3a1452f0),
	.w3(32'hbbaf5512),
	.w4(32'hbb3918c9),
	.w5(32'h3a231fc2),
	.w6(32'hbc0ffb68),
	.w7(32'hbb5611bb),
	.w8(32'h3bad9fa0),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38538d37),
	.w1(32'h397ae10b),
	.w2(32'h3944d0e1),
	.w3(32'h3883cc82),
	.w4(32'h398f945f),
	.w5(32'h398e582d),
	.w6(32'hb80aa3d9),
	.w7(32'h393a2cb7),
	.w8(32'hb8081581),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb799e166),
	.w1(32'h37e1d9c0),
	.w2(32'h37a695d0),
	.w3(32'hb80ef92f),
	.w4(32'h3787f46f),
	.w5(32'h36fed269),
	.w6(32'hb83167d6),
	.w7(32'h36b401ca),
	.w8(32'h362015e1),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d5bfb),
	.w1(32'hb8172c2d),
	.w2(32'h38e8d513),
	.w3(32'hb61038eb),
	.w4(32'h3815f0a4),
	.w5(32'h38bd7c21),
	.w6(32'hb8414570),
	.w7(32'h37a41898),
	.w8(32'h37a3aafd),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233983),
	.w1(32'hbb09e103),
	.w2(32'hb97d07f8),
	.w3(32'hbb4f26f8),
	.w4(32'hbb04d1fa),
	.w5(32'h3a0e62a6),
	.w6(32'hbb876239),
	.w7(32'hbb11ecd7),
	.w8(32'h3982ab62),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7cd41),
	.w1(32'h3b1c3888),
	.w2(32'h3b06182e),
	.w3(32'h3ade53ef),
	.w4(32'h3adc203d),
	.w5(32'h3af1dcf7),
	.w6(32'h3a5b8c42),
	.w7(32'h3a5d5726),
	.w8(32'h3adc2c1d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9001a00),
	.w1(32'hba85135d),
	.w2(32'hba4d8cd1),
	.w3(32'hb9bc2905),
	.w4(32'hba84ef68),
	.w5(32'hba4aa139),
	.w6(32'hbaa35849),
	.w7(32'hbb0f3c5b),
	.w8(32'hbacb7b31),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377842d4),
	.w1(32'hbaf43b50),
	.w2(32'hbadf941e),
	.w3(32'h3a019d37),
	.w4(32'hba700748),
	.w5(32'hb9952479),
	.w6(32'h39e1082e),
	.w7(32'h3b1a9ae5),
	.w8(32'h3b1a8e85),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fd5ad),
	.w1(32'h3993fd92),
	.w2(32'h3b30d7c6),
	.w3(32'h39e0665f),
	.w4(32'h3b04143c),
	.w5(32'h3b93a0eb),
	.w6(32'hb8ea2944),
	.w7(32'h3ab6e52d),
	.w8(32'h3b68456c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942a314),
	.w1(32'h398046a5),
	.w2(32'h3ad605ca),
	.w3(32'h38cf475f),
	.w4(32'h39a5a616),
	.w5(32'h3ad15cf9),
	.w6(32'hb9f0920f),
	.w7(32'h37c18978),
	.w8(32'h39f22334),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfea09),
	.w1(32'hbb07c2b5),
	.w2(32'h3ac54117),
	.w3(32'hbaeca9ca),
	.w4(32'h396380cf),
	.w5(32'h3b598efd),
	.w6(32'hbb8f73da),
	.w7(32'hbb54f925),
	.w8(32'hbac23742),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1351c4),
	.w1(32'hbc147f2f),
	.w2(32'hba4bacaf),
	.w3(32'hbbccc610),
	.w4(32'hbb819bd2),
	.w5(32'h3b8d9e84),
	.w6(32'hbbdfa164),
	.w7(32'hb9124c74),
	.w8(32'h3bbb7d3f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79707e3),
	.w1(32'h37c67642),
	.w2(32'h37bc0635),
	.w3(32'h37292634),
	.w4(32'h381d7450),
	.w5(32'h37ab8f2a),
	.w6(32'hb65da72d),
	.w7(32'h3806ad1f),
	.w8(32'h342d5a0a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c4313),
	.w1(32'hb78c82fe),
	.w2(32'hb9287608),
	.w3(32'hb91f580e),
	.w4(32'hb7c46f06),
	.w5(32'hb92d9ee9),
	.w6(32'hb945cb3b),
	.w7(32'hb845d00d),
	.w8(32'hb930345a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1f2e4),
	.w1(32'h38928dee),
	.w2(32'h3782b786),
	.w3(32'hb84dae70),
	.w4(32'h383f0bd0),
	.w5(32'h3593e654),
	.w6(32'hb8a6c344),
	.w7(32'h37fc0c4b),
	.w8(32'h36c61ebf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed5fd0),
	.w1(32'h39cd1cd2),
	.w2(32'h39df3bc2),
	.w3(32'h3a26ca02),
	.w4(32'h3958b963),
	.w5(32'h3953aaac),
	.w6(32'h39bc61ba),
	.w7(32'h396b961b),
	.w8(32'h399b684e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a704d),
	.w1(32'h3b4c65a2),
	.w2(32'h3b4359c7),
	.w3(32'h3b1fe052),
	.w4(32'h3b2a7c11),
	.w5(32'h3b27c8cb),
	.w6(32'hb923fd70),
	.w7(32'h39dfeea3),
	.w8(32'h3a1250dd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea90d6),
	.w1(32'h39195a63),
	.w2(32'h3a8237b9),
	.w3(32'h3910bb0e),
	.w4(32'h3a483817),
	.w5(32'h3a6c8f1d),
	.w6(32'hbb17a472),
	.w7(32'hbaa2dc42),
	.w8(32'hba782309),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f8f8),
	.w1(32'h3b49aa26),
	.w2(32'h3b5835d1),
	.w3(32'h3b1c418f),
	.w4(32'h3a39cbde),
	.w5(32'h39ce4618),
	.w6(32'h3ba5b8ce),
	.w7(32'h3c1c3b08),
	.w8(32'h3bcccb5b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380788c8),
	.w1(32'h3936cdde),
	.w2(32'hb98999a0),
	.w3(32'h3a47e5f0),
	.w4(32'hb8b41392),
	.w5(32'hba93a4d2),
	.w6(32'h3aa7c0b8),
	.w7(32'h39dd7b9d),
	.w8(32'hba4005f1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a731d9e),
	.w1(32'hbb818dc2),
	.w2(32'hbb61dbe4),
	.w3(32'hbb4743bb),
	.w4(32'hbbab2f8f),
	.w5(32'h3b1f7e3d),
	.w6(32'hbb847ad2),
	.w7(32'hba1890c8),
	.w8(32'h3bb96f7a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa4ec6),
	.w1(32'hbb0a08c0),
	.w2(32'hba2a0f27),
	.w3(32'hbc12930b),
	.w4(32'hbb5796ed),
	.w5(32'hbac4fa0e),
	.w6(32'h3af6b814),
	.w7(32'hbb2f03bb),
	.w8(32'h3ad5a58e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2a31e),
	.w1(32'hbb3e7476),
	.w2(32'hba8ec1dd),
	.w3(32'h3a60ca72),
	.w4(32'hb990b174),
	.w5(32'h39e15d8d),
	.w6(32'hba8ace78),
	.w7(32'hb9539ee3),
	.w8(32'h3b110a7e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a918c5a),
	.w1(32'hb6b67751),
	.w2(32'h3a3d1f66),
	.w3(32'h3a82c048),
	.w4(32'hb9cc89c1),
	.w5(32'h381dce32),
	.w6(32'hb8b8a60a),
	.w7(32'hba845ead),
	.w8(32'hbad8bf66),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7eca7),
	.w1(32'h3b2ad139),
	.w2(32'h3b5b5dd4),
	.w3(32'h3b9a02af),
	.w4(32'h3bb3db04),
	.w5(32'h3bbaabc8),
	.w6(32'hba917bf3),
	.w7(32'h3b2ac6da),
	.w8(32'h3b8ef7b2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd737),
	.w1(32'hbc17376b),
	.w2(32'hbbf51ae0),
	.w3(32'hba92f1d0),
	.w4(32'hbb41090e),
	.w5(32'hbabf9e1a),
	.w6(32'hba863dcc),
	.w7(32'hbb4f5f3b),
	.w8(32'hbb294abe),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c83cc),
	.w1(32'h3a8f1166),
	.w2(32'h3b25fc18),
	.w3(32'h3afbcf0c),
	.w4(32'h3af7bce3),
	.w5(32'h3b876d5b),
	.w6(32'h3b54ef96),
	.w7(32'h3a8bc7ff),
	.w8(32'h3b2af19a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12aa33),
	.w1(32'hbac41dbd),
	.w2(32'hba7e388f),
	.w3(32'h398fcc5c),
	.w4(32'hbb01b66e),
	.w5(32'hba0b0f16),
	.w6(32'h3b91f2f5),
	.w7(32'h3a849267),
	.w8(32'hba33a26d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad03a27),
	.w1(32'h3a615b20),
	.w2(32'h3a812e41),
	.w3(32'h3ace6e35),
	.w4(32'h3a7e380c),
	.w5(32'h3a740eb4),
	.w6(32'hb8f8f661),
	.w7(32'h3a2317c3),
	.w8(32'h3a1ecf2e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399080e3),
	.w1(32'hb968a0dd),
	.w2(32'h3a34b2e3),
	.w3(32'h3a92b8e1),
	.w4(32'h3aa5d19a),
	.w5(32'h3a9668c5),
	.w6(32'hb900ac7e),
	.w7(32'h39aea302),
	.w8(32'h3aabc9d4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce992a),
	.w1(32'hbb02a487),
	.w2(32'hba731f10),
	.w3(32'hb819c75d),
	.w4(32'hba299ba0),
	.w5(32'hba8b3b6e),
	.w6(32'hbb777c06),
	.w7(32'hbb5cd01d),
	.w8(32'hbbc56a4d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba955723),
	.w1(32'hba7e7608),
	.w2(32'hbb82a248),
	.w3(32'h3ad94886),
	.w4(32'hba2e85cf),
	.w5(32'hbbac0eaa),
	.w6(32'h3b21e9e9),
	.w7(32'h39e03a7f),
	.w8(32'h3abf8720),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac752e0),
	.w1(32'hb99018a9),
	.w2(32'h3a69acc3),
	.w3(32'h3b02dc97),
	.w4(32'h3a61561d),
	.w5(32'h3badcf07),
	.w6(32'h3a3d70df),
	.w7(32'h39a4d91b),
	.w8(32'h3b5c143a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a966f71),
	.w1(32'hba96828a),
	.w2(32'hbbd80d9c),
	.w3(32'hb9c130a8),
	.w4(32'hbb039795),
	.w5(32'hbb9fcefa),
	.w6(32'h3b850497),
	.w7(32'hbb0964a5),
	.w8(32'hb9a827b6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc0ed8),
	.w1(32'h3b1473d8),
	.w2(32'hbb13c5bf),
	.w3(32'hba8a327d),
	.w4(32'hbb8b417a),
	.w5(32'hbb8667bb),
	.w6(32'h38cc2864),
	.w7(32'hbadcafee),
	.w8(32'hbaa96eeb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c632c),
	.w1(32'h3b1c4231),
	.w2(32'h3b4a5f85),
	.w3(32'h3a9832d9),
	.w4(32'hbb071c49),
	.w5(32'hbb9a5d94),
	.w6(32'hbb884f54),
	.w7(32'hbb61c34a),
	.w8(32'h39658e99),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b718),
	.w1(32'h3b474a85),
	.w2(32'h3bc07152),
	.w3(32'hbbc97cd2),
	.w4(32'hbaeb9aa4),
	.w5(32'h3b9dadc9),
	.w6(32'hbb6b58e9),
	.w7(32'hbb553f1f),
	.w8(32'h3b2e3bcf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39afcb36),
	.w1(32'h3a9f6bbc),
	.w2(32'h3b02ed6c),
	.w3(32'h397e45a2),
	.w4(32'h3aff55b6),
	.w5(32'h3b2e1a13),
	.w6(32'h3b2b6352),
	.w7(32'h3b8004c3),
	.w8(32'hbb85a26f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ab0a),
	.w1(32'hbb21796f),
	.w2(32'hbb2ca6d0),
	.w3(32'hbaab6a45),
	.w4(32'hb942ee06),
	.w5(32'hbaffec0c),
	.w6(32'hbba2903b),
	.w7(32'hbbbeb2e6),
	.w8(32'hbadb05a9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b63d8f),
	.w1(32'hb98b086d),
	.w2(32'hb84d24e9),
	.w3(32'hba60fdad),
	.w4(32'hba8385df),
	.w5(32'hbbbea338),
	.w6(32'h3b021161),
	.w7(32'h3a8dc1d6),
	.w8(32'h37424999),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43bcb9),
	.w1(32'hb9d7795f),
	.w2(32'h3842561f),
	.w3(32'h3b2484f3),
	.w4(32'hb9b96468),
	.w5(32'h39ebc9ef),
	.w6(32'h3a6c60cb),
	.w7(32'hb9d386e4),
	.w8(32'h3ab6a017),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399274c1),
	.w1(32'h3a8394c8),
	.w2(32'h3b8376c4),
	.w3(32'h3a43499a),
	.w4(32'h3a9b5e8d),
	.w5(32'h3b234de5),
	.w6(32'hba526d78),
	.w7(32'h3a803ddc),
	.w8(32'h3ac6ea71),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ead01),
	.w1(32'hbb31818f),
	.w2(32'h3b8fa057),
	.w3(32'hbb348be6),
	.w4(32'hbb34c766),
	.w5(32'h3bdc520e),
	.w6(32'hba153416),
	.w7(32'hbadbac05),
	.w8(32'hb9e02bcc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule