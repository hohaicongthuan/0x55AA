module layer_6_featuremap_110(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01270b),
	.w1(32'hbb8ee4a5),
	.w2(32'hba1c34c8),
	.w3(32'hba4dd859),
	.w4(32'h3b910bb8),
	.w5(32'h3b742a11),
	.w6(32'hbb35ccd7),
	.w7(32'h3808b2f6),
	.w8(32'hba674ea7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8be54),
	.w1(32'h3a710071),
	.w2(32'hba0ae652),
	.w3(32'h39fef63b),
	.w4(32'hbb8f2c4c),
	.w5(32'h39e352b3),
	.w6(32'hbbaec105),
	.w7(32'hbbb13c9f),
	.w8(32'hbc039569),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d6999),
	.w1(32'h3b96d53f),
	.w2(32'h3c5a2f8d),
	.w3(32'hbac11fbd),
	.w4(32'h3acbc77c),
	.w5(32'h3beb6618),
	.w6(32'h3b0c6bf4),
	.w7(32'h3becc45e),
	.w8(32'hbbb33fbc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf32b9f),
	.w1(32'hbbc48f6f),
	.w2(32'h39a61379),
	.w3(32'h3b11a3cb),
	.w4(32'hba7cd40d),
	.w5(32'h3b0ab133),
	.w6(32'h3bda4552),
	.w7(32'h3bc776c8),
	.w8(32'h3be8b794),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d9f1),
	.w1(32'h3c67c19f),
	.w2(32'h3cca6846),
	.w3(32'hbc353821),
	.w4(32'h3b3dda97),
	.w5(32'hbbeafcf4),
	.w6(32'hbc113d30),
	.w7(32'h3cc1ec44),
	.w8(32'hbd8d5a5f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd398e9d),
	.w1(32'h39e93e46),
	.w2(32'hba97ef1c),
	.w3(32'hbaa90924),
	.w4(32'h3a7b6820),
	.w5(32'h3b484c68),
	.w6(32'hbad49211),
	.w7(32'hbaa637be),
	.w8(32'h3aee1a6b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5c477),
	.w1(32'h3bb0b413),
	.w2(32'h3b2d29f4),
	.w3(32'hba3bfd89),
	.w4(32'hbb7cc8b0),
	.w5(32'hbb873db4),
	.w6(32'hbb3df419),
	.w7(32'hbc199097),
	.w8(32'hba9517ac),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd2a67),
	.w1(32'h3c650a0c),
	.w2(32'hbc0bf030),
	.w3(32'h3b8205de),
	.w4(32'hbc6ab49c),
	.w5(32'h3c76a23e),
	.w6(32'hba810d8c),
	.w7(32'hbcf9f98b),
	.w8(32'h3c5f07ad),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd798e),
	.w1(32'h3bfe6548),
	.w2(32'hbc832788),
	.w3(32'hbc59c29c),
	.w4(32'h3c4f5faa),
	.w5(32'hbc383011),
	.w6(32'hba1b6437),
	.w7(32'h3cad188d),
	.w8(32'hbcfe387f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbea3fa),
	.w1(32'hbb85953a),
	.w2(32'hbb297a7a),
	.w3(32'hb910690a),
	.w4(32'h3bc42c42),
	.w5(32'h3b51bf2e),
	.w6(32'hbbbca075),
	.w7(32'h3a2005b6),
	.w8(32'hbb53f61c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e146ad),
	.w1(32'h3c56d978),
	.w2(32'hbb959744),
	.w3(32'h3b26f1b2),
	.w4(32'hbbf5a34b),
	.w5(32'hbca60e6e),
	.w6(32'hb8070327),
	.w7(32'hbc273784),
	.w8(32'hbd1e27e8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca08f74),
	.w1(32'hba5d6bc0),
	.w2(32'h3c0a52db),
	.w3(32'hbaac2ee4),
	.w4(32'h3bc35c56),
	.w5(32'h3b95fe51),
	.w6(32'hbb3dab9e),
	.w7(32'h3c08bc03),
	.w8(32'hbac05919),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060178),
	.w1(32'h3ac7a411),
	.w2(32'h3c1f1793),
	.w3(32'hbb51fb4a),
	.w4(32'h3c38dc75),
	.w5(32'hbb4abebd),
	.w6(32'h39ff0e17),
	.w7(32'h3c2a6e31),
	.w8(32'h395255d2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42837),
	.w1(32'hbb0b3efa),
	.w2(32'hbb6cfbe8),
	.w3(32'hbbc60710),
	.w4(32'hbc44979b),
	.w5(32'hbb840ce7),
	.w6(32'hbc16a8e6),
	.w7(32'hbc5167bf),
	.w8(32'hbacdb4da),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63274d),
	.w1(32'h3b72c990),
	.w2(32'h39476a0a),
	.w3(32'hbb582441),
	.w4(32'hbb2ed505),
	.w5(32'hb97801f3),
	.w6(32'h3a64957f),
	.w7(32'hbaefce66),
	.w8(32'hba8cba0f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac16e40),
	.w1(32'hba2e38dc),
	.w2(32'hb9bf405c),
	.w3(32'h3b398aee),
	.w4(32'h3708face),
	.w5(32'h3ba041d5),
	.w6(32'h3b3ff8f6),
	.w7(32'hbae25ec2),
	.w8(32'h3b9e92af),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb821f70),
	.w1(32'hbc392548),
	.w2(32'h3b91ecee),
	.w3(32'h391b1486),
	.w4(32'h3bb256a3),
	.w5(32'h3be17b07),
	.w6(32'hbc26cf96),
	.w7(32'h3be99b4a),
	.w8(32'h3c3a5015),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca29c6c),
	.w1(32'hb9cac4e9),
	.w2(32'hb9ac6946),
	.w3(32'hb9d598ac),
	.w4(32'hba8a44e2),
	.w5(32'hbb3ed69a),
	.w6(32'h3aba72f7),
	.w7(32'hbb373830),
	.w8(32'h375e3130),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadea9f8),
	.w1(32'h3b4a4a8b),
	.w2(32'h3b5fbd6b),
	.w3(32'h3bb48b40),
	.w4(32'h3bf6c300),
	.w5(32'h3bc899fa),
	.w6(32'h3bc8e59f),
	.w7(32'h3b8ef14d),
	.w8(32'h3b2e9aaa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc4c1b),
	.w1(32'h3c57e827),
	.w2(32'h3b568986),
	.w3(32'hbc835b3e),
	.w4(32'h3d3473d4),
	.w5(32'hbb8c5d51),
	.w6(32'hbbb43d32),
	.w7(32'h3d5c9c00),
	.w8(32'hbc5366d7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3f508),
	.w1(32'h3a688f27),
	.w2(32'h3a477746),
	.w3(32'h39a15d8b),
	.w4(32'hbaea0438),
	.w5(32'hbb1725ac),
	.w6(32'hbaaa0ee0),
	.w7(32'hbac6f39c),
	.w8(32'hbab36a63),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf59aaa),
	.w1(32'hbc497e07),
	.w2(32'hbaf308f2),
	.w3(32'h3b4211b1),
	.w4(32'h3b3fc81d),
	.w5(32'hba769c92),
	.w6(32'h38cfbe70),
	.w7(32'h3c0485ce),
	.w8(32'hbb8cb1e3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0add2b),
	.w1(32'hbc3f5a8e),
	.w2(32'h3b1c9878),
	.w3(32'h3ae9c244),
	.w4(32'hbb38e981),
	.w5(32'h3c922b60),
	.w6(32'hbbd7f39f),
	.w7(32'hbae97b5c),
	.w8(32'h3b6a4423),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d3d53),
	.w1(32'h3c138a13),
	.w2(32'h39ce127b),
	.w3(32'h3b7af0ab),
	.w4(32'h3d0b0941),
	.w5(32'h3c229d17),
	.w6(32'h3b1678e4),
	.w7(32'hb91094ad),
	.w8(32'h3b5b4f2a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8ffa5),
	.w1(32'hbc44281d),
	.w2(32'hbc63768c),
	.w3(32'h3c62113c),
	.w4(32'hbc1b2645),
	.w5(32'hbc1b68c8),
	.w6(32'h3c907624),
	.w7(32'hbbee13fc),
	.w8(32'hbbc79c82),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7d49b),
	.w1(32'hbc843e2d),
	.w2(32'hbb5c2553),
	.w3(32'hbc8d88f1),
	.w4(32'hbb0b397b),
	.w5(32'hbb8d62fc),
	.w6(32'hbc535972),
	.w7(32'h3b273b7f),
	.w8(32'hbae70877),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe35897),
	.w1(32'hba7940b9),
	.w2(32'h3af342c2),
	.w3(32'h3aa51e46),
	.w4(32'hba0424be),
	.w5(32'hbb8dfbfe),
	.w6(32'h3b706aee),
	.w7(32'hbbbb07e3),
	.w8(32'hbbd71760),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6145),
	.w1(32'hbab47d81),
	.w2(32'h39f400e5),
	.w3(32'hbb718c7b),
	.w4(32'hba7cfe6b),
	.w5(32'hbb9ef3a3),
	.w6(32'hba88a631),
	.w7(32'hbb94e1fe),
	.w8(32'hbb50ec5f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87d8f5),
	.w1(32'h3978f131),
	.w2(32'h39cb761c),
	.w3(32'h3b869d3b),
	.w4(32'h39ba5aec),
	.w5(32'hbb6bf415),
	.w6(32'h3b04a074),
	.w7(32'h3865f983),
	.w8(32'hbb4381ca),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd050ab),
	.w1(32'hbd1718cf),
	.w2(32'hbd1a0058),
	.w3(32'hbce5e2f2),
	.w4(32'hbc9f44a3),
	.w5(32'hbcfb2d1d),
	.w6(32'hb9814e51),
	.w7(32'hbbbf1cc6),
	.w8(32'h3c49daed),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c948f70),
	.w1(32'hbc178524),
	.w2(32'h3c468bc1),
	.w3(32'hbbf4c91e),
	.w4(32'hbbfcc599),
	.w5(32'hbc466834),
	.w6(32'hbbcb160d),
	.w7(32'h3c6f6f7e),
	.w8(32'hbd01e33f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc809744),
	.w1(32'hbc691ce2),
	.w2(32'h3c810316),
	.w3(32'h3be0db3e),
	.w4(32'hbc73f8bb),
	.w5(32'hbc2d6ee1),
	.w6(32'hba9eae64),
	.w7(32'hbb610ced),
	.w8(32'hbc759ed8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ba0e0),
	.w1(32'hbbe6afb5),
	.w2(32'hbc994203),
	.w3(32'hbc030894),
	.w4(32'hbc1f1aa2),
	.w5(32'h3ca665e6),
	.w6(32'hba7464aa),
	.w7(32'hbcf02172),
	.w8(32'h3d24b3ec),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fceb3),
	.w1(32'hbb6eceaf),
	.w2(32'h3d1544dc),
	.w3(32'hbb1de8dd),
	.w4(32'h3d177b09),
	.w5(32'h3cce7120),
	.w6(32'hbca7b066),
	.w7(32'h3d8d4743),
	.w8(32'h3d580f00),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed79b6),
	.w1(32'h3a58c00b),
	.w2(32'h3ba65fff),
	.w3(32'h3b38c5e7),
	.w4(32'h3c0071ce),
	.w5(32'h3b80ef07),
	.w6(32'h3a9be8f9),
	.w7(32'h3bf8ce25),
	.w8(32'h37c736c6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5dec6),
	.w1(32'hbb972a27),
	.w2(32'hbb8262e4),
	.w3(32'hbb01173a),
	.w4(32'hbbff18ad),
	.w5(32'h3c4bb712),
	.w6(32'hba8c734f),
	.w7(32'h3b205850),
	.w8(32'h3c445a1f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a73d8),
	.w1(32'h3b00d0d6),
	.w2(32'h3b7e96ba),
	.w3(32'hbb8fb1a7),
	.w4(32'h3bd2eaf6),
	.w5(32'h3ad34245),
	.w6(32'hbb6e4421),
	.w7(32'h3b14efe4),
	.w8(32'hbbad28f3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1765f6),
	.w1(32'hbb0a494c),
	.w2(32'h3a5827e6),
	.w3(32'hb9d34681),
	.w4(32'h3aa3b4a0),
	.w5(32'hbb17be35),
	.w6(32'h3af87b9d),
	.w7(32'h3b99fa9f),
	.w8(32'hbb97d469),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167798),
	.w1(32'h3b78b93f),
	.w2(32'hbc585c05),
	.w3(32'hbb11020a),
	.w4(32'h3ab94cf8),
	.w5(32'hbac859cb),
	.w6(32'hb9e9bb43),
	.w7(32'h3b80896d),
	.w8(32'hbc4e872d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb5242),
	.w1(32'h3ca5ddbd),
	.w2(32'hbcc1ef2e),
	.w3(32'h3c01f4aa),
	.w4(32'h3d7b93f5),
	.w5(32'hbd13d948),
	.w6(32'h3c54d5fc),
	.w7(32'h3c346c89),
	.w8(32'hbc2bc41d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d883119),
	.w1(32'hbaecf51b),
	.w2(32'h3cbbc2b7),
	.w3(32'h3c34a5e8),
	.w4(32'hbc4b8966),
	.w5(32'hbbe607d5),
	.w6(32'h3bc5fcb5),
	.w7(32'h3c04c657),
	.w8(32'hbca215fe),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd24463e),
	.w1(32'hb9133f8c),
	.w2(32'h3a404ad4),
	.w3(32'h3a89850c),
	.w4(32'h3a404914),
	.w5(32'hb99b0cdd),
	.w6(32'h3b3ac214),
	.w7(32'h3a9df222),
	.w8(32'h3a7b2142),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93dd446),
	.w1(32'hb90a8f73),
	.w2(32'h3a487d62),
	.w3(32'h3a3e3b62),
	.w4(32'h3a9d0f19),
	.w5(32'h3b9423f2),
	.w6(32'hbbd48323),
	.w7(32'h3afc3efb),
	.w8(32'hbaef8349),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc1daa),
	.w1(32'hbc0c0fcd),
	.w2(32'hbc875ef1),
	.w3(32'hbc590092),
	.w4(32'hbc59d07d),
	.w5(32'hbbd35454),
	.w6(32'h3bfc4a38),
	.w7(32'h3bf539b8),
	.w8(32'h38c98ac8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bee0),
	.w1(32'h39c45c0d),
	.w2(32'h3b0fbc9d),
	.w3(32'h3ba40cac),
	.w4(32'h3bb0a30b),
	.w5(32'h3ae14dfe),
	.w6(32'h3b424fe1),
	.w7(32'hb9a97bde),
	.w8(32'hba87a08f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca68df),
	.w1(32'h3b42177d),
	.w2(32'hbcd9f4df),
	.w3(32'h38c756c4),
	.w4(32'hbc7650f5),
	.w5(32'hbca68cf8),
	.w6(32'hbaa428ee),
	.w7(32'hbccb5d24),
	.w8(32'hbd037d86),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbafc7d),
	.w1(32'h3bb3cda5),
	.w2(32'hbbb86b9f),
	.w3(32'hbbdabf55),
	.w4(32'hbb9a5f8e),
	.w5(32'hbc7e620f),
	.w6(32'hbb0c71e1),
	.w7(32'hbc3f150a),
	.w8(32'hbbb9a2d5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf55903),
	.w1(32'hba7c950f),
	.w2(32'hbc99a859),
	.w3(32'hbc80dc4b),
	.w4(32'h3d022ad2),
	.w5(32'hbc566d32),
	.w6(32'hbb01b693),
	.w7(32'h3d05f4c8),
	.w8(32'h3c924a8b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1bc572),
	.w1(32'h3b642249),
	.w2(32'hbaea425e),
	.w3(32'hba850b08),
	.w4(32'hbb47b940),
	.w5(32'hba83ff61),
	.w6(32'h3ab74dae),
	.w7(32'hbb0f50ca),
	.w8(32'hbb48ff09),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ab4d),
	.w1(32'hbb9fbb01),
	.w2(32'hbbf38563),
	.w3(32'h3b91b1ab),
	.w4(32'hbc3dbe7f),
	.w5(32'h3d1e7d1e),
	.w6(32'h3b7c999a),
	.w7(32'hbcb473d2),
	.w8(32'h3d4d0fe6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0218b0),
	.w1(32'h3be85e63),
	.w2(32'h3bac7f1d),
	.w3(32'h3b7e7d5b),
	.w4(32'h3b904867),
	.w5(32'hb9482590),
	.w6(32'h3bb188f0),
	.w7(32'h3a8d1b68),
	.w8(32'h3ad52168),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2f70d),
	.w1(32'h3c84a518),
	.w2(32'h3b4735ca),
	.w3(32'h3c1021d9),
	.w4(32'h3be07faf),
	.w5(32'h3b99ab74),
	.w6(32'h3c1ad343),
	.w7(32'hb93f0f23),
	.w8(32'h3ab3da5c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e201e),
	.w1(32'h3bbc0759),
	.w2(32'h3b998eb0),
	.w3(32'h3c56924a),
	.w4(32'h3bdf7c2e),
	.w5(32'h3c0ba47c),
	.w6(32'h3c8fe1e1),
	.w7(32'h3c11003d),
	.w8(32'h3c0b2d02),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be586ac),
	.w1(32'h3ba736b6),
	.w2(32'h3b6ed95a),
	.w3(32'h3c233e0a),
	.w4(32'h3bcce647),
	.w5(32'h3a539ea0),
	.w6(32'h3c242873),
	.w7(32'h3b8d295c),
	.w8(32'h3acd4ca4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf61f1b),
	.w1(32'h3c25a269),
	.w2(32'h3be136f1),
	.w3(32'h3c4d3b0c),
	.w4(32'h3c383291),
	.w5(32'h3bd6bdfa),
	.w6(32'h3c018d15),
	.w7(32'h3bd49248),
	.w8(32'h3bf1962b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde68fb),
	.w1(32'hbc1bc197),
	.w2(32'h3abb3750),
	.w3(32'hbb2b5198),
	.w4(32'hbc83391b),
	.w5(32'hbcc783df),
	.w6(32'h3c94d6e5),
	.w7(32'h3c448784),
	.w8(32'hbb4d290c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06393b),
	.w1(32'h3b57de90),
	.w2(32'h3b9c0c3c),
	.w3(32'h3b8ca3e6),
	.w4(32'h3c296fe0),
	.w5(32'h3bef7b48),
	.w6(32'hbb83639c),
	.w7(32'hb99aa413),
	.w8(32'h3b43f2c5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c1f2b),
	.w1(32'h3c0f69db),
	.w2(32'h3cd4e24f),
	.w3(32'hbb6d6036),
	.w4(32'hbc7e47c1),
	.w5(32'hbba160fd),
	.w6(32'h3cc09876),
	.w7(32'h3d1db75a),
	.w8(32'h3c679a7a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49a769),
	.w1(32'hba908ad7),
	.w2(32'h3a89c033),
	.w3(32'hbac78360),
	.w4(32'hbb7f658b),
	.w5(32'hbb993128),
	.w6(32'h3b59082d),
	.w7(32'h3b3083b8),
	.w8(32'hb84ca447),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8549eb),
	.w1(32'hbd0613a1),
	.w2(32'hbd019000),
	.w3(32'h3c88e2eb),
	.w4(32'h3d0d57c9),
	.w5(32'h3cb637c7),
	.w6(32'h3bc0f096),
	.w7(32'h3cdc5afb),
	.w8(32'h3cc85c90),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826895),
	.w1(32'h3bb60d3a),
	.w2(32'h3b1066a9),
	.w3(32'hb9793e2d),
	.w4(32'hbb6e2196),
	.w5(32'hbb9c4ade),
	.w6(32'h3b55556f),
	.w7(32'h3af18542),
	.w8(32'h3a42d36c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddf70a),
	.w1(32'hbcd1e24f),
	.w2(32'hbca860d5),
	.w3(32'hbc98c6d1),
	.w4(32'hbcc78686),
	.w5(32'hbc35da82),
	.w6(32'h3aa5bbf2),
	.w7(32'h3c69b06d),
	.w8(32'h3c6aa203),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e8f16),
	.w1(32'hbbc22c4b),
	.w2(32'h3c124bdf),
	.w3(32'hbc9be578),
	.w4(32'hbbad3cbd),
	.w5(32'h3caaee2d),
	.w6(32'hbd386dc7),
	.w7(32'hbd42b524),
	.w8(32'hbd03571e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33df62),
	.w1(32'hbbe8d804),
	.w2(32'hbb179e9a),
	.w3(32'hbb8667fe),
	.w4(32'hbbe94334),
	.w5(32'hbb99b747),
	.w6(32'hb98344f6),
	.w7(32'h3bcb0915),
	.w8(32'h3b47084d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule