module layer_6_featuremap_18(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d5c8b),
	.w1(32'h3cce1271),
	.w2(32'h3d050464),
	.w3(32'hbd085ff3),
	.w4(32'h3c90a951),
	.w5(32'h3c9a652f),
	.w6(32'hbb85d3e1),
	.w7(32'h3c5c1729),
	.w8(32'hbd045628),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf4329),
	.w1(32'hbcf8d8d9),
	.w2(32'hbd0b8d09),
	.w3(32'hbb1fac1f),
	.w4(32'hbc99951c),
	.w5(32'hbca7e360),
	.w6(32'hbc28a3c4),
	.w7(32'hbc8e391b),
	.w8(32'hbb92a3ab),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b0d7b),
	.w1(32'hbd78e5ca),
	.w2(32'hbd8f8b29),
	.w3(32'hbc144e39),
	.w4(32'hbc35738a),
	.w5(32'hbc1f6fad),
	.w6(32'h3c4ce16b),
	.w7(32'h3cb46235),
	.w8(32'h3ca2ab2e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf746),
	.w1(32'h3ccfc173),
	.w2(32'h3c4c9410),
	.w3(32'hbc00f942),
	.w4(32'hbc5bd5cc),
	.w5(32'hbd188d1f),
	.w6(32'h3c56c521),
	.w7(32'hbc4f8b5e),
	.w8(32'hbc726bd4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0b63e5),
	.w1(32'h3b3c5fcf),
	.w2(32'hbc561983),
	.w3(32'hba20b877),
	.w4(32'h3ba3b73b),
	.w5(32'hbbd974e1),
	.w6(32'h3c96c35b),
	.w7(32'h3b8de7fd),
	.w8(32'hbabf40d4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9555c0),
	.w1(32'hbb0444fd),
	.w2(32'hbd45c4fc),
	.w3(32'hbbe5bfcb),
	.w4(32'h3c944583),
	.w5(32'h3c9eef4e),
	.w6(32'h3ce555dd),
	.w7(32'h3cb0ea85),
	.w8(32'hbb159ab8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b09ac),
	.w1(32'h3c06d316),
	.w2(32'h3c5f93cd),
	.w3(32'h3bc965b5),
	.w4(32'h3aa1c7e0),
	.w5(32'hbafa885b),
	.w6(32'hbb98f70d),
	.w7(32'h3bf48ac2),
	.w8(32'h3b12a499),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe3d52),
	.w1(32'h3c635c3f),
	.w2(32'h38c5576c),
	.w3(32'hbbea506c),
	.w4(32'h3c2ec2e3),
	.w5(32'h3bf866ec),
	.w6(32'h3be88b10),
	.w7(32'hbb9f47ac),
	.w8(32'h3c3a15ca),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964265b),
	.w1(32'hbcee6ebc),
	.w2(32'hbd249f3e),
	.w3(32'hbc51a3a6),
	.w4(32'hbc36143e),
	.w5(32'hbc99484a),
	.w6(32'h3c49717f),
	.w7(32'hbc3d5ac9),
	.w8(32'hbc0bddde),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc34514),
	.w1(32'h3be22ffb),
	.w2(32'h3b764468),
	.w3(32'h3cb578db),
	.w4(32'hb9d51c59),
	.w5(32'hbc067362),
	.w6(32'h3ac7dadb),
	.w7(32'h3c03cc6b),
	.w8(32'h3ab42631),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6681de),
	.w1(32'h39b07eb3),
	.w2(32'hbcfeefd9),
	.w3(32'hbbadcd33),
	.w4(32'h3aa1d96c),
	.w5(32'hbb4bc1e6),
	.w6(32'h3c0632ea),
	.w7(32'h3c2b1d0b),
	.w8(32'h3c942bb0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb108),
	.w1(32'hbd768c17),
	.w2(32'hbe48449f),
	.w3(32'h388d122a),
	.w4(32'hbcc82526),
	.w5(32'h3ddf696b),
	.w6(32'h3b74c644),
	.w7(32'hbcd8148f),
	.w8(32'hbd4f5120),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e3f1c29),
	.w1(32'h3c66a737),
	.w2(32'hbda845f4),
	.w3(32'hbca718de),
	.w4(32'h3bc7f6c7),
	.w5(32'h3ae34ae6),
	.w6(32'h3c807660),
	.w7(32'hbbf692e8),
	.w8(32'hbbde30a4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c4e3f),
	.w1(32'hbc5923cb),
	.w2(32'hbd399901),
	.w3(32'hbd4ca863),
	.w4(32'h3c80ab5e),
	.w5(32'h3c84c21f),
	.w6(32'h3b7458d2),
	.w7(32'h3c7ca962),
	.w8(32'hbca423d3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eb2a2),
	.w1(32'h3c822503),
	.w2(32'hbd645628),
	.w3(32'h3d24df0a),
	.w4(32'h3d075196),
	.w5(32'hbc6319d7),
	.w6(32'h3bc51b1d),
	.w7(32'hbc92b1d0),
	.w8(32'hbc000311),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd097a31),
	.w1(32'h3c40bfa7),
	.w2(32'hbcd48ef4),
	.w3(32'hbd425538),
	.w4(32'h3c5a71fb),
	.w5(32'hbc289f9d),
	.w6(32'h3ca8cb5f),
	.w7(32'h3d3e12a4),
	.w8(32'h3cfc8054),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd09ae7d),
	.w1(32'hbcffa466),
	.w2(32'h3bf39dfe),
	.w3(32'hbd04dbd2),
	.w4(32'hbd561eba),
	.w5(32'h3c3278d7),
	.w6(32'h3cebbdc5),
	.w7(32'h3d5ff47e),
	.w8(32'h3cf96afb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d6c59),
	.w1(32'hbbe9ce0d),
	.w2(32'h3c4be52f),
	.w3(32'h3b97f036),
	.w4(32'h3c884722),
	.w5(32'h3cd84f67),
	.w6(32'hbc8ce0d6),
	.w7(32'hbc4c5d87),
	.w8(32'hbca22b88),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12a75c),
	.w1(32'h3c342b13),
	.w2(32'hbc89dda7),
	.w3(32'h3b806715),
	.w4(32'hbbd79860),
	.w5(32'hbb718bbb),
	.w6(32'h3be1fd8f),
	.w7(32'hbc91c8c3),
	.w8(32'hbbbcae98),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3affc0aa),
	.w1(32'hbc2efbc5),
	.w2(32'hbc2ca2b1),
	.w3(32'h3addf3e6),
	.w4(32'hbc938c98),
	.w5(32'hbcbbed64),
	.w6(32'h3c0dc64f),
	.w7(32'h3d0ab2a8),
	.w8(32'h3c23f078),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b9d7b),
	.w1(32'h3bc60bbe),
	.w2(32'h3b835792),
	.w3(32'hbcb46dc9),
	.w4(32'hbbbd2825),
	.w5(32'h3b7c55c7),
	.w6(32'h3ba4502e),
	.w7(32'h3cf72e0f),
	.w8(32'hbc3cbc79),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1548cc),
	.w1(32'hbd0e6712),
	.w2(32'hbd1db852),
	.w3(32'hbcba3c14),
	.w4(32'hbcf88da7),
	.w5(32'hbcc188ab),
	.w6(32'h3c3df167),
	.w7(32'hbb9a0eb5),
	.w8(32'hbc225e02),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3ab0ea),
	.w1(32'hbbe6dea9),
	.w2(32'hbd0479cc),
	.w3(32'h3b72372d),
	.w4(32'hbc0dd880),
	.w5(32'h3bf27870),
	.w6(32'hbad9fb84),
	.w7(32'hbb8f8eb7),
	.w8(32'hbba5bd44),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f2b38),
	.w1(32'hbd186a18),
	.w2(32'hbe00b09b),
	.w3(32'hbcedf158),
	.w4(32'h3b17ee0a),
	.w5(32'hbd7ad778),
	.w6(32'hbd021b78),
	.w7(32'hbc284669),
	.w8(32'hbc4972dc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37dcec),
	.w1(32'hbcb6475d),
	.w2(32'hbbf4e8da),
	.w3(32'hbd75def1),
	.w4(32'hbdb50c62),
	.w5(32'hbda48c0b),
	.w6(32'hbc8ee563),
	.w7(32'hbd185f86),
	.w8(32'hbd8ce939),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb0b8c),
	.w1(32'h3d3d3470),
	.w2(32'hbe7423a9),
	.w3(32'hbaf4838c),
	.w4(32'hbe1d2598),
	.w5(32'hbda039d4),
	.w6(32'h3d1e531e),
	.w7(32'hbd61bc40),
	.w8(32'hbe3089d5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd18d9d),
	.w1(32'h3c4d1b4b),
	.w2(32'hbda07846),
	.w3(32'hbd9c8a7e),
	.w4(32'h3ce3b753),
	.w5(32'hbbc0a361),
	.w6(32'h3caa8b8d),
	.w7(32'hbcae10ae),
	.w8(32'hbc59885f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd59bce8),
	.w1(32'hbc57a322),
	.w2(32'hbd2c5a20),
	.w3(32'hbcc3e772),
	.w4(32'h3b160f23),
	.w5(32'hbd091eab),
	.w6(32'h3cf38516),
	.w7(32'h3cd71307),
	.w8(32'hbb48d48d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30dc79),
	.w1(32'h3ca8a6cd),
	.w2(32'hbd2d8c2b),
	.w3(32'hbcb36d9a),
	.w4(32'h3d212386),
	.w5(32'h3cac67ba),
	.w6(32'h3c487272),
	.w7(32'hbc3ac1cb),
	.w8(32'h3b0d7dc9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe0258a2),
	.w1(32'h3da91f11),
	.w2(32'h3d238edf),
	.w3(32'h3ceee861),
	.w4(32'h3daec48e),
	.w5(32'h3c77d18f),
	.w6(32'h3d0427db),
	.w7(32'hbe519d44),
	.w8(32'hbddff6ba),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef444),
	.w1(32'h3bd83898),
	.w2(32'h3b89cdb8),
	.w3(32'h3c189929),
	.w4(32'h3b8ac261),
	.w5(32'h3b376287),
	.w6(32'h3c40c10b),
	.w7(32'h3be2b0ca),
	.w8(32'h3bbdeb57),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1102d7),
	.w1(32'hbc42ccdb),
	.w2(32'hbb0e1782),
	.w3(32'hbc4f09c0),
	.w4(32'hbc774b45),
	.w5(32'hbb304aff),
	.w6(32'hba9c2eb0),
	.w7(32'hbb18190d),
	.w8(32'hba176c7c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8a95d),
	.w1(32'hbb960ff0),
	.w2(32'hbbe908a3),
	.w3(32'hbbcbb7d5),
	.w4(32'hba8f5c62),
	.w5(32'hbc27a232),
	.w6(32'hbacfe381),
	.w7(32'h3aea7a33),
	.w8(32'hbb98d3a6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ecfde),
	.w1(32'hbb636870),
	.w2(32'hbb158e35),
	.w3(32'hbc049d59),
	.w4(32'hbb5c60cc),
	.w5(32'hbb053cfa),
	.w6(32'hbac9c76e),
	.w7(32'h39eabfcb),
	.w8(32'h3ad2db08),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b8a19),
	.w1(32'hba4cfb8d),
	.w2(32'hbbaf11cf),
	.w3(32'hbb024e40),
	.w4(32'hba4d69a2),
	.w5(32'hbb87e566),
	.w6(32'hbaa126f0),
	.w7(32'hbb7d19e6),
	.w8(32'h3b2bd0e9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc941de2),
	.w1(32'h3b8dbab7),
	.w2(32'hbc1899c1),
	.w3(32'hba93754b),
	.w4(32'hbc2db25e),
	.w5(32'hbb059e56),
	.w6(32'h3c096f72),
	.w7(32'hbd2aee39),
	.w8(32'hbd52ada1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266443),
	.w1(32'h3bbfc194),
	.w2(32'hb7ddf235),
	.w3(32'h3c0ed910),
	.w4(32'h3b77b08e),
	.w5(32'h3b9eb718),
	.w6(32'h3b84958e),
	.w7(32'hbb30edbf),
	.w8(32'hba64cd40),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c249404),
	.w1(32'h3c37ef50),
	.w2(32'h3c5a1cf9),
	.w3(32'h3c89416f),
	.w4(32'h3c26216c),
	.w5(32'h3cb7c12d),
	.w6(32'h3c200d59),
	.w7(32'hbb4c62b6),
	.w8(32'hbc0fecfa),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d10c0),
	.w1(32'hbb9e9901),
	.w2(32'hbb51bc00),
	.w3(32'h3a2200a2),
	.w4(32'hbbd30a41),
	.w5(32'hbbacb379),
	.w6(32'hbb9d962a),
	.w7(32'hbb641ffa),
	.w8(32'hbb86c84d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2241dd),
	.w1(32'hbd9794d1),
	.w2(32'h3bc44a16),
	.w3(32'hbcd8dc55),
	.w4(32'hbc83f8e3),
	.w5(32'h3c9b19df),
	.w6(32'h3d2d933c),
	.w7(32'h3dadd592),
	.w8(32'h3d4b1bc4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf2e4f5),
	.w1(32'h3d1fbe0e),
	.w2(32'h3cbf6a8b),
	.w3(32'h3cb3100c),
	.w4(32'h3c934b4d),
	.w5(32'h3c04f096),
	.w6(32'h3cdba278),
	.w7(32'h3cee3966),
	.w8(32'h3c641a80),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c635317),
	.w1(32'h3c87bea2),
	.w2(32'h3bea3eef),
	.w3(32'h3c431007),
	.w4(32'hba8419d1),
	.w5(32'h3b717884),
	.w6(32'hbc1978e0),
	.w7(32'hbccd1b0a),
	.w8(32'hbc7b3457),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac06987),
	.w1(32'hbbcce4a0),
	.w2(32'hbc1d394f),
	.w3(32'hbaf7d8e0),
	.w4(32'hbb835c9e),
	.w5(32'hbb4d61cd),
	.w6(32'hbbb380d9),
	.w7(32'hbc2070c8),
	.w8(32'hbb61954f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd146ba0),
	.w1(32'h3dc346e0),
	.w2(32'h3d8437e6),
	.w3(32'h3d5033fe),
	.w4(32'h3d740d21),
	.w5(32'h3d542455),
	.w6(32'h3d6789ee),
	.w7(32'hbe0e08b8),
	.w8(32'hbe072bf4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd16e4a0),
	.w1(32'hbd7c42b8),
	.w2(32'hbcf31b53),
	.w3(32'hbcdaa29a),
	.w4(32'hbd173df6),
	.w5(32'hbc88c50f),
	.w6(32'h3bcf7bb1),
	.w7(32'h3cd20ba6),
	.w8(32'h3cc600c0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb257708),
	.w1(32'hbc0b460d),
	.w2(32'hbc0b48eb),
	.w3(32'hbb751e7b),
	.w4(32'hbc185352),
	.w5(32'hbc3b6607),
	.w6(32'hbc0d2196),
	.w7(32'hbc390655),
	.w8(32'hbc41a09f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1016d1),
	.w1(32'hbab8c1c9),
	.w2(32'hba987e37),
	.w3(32'hbc1c6fa9),
	.w4(32'hbc0a4dae),
	.w5(32'hbc088255),
	.w6(32'hba166be6),
	.w7(32'h3adb6506),
	.w8(32'hba9af1a9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf7baa4),
	.w1(32'hbcb5c8c5),
	.w2(32'hbc709aa7),
	.w3(32'hbd3f3110),
	.w4(32'hbd3587c7),
	.w5(32'hbcb8d7f1),
	.w6(32'hbcd99eaa),
	.w7(32'hbd6bde5b),
	.w8(32'hbd0c41e3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b925875),
	.w1(32'h3c901938),
	.w2(32'h3cce4a54),
	.w3(32'h3be91a19),
	.w4(32'h3cc24e09),
	.w5(32'h3cd02531),
	.w6(32'h3ca11301),
	.w7(32'h3cd9bd65),
	.w8(32'h3c761a1b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3332),
	.w1(32'hbca0545d),
	.w2(32'hbcc99f96),
	.w3(32'hbb0ef1db),
	.w4(32'hbb7e0576),
	.w5(32'hbcb89e09),
	.w6(32'h3ca0776b),
	.w7(32'h3bbfdb92),
	.w8(32'h3af3446c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813ec1),
	.w1(32'h3c58690d),
	.w2(32'h3c329787),
	.w3(32'h3b1531ce),
	.w4(32'hbc0fd392),
	.w5(32'hbbb82a64),
	.w6(32'h3c3f68b8),
	.w7(32'h3b64023a),
	.w8(32'h3ad89375),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2be457),
	.w1(32'h3c89efd2),
	.w2(32'h3b1cd79d),
	.w3(32'h3d1116b5),
	.w4(32'h3b973bc2),
	.w5(32'hbb2d45a4),
	.w6(32'h3c143764),
	.w7(32'h3c32037b),
	.w8(32'hbbd6ab2a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2b7973),
	.w1(32'hbd7c66b5),
	.w2(32'hbd01f868),
	.w3(32'hbd8f2fbb),
	.w4(32'hbd819b33),
	.w5(32'hbca22483),
	.w6(32'hbccc2d5a),
	.w7(32'h3ca399dc),
	.w8(32'h3c3d482c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2a41b),
	.w1(32'h3d2a6ce8),
	.w2(32'h3d07ba18),
	.w3(32'h3cfc9e16),
	.w4(32'h3d2ea262),
	.w5(32'h3d1bd945),
	.w6(32'h3d5753c0),
	.w7(32'h3d40e576),
	.w8(32'h3d4c3a9b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca52356),
	.w1(32'hbb4b5297),
	.w2(32'hbb90c5d8),
	.w3(32'h3cc980aa),
	.w4(32'h3b188d72),
	.w5(32'hbb96025f),
	.w6(32'h3b6694ca),
	.w7(32'h3b466015),
	.w8(32'h3be10037),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bcba7),
	.w1(32'h3c8a2634),
	.w2(32'h3baad6ab),
	.w3(32'hbc8e425d),
	.w4(32'hbca8a464),
	.w5(32'hbc8f731c),
	.w6(32'hbc232f35),
	.w7(32'hbd10cf68),
	.w8(32'hbd0505ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbc50e),
	.w1(32'h3bcb9234),
	.w2(32'h3b8f049a),
	.w3(32'h3b8588b6),
	.w4(32'h3c0862f9),
	.w5(32'h3c356c3e),
	.w6(32'h3b86aad1),
	.w7(32'h3c169156),
	.w8(32'h3bf299d8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f349b),
	.w1(32'h3b047989),
	.w2(32'h3b90cbd1),
	.w3(32'h3812b1f8),
	.w4(32'hba673aee),
	.w5(32'h3ba56d57),
	.w6(32'hbb610cf1),
	.w7(32'hbb936bad),
	.w8(32'hbae7b8d2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c782e3e),
	.w1(32'h3bff325d),
	.w2(32'h3c08847e),
	.w3(32'h3cb69f66),
	.w4(32'h3bd2c029),
	.w5(32'h3bd0fe9d),
	.w6(32'h3bbfd248),
	.w7(32'h3c6ce75c),
	.w8(32'h3bfaaafc),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c1329),
	.w1(32'hbd329814),
	.w2(32'hbd514fde),
	.w3(32'hbc8a79b5),
	.w4(32'hbd4d0dcf),
	.w5(32'hbd896616),
	.w6(32'h3b7670ee),
	.w7(32'h3cbe21d2),
	.w8(32'hbc6cfa98),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb452a3),
	.w1(32'hbbe4a9a2),
	.w2(32'hbc768f2f),
	.w3(32'hbbe6d230),
	.w4(32'hbc8fbdc5),
	.w5(32'hbcab9af0),
	.w6(32'h3af251ef),
	.w7(32'hbbc4b790),
	.w8(32'hbc13bb38),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ee9d1),
	.w1(32'h3c2ebfe6),
	.w2(32'h3ba77acd),
	.w3(32'hbcb72e90),
	.w4(32'hbce8e83c),
	.w5(32'hbcbf3fa2),
	.w6(32'h3b3b2d5a),
	.w7(32'hbb37a34b),
	.w8(32'hbc9a639a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca86f3d),
	.w1(32'h3d3ce76b),
	.w2(32'hbd2d7909),
	.w3(32'h3d7c2203),
	.w4(32'h3dc55245),
	.w5(32'h3cf17ed7),
	.w6(32'h3d81e385),
	.w7(32'hbdfe0641),
	.w8(32'hbdffa39c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d94e),
	.w1(32'hba6c9109),
	.w2(32'hba6537c9),
	.w3(32'h3c0b5494),
	.w4(32'h3bf08c20),
	.w5(32'h3b738224),
	.w6(32'hba49931b),
	.w7(32'hbb424023),
	.w8(32'hbb32e9e5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule