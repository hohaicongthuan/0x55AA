module layer_10_featuremap_428(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30e7dd),
	.w1(32'hb9d6e8f2),
	.w2(32'hba13ffb1),
	.w3(32'h3940da26),
	.w4(32'hba334db1),
	.w5(32'h3844280d),
	.w6(32'h399b40cd),
	.w7(32'h39c64241),
	.w8(32'h39ef0322),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccbfd3),
	.w1(32'h3ac44139),
	.w2(32'h3b2a8956),
	.w3(32'h3a26e78e),
	.w4(32'h3b8b7729),
	.w5(32'h3b40031d),
	.w6(32'h3b2b8cd8),
	.w7(32'h3b77410b),
	.w8(32'h3b0986d3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c4fd1),
	.w1(32'hb9d0540a),
	.w2(32'hb9e26815),
	.w3(32'hba1ec2cb),
	.w4(32'h39d0360f),
	.w5(32'h3a57c707),
	.w6(32'hb91e9089),
	.w7(32'h390d3448),
	.w8(32'h38293088),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba157be1),
	.w1(32'hba174046),
	.w2(32'hbaa69299),
	.w3(32'h39bb9f04),
	.w4(32'hb8b4b1a9),
	.w5(32'hba2e6955),
	.w6(32'h39dab7be),
	.w7(32'h3a281a18),
	.w8(32'hba864903),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e2636),
	.w1(32'h3a066112),
	.w2(32'h39381ce2),
	.w3(32'hb8c321d6),
	.w4(32'h3a12a62c),
	.w5(32'h39ac69d4),
	.w6(32'hb9a21bf2),
	.w7(32'h3a054bf9),
	.w8(32'h3a090f49),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3844ceac),
	.w1(32'hba442be8),
	.w2(32'hb9a12e7d),
	.w3(32'h399bd9ac),
	.w4(32'hb9c0b725),
	.w5(32'hbaa2aff7),
	.w6(32'h39446d86),
	.w7(32'hba70817a),
	.w8(32'hba1b81dc),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f22c7),
	.w1(32'h3b56b642),
	.w2(32'h39c8a41b),
	.w3(32'h3b82a755),
	.w4(32'h3ab2dc9a),
	.w5(32'h39a2e3e3),
	.w6(32'h3b03a867),
	.w7(32'hba8191c8),
	.w8(32'hba9bbda4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87169c),
	.w1(32'hbb9bd1b4),
	.w2(32'hbc031949),
	.w3(32'hbc8836a2),
	.w4(32'hbc41b446),
	.w5(32'hbbe23573),
	.w6(32'hbbb2a343),
	.w7(32'hbc8a1a4e),
	.w8(32'hbc605158),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38922af1),
	.w1(32'hb9edaa10),
	.w2(32'hba80a56c),
	.w3(32'h3a4dc8d2),
	.w4(32'h3a444e10),
	.w5(32'hba81135c),
	.w6(32'h3ab6dc3e),
	.w7(32'h398bd58c),
	.w8(32'hba96bb21),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c174d9d),
	.w1(32'h3b635921),
	.w2(32'h3bdf5c63),
	.w3(32'h3ab90412),
	.w4(32'hba1d7008),
	.w5(32'h3b0872b1),
	.w6(32'hbb31d17e),
	.w7(32'hbbaba628),
	.w8(32'hbb13408e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61d290a),
	.w1(32'hb96428e2),
	.w2(32'hba29a48b),
	.w3(32'h381bdbb6),
	.w4(32'hba07719e),
	.w5(32'hba9009ca),
	.w6(32'hba006245),
	.w7(32'hba65521b),
	.w8(32'hba93977a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25dfbc),
	.w1(32'h3b8b2bee),
	.w2(32'hbb498513),
	.w3(32'h3af32ba9),
	.w4(32'h3a795ca7),
	.w5(32'hb9d9516d),
	.w6(32'h3b42afab),
	.w7(32'h3a7c149f),
	.w8(32'hbb0dcba3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5eafa8),
	.w1(32'h3baa01c8),
	.w2(32'h3c044874),
	.w3(32'hba2b6ebc),
	.w4(32'hbb99f395),
	.w5(32'hbb896e20),
	.w6(32'hbbf3d8b6),
	.w7(32'hbc80c4f9),
	.w8(32'hbc26ec6d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2db6c7),
	.w1(32'h3b31248a),
	.w2(32'h3a179102),
	.w3(32'h3b172816),
	.w4(32'h3b3df040),
	.w5(32'h3b1fe0db),
	.w6(32'h3aa998d6),
	.w7(32'h3a80ea0e),
	.w8(32'h3a26d475),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0f6f),
	.w1(32'h3b295b45),
	.w2(32'h3b51f768),
	.w3(32'h39b69162),
	.w4(32'h3b235b55),
	.w5(32'h3adece8c),
	.w6(32'h3b111bb8),
	.w7(32'h3b2f5458),
	.w8(32'h3a452766),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207d24),
	.w1(32'h3ab3d750),
	.w2(32'h3b2c7d3c),
	.w3(32'h3abe162c),
	.w4(32'hbb0da144),
	.w5(32'hba680347),
	.w6(32'hbb1260b0),
	.w7(32'hbb9d0c11),
	.w8(32'hbb8163d9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5ce2e),
	.w1(32'h3a701518),
	.w2(32'h39fe4262),
	.w3(32'h39825310),
	.w4(32'h3a5a14ee),
	.w5(32'hb8d0201a),
	.w6(32'h39294757),
	.w7(32'h3a44ee71),
	.w8(32'h3a119004),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc26154),
	.w1(32'hbbad772b),
	.w2(32'hbc091d3b),
	.w3(32'hbc09bcbe),
	.w4(32'hbc6eb782),
	.w5(32'hbc4595d1),
	.w6(32'hbc4153bf),
	.w7(32'hbcaf72e5),
	.w8(32'hbc8b4f15),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70fb0b),
	.w1(32'hbb482184),
	.w2(32'hbb3de2f4),
	.w3(32'hbb2921ee),
	.w4(32'hbbad75d6),
	.w5(32'hbbba857f),
	.w6(32'hbbd272a8),
	.w7(32'hbc592ed9),
	.w8(32'hbbfdf06e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba033f82),
	.w1(32'hb99855d4),
	.w2(32'h3a738a39),
	.w3(32'hb9a95ef0),
	.w4(32'hb9d3b746),
	.w5(32'h3866c7e9),
	.w6(32'hb85b06cc),
	.w7(32'h39ef6491),
	.w8(32'h3aa5036d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c028c),
	.w1(32'hba0598ee),
	.w2(32'h3980dabb),
	.w3(32'h392f8a50),
	.w4(32'h3915e806),
	.w5(32'h3a2c531d),
	.w6(32'h3a09f7cd),
	.w7(32'h39db1903),
	.w8(32'hb8d0e58b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1b2f5),
	.w1(32'h3981d9cf),
	.w2(32'h3aad263c),
	.w3(32'h3a85c79a),
	.w4(32'h3a5a19af),
	.w5(32'h3a18c364),
	.w6(32'hba1331bf),
	.w7(32'h3ae0288c),
	.w8(32'h3a86635e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83c81f),
	.w1(32'h3a0feef4),
	.w2(32'hb9bda5f4),
	.w3(32'h3b66686e),
	.w4(32'hbc483dad),
	.w5(32'hbc468c73),
	.w6(32'hbc4d892c),
	.w7(32'hbbd61c8a),
	.w8(32'hbc01dd08),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec44c8),
	.w1(32'h3bb6ab6f),
	.w2(32'h3c073c8a),
	.w3(32'h3b29d13a),
	.w4(32'h39a6e762),
	.w5(32'h3b511664),
	.w6(32'hba069781),
	.w7(32'h39f51e8b),
	.w8(32'h3b19fe0f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf4565),
	.w1(32'h3be1676a),
	.w2(32'h3c317977),
	.w3(32'hbb17b264),
	.w4(32'hba4886d5),
	.w5(32'h3bca07b8),
	.w6(32'h3abb077f),
	.w7(32'h3b862057),
	.w8(32'h3b8d957c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d5abd),
	.w1(32'hb9888240),
	.w2(32'h3a239a89),
	.w3(32'hba87f69c),
	.w4(32'hb9d3c691),
	.w5(32'hb8d4353b),
	.w6(32'hba96476a),
	.w7(32'h399f4c4f),
	.w8(32'h39c00f90),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba158d13),
	.w1(32'hba5e714c),
	.w2(32'hba5a8006),
	.w3(32'hb9ffdaa2),
	.w4(32'hba7040c6),
	.w5(32'hb8419bde),
	.w6(32'hb7b2c327),
	.w7(32'hba776efc),
	.w8(32'hb983802f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac71fc3),
	.w1(32'hbaeafc96),
	.w2(32'h3afff671),
	.w3(32'h3ae8ffda),
	.w4(32'hba4cc83b),
	.w5(32'h3a667dd9),
	.w6(32'h3a44cf5b),
	.w7(32'h3ab3acde),
	.w8(32'h3aa6f8fb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60ebe6),
	.w1(32'h382c1d96),
	.w2(32'h3b16e472),
	.w3(32'hba42bf42),
	.w4(32'h39814cfa),
	.w5(32'h39a08c07),
	.w6(32'hba5f9924),
	.w7(32'h3a4bf6b6),
	.w8(32'h3aaa54f8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7aeb4),
	.w1(32'h3ba6f522),
	.w2(32'h3c02d180),
	.w3(32'h3b38eedd),
	.w4(32'h3b49bd00),
	.w5(32'h3b94e600),
	.w6(32'h3b845b87),
	.w7(32'h3ba0d95b),
	.w8(32'h3b9188c6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96f9b3a),
	.w1(32'h3a1d724d),
	.w2(32'h39bdb8c1),
	.w3(32'h37ea019d),
	.w4(32'h3994b458),
	.w5(32'hb98bfaa2),
	.w6(32'hba3ff857),
	.w7(32'hb98280f6),
	.w8(32'h3888474d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b8f98),
	.w1(32'hb9b3f849),
	.w2(32'hba0578f3),
	.w3(32'h3a4ffc82),
	.w4(32'hb8814092),
	.w5(32'hb883eb56),
	.w6(32'hb952c61a),
	.w7(32'hb9c2b95c),
	.w8(32'h3963b389),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b324ebe),
	.w1(32'h3a7ffa30),
	.w2(32'h3a6e6fe2),
	.w3(32'h399bacc3),
	.w4(32'hba8f4aa2),
	.w5(32'h3a0cbd39),
	.w6(32'hba983ac0),
	.w7(32'hbb0d9c06),
	.w8(32'hba908246),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944437b),
	.w1(32'h3af65865),
	.w2(32'h3b12392b),
	.w3(32'h388f26e9),
	.w4(32'h3aab0daf),
	.w5(32'h3ab697a6),
	.w6(32'h3aacd0de),
	.w7(32'h3b25d914),
	.w8(32'h3acd7af6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9351885),
	.w1(32'hb9a0c244),
	.w2(32'hb9bf9cc8),
	.w3(32'h3a6ba38c),
	.w4(32'h3a05d6d8),
	.w5(32'hba14671d),
	.w6(32'h3a16eda8),
	.w7(32'h3a194ac3),
	.w8(32'h399053e6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853255),
	.w1(32'h3a884848),
	.w2(32'h39dad92d),
	.w3(32'hb9b98dff),
	.w4(32'hba1e93cd),
	.w5(32'hba56f238),
	.w6(32'hba3ffdd0),
	.w7(32'hbb3c8f34),
	.w8(32'hbb5cd5f9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea3a01),
	.w1(32'h3aaad40f),
	.w2(32'hbbc2b352),
	.w3(32'h3b854091),
	.w4(32'h3b162397),
	.w5(32'h3aa1b9a9),
	.w6(32'h3bcf3335),
	.w7(32'hba639013),
	.w8(32'hbb8229b7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a136970),
	.w1(32'h3c2af816),
	.w2(32'h3c7da0fd),
	.w3(32'h3b18239d),
	.w4(32'h3c4cd171),
	.w5(32'h3c52f3d5),
	.w6(32'h3bdc2992),
	.w7(32'h3c5ec32c),
	.w8(32'h3c6a1c78),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0299ed),
	.w1(32'h3c047cb1),
	.w2(32'h3c605999),
	.w3(32'h3b81e5ca),
	.w4(32'h3c175d85),
	.w5(32'h3c20f815),
	.w6(32'h3c052987),
	.w7(32'h3c4e584a),
	.w8(32'h3c4d41cd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e269),
	.w1(32'h3add8f8a),
	.w2(32'h3b12609e),
	.w3(32'h3ab11152),
	.w4(32'h3a413284),
	.w5(32'h3af5744f),
	.w6(32'h3b011e69),
	.w7(32'h39ec1c36),
	.w8(32'h3962234a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91263b3),
	.w1(32'h3a019939),
	.w2(32'h3949a04b),
	.w3(32'hb9c14bfd),
	.w4(32'hb8201056),
	.w5(32'h39e768e4),
	.w6(32'hb8af8c3f),
	.w7(32'h3910f4d5),
	.w8(32'h3a80ac30),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfc6e0),
	.w1(32'h39b3f317),
	.w2(32'hb99a726b),
	.w3(32'h3a8c61f6),
	.w4(32'hb9518897),
	.w5(32'hb7546784),
	.w6(32'h3aa3493a),
	.w7(32'hb94cdaa2),
	.w8(32'hb9ba56ae),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14b8a1),
	.w1(32'h3a00ef73),
	.w2(32'hb9a56087),
	.w3(32'hb97f5bfc),
	.w4(32'h39c1ac14),
	.w5(32'hb7147253),
	.w6(32'h3a16fd87),
	.w7(32'h3a150e7a),
	.w8(32'hb9b2a3b4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd9d7d),
	.w1(32'h3b221e8f),
	.w2(32'h3c09807f),
	.w3(32'hba7bcfae),
	.w4(32'hbbf9b17d),
	.w5(32'hbb8c0884),
	.w6(32'hbbe05624),
	.w7(32'hbc450843),
	.w8(32'hbb8b1bec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9694b0),
	.w1(32'h3bc72b13),
	.w2(32'h3c00355b),
	.w3(32'hb99bdd3b),
	.w4(32'h3b2b96c2),
	.w5(32'h3b9817c1),
	.w6(32'h3a31b55b),
	.w7(32'h3b8cb332),
	.w8(32'h3b8490ca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b3b2),
	.w1(32'h3bd4807d),
	.w2(32'h3c1e5450),
	.w3(32'h3ab3272a),
	.w4(32'hba8f986a),
	.w5(32'h3b7c640a),
	.w6(32'h3aa0b9dd),
	.w7(32'h3a2fd0d7),
	.w8(32'h3b2a7a92),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94e322),
	.w1(32'h3bbb9822),
	.w2(32'h3b9ac554),
	.w3(32'h3b123383),
	.w4(32'h3a1384d2),
	.w5(32'h3b24b1e6),
	.w6(32'h3ab00334),
	.w7(32'h3a097767),
	.w8(32'h3a27f323),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6349ed),
	.w1(32'hbb78f0a6),
	.w2(32'hbc237218),
	.w3(32'hbb910959),
	.w4(32'hbc73daf0),
	.w5(32'hbc84d4c1),
	.w6(32'hbc62f070),
	.w7(32'hbcdcf51f),
	.w8(32'hbca8b4bb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a84df),
	.w1(32'hb9b21752),
	.w2(32'h3a237b7a),
	.w3(32'hb9f0e439),
	.w4(32'hba035838),
	.w5(32'h34f7e45c),
	.w6(32'hb907701e),
	.w7(32'hba3da7a5),
	.w8(32'hba8de762),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a729ff),
	.w1(32'hb9fd626e),
	.w2(32'hba9b7b04),
	.w3(32'hba7a967a),
	.w4(32'hb94bdfcb),
	.w5(32'hb9fb8e32),
	.w6(32'hba5cc70d),
	.w7(32'hba37122a),
	.w8(32'hbaa90c05),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49e886),
	.w1(32'h39cf3b07),
	.w2(32'h3847e320),
	.w3(32'hba623471),
	.w4(32'h396cbf91),
	.w5(32'hba236b06),
	.w6(32'hba468e29),
	.w7(32'hb98f0195),
	.w8(32'hb9849aec),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01bce3),
	.w1(32'h3a6dc2d8),
	.w2(32'h3b2e3c47),
	.w3(32'hbabd830f),
	.w4(32'hbb5d6c11),
	.w5(32'hbb0f2a65),
	.w6(32'hba903b78),
	.w7(32'hbb657554),
	.w8(32'hbafcc544),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a2148),
	.w1(32'hb9d3641c),
	.w2(32'hba61713b),
	.w3(32'hb9e6a462),
	.w4(32'hba822074),
	.w5(32'hbaaa2493),
	.w6(32'hb9a477a1),
	.w7(32'hbb04fbfc),
	.w8(32'hbadfe3af),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e693a),
	.w1(32'hbb0e1ff6),
	.w2(32'hbbaa6ef7),
	.w3(32'hbb884b9d),
	.w4(32'hbc381d19),
	.w5(32'hbbbb944c),
	.w6(32'hbc0eaa31),
	.w7(32'hbc76590a),
	.w8(32'hbbe5765c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992256f),
	.w1(32'hba52f6ed),
	.w2(32'h395caf02),
	.w3(32'hbad4ff45),
	.w4(32'hbae39173),
	.w5(32'hba985d5b),
	.w6(32'hb902b3aa),
	.w7(32'hba52df99),
	.w8(32'hba859f96),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39345ff2),
	.w1(32'h39b81cbf),
	.w2(32'hb922191a),
	.w3(32'h3900da07),
	.w4(32'hb8a2fdde),
	.w5(32'h3a033fa1),
	.w6(32'h38c22c16),
	.w7(32'h39bf44fb),
	.w8(32'h3a8aff6a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c4e8d),
	.w1(32'h39bfd941),
	.w2(32'h38963ae0),
	.w3(32'hb91551d8),
	.w4(32'h3978c7bb),
	.w5(32'hb92dd1b3),
	.w6(32'h39c50ba0),
	.w7(32'hb73a8c08),
	.w8(32'h3904cafb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c60123),
	.w1(32'h39684624),
	.w2(32'h3a60c711),
	.w3(32'hb865613d),
	.w4(32'hb8a30a7d),
	.w5(32'h394708d8),
	.w6(32'hb9ff72c0),
	.w7(32'h38e7b318),
	.w8(32'h3a05df0b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dc3d2),
	.w1(32'h3a583dbb),
	.w2(32'hb920ab76),
	.w3(32'h39e5ec13),
	.w4(32'h3a23cf3a),
	.w5(32'hba4d1126),
	.w6(32'h3a89de2b),
	.w7(32'h3a945d22),
	.w8(32'hb9f4a69d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82c4d01),
	.w1(32'h3970158f),
	.w2(32'hb9c2474f),
	.w3(32'h3a19d555),
	.w4(32'h3a3409b8),
	.w5(32'hb95260a7),
	.w6(32'h38e15f59),
	.w7(32'h378420fc),
	.w8(32'hb907b1e8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770d1f),
	.w1(32'hbaa22674),
	.w2(32'hbac63d71),
	.w3(32'hbb72c975),
	.w4(32'hbbf78ac3),
	.w5(32'hbb485edd),
	.w6(32'hbc0838b9),
	.w7(32'hbc37bf9a),
	.w8(32'hbbefa4d8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb321a8a),
	.w1(32'hbb153c0d),
	.w2(32'hbaaa1f5c),
	.w3(32'hba410c00),
	.w4(32'hbba82212),
	.w5(32'hbb97d69b),
	.w6(32'hbb6a53d2),
	.w7(32'hbb283bf2),
	.w8(32'hbb858485),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c38c8),
	.w1(32'hb9f161f2),
	.w2(32'hba98448a),
	.w3(32'hb9a9d5cb),
	.w4(32'hba1dc8bc),
	.w5(32'hba0b1055),
	.w6(32'hb806c1e7),
	.w7(32'hb9d8884f),
	.w8(32'hb909214e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba031549),
	.w1(32'h3997fcf8),
	.w2(32'hba0a6252),
	.w3(32'hba7bb5e5),
	.w4(32'hb9498805),
	.w5(32'hb992d622),
	.w6(32'hba177d37),
	.w7(32'h38b7ff0b),
	.w8(32'hb96400c0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17788a),
	.w1(32'h39e3249a),
	.w2(32'h38f32079),
	.w3(32'hb9a919ee),
	.w4(32'h3901c52c),
	.w5(32'h34e2a44a),
	.w6(32'h390d8b3c),
	.w7(32'h3930f86b),
	.w8(32'hb7b1fca3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399efafe),
	.w1(32'hb8733df8),
	.w2(32'hba0eb0fd),
	.w3(32'hb9b007fe),
	.w4(32'hb96048e9),
	.w5(32'h390b245b),
	.w6(32'hb9d9cfa8),
	.w7(32'hb9708e33),
	.w8(32'hb979804a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02283a),
	.w1(32'hbbcc2206),
	.w2(32'hbb3759a8),
	.w3(32'h3b367b3f),
	.w4(32'h3a18bc2d),
	.w5(32'h3b148eae),
	.w6(32'hbaf2b6f4),
	.w7(32'hbb9607d4),
	.w8(32'hb8b4f036),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50e37d),
	.w1(32'h3b8c2eee),
	.w2(32'h3c0e302e),
	.w3(32'h39852ce0),
	.w4(32'hb9cd7fc0),
	.w5(32'h3b9d6292),
	.w6(32'h3ba2e7b1),
	.w7(32'h3b78aaaa),
	.w8(32'hba7ce073),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf99e40),
	.w1(32'hbadaabff),
	.w2(32'hba9aceb2),
	.w3(32'hbbb207da),
	.w4(32'hbc087b6b),
	.w5(32'hbbc752f8),
	.w6(32'hbba07128),
	.w7(32'hbbe1df4b),
	.w8(32'hbbe2b6a2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24897a),
	.w1(32'h3c4ff9c4),
	.w2(32'h3c0a273d),
	.w3(32'hb9ca4351),
	.w4(32'h3be0bb78),
	.w5(32'h3b8901a8),
	.w6(32'h3b842c31),
	.w7(32'h3c4cd7a2),
	.w8(32'hbb6dd37f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda0c1f),
	.w1(32'h3b12763b),
	.w2(32'h3a6ffee6),
	.w3(32'hbcac8be1),
	.w4(32'hbc01f12e),
	.w5(32'hbb4534a4),
	.w6(32'hbc1967c3),
	.w7(32'hbc03dbe1),
	.w8(32'hbc360884),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34ff8b),
	.w1(32'hbbd44217),
	.w2(32'hbabcd106),
	.w3(32'h3c1b9b70),
	.w4(32'hbc848902),
	.w5(32'hbc4700a7),
	.w6(32'h3aeb5006),
	.w7(32'hbb3180b2),
	.w8(32'h3bb6da28),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc84d3c),
	.w1(32'h3aa57c86),
	.w2(32'h3b086e51),
	.w3(32'h3bffdabe),
	.w4(32'h3bf8eba9),
	.w5(32'h3c7063dd),
	.w6(32'h3c1d410a),
	.w7(32'h3b8ef1c6),
	.w8(32'h3c2f3000),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0e72),
	.w1(32'hbb99c124),
	.w2(32'hbb4a40a1),
	.w3(32'hba61ba78),
	.w4(32'h3b334fc9),
	.w5(32'hbb8bb16d),
	.w6(32'h3b0e0998),
	.w7(32'hbbfd8fca),
	.w8(32'hbb734032),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d75f),
	.w1(32'hbbcc97b7),
	.w2(32'hbc132091),
	.w3(32'hba9f5cb4),
	.w4(32'hbbb05b86),
	.w5(32'hbc4afab7),
	.w6(32'h3ba09868),
	.w7(32'h3b78dc28),
	.w8(32'h3bb18ce0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26144a),
	.w1(32'hbaa7c1da),
	.w2(32'hbc0ec64c),
	.w3(32'hbc10c118),
	.w4(32'hbbba8c45),
	.w5(32'hbbad9d3f),
	.w6(32'hbb8a28a5),
	.w7(32'hbc9436d2),
	.w8(32'hbc1bde48),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b733485),
	.w1(32'hbbf9a527),
	.w2(32'hbb50285a),
	.w3(32'hbc5f7b6a),
	.w4(32'hbce0b78d),
	.w5(32'hbc5e5a75),
	.w6(32'hbc1cf324),
	.w7(32'hbd03af39),
	.w8(32'hbc7c0c42),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce739e8),
	.w1(32'h3b10d901),
	.w2(32'h3c0b848e),
	.w3(32'h3d0cab20),
	.w4(32'h3a3474c1),
	.w5(32'h3c8c1341),
	.w6(32'h3c8c63ec),
	.w7(32'hbb2aedb2),
	.w8(32'hbb883793),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed390f),
	.w1(32'hba84972a),
	.w2(32'h3ba00b78),
	.w3(32'h3c110ad8),
	.w4(32'hbb80dede),
	.w5(32'h3bca29e4),
	.w6(32'h3b2283a3),
	.w7(32'hbc064c09),
	.w8(32'h3977de60),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc1709),
	.w1(32'hbc514b74),
	.w2(32'hbbe6094c),
	.w3(32'hbb003c8d),
	.w4(32'hbc8d7fe3),
	.w5(32'hbbbc716a),
	.w6(32'hbb288be1),
	.w7(32'hbbd379cc),
	.w8(32'hbc2d11a3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c270a3d),
	.w1(32'h3b20799c),
	.w2(32'h3c15b492),
	.w3(32'h3beb4184),
	.w4(32'h3b52b0ff),
	.w5(32'h3a5b739c),
	.w6(32'h3b048ea5),
	.w7(32'h3b9a3517),
	.w8(32'h3c282613),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c666621),
	.w1(32'hbb8cd0e4),
	.w2(32'h3b0ff2ed),
	.w3(32'h3c408756),
	.w4(32'h3b18442d),
	.w5(32'h3c2bcdda),
	.w6(32'h3c82e9c3),
	.w7(32'hbbb442b9),
	.w8(32'h3b8e848b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5ba8c),
	.w1(32'h3b1e405f),
	.w2(32'hb937bd96),
	.w3(32'h3cb0ad87),
	.w4(32'h3c3a1af8),
	.w5(32'h3a98ea48),
	.w6(32'h3c3523ae),
	.w7(32'h3b25b285),
	.w8(32'hbbe2733f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7dd2a),
	.w1(32'hbb3b8532),
	.w2(32'hba8fdced),
	.w3(32'hbace1998),
	.w4(32'hbb2671f1),
	.w5(32'h3a08ffcb),
	.w6(32'hbb1c0f48),
	.w7(32'hbad7d38c),
	.w8(32'h3b1983ab),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63ae81),
	.w1(32'hbbc4779b),
	.w2(32'h3ba05158),
	.w3(32'h3b937093),
	.w4(32'hbbe95b44),
	.w5(32'h3c28e2fa),
	.w6(32'hbbbc1bbe),
	.w7(32'hbb0c19a0),
	.w8(32'h3c4cdad5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13f459),
	.w1(32'h3bd65015),
	.w2(32'h3b9434cf),
	.w3(32'h3c1b08c8),
	.w4(32'h3a9983af),
	.w5(32'h3c5cc0a7),
	.w6(32'h3b6296de),
	.w7(32'hbb28ca86),
	.w8(32'hbc92730c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eb191),
	.w1(32'hb9260790),
	.w2(32'h3c1a2d5a),
	.w3(32'hbc2f3dc1),
	.w4(32'hbbd5584d),
	.w5(32'h3c09d657),
	.w6(32'hbc387bd5),
	.w7(32'hbab10c39),
	.w8(32'h3ad8742e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09118c),
	.w1(32'h3b830fac),
	.w2(32'hbba22dd3),
	.w3(32'h3c207034),
	.w4(32'hbb031ec1),
	.w5(32'hbc034f34),
	.w6(32'h3c00f0c1),
	.w7(32'hbb9a7f80),
	.w8(32'hbbac2577),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0741ae),
	.w1(32'hbb6f843f),
	.w2(32'hbb1e3ff7),
	.w3(32'hbba6b49c),
	.w4(32'hbc25236b),
	.w5(32'hbb815db6),
	.w6(32'h3be8cca7),
	.w7(32'hbc041860),
	.w8(32'h3baaceb1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24bc76),
	.w1(32'hbafa238a),
	.w2(32'hbb0ffe6b),
	.w3(32'h3c2681c6),
	.w4(32'hb52ddc64),
	.w5(32'h3bbf76b0),
	.w6(32'hbc9ea0f8),
	.w7(32'hbc74aa4a),
	.w8(32'hb9a280af),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05414c),
	.w1(32'h3be02afe),
	.w2(32'h3b9984c5),
	.w3(32'hbc8e55d6),
	.w4(32'h3bba7f4b),
	.w5(32'hba230861),
	.w6(32'hbbcbeb75),
	.w7(32'h3b438166),
	.w8(32'hbb0e8a47),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96942d),
	.w1(32'hbb2040ea),
	.w2(32'h3c2cdcbd),
	.w3(32'h3c4b8f76),
	.w4(32'h3b90eae4),
	.w5(32'h3c5abe8c),
	.w6(32'h3b90cbfc),
	.w7(32'h3cbd98ef),
	.w8(32'h3be34cff),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97f1cf),
	.w1(32'h3ba8ed60),
	.w2(32'hbabd860e),
	.w3(32'hba51fa9d),
	.w4(32'h3bde5135),
	.w5(32'hbb3f427e),
	.w6(32'hbc1b9f7e),
	.w7(32'h3b523f22),
	.w8(32'h3b7afbda),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf77abc),
	.w1(32'h3bb4a853),
	.w2(32'hbb68b855),
	.w3(32'hbc7c2966),
	.w4(32'h3be409c3),
	.w5(32'h3b4b8465),
	.w6(32'hba967363),
	.w7(32'hba4c6655),
	.w8(32'hba4da0cb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc419a71),
	.w1(32'hbba91ec9),
	.w2(32'h3c0b9baa),
	.w3(32'hbc154ff3),
	.w4(32'hbc221cf3),
	.w5(32'h3c5c9eca),
	.w6(32'hbaf6f512),
	.w7(32'hbb75e521),
	.w8(32'h3ba9f84e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c65f3),
	.w1(32'h3b3dae6a),
	.w2(32'h3bd93b58),
	.w3(32'h3c5ea7b3),
	.w4(32'hbb6b947d),
	.w5(32'h3bbfcaed),
	.w6(32'hb91d8bcc),
	.w7(32'hbbb16e70),
	.w8(32'hb92515ba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52187),
	.w1(32'hba051a61),
	.w2(32'hbad6cd01),
	.w3(32'hbc275c78),
	.w4(32'hbb97e170),
	.w5(32'h3c491b81),
	.w6(32'hbb834dd9),
	.w7(32'hbb5a4dd9),
	.w8(32'h3b9feadf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3db42a),
	.w1(32'h3b95c850),
	.w2(32'h3bf76c93),
	.w3(32'h3c3324b8),
	.w4(32'h3c45401a),
	.w5(32'h3c9fc7ad),
	.w6(32'h3b9648dd),
	.w7(32'h3bb37855),
	.w8(32'h3c412c67),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a54c7),
	.w1(32'hbba32077),
	.w2(32'h3b7e0025),
	.w3(32'h3a563346),
	.w4(32'h3c21d87a),
	.w5(32'h3c6ceea8),
	.w6(32'h3b6ad0d2),
	.w7(32'h3bb0f408),
	.w8(32'h3c39fd7a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11aa32),
	.w1(32'h3c4ef78c),
	.w2(32'hbbc4ef31),
	.w3(32'h3b47e141),
	.w4(32'h3c816bd7),
	.w5(32'h3c52179e),
	.w6(32'h3a99f854),
	.w7(32'hbc84a642),
	.w8(32'hbbba1f22),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8740e8),
	.w1(32'h3b344260),
	.w2(32'h3b79ea04),
	.w3(32'hbc89cbff),
	.w4(32'hbb5e57fa),
	.w5(32'h3bacdea0),
	.w6(32'h3c6a2729),
	.w7(32'hbb4c5f27),
	.w8(32'h3bc10b11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2ef50),
	.w1(32'hba574c65),
	.w2(32'h3c197533),
	.w3(32'h3bc852ab),
	.w4(32'h3af56e1e),
	.w5(32'h3cdfeff3),
	.w6(32'h3bbf0898),
	.w7(32'h3b25533b),
	.w8(32'h3bbfbc36),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4293c),
	.w1(32'h3aeeed11),
	.w2(32'hbbd0012a),
	.w3(32'h3b17bcf3),
	.w4(32'h3a925a71),
	.w5(32'hba9682da),
	.w6(32'h3b6a0c45),
	.w7(32'hbb75dc8a),
	.w8(32'hbbeb656f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe497a),
	.w1(32'hba9d152a),
	.w2(32'h3c01b1b3),
	.w3(32'hbbe2b689),
	.w4(32'h3a12e675),
	.w5(32'h3cc55862),
	.w6(32'hbc262323),
	.w7(32'hbc0d2c0d),
	.w8(32'h3af9e42b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3214f2),
	.w1(32'hbb98f4d2),
	.w2(32'hbc5a96c4),
	.w3(32'h39f30f7f),
	.w4(32'hbca808e4),
	.w5(32'hbc5712ba),
	.w6(32'hbc3743c7),
	.w7(32'hbce43367),
	.w8(32'hbc0557fd),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacebcb),
	.w1(32'h3b37cc73),
	.w2(32'h3a5292b9),
	.w3(32'h3b423b66),
	.w4(32'hbadeebc5),
	.w5(32'h3b741c1f),
	.w6(32'h3bdf9d61),
	.w7(32'hb92aff79),
	.w8(32'hba6e136b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b785336),
	.w1(32'h3bdbf671),
	.w2(32'h3b6e9d6b),
	.w3(32'h3bc3ee3c),
	.w4(32'h3c865983),
	.w5(32'h3c517484),
	.w6(32'h3b01f35a),
	.w7(32'h3bf8c204),
	.w8(32'h3af163d6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc89262),
	.w1(32'h39ea6eab),
	.w2(32'hbae8742d),
	.w3(32'h3b2ffbcc),
	.w4(32'hba9d9271),
	.w5(32'h3b5ff407),
	.w6(32'hbc061403),
	.w7(32'h3b32bdd0),
	.w8(32'hbbe5785a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c680b),
	.w1(32'hbb1eb799),
	.w2(32'hbb1773ee),
	.w3(32'hbc565cbf),
	.w4(32'hba6c8998),
	.w5(32'hbc2b6f4f),
	.w6(32'hbc4901a2),
	.w7(32'hbc242fb5),
	.w8(32'hbc0ebaa4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5048b),
	.w1(32'hbb07534a),
	.w2(32'h3b2c864e),
	.w3(32'hbc0253bb),
	.w4(32'hbc0e9a59),
	.w5(32'hb9a282c5),
	.w6(32'h3a4cf0eb),
	.w7(32'h3a9fa3a4),
	.w8(32'h3b2ef873),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a5c2a),
	.w1(32'hbb8336f4),
	.w2(32'h3c8fa041),
	.w3(32'hbc07f4c6),
	.w4(32'h3c349086),
	.w5(32'h3c1808ee),
	.w6(32'hbbbde3c1),
	.w7(32'h3c310a3a),
	.w8(32'h3c10ae35),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5371a7),
	.w1(32'hbbcba4fd),
	.w2(32'h3c0d21a3),
	.w3(32'hbc08b409),
	.w4(32'h3bd88c86),
	.w5(32'h3d0a2ba3),
	.w6(32'h3b74432b),
	.w7(32'h3b6b7d99),
	.w8(32'h3c6517df),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3dbe8),
	.w1(32'hbc047791),
	.w2(32'hbb1afe52),
	.w3(32'h3c1b97bf),
	.w4(32'hbbd23a20),
	.w5(32'h3b059fdf),
	.w6(32'h3c0058ee),
	.w7(32'h3bac61d5),
	.w8(32'hbac6be04),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dbcb9),
	.w1(32'h3bb612cd),
	.w2(32'h39ca3296),
	.w3(32'h3bd0d206),
	.w4(32'h3b23712e),
	.w5(32'hbbd9e11d),
	.w6(32'h3aa8c6e0),
	.w7(32'h3a835181),
	.w8(32'hbb172a4a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4cc3c),
	.w1(32'h3bb17569),
	.w2(32'hbbe00d06),
	.w3(32'h3aaed935),
	.w4(32'h3c389608),
	.w5(32'hbc2e5064),
	.w6(32'hbafcfa9f),
	.w7(32'h3c22900a),
	.w8(32'h391a6aa2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6f391),
	.w1(32'h3bcbac54),
	.w2(32'hbb5c3c45),
	.w3(32'hbc9e8866),
	.w4(32'h3b2ee64b),
	.w5(32'h3ba0e612),
	.w6(32'hbc17e39d),
	.w7(32'h3a3006bd),
	.w8(32'h3a7da6b6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b654f9f),
	.w1(32'h3ba6743c),
	.w2(32'hbc0bbcab),
	.w3(32'h3bf5011c),
	.w4(32'h3c7096cf),
	.w5(32'hbba92491),
	.w6(32'h3be1cf17),
	.w7(32'h3bde5a7f),
	.w8(32'hbaaccf7b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cff8c),
	.w1(32'hbb009418),
	.w2(32'hbc23b6e2),
	.w3(32'hbc3d673e),
	.w4(32'h3c20f5ac),
	.w5(32'hbbec0b2d),
	.w6(32'hbb94c34f),
	.w7(32'h3c11855f),
	.w8(32'hbab7e285),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e11b0),
	.w1(32'hbbdab264),
	.w2(32'hbbd39d7b),
	.w3(32'h3ac4f5ea),
	.w4(32'hbc0933ef),
	.w5(32'hbc3bd3f2),
	.w6(32'h3bd0ea35),
	.w7(32'hbba0e1e7),
	.w8(32'hbb562f79),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b3fc5),
	.w1(32'hbb1f0da0),
	.w2(32'h3bfeb6b2),
	.w3(32'hbb9d71d7),
	.w4(32'hbc2eb0b2),
	.w5(32'h3cc32d47),
	.w6(32'hbb30b22f),
	.w7(32'hbbb7667b),
	.w8(32'h3b86ff63),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8c290),
	.w1(32'hbc2e1b27),
	.w2(32'hbb0afc55),
	.w3(32'h3acefbdc),
	.w4(32'hbbdafde5),
	.w5(32'hbbb76928),
	.w6(32'hbab8a137),
	.w7(32'hbbd84e27),
	.w8(32'h3ac7214f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2779bb),
	.w1(32'hbb50067e),
	.w2(32'hbc221d6e),
	.w3(32'h3cb09f30),
	.w4(32'h3b2f474b),
	.w5(32'hbba2e52f),
	.w6(32'h3b7f5136),
	.w7(32'hbc05dc93),
	.w8(32'hbc38c266),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e97e9),
	.w1(32'h3be56e6a),
	.w2(32'hbb1584db),
	.w3(32'hbc5c99e7),
	.w4(32'hba99384a),
	.w5(32'hbb11c463),
	.w6(32'hbbb60802),
	.w7(32'hbb3633af),
	.w8(32'hbc1580ed),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be075),
	.w1(32'h3bf3a192),
	.w2(32'h3c5217e7),
	.w3(32'h3c54c502),
	.w4(32'h3c49ac57),
	.w5(32'h3cbb48aa),
	.w6(32'h3b282c3d),
	.w7(32'h3c717a48),
	.w8(32'h3c8808f7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24e678),
	.w1(32'hbba9986e),
	.w2(32'hbb331cc5),
	.w3(32'hbc76de3a),
	.w4(32'hbbff484d),
	.w5(32'hbbe02c2b),
	.w6(32'h39efade8),
	.w7(32'h39c8bad3),
	.w8(32'hbad7c3b9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c195442),
	.w1(32'hbbcb4bad),
	.w2(32'hbb8bdce5),
	.w3(32'h3aa1c03e),
	.w4(32'hbb18e239),
	.w5(32'hbb4095e0),
	.w6(32'hbae8c24a),
	.w7(32'h3b8836e4),
	.w8(32'hba7dec67),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f8dcd),
	.w1(32'h3bc94534),
	.w2(32'hbb06c6be),
	.w3(32'hbb6fa764),
	.w4(32'h39dedcde),
	.w5(32'h3bd8efd4),
	.w6(32'hba88edbb),
	.w7(32'h3bee0eb5),
	.w8(32'hbbf3d5f5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33a22c),
	.w1(32'h3be9b101),
	.w2(32'hba205bcd),
	.w3(32'h3b8937b2),
	.w4(32'hbb8fcff8),
	.w5(32'hbb953616),
	.w6(32'hbc4a8dd8),
	.w7(32'hbbd6acab),
	.w8(32'hbbf3f8c0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d6b7),
	.w1(32'hba2011e4),
	.w2(32'h3aafee1d),
	.w3(32'hbb2c9b59),
	.w4(32'hbc275a51),
	.w5(32'hbc000f6d),
	.w6(32'hbbaa0d75),
	.w7(32'hbbde58a9),
	.w8(32'hbb159b16),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc497ba),
	.w1(32'h3b27db41),
	.w2(32'hb9e43d87),
	.w3(32'h3a10af87),
	.w4(32'hba941ad7),
	.w5(32'h3cae9902),
	.w6(32'h3b8cfee8),
	.w7(32'hbb3dbc69),
	.w8(32'h3ba06682),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7adf74),
	.w1(32'hbbd87d69),
	.w2(32'hbb1645fa),
	.w3(32'h3bff2e9e),
	.w4(32'hb9583718),
	.w5(32'h3bef2fb5),
	.w6(32'h3c0fe0ff),
	.w7(32'hbc54d4f9),
	.w8(32'hbb832209),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb775bbc),
	.w1(32'h3c18a650),
	.w2(32'h3b13a2d0),
	.w3(32'hbb5967f9),
	.w4(32'h3bedfdf1),
	.w5(32'h3b96d044),
	.w6(32'hbc0db710),
	.w7(32'h3b66f898),
	.w8(32'h3c467ddc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd79c6),
	.w1(32'hbaa358c5),
	.w2(32'hbaf0c388),
	.w3(32'hbb68f048),
	.w4(32'h3be400c1),
	.w5(32'h3b96ef8a),
	.w6(32'h3b418692),
	.w7(32'hbb40b712),
	.w8(32'hb9076388),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccec64),
	.w1(32'h3c15c76d),
	.w2(32'hbbb00bc2),
	.w3(32'hbc4c39b7),
	.w4(32'h3d060fb5),
	.w5(32'h3a9814ea),
	.w6(32'hbbc563d3),
	.w7(32'h3ccfddb7),
	.w8(32'h3bbe44eb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe78930),
	.w1(32'hbb921d23),
	.w2(32'hbb9590fa),
	.w3(32'hbc8ee34f),
	.w4(32'hbc85044b),
	.w5(32'hbc6516b2),
	.w6(32'hbc8882b0),
	.w7(32'hbc999402),
	.w8(32'hbc1ba510),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb94a74),
	.w1(32'h3c0f8bfd),
	.w2(32'hba3d6f7f),
	.w3(32'hb92d05bf),
	.w4(32'h3c8fe086),
	.w5(32'h3b14f952),
	.w6(32'h3a62fc21),
	.w7(32'h3c7b9cf4),
	.w8(32'h3bfe4da8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fdb96),
	.w1(32'hbb5e5329),
	.w2(32'h3b8d40ae),
	.w3(32'hbb3e8462),
	.w4(32'h3b1e5c34),
	.w5(32'h3cc73eaf),
	.w6(32'hbc180e7f),
	.w7(32'hbb88cd68),
	.w8(32'h3b696e22),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b8fc),
	.w1(32'hbbc9089c),
	.w2(32'h3b766d27),
	.w3(32'h39b68f6d),
	.w4(32'hbaae4dd1),
	.w5(32'hbb5ce494),
	.w6(32'hbb33b645),
	.w7(32'hbc151ab7),
	.w8(32'hbba984bc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae92977),
	.w1(32'h37e19f8a),
	.w2(32'h3b4d1c86),
	.w3(32'hbc304fb3),
	.w4(32'hbb8f4645),
	.w5(32'h3a8f8860),
	.w6(32'hbb01f8c5),
	.w7(32'h3b981b6b),
	.w8(32'h3b814425),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a953eee),
	.w1(32'hbc626b1e),
	.w2(32'h3c0523a0),
	.w3(32'hbc003c3a),
	.w4(32'hbc8fcba7),
	.w5(32'h3bc6fccc),
	.w6(32'hbb75ff1b),
	.w7(32'hbc8a442e),
	.w8(32'h3b8a06d5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca02b65),
	.w1(32'hba945054),
	.w2(32'h3b156fb6),
	.w3(32'h3d22c430),
	.w4(32'hbba2574c),
	.w5(32'h3cd7e6bd),
	.w6(32'h3c3b0559),
	.w7(32'hbc031e35),
	.w8(32'h3b147bc2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344d93),
	.w1(32'hba95348c),
	.w2(32'h3b7e269b),
	.w3(32'h3ce8744e),
	.w4(32'h3b0c3475),
	.w5(32'h3c1c8fd6),
	.w6(32'h3c21ffed),
	.w7(32'h3a409625),
	.w8(32'h3bd72339),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d7739),
	.w1(32'h3b2128cf),
	.w2(32'h3acb39c9),
	.w3(32'hbbf9846b),
	.w4(32'hbab4a031),
	.w5(32'h3c8b8d15),
	.w6(32'hbc0aeaec),
	.w7(32'h3be785ce),
	.w8(32'h3ae608fd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7702f8),
	.w1(32'hbbfaacb6),
	.w2(32'hbb013ee2),
	.w3(32'h3c043b49),
	.w4(32'hbb705239),
	.w5(32'h3a948900),
	.w6(32'h3bba1d5e),
	.w7(32'hbba9cd89),
	.w8(32'hb84a8918),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32c0ac),
	.w1(32'hbbd0e967),
	.w2(32'h3c1f4aa9),
	.w3(32'h3cd5e1b0),
	.w4(32'hbbb2e1b5),
	.w5(32'h3bc6c12b),
	.w6(32'h3c171706),
	.w7(32'h3c022114),
	.w8(32'h3c347fce),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60dbc),
	.w1(32'h3bd8b85b),
	.w2(32'hba50a3e3),
	.w3(32'h3ca2cc06),
	.w4(32'hbb9640c0),
	.w5(32'hbc67ccee),
	.w6(32'h3b7a6908),
	.w7(32'hbb99bc39),
	.w8(32'hbc3fd36b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dcf21),
	.w1(32'h3abdc9b4),
	.w2(32'h3a8c85a9),
	.w3(32'hbb8a4721),
	.w4(32'h3a101581),
	.w5(32'h3c1a42a2),
	.w6(32'hbbf2dca8),
	.w7(32'hbb778488),
	.w8(32'h3b6e93b4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd1ce49),
	.w1(32'hbb10a529),
	.w2(32'h3c5903b2),
	.w3(32'h3cd0374b),
	.w4(32'hbc42e704),
	.w5(32'h3b8cc0cd),
	.w6(32'h3bc20135),
	.w7(32'hbc84f22a),
	.w8(32'hbc6c823a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bb0e1),
	.w1(32'h3c2e0bba),
	.w2(32'h3b0911bd),
	.w3(32'h3ca7be1e),
	.w4(32'h3cb25ca4),
	.w5(32'h3bbedfee),
	.w6(32'h3c3e6831),
	.w7(32'h3be4b80e),
	.w8(32'h3c2404ae),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae69ee0),
	.w1(32'h3c3bca4b),
	.w2(32'h3b8e72bd),
	.w3(32'hbb8dc5c2),
	.w4(32'h3c4e14ad),
	.w5(32'h3c85e8ec),
	.w6(32'hbbddd606),
	.w7(32'h3c2a8833),
	.w8(32'h3c9b5d62),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33bff3),
	.w1(32'h3c802309),
	.w2(32'h3bf343bd),
	.w3(32'h3bd3c77b),
	.w4(32'h3c692a54),
	.w5(32'hbb6f57d0),
	.w6(32'h3a3e6a85),
	.w7(32'h3b7933c9),
	.w8(32'hbb0b259f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a2610),
	.w1(32'hbb8540c8),
	.w2(32'hbbbeb6c8),
	.w3(32'hbc4f11db),
	.w4(32'hbc2b366b),
	.w5(32'hbc2d9e92),
	.w6(32'hba87ed1a),
	.w7(32'hbb99dcbf),
	.w8(32'hbb84a68a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3fa32),
	.w1(32'hbb230d07),
	.w2(32'hbbba970f),
	.w3(32'hbb579945),
	.w4(32'h3a95ae07),
	.w5(32'hbc3bbcd0),
	.w6(32'h3ae3ea38),
	.w7(32'h3bafc13f),
	.w8(32'hbc3c4ec9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc695690),
	.w1(32'h3cc581d4),
	.w2(32'h3c1fe5f4),
	.w3(32'hbcc32070),
	.w4(32'h3d2d1c0f),
	.w5(32'h3c027ab1),
	.w6(32'hbcbdd0d0),
	.w7(32'h3ce162a5),
	.w8(32'h3c15be40),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95b327),
	.w1(32'h3996d8a6),
	.w2(32'hbb5a69c1),
	.w3(32'hbcedd9ba),
	.w4(32'h3b3908a4),
	.w5(32'hbb720937),
	.w6(32'hbc2b129c),
	.w7(32'h3b2042d0),
	.w8(32'hbadf0098),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9c346),
	.w1(32'h3bc16d2f),
	.w2(32'h3aefae1c),
	.w3(32'hbb36c0e2),
	.w4(32'h3b4d23e2),
	.w5(32'h38b052e1),
	.w6(32'hbba47387),
	.w7(32'h3b9060d7),
	.w8(32'hbb9ef740),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5882e),
	.w1(32'hba902fde),
	.w2(32'h3b1133a2),
	.w3(32'hbc2de098),
	.w4(32'hbb8427b8),
	.w5(32'hbb50ac0b),
	.w6(32'h3a308c9c),
	.w7(32'h3a59d24d),
	.w8(32'hbabefbac),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae42198),
	.w1(32'h3a381932),
	.w2(32'h3c972f7c),
	.w3(32'h3c524e7c),
	.w4(32'h3c7d302b),
	.w5(32'h3c953b69),
	.w6(32'h3c1a3575),
	.w7(32'h3bccb01d),
	.w8(32'h3c9be561),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847e01),
	.w1(32'hbaae5a70),
	.w2(32'h3bf80b19),
	.w3(32'h3b6cc524),
	.w4(32'hbc12063d),
	.w5(32'h3a0dda2e),
	.w6(32'hbb20e64d),
	.w7(32'hbc3d0fea),
	.w8(32'hbb1a9767),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf903c8),
	.w1(32'hbbb51a66),
	.w2(32'h3bb62218),
	.w3(32'h3c921b10),
	.w4(32'hbb8bb26b),
	.w5(32'h3cdcf511),
	.w6(32'h3c0ffc01),
	.w7(32'hbb068b30),
	.w8(32'h3c23534c),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0e63),
	.w1(32'h3b2e1637),
	.w2(32'h3b6462e5),
	.w3(32'h3b2fce93),
	.w4(32'h3c463d73),
	.w5(32'h3b8d3c2e),
	.w6(32'hbaa08f82),
	.w7(32'hba7cfd5e),
	.w8(32'hbb9450d3),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0be34),
	.w1(32'hbb43d98d),
	.w2(32'hbad2c92e),
	.w3(32'hb9c1eb41),
	.w4(32'h3c293c96),
	.w5(32'h38c071a6),
	.w6(32'h3c241feb),
	.w7(32'h3be47503),
	.w8(32'hbb838fc9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2736),
	.w1(32'hbb679675),
	.w2(32'hbb0a2736),
	.w3(32'hbc62383c),
	.w4(32'h3c22be6c),
	.w5(32'hbb1a40d8),
	.w6(32'hbb8edca6),
	.w7(32'h3be07a93),
	.w8(32'h3b3cd3de),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82ee09),
	.w1(32'hbc19a787),
	.w2(32'hbbceb937),
	.w3(32'hbbbc4f51),
	.w4(32'hbc80e3c6),
	.w5(32'hbc84115c),
	.w6(32'hbc190d35),
	.w7(32'hbc307396),
	.w8(32'hbc332897),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c38c),
	.w1(32'h3bd120a4),
	.w2(32'h39e3be0d),
	.w3(32'h3b937a8e),
	.w4(32'h3a39aeaa),
	.w5(32'h3bdf0e49),
	.w6(32'hbbc04406),
	.w7(32'h389f28aa),
	.w8(32'h3a9e4fef),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2df0),
	.w1(32'hbb1f23c6),
	.w2(32'h3bd4809f),
	.w3(32'hbbcac9d8),
	.w4(32'hbba6957b),
	.w5(32'h3cfc0e75),
	.w6(32'h3a6c6ebb),
	.w7(32'hbb2f32be),
	.w8(32'h3c2f9577),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cd087),
	.w1(32'hbb9107f6),
	.w2(32'hb9c04acb),
	.w3(32'h3c8feeda),
	.w4(32'hbc68223c),
	.w5(32'h3ade1206),
	.w6(32'h3b6a914e),
	.w7(32'hbbcec355),
	.w8(32'h3ab191cb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fc620),
	.w1(32'h3c1af0eb),
	.w2(32'h3b195793),
	.w3(32'h3b03c8d0),
	.w4(32'h3c1335a8),
	.w5(32'h3bf822af),
	.w6(32'h3bed1be2),
	.w7(32'h3c1c78fa),
	.w8(32'h3be8e4fb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2bced),
	.w1(32'h39e443d4),
	.w2(32'hbbe260c5),
	.w3(32'hbc2c61a1),
	.w4(32'hbbdb679e),
	.w5(32'hbc88866c),
	.w6(32'hbacbfe1e),
	.w7(32'hbb7071eb),
	.w8(32'hbbdee3c6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9e31b),
	.w1(32'h3c1ed3c0),
	.w2(32'h3b9b7e91),
	.w3(32'h3c17617a),
	.w4(32'h3bf9f8b5),
	.w5(32'h3ca4563a),
	.w6(32'h3b8fa6fc),
	.w7(32'h3c3a073c),
	.w8(32'h3b259877),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0dce),
	.w1(32'h3be506d7),
	.w2(32'h3a46ddba),
	.w3(32'h3c4c382e),
	.w4(32'h3abd6682),
	.w5(32'h3c4e9522),
	.w6(32'h3bcfabee),
	.w7(32'h3b87d3f5),
	.w8(32'h3b661f1e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ac68),
	.w1(32'h3c21ce97),
	.w2(32'h3bba1d4c),
	.w3(32'hbc1a610b),
	.w4(32'h3c369576),
	.w5(32'hba5632cd),
	.w6(32'hba92480d),
	.w7(32'h3bea2075),
	.w8(32'h3c09e67f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb71af9),
	.w1(32'h3c5900be),
	.w2(32'h3c8c4f95),
	.w3(32'h3bc40fdd),
	.w4(32'hbac25dd0),
	.w5(32'h3c01e9f8),
	.w6(32'h3aa1811f),
	.w7(32'hbc5ec7bf),
	.w8(32'hbb295b5a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add7c7e),
	.w1(32'hbc35d6c4),
	.w2(32'h3af458e6),
	.w3(32'hbb1cdce8),
	.w4(32'hbc8d4e0c),
	.w5(32'h3b924ed9),
	.w6(32'h3b748519),
	.w7(32'hbc826745),
	.w8(32'hb996c2dc),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55d671),
	.w1(32'h3bc9bcf3),
	.w2(32'h3b73f773),
	.w3(32'h3c9e10fa),
	.w4(32'hbbf9a36d),
	.w5(32'hbbab615e),
	.w6(32'h3c09bc5e),
	.w7(32'hbc3f3c99),
	.w8(32'hbc3ac912),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c32b4),
	.w1(32'hbc4a1986),
	.w2(32'h3bbd3788),
	.w3(32'hbc2030f4),
	.w4(32'hbc8c1065),
	.w5(32'h3c3e7201),
	.w6(32'hbc2b79e2),
	.w7(32'hbc2a305c),
	.w8(32'h3bf2e894),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0185df),
	.w1(32'h3bca4edc),
	.w2(32'h3bf15ea0),
	.w3(32'h3c17fe2b),
	.w4(32'h3b517e4e),
	.w5(32'hba932202),
	.w6(32'h3bdde226),
	.w7(32'hbad0c8c5),
	.w8(32'h3ba07407),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa5cdb),
	.w1(32'hbb2a6723),
	.w2(32'hbb8328e9),
	.w3(32'hbc15666f),
	.w4(32'hba5718f8),
	.w5(32'hbbc388f9),
	.w6(32'hbc3ba105),
	.w7(32'hbb05aaba),
	.w8(32'hbb51e944),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58ad36),
	.w1(32'hbc6ff21f),
	.w2(32'hbb16d29b),
	.w3(32'hbc063b91),
	.w4(32'hbc552608),
	.w5(32'hb8a7bb44),
	.w6(32'hbc3d8701),
	.w7(32'hbc162e26),
	.w8(32'hbc3dfc0a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c415450),
	.w1(32'h3a111775),
	.w2(32'hbbc023b7),
	.w3(32'h3cb47b56),
	.w4(32'hbb95f3f2),
	.w5(32'hbbaa6b37),
	.w6(32'h3c2372da),
	.w7(32'h39f471da),
	.w8(32'hbbc411f7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff105),
	.w1(32'h3bbed93c),
	.w2(32'h3ae0f378),
	.w3(32'h3c37e547),
	.w4(32'h3c2057b0),
	.w5(32'hbb9d817e),
	.w6(32'h3a04690f),
	.w7(32'h3c0f6f10),
	.w8(32'h3b58b972),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc236508),
	.w1(32'h3b17cb46),
	.w2(32'hbc252844),
	.w3(32'hbc7ab359),
	.w4(32'h3c0d9eaf),
	.w5(32'hbc0945fc),
	.w6(32'hbbecddd0),
	.w7(32'h3bc7b05e),
	.w8(32'hbbb7a081),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ab846),
	.w1(32'hbb31cc7d),
	.w2(32'hbc15751a),
	.w3(32'hbc0e7fe3),
	.w4(32'h3b8439d0),
	.w5(32'h3bfe09d4),
	.w6(32'hbc6e4270),
	.w7(32'h3bdd5bdb),
	.w8(32'hbacdadd1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc8095),
	.w1(32'h3ba6048b),
	.w2(32'hbb89787c),
	.w3(32'hba78ac1b),
	.w4(32'h3a59413b),
	.w5(32'h3cc4b5c2),
	.w6(32'hbb7f43d8),
	.w7(32'hbbb659ee),
	.w8(32'hbb2621f2),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3911d6),
	.w1(32'hbc23c6a5),
	.w2(32'hbb319205),
	.w3(32'hbac22444),
	.w4(32'hbb83a1af),
	.w5(32'hbbb6a95b),
	.w6(32'hba53f14e),
	.w7(32'h3a5e6e41),
	.w8(32'hbc0bf16a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37bcac),
	.w1(32'h3c5a9a53),
	.w2(32'hbb2c6883),
	.w3(32'h3a32d218),
	.w4(32'h3d01210b),
	.w5(32'h3c8b26e6),
	.w6(32'hbb9cadce),
	.w7(32'h39d00cfd),
	.w8(32'h3bab69a6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298c60),
	.w1(32'hbb8a1995),
	.w2(32'hbcd2790a),
	.w3(32'hbc0d6cd0),
	.w4(32'hbc02a366),
	.w5(32'hbcb748c1),
	.w6(32'hbb08444c),
	.w7(32'hbb70febe),
	.w8(32'hbcd5fb8e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90d16c),
	.w1(32'h3c2f18bb),
	.w2(32'hbb7224c2),
	.w3(32'hbc8a3425),
	.w4(32'hbca5ad73),
	.w5(32'hbc5fe4aa),
	.w6(32'hbd229c95),
	.w7(32'hbd0f05bb),
	.w8(32'hbd18967a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39411f),
	.w1(32'h3c1b4ae2),
	.w2(32'h3c665f2b),
	.w3(32'hbc509d6e),
	.w4(32'h3ce2d0a1),
	.w5(32'h3c97846c),
	.w6(32'hbba30b6c),
	.w7(32'h3c89454b),
	.w8(32'h3c76dff2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a32b4),
	.w1(32'hba1c1ed9),
	.w2(32'hbb8d85b1),
	.w3(32'hbc8fc07b),
	.w4(32'hbbb7f417),
	.w5(32'h3bc82b9a),
	.w6(32'hbbdc21b6),
	.w7(32'hbbba78f9),
	.w8(32'hbacb94be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a860105),
	.w1(32'hbb537d9d),
	.w2(32'h3b789a15),
	.w3(32'hbb8002f6),
	.w4(32'hbb81281a),
	.w5(32'h3c2dd9d4),
	.w6(32'hb9372112),
	.w7(32'hbc01ed72),
	.w8(32'hbb884167),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e29ca),
	.w1(32'hbbb74bfb),
	.w2(32'hbaf20259),
	.w3(32'hbb3f6e13),
	.w4(32'hbc07e9b2),
	.w5(32'hba832a5d),
	.w6(32'hbb8e8849),
	.w7(32'hbc39f85e),
	.w8(32'h3abcc92a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed238d),
	.w1(32'h3b2dbf3a),
	.w2(32'h3bd59350),
	.w3(32'h3cb6e1cb),
	.w4(32'h3c10f10b),
	.w5(32'h3ae84e15),
	.w6(32'h3c508faf),
	.w7(32'h3bb7533d),
	.w8(32'h3bd34f99),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb49588),
	.w1(32'hbb1c130d),
	.w2(32'hbc03e025),
	.w3(32'h3c47e57f),
	.w4(32'hbc14d69a),
	.w5(32'hbba39fae),
	.w6(32'h3c5999c1),
	.w7(32'hbc0cad4b),
	.w8(32'hbc19a325),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8060),
	.w1(32'hbbea465c),
	.w2(32'h3bb0f6bd),
	.w3(32'hbc274ab9),
	.w4(32'hbc2278bb),
	.w5(32'h3b6e2df6),
	.w6(32'hbbca6e94),
	.w7(32'hbc173a50),
	.w8(32'h39b0e748),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93cc8c),
	.w1(32'h3ba766c1),
	.w2(32'h3bd6a968),
	.w3(32'h3c65a18d),
	.w4(32'hbc3f7ada),
	.w5(32'h3a9fbbb3),
	.w6(32'hbaf0718d),
	.w7(32'hbc2135be),
	.w8(32'hbb9d0ac8),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c758d),
	.w1(32'hbc19b676),
	.w2(32'h3aefa050),
	.w3(32'h3abd3b85),
	.w4(32'hbc8587f1),
	.w5(32'h3c28842a),
	.w6(32'h3b039cc7),
	.w7(32'hbad8d759),
	.w8(32'h3b4e5ce4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc57b01),
	.w1(32'h3b72c7fd),
	.w2(32'h3bb3e4b0),
	.w3(32'h3b89d38d),
	.w4(32'hba9c6bc7),
	.w5(32'h370043e6),
	.w6(32'hb955adec),
	.w7(32'hbbb1c8fd),
	.w8(32'hba9eb612),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c073ede),
	.w1(32'hba06a57c),
	.w2(32'hbaf83b3a),
	.w3(32'h3bec2fad),
	.w4(32'hbb5df6ab),
	.w5(32'hbb0277d4),
	.w6(32'h3bc88c71),
	.w7(32'hb9d63159),
	.w8(32'h3b73c904),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bd51e),
	.w1(32'h3baf2ed4),
	.w2(32'hbbf66d75),
	.w3(32'hba9cd938),
	.w4(32'h3c649a55),
	.w5(32'hbc543153),
	.w6(32'h3b0d3214),
	.w7(32'hbb41f15f),
	.w8(32'hbb23d587),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe461e4),
	.w1(32'hbb3a7ba5),
	.w2(32'hbb22ed5c),
	.w3(32'hbc42df23),
	.w4(32'hb98f0c10),
	.w5(32'hbbac58c5),
	.w6(32'h3b05d0ed),
	.w7(32'h39d4aa82),
	.w8(32'h3b57aa95),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a818),
	.w1(32'hbb56ee6f),
	.w2(32'h3c5fdefb),
	.w3(32'hbae24db9),
	.w4(32'hb8e90475),
	.w5(32'h3925baa3),
	.w6(32'h3bb75b52),
	.w7(32'h3c289db0),
	.w8(32'hbc220ef9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5a205),
	.w1(32'h3bf6156d),
	.w2(32'h3b8792d2),
	.w3(32'hbc5ad6d7),
	.w4(32'hbb2de4b1),
	.w5(32'hbb4c725c),
	.w6(32'hbb1c8640),
	.w7(32'hbbcf734e),
	.w8(32'hba5eca7c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1353),
	.w1(32'hbc3d7f98),
	.w2(32'h3c864c0b),
	.w3(32'h3b41c1ae),
	.w4(32'h3b4e14d9),
	.w5(32'hbb139112),
	.w6(32'h3bd6a8c6),
	.w7(32'hbb8df732),
	.w8(32'h3a06e663),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef00fc),
	.w1(32'h3c1d2390),
	.w2(32'h3c002229),
	.w3(32'hbc0a9315),
	.w4(32'h3b8b955a),
	.w5(32'h3b938628),
	.w6(32'h3ba2f2ea),
	.w7(32'h3c00829b),
	.w8(32'h3bc622c9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90e3fb),
	.w1(32'hba47461f),
	.w2(32'hb9ae0506),
	.w3(32'h3b519160),
	.w4(32'hbc1b9829),
	.w5(32'h3cebefa6),
	.w6(32'h3b861b6e),
	.w7(32'h3ad320c7),
	.w8(32'hbc4743a5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cc2ce),
	.w1(32'h3be126a4),
	.w2(32'h3cd57da9),
	.w3(32'h3c540e9f),
	.w4(32'hbaddbe2f),
	.w5(32'h3d061c60),
	.w6(32'h3c297a39),
	.w7(32'h3ab53edd),
	.w8(32'hbcb1298a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cff517),
	.w1(32'hbac97b3f),
	.w2(32'hbbc059e8),
	.w3(32'hbbcf24d4),
	.w4(32'hbc03c391),
	.w5(32'hbc017f55),
	.w6(32'h3c1c8936),
	.w7(32'hbbc8fdf2),
	.w8(32'hbb051dee),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a3901),
	.w1(32'h3ba49c2b),
	.w2(32'h3b41420b),
	.w3(32'hbbf17429),
	.w4(32'hbc36ee72),
	.w5(32'hbb8b87ce),
	.w6(32'hbbb40ba4),
	.w7(32'hbc33ca82),
	.w8(32'hbbb2ee61),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb854870),
	.w1(32'hbb9ff2cc),
	.w2(32'hbb958367),
	.w3(32'h3a0a16f1),
	.w4(32'hbb7d916c),
	.w5(32'hbb329ae8),
	.w6(32'h3be58d52),
	.w7(32'h3b5c2614),
	.w8(32'h3b3877c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba936be5),
	.w1(32'h3b4f5d8a),
	.w2(32'hbc8ec86f),
	.w3(32'hbae004d6),
	.w4(32'hbc40f0c1),
	.w5(32'hbb447f6e),
	.w6(32'hbb08f63a),
	.w7(32'hba7fb636),
	.w8(32'h3bb0497c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b167bc1),
	.w1(32'h3a4d5321),
	.w2(32'h3c11f484),
	.w3(32'h3c05d436),
	.w4(32'hbbe50012),
	.w5(32'hbc1651b7),
	.w6(32'h3a9b9741),
	.w7(32'h3b88b1d5),
	.w8(32'hbb7973eb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7429b),
	.w1(32'h3b56c1ab),
	.w2(32'h3b839360),
	.w3(32'hbc194145),
	.w4(32'hbc45e97c),
	.w5(32'hbbb8d004),
	.w6(32'hbb147562),
	.w7(32'hbb71d7a6),
	.w8(32'h3a2b5bb3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd896f),
	.w1(32'h3b81e3b6),
	.w2(32'h3946b5cb),
	.w3(32'h3a3946df),
	.w4(32'hbadc9284),
	.w5(32'h3aa7ee69),
	.w6(32'h3b9e3879),
	.w7(32'h39283c93),
	.w8(32'h3affef1b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ced069),
	.w1(32'h3c20d000),
	.w2(32'hbb842507),
	.w3(32'h3b8ebb2a),
	.w4(32'hbae79016),
	.w5(32'h3cea9fc5),
	.w6(32'hbbc5368d),
	.w7(32'h3bb97e75),
	.w8(32'hbc5f3645),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c0fb41),
	.w1(32'h3ba79b57),
	.w2(32'hbbd7bb4b),
	.w3(32'h3b3adc25),
	.w4(32'hbc3917f9),
	.w5(32'h3c6a5ba7),
	.w6(32'h3c392d79),
	.w7(32'h3aaf634f),
	.w8(32'h3c3191c2),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a18f6),
	.w1(32'hbb5944d0),
	.w2(32'hbb897c70),
	.w3(32'h3c826e68),
	.w4(32'hbbfc0795),
	.w5(32'hbba46e9c),
	.w6(32'h3bce5d15),
	.w7(32'hba60d6e0),
	.w8(32'h3a8b8496),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd990d3),
	.w1(32'h3b864b0c),
	.w2(32'h3bc1f10f),
	.w3(32'h3aa69bae),
	.w4(32'hbb8d2e19),
	.w5(32'h3c0acad4),
	.w6(32'h394c7f27),
	.w7(32'hbbb0afcb),
	.w8(32'hbc80db84),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d965c),
	.w1(32'h3a8e051d),
	.w2(32'hba01855f),
	.w3(32'hbb17ad6e),
	.w4(32'hbc52cf8b),
	.w5(32'hbc056de5),
	.w6(32'hbc76df07),
	.w7(32'hbc8a39a5),
	.w8(32'hbc8c8c11),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3898ee),
	.w1(32'h3ada44d5),
	.w2(32'hbbc6f015),
	.w3(32'h3b8f6846),
	.w4(32'hbba4508a),
	.w5(32'hbbb5bbb1),
	.w6(32'h3c04e77a),
	.w7(32'hbc474e54),
	.w8(32'hbc768222),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4b9b8),
	.w1(32'hbb283a45),
	.w2(32'h3bb457df),
	.w3(32'hbb30e7c3),
	.w4(32'h3c659511),
	.w5(32'hbbfa38a3),
	.w6(32'hbbaa6e32),
	.w7(32'h3bef8a23),
	.w8(32'h3bf4c212),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e930a0),
	.w1(32'hbb8d5f4f),
	.w2(32'h3bfe7c9d),
	.w3(32'hbc60dfe8),
	.w4(32'h3cb95fed),
	.w5(32'hbc80e5cc),
	.w6(32'hbb679cc8),
	.w7(32'h3c2d4e0b),
	.w8(32'h3b3f9ab8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7d523),
	.w1(32'h3baee25f),
	.w2(32'hbb31386c),
	.w3(32'hbcae57eb),
	.w4(32'h3b96ff42),
	.w5(32'hbc33552e),
	.w6(32'hbaead083),
	.w7(32'hb9d5c7e3),
	.w8(32'hbb5796c4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc52a20),
	.w1(32'h3bb75c8b),
	.w2(32'h3b8a6267),
	.w3(32'hbb2c9470),
	.w4(32'h3b1ee241),
	.w5(32'hbb69bd0f),
	.w6(32'hbb33ff54),
	.w7(32'hbb7f7eba),
	.w8(32'h3cc7c371),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0baaa7),
	.w1(32'hbc0f8bab),
	.w2(32'hbb120d85),
	.w3(32'h3c858f1a),
	.w4(32'hbb73d140),
	.w5(32'hbb99f667),
	.w6(32'hbbc6eaaf),
	.w7(32'hbb72344a),
	.w8(32'h3beb2848),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01d197),
	.w1(32'h3b24efbd),
	.w2(32'h3b573f62),
	.w3(32'hbb3ac05a),
	.w4(32'h3af8877f),
	.w5(32'hb9c4bae2),
	.w6(32'h39b6e317),
	.w7(32'h3a600e5f),
	.w8(32'h3a95f6a9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1afe62),
	.w1(32'hbb29cae8),
	.w2(32'h3b3027ee),
	.w3(32'hbb87e0bf),
	.w4(32'h3bcb63a2),
	.w5(32'h3c439ab7),
	.w6(32'hbbf2e4da),
	.w7(32'hbae9562e),
	.w8(32'h3ba93d29),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cf83f),
	.w1(32'h3b8ed02f),
	.w2(32'h3b684994),
	.w3(32'h3b80ce35),
	.w4(32'hbb3aa373),
	.w5(32'hbbca2305),
	.w6(32'h3bb25572),
	.w7(32'hbaa05878),
	.w8(32'hbbce2903),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ecea4),
	.w1(32'hbb559f5f),
	.w2(32'h3c033fa7),
	.w3(32'hbc0a0a4a),
	.w4(32'h3b9d81ec),
	.w5(32'hbba6340d),
	.w6(32'hb9cdf3b2),
	.w7(32'h3b9e5b5e),
	.w8(32'h3aee4d95),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61166f),
	.w1(32'h3adbafce),
	.w2(32'hba9e7826),
	.w3(32'hbbd53046),
	.w4(32'hbb4d5101),
	.w5(32'hbc1937d0),
	.w6(32'h3bb0e4f7),
	.w7(32'hbbdea329),
	.w8(32'h3bc5f59a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ef90),
	.w1(32'h3caaadd7),
	.w2(32'hbc2f6b4c),
	.w3(32'hbbd84bdc),
	.w4(32'hbca958ff),
	.w5(32'h3af7b184),
	.w6(32'hbae45c58),
	.w7(32'hbce7dc47),
	.w8(32'h3c434f86),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f653),
	.w1(32'hbb9db558),
	.w2(32'h3c3ec4b9),
	.w3(32'h3cc78f4a),
	.w4(32'hbc944f0f),
	.w5(32'h3cd62160),
	.w6(32'hbc0dbb79),
	.w7(32'hbbc1062a),
	.w8(32'hbce9faf2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7c7950),
	.w1(32'hbb3edb80),
	.w2(32'h3ba292c6),
	.w3(32'hbc383160),
	.w4(32'h3c4b3eea),
	.w5(32'hbb8af91f),
	.w6(32'h3ba6f238),
	.w7(32'hbb1dfc33),
	.w8(32'hba5b95db),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b014c5a),
	.w1(32'h3a36ece5),
	.w2(32'h3b39690a),
	.w3(32'hbc026cbc),
	.w4(32'h3b1a5a66),
	.w5(32'h3b2f934d),
	.w6(32'h39e2f04a),
	.w7(32'hbb02f389),
	.w8(32'h3b6ed3d2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa063f),
	.w1(32'hbb34f3ba),
	.w2(32'h3bee4be3),
	.w3(32'h3b3c9c3b),
	.w4(32'hba3298e4),
	.w5(32'h3b8bc176),
	.w6(32'h3b3f560d),
	.w7(32'h3a80d23a),
	.w8(32'hbc35e50b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9498a),
	.w1(32'hbaf47df2),
	.w2(32'hbb807703),
	.w3(32'hbbcf911b),
	.w4(32'h3c4247a0),
	.w5(32'hbbd1e7f7),
	.w6(32'hbb5cea02),
	.w7(32'h3b776402),
	.w8(32'h3c4df131),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0935ad),
	.w1(32'hbb75071b),
	.w2(32'h3b107b05),
	.w3(32'h3bea7171),
	.w4(32'h3bc38bf0),
	.w5(32'hbc664de8),
	.w6(32'hbab025c5),
	.w7(32'hbbf6fad8),
	.w8(32'hb9c693c2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41e863),
	.w1(32'h3a3b63d2),
	.w2(32'h3c0f7581),
	.w3(32'hbb576078),
	.w4(32'h3c400ae9),
	.w5(32'hbc4f2671),
	.w6(32'hbba2e124),
	.w7(32'hbc85428f),
	.w8(32'h3bf64b4d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97934b),
	.w1(32'hb995a626),
	.w2(32'h3bdbe278),
	.w3(32'h3baaf4ec),
	.w4(32'h3b910df5),
	.w5(32'hbb63a6df),
	.w6(32'h3b134957),
	.w7(32'hbb1fbdd6),
	.w8(32'h3b13e76a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8821d8),
	.w1(32'hb978398b),
	.w2(32'h3aeb60d9),
	.w3(32'hbbc12028),
	.w4(32'h3ae588c8),
	.w5(32'hbaa9005e),
	.w6(32'hbaa1425f),
	.w7(32'h3bcd70d2),
	.w8(32'h3c40958a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b549f55),
	.w1(32'h3c1b9700),
	.w2(32'hbc26860f),
	.w3(32'h3aaba0ed),
	.w4(32'hbb1469ff),
	.w5(32'h3b4ac401),
	.w6(32'hbb626828),
	.w7(32'h3aceecf1),
	.w8(32'h3ce6b067),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e713),
	.w1(32'hbcab9e14),
	.w2(32'h3cfa13af),
	.w3(32'h3cef627a),
	.w4(32'hbc2f0ecf),
	.w5(32'h3ca8a7f9),
	.w6(32'hbc1c4f95),
	.w7(32'h3ba15f41),
	.w8(32'hbcee9d55),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d48b),
	.w1(32'hbb9fc55d),
	.w2(32'h3b1b6e89),
	.w3(32'hba8daf76),
	.w4(32'h3a88645a),
	.w5(32'h3c27ff3b),
	.w6(32'h3c5bdbc7),
	.w7(32'hbb314cad),
	.w8(32'hbc20e5d1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa05513),
	.w1(32'h3b7ae1aa),
	.w2(32'hbbf6cfa8),
	.w3(32'hbbef8783),
	.w4(32'hba66a943),
	.w5(32'hbaf87075),
	.w6(32'hbb00aedc),
	.w7(32'hba83743b),
	.w8(32'hba7368df),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990179e),
	.w1(32'h3b49ef3f),
	.w2(32'h3b8d7657),
	.w3(32'hbb4b9a33),
	.w4(32'h3bce4e10),
	.w5(32'hbc4e7d99),
	.w6(32'hbb12349c),
	.w7(32'h3b1e3d31),
	.w8(32'h3c2e1aef),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18924),
	.w1(32'hbc60a6c4),
	.w2(32'h3c335039),
	.w3(32'h3c4aef38),
	.w4(32'h3cd5f335),
	.w5(32'hbc57c367),
	.w6(32'hbbeac9bc),
	.w7(32'h3c00323d),
	.w8(32'hbbe2a897),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4d5b4),
	.w1(32'hbb6f74a3),
	.w2(32'hbb02bdf2),
	.w3(32'hbccf1fa9),
	.w4(32'hbc2a956e),
	.w5(32'h3c18ffef),
	.w6(32'h3baa1b0d),
	.w7(32'hbb4f9d0a),
	.w8(32'h3c6bfe2d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dd4ad),
	.w1(32'h3b7ff57d),
	.w2(32'hbc8ffdc5),
	.w3(32'h3c393513),
	.w4(32'h3c1db3f5),
	.w5(32'hbc794d59),
	.w6(32'h3c1a225c),
	.w7(32'hbb607f63),
	.w8(32'h3cb2f0e2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c478650),
	.w1(32'h3b0c52ac),
	.w2(32'h3bca4e41),
	.w3(32'h3ca5034f),
	.w4(32'hb9cbc37f),
	.w5(32'h3b5f92ab),
	.w6(32'hbca2954e),
	.w7(32'h3af7b711),
	.w8(32'hb8b12f28),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad907f3),
	.w1(32'hbb8f503c),
	.w2(32'hbb82f5d1),
	.w3(32'hbb413724),
	.w4(32'hbb4dca70),
	.w5(32'hbb3500d1),
	.w6(32'h3b17bfa9),
	.w7(32'hba2b44db),
	.w8(32'h39e3e700),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676dfa),
	.w1(32'h3ba0124c),
	.w2(32'hbc75cffe),
	.w3(32'h3c013e18),
	.w4(32'hbc2bb451),
	.w5(32'hbb4788e9),
	.w6(32'h3adc4f1d),
	.w7(32'hbaed5c6d),
	.w8(32'h3c8a797d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f0f8a),
	.w1(32'h3959611a),
	.w2(32'hbc65670e),
	.w3(32'h3ca04c94),
	.w4(32'hbad26fe9),
	.w5(32'hbce0a32c),
	.w6(32'hbc1d26e9),
	.w7(32'hbbff3faf),
	.w8(32'h3c8e2d85),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338492),
	.w1(32'hbba97abf),
	.w2(32'h3c15f679),
	.w3(32'h3c47f4f7),
	.w4(32'h3cbbf3fe),
	.w5(32'hbc755a78),
	.w6(32'hbc1fdcc5),
	.w7(32'hba7d67aa),
	.w8(32'h3c818b85),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6f234),
	.w1(32'hbc31f844),
	.w2(32'h3c90388d),
	.w3(32'h3a0f144a),
	.w4(32'h3c26e500),
	.w5(32'h3cadf777),
	.w6(32'hbb3ad490),
	.w7(32'hbb8397e4),
	.w8(32'hbbf52d82),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0557f7),
	.w1(32'hbbec9edc),
	.w2(32'hbc19513e),
	.w3(32'h3b9db4cd),
	.w4(32'hbbc899ec),
	.w5(32'hbc03dac5),
	.w6(32'h3c9cca00),
	.w7(32'hbc094261),
	.w8(32'hbba354b6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05c29b),
	.w1(32'h3b351f79),
	.w2(32'h39c57dec),
	.w3(32'hbc55cf16),
	.w4(32'hbb972361),
	.w5(32'hbc04335f),
	.w6(32'hbb856deb),
	.w7(32'h3a714f39),
	.w8(32'hbaaeb7c5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule