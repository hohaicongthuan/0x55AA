module layer_6_featuremap_5(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c050621),
	.w1(32'h3bf3516f),
	.w2(32'h3b8ad235),
	.w3(32'h3be6b26f),
	.w4(32'h3c066795),
	.w5(32'h3b2426fd),
	.w6(32'h3be3664a),
	.w7(32'h3c06d958),
	.w8(32'h3b4c834c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a045f57),
	.w1(32'h39a7e7d7),
	.w2(32'hb8d74552),
	.w3(32'h396a5618),
	.w4(32'h38e68193),
	.w5(32'hb8c9b53c),
	.w6(32'h38db0546),
	.w7(32'hb586f417),
	.w8(32'hb9204c0a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2414fe),
	.w1(32'hbc3f705c),
	.w2(32'hb99eb17c),
	.w3(32'h3a22a0a1),
	.w4(32'hbbc2858c),
	.w5(32'h3bf253bd),
	.w6(32'h3aa56cf0),
	.w7(32'hbc109ba2),
	.w8(32'h39dda51d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c160b68),
	.w1(32'h3b9c2f24),
	.w2(32'h3b9d5477),
	.w3(32'h3b620b5d),
	.w4(32'h3a6d9569),
	.w5(32'h3bd5f8d7),
	.w6(32'h3bae2b60),
	.w7(32'h3ac93e2a),
	.w8(32'h3b9c57b9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f63e4c),
	.w1(32'hb9cda62e),
	.w2(32'h39b71915),
	.w3(32'hba23746d),
	.w4(32'h3a67fd91),
	.w5(32'hba24414e),
	.w6(32'h3a174fac),
	.w7(32'h3aa827d7),
	.w8(32'hba728203),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a824a47),
	.w1(32'h3993f9f4),
	.w2(32'h39898586),
	.w3(32'h3a58eb90),
	.w4(32'h39cdf98a),
	.w5(32'h39aedb61),
	.w6(32'h3a554e87),
	.w7(32'h3a590014),
	.w8(32'h398fcf30),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914fa8),
	.w1(32'h3bb00cac),
	.w2(32'h3bfb0bb1),
	.w3(32'h3c08dc1f),
	.w4(32'h3c00340a),
	.w5(32'h3c0ee3f3),
	.w6(32'h3c0ffc06),
	.w7(32'h3c1191d9),
	.w8(32'h3c183fd7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb29f0),
	.w1(32'hba32950d),
	.w2(32'hb97324a4),
	.w3(32'hba2896b7),
	.w4(32'h38f696c0),
	.w5(32'h39aa22f7),
	.w6(32'hbaa9665a),
	.w7(32'hb98b1c9b),
	.w8(32'hb9106de8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27b640),
	.w1(32'hbc33d91e),
	.w2(32'hbb03d45a),
	.w3(32'hbbffe872),
	.w4(32'hbc13f511),
	.w5(32'hbb396812),
	.w6(32'hbbfcd01b),
	.w7(32'hbc109f59),
	.w8(32'hba87242a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3df6e2),
	.w1(32'h39917c49),
	.w2(32'hba77a0cf),
	.w3(32'h3b17ff1e),
	.w4(32'h3a51b3fd),
	.w5(32'h3ac1c80a),
	.w6(32'h3b78c404),
	.w7(32'h3b0ecf6e),
	.w8(32'h3b198342),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9990b0),
	.w1(32'hbc962337),
	.w2(32'hbbb44618),
	.w3(32'hbc66e13b),
	.w4(32'hbc741db3),
	.w5(32'hbc08293a),
	.w6(32'hbc716375),
	.w7(32'hbc77bacd),
	.w8(32'hbc54e11d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38abf97e),
	.w1(32'h3a01571b),
	.w2(32'h3a58359a),
	.w3(32'h39191535),
	.w4(32'h39900690),
	.w5(32'h3a053903),
	.w6(32'h391ee2ad),
	.w7(32'h3844c2e2),
	.w8(32'h3979ea8a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f789a9),
	.w1(32'hb6247204),
	.w2(32'hb5f9a50a),
	.w3(32'h389b38fe),
	.w4(32'h3823cf64),
	.w5(32'h37dbd6e5),
	.w6(32'h3830860f),
	.w7(32'h3823b21c),
	.w8(32'h37f6e0a7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb55bd6),
	.w1(32'hbcca570d),
	.w2(32'hbbed20bb),
	.w3(32'hbc9a484e),
	.w4(32'hbcadbb5c),
	.w5(32'hbc186cd2),
	.w6(32'hbca08c0d),
	.w7(32'hbcaa1e77),
	.w8(32'hbc6508f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c8e41),
	.w1(32'hbb46d216),
	.w2(32'hbb1d00e2),
	.w3(32'hbb216ded),
	.w4(32'hbb6fadd1),
	.w5(32'hba9c29a3),
	.w6(32'hba83ffb9),
	.w7(32'hbb5b17e6),
	.w8(32'hbab411fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ecc16),
	.w1(32'hbb99e73e),
	.w2(32'hbb5b0d76),
	.w3(32'hbbb810b2),
	.w4(32'hbb8c4a2c),
	.w5(32'hb71ae85e),
	.w6(32'hbbb219b5),
	.w7(32'hbba18a0c),
	.w8(32'h360a8a87),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097b58),
	.w1(32'hbc51556c),
	.w2(32'h3bd18ee3),
	.w3(32'hbc3be921),
	.w4(32'hbc41f2f9),
	.w5(32'h3c8947f5),
	.w6(32'hbbd0f483),
	.w7(32'hbc25ce7b),
	.w8(32'h3c884452),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381c3957),
	.w1(32'h381be23a),
	.w2(32'hb7c50ded),
	.w3(32'hb5cbd908),
	.w4(32'h36ce8726),
	.w5(32'hb8633c5c),
	.w6(32'hb7366032),
	.w7(32'hb78f024f),
	.w8(32'hb8a14385),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba929b),
	.w1(32'h3928b72a),
	.w2(32'hbb3dc466),
	.w3(32'h3b942e38),
	.w4(32'h3a3c4d18),
	.w5(32'hb9fdd5c0),
	.w6(32'h3ba85293),
	.w7(32'h3a929703),
	.w8(32'h3a0b4781),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86a509),
	.w1(32'hbb21ffef),
	.w2(32'hb92c3316),
	.w3(32'hba9229b7),
	.w4(32'hbadcf867),
	.w5(32'h3aae6663),
	.w6(32'h38198fa8),
	.w7(32'hba826450),
	.w8(32'h3b13f54d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801ba1),
	.w1(32'h3a921ae6),
	.w2(32'h3adc0844),
	.w3(32'h39d004cb),
	.w4(32'hb9b696b8),
	.w5(32'h39f3dde6),
	.w6(32'h3a5e8a75),
	.w7(32'hba827f48),
	.w8(32'hba5261aa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde81ff),
	.w1(32'hbcdb8e26),
	.w2(32'hbc21bac7),
	.w3(32'hbcd2be38),
	.w4(32'hbccd198b),
	.w5(32'hbc2bbd71),
	.w6(32'hbcaab513),
	.w7(32'hbcc28f54),
	.w8(32'hbc5c4a9c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265737),
	.w1(32'hba98bf73),
	.w2(32'hba367591),
	.w3(32'hba9ccb93),
	.w4(32'hb9453f13),
	.w5(32'hb80812a0),
	.w6(32'hbad27198),
	.w7(32'hba454dba),
	.w8(32'hb9abc2cc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd22855c),
	.w1(32'hbd39c873),
	.w2(32'hbd12664b),
	.w3(32'hbd0efeaa),
	.w4(32'hbd300301),
	.w5(32'hbd2590b3),
	.w6(32'hbcfde4a6),
	.w7(32'hbd0e9e73),
	.w8(32'hbd2b2d1a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf836d8),
	.w1(32'h3c824904),
	.w2(32'h3c63eed5),
	.w3(32'h3c81194d),
	.w4(32'h3c15eafb),
	.w5(32'h3cc2a37d),
	.w6(32'h3cca528f),
	.w7(32'h3c635ca7),
	.w8(32'h3c951892),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bc2ad),
	.w1(32'hbba25849),
	.w2(32'hb7f30cfc),
	.w3(32'hbb14825b),
	.w4(32'hbc5ec166),
	.w5(32'h3c04753c),
	.w6(32'h3bad0a08),
	.w7(32'hbbfb4489),
	.w8(32'h3beef335),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc340ad7),
	.w1(32'hbc916491),
	.w2(32'hbc6bd513),
	.w3(32'hbc2a7515),
	.w4(32'hbc908fc7),
	.w5(32'hbca38f18),
	.w6(32'hbc6879e8),
	.w7(32'hbc9fe8e0),
	.w8(32'hbca0206b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3597b1),
	.w1(32'hbb8007bb),
	.w2(32'h393bce74),
	.w3(32'hbb76a8c6),
	.w4(32'hbb08b237),
	.w5(32'h38c81dcd),
	.w6(32'hbb46a13c),
	.w7(32'hba8d7b2c),
	.w8(32'h3a1ad2c2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb781ef5),
	.w1(32'hbb43787a),
	.w2(32'hbad9b97c),
	.w3(32'hbb773fb0),
	.w4(32'hbb544e74),
	.w5(32'hbafe10a2),
	.w6(32'hbb7541d8),
	.w7(32'hbb42809d),
	.w8(32'hbb11db8b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d505e2d),
	.w1(32'hbc4a1ce2),
	.w2(32'hbd84aae1),
	.w3(32'hbb5010d2),
	.w4(32'hbd23d9c6),
	.w5(32'hbd06c516),
	.w6(32'h3b63bf9d),
	.w7(32'hbd1e1c82),
	.w8(32'hbc0f9067),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3884ea67),
	.w1(32'hbbe4d277),
	.w2(32'hbc8a7a73),
	.w3(32'h386fa205),
	.w4(32'h3c2c1c17),
	.w5(32'h3c8b6ee8),
	.w6(32'hb98161d8),
	.w7(32'hbbd264a6),
	.w8(32'h3cccee9e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3801d1),
	.w1(32'hbd45e35d),
	.w2(32'h3db71c5f),
	.w3(32'hbd0093ee),
	.w4(32'hbd008477),
	.w5(32'hbd494db7),
	.w6(32'hbd23bff1),
	.w7(32'hbd5e43db),
	.w8(32'hbd04b89d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7a6eb4),
	.w1(32'hbd185773),
	.w2(32'h3df5ac87),
	.w3(32'hbce6fc21),
	.w4(32'h3c0c6354),
	.w5(32'hbd1e8013),
	.w6(32'h3c9f0486),
	.w7(32'hbd141fd1),
	.w8(32'hbcbf642e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd62a7dd),
	.w1(32'h3bdcdfa1),
	.w2(32'hbb7f588c),
	.w3(32'h3cd699ee),
	.w4(32'hba3681a8),
	.w5(32'h3aa3a6f2),
	.w6(32'h3c803cbb),
	.w7(32'hbc719ac0),
	.w8(32'h3b1b710d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf41c85),
	.w1(32'h3c1579d4),
	.w2(32'hbcf430aa),
	.w3(32'h3be7dbc4),
	.w4(32'h3b99ac76),
	.w5(32'hbc8eeab2),
	.w6(32'h3c7125c3),
	.w7(32'h3c20a4bd),
	.w8(32'hbabc592a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc4a7c),
	.w1(32'h3d11130d),
	.w2(32'hbe20c5a4),
	.w3(32'hbcb7a7d3),
	.w4(32'hbd0d78f8),
	.w5(32'h3caafcbc),
	.w6(32'hbd277ef0),
	.w7(32'h3b379c46),
	.w8(32'hbcdd19b9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d161531),
	.w1(32'h3c16a476),
	.w2(32'hbbdedb88),
	.w3(32'hbc28e00a),
	.w4(32'h3b59dc55),
	.w5(32'h3a99fb1d),
	.w6(32'h3b04048a),
	.w7(32'hbb4762ce),
	.w8(32'hbbd83abe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf98af5),
	.w1(32'hbca235b5),
	.w2(32'hbd41fbf4),
	.w3(32'hba7d7732),
	.w4(32'hbb484dc7),
	.w5(32'hbb3d29dd),
	.w6(32'hbc006899),
	.w7(32'hbc56af4e),
	.w8(32'h3bac0816),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb31d40),
	.w1(32'h3a79727f),
	.w2(32'h3aaf9777),
	.w3(32'hbc456d4c),
	.w4(32'hbb0d18ab),
	.w5(32'hbb7e8e54),
	.w6(32'hbbb73d07),
	.w7(32'hbbbfe956),
	.w8(32'h3ac8d966),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce29ec0),
	.w1(32'hbd1b08df),
	.w2(32'h3c5cd40b),
	.w3(32'hbc51b360),
	.w4(32'hbc898352),
	.w5(32'h3a381753),
	.w6(32'hbcf129cc),
	.w7(32'hbd2e08a4),
	.w8(32'hbb3ad73b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6db627),
	.w1(32'hbb90f49d),
	.w2(32'hbb321243),
	.w3(32'hbc66e04b),
	.w4(32'hbbc2af4a),
	.w5(32'hbc04bf09),
	.w6(32'hbb8edf5b),
	.w7(32'hbc936f91),
	.w8(32'h3bd86875),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aee83),
	.w1(32'h3a6a5630),
	.w2(32'hbb20bc2d),
	.w3(32'h3c13ad0e),
	.w4(32'hbbe15128),
	.w5(32'h3b82b8fe),
	.w6(32'hbb59beb4),
	.w7(32'hbc0f722d),
	.w8(32'h3aeb5496),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935bee1),
	.w1(32'h3c25f0b8),
	.w2(32'hbcfddeba),
	.w3(32'h3af630ef),
	.w4(32'hbbfa79d1),
	.w5(32'h39b0a6b4),
	.w6(32'h3bc44fb6),
	.w7(32'h3c5f3608),
	.w8(32'h3ba6c114),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8969c7),
	.w1(32'h3c6e22e1),
	.w2(32'hbd3143cf),
	.w3(32'h3c4e2914),
	.w4(32'hbd155122),
	.w5(32'h3c379bb5),
	.w6(32'hbce95101),
	.w7(32'hbc93c3b9),
	.w8(32'h3d08f4a5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd299806),
	.w1(32'hbd499c50),
	.w2(32'h3b4a625d),
	.w3(32'hbcd7cba5),
	.w4(32'hbd33c2fe),
	.w5(32'hbbfe54ac),
	.w6(32'hbc8160a4),
	.w7(32'h3bdd2344),
	.w8(32'hbce2dcad),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17d11e),
	.w1(32'hbba80f8c),
	.w2(32'h3cf34969),
	.w3(32'h3bc2cffe),
	.w4(32'h3c8c0b61),
	.w5(32'h3b26e1ca),
	.w6(32'h3c1e0947),
	.w7(32'hbc49b0bf),
	.w8(32'h3c16d28f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fbb2b),
	.w1(32'hbd0ff491),
	.w2(32'h3c5b54b0),
	.w3(32'h3bb00606),
	.w4(32'h3c253207),
	.w5(32'hbd556681),
	.w6(32'h3bd31690),
	.w7(32'hbd2b8986),
	.w8(32'hbc99aa7c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd80421),
	.w1(32'h3bea2cc2),
	.w2(32'hbc269937),
	.w3(32'hbb878635),
	.w4(32'h3b0e531b),
	.w5(32'hbcbcbffd),
	.w6(32'hba9c1b49),
	.w7(32'h3c6bca6e),
	.w8(32'h3c3f662f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e8a7d),
	.w1(32'hbda6e8eb),
	.w2(32'hbca67231),
	.w3(32'hbaf37642),
	.w4(32'h3d40752d),
	.w5(32'hbd9909e5),
	.w6(32'hbc2af3b5),
	.w7(32'h3db2e446),
	.w8(32'hbd8af0a8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dc79f94),
	.w1(32'hbd1a2ad5),
	.w2(32'h3c889992),
	.w3(32'h3c4bc4e0),
	.w4(32'h3c0e34b3),
	.w5(32'hbcb93073),
	.w6(32'h3c4d3e8c),
	.w7(32'hbc4d72e1),
	.w8(32'hbb9a2905),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d379163),
	.w1(32'h3c4bab94),
	.w2(32'h3c243c70),
	.w3(32'hbba81e0a),
	.w4(32'h3ba61eee),
	.w5(32'h3c5a684a),
	.w6(32'h3c1cdd1f),
	.w7(32'hba17167c),
	.w8(32'h3c4c50a1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8639d0),
	.w1(32'hbd8961ae),
	.w2(32'h3df70baa),
	.w3(32'h3c0a0a97),
	.w4(32'hbc52b4ec),
	.w5(32'hbd1980a3),
	.w6(32'h3d131beb),
	.w7(32'hbc3a0a8c),
	.w8(32'hbbb031b3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc6d2b8),
	.w1(32'hbcea324d),
	.w2(32'hbcacaa56),
	.w3(32'h3c5c9912),
	.w4(32'hbc776015),
	.w5(32'hbc156473),
	.w6(32'hbc02c1a9),
	.w7(32'hbd1932ff),
	.w8(32'h3cac600b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceab15),
	.w1(32'h3cd9f0eb),
	.w2(32'h3a381616),
	.w3(32'h3b1a3c80),
	.w4(32'h3c9d3b4c),
	.w5(32'h3913030d),
	.w6(32'h3c731eed),
	.w7(32'h3ca98aee),
	.w8(32'h3c592a62),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f8d28),
	.w1(32'hbc8a1183),
	.w2(32'hbc82f856),
	.w3(32'hbb59b337),
	.w4(32'h3c4afe9d),
	.w5(32'hbcbf597a),
	.w6(32'h3b862960),
	.w7(32'h3ba3d692),
	.w8(32'h3c3a7e95),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0580),
	.w1(32'h3d2aa501),
	.w2(32'h3cd33bff),
	.w3(32'h3a88a879),
	.w4(32'hbcad95d5),
	.w5(32'h3d03dc55),
	.w6(32'hbc0e2409),
	.w7(32'hbd49a61e),
	.w8(32'h3af9ca6c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9b5c27),
	.w1(32'h3cc78cd6),
	.w2(32'h3c819f87),
	.w3(32'hb9120f5f),
	.w4(32'hbd55724a),
	.w5(32'h3ca1dfde),
	.w6(32'hbc709bb4),
	.w7(32'hbc2a84d2),
	.w8(32'h3c34fd29),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca75df0),
	.w1(32'hbc884574),
	.w2(32'h3cc51133),
	.w3(32'h3c3d56b5),
	.w4(32'h3ad7c4b4),
	.w5(32'h396de2ff),
	.w6(32'hbbad972a),
	.w7(32'h3b67a82a),
	.w8(32'hbc0bb3b0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ef4b4),
	.w1(32'hbd1fc3bd),
	.w2(32'hbce96157),
	.w3(32'hbc1074fa),
	.w4(32'hbae1be8e),
	.w5(32'hbc331399),
	.w6(32'hbc2011cb),
	.w7(32'h39053d7a),
	.w8(32'h3b4d9fd0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae32a74),
	.w1(32'hbd054343),
	.w2(32'hbbc52a38),
	.w3(32'hbb9f4d68),
	.w4(32'hbd07fe23),
	.w5(32'h3b5efe22),
	.w6(32'h3d0fc204),
	.w7(32'hbd42dd3d),
	.w8(32'h3cb62c06),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1a8e),
	.w1(32'hbcebf603),
	.w2(32'hbc90d0c9),
	.w3(32'hbcff5cc9),
	.w4(32'hbd17b2f9),
	.w5(32'hbc4b7e25),
	.w6(32'h3c280f78),
	.w7(32'h3c35a91e),
	.w8(32'hba8870f1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9306e),
	.w1(32'h3cd6b4ff),
	.w2(32'hbcaae22d),
	.w3(32'hbc7fef44),
	.w4(32'hbc7b4715),
	.w5(32'h3c87c3ff),
	.w6(32'hbc9e9812),
	.w7(32'h3cbbc53a),
	.w8(32'h3c3d3360),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc011a52),
	.w1(32'h3c420b6a),
	.w2(32'hbcffa68c),
	.w3(32'h3c226269),
	.w4(32'h3c73fb95),
	.w5(32'hbcac8838),
	.w6(32'hba280559),
	.w7(32'hbbbc293a),
	.w8(32'hbc350374),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe610c7),
	.w1(32'hbc0eaf82),
	.w2(32'h3b88b590),
	.w3(32'hbba7c1de),
	.w4(32'hbb9216a9),
	.w5(32'h3999beba),
	.w6(32'hbad68bd0),
	.w7(32'hbb00291f),
	.w8(32'hbb75f355),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule