module layer_8_featuremap_220(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8ec0a),
	.w1(32'hbc89e5c9),
	.w2(32'hbd081046),
	.w3(32'hbc35410e),
	.w4(32'h3cea02c5),
	.w5(32'hbbfa7d31),
	.w6(32'hbbabf178),
	.w7(32'hbaf73bbd),
	.w8(32'h3a8ddb8b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844f3d),
	.w1(32'h3b60ea66),
	.w2(32'h3ae820c1),
	.w3(32'hbc59922f),
	.w4(32'h3b072ec1),
	.w5(32'h3a15dcbd),
	.w6(32'h3b57d4c7),
	.w7(32'h3b1babd1),
	.w8(32'hb9a2c453),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9feafac),
	.w1(32'hbb23daf4),
	.w2(32'h3b74d278),
	.w3(32'h3b6780ed),
	.w4(32'h3b5fc4c8),
	.w5(32'hbb4ffc19),
	.w6(32'h3b4554c3),
	.w7(32'h3bf9b629),
	.w8(32'h3ad10a53),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a45d6),
	.w1(32'hbc929838),
	.w2(32'hbc0af3f2),
	.w3(32'hbc00858e),
	.w4(32'h3cade2d0),
	.w5(32'hbc122d9e),
	.w6(32'hbbb794b7),
	.w7(32'h3c2872a6),
	.w8(32'hbc69f611),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03182a),
	.w1(32'hbb12ce79),
	.w2(32'hbb470e6e),
	.w3(32'hbbeeb5ee),
	.w4(32'h3a4595ee),
	.w5(32'hbaf5dbc0),
	.w6(32'h398975e5),
	.w7(32'h3963e1d9),
	.w8(32'h3a18488b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc307488),
	.w1(32'hbbb3f521),
	.w2(32'h3b0fc641),
	.w3(32'hbb9d8ec8),
	.w4(32'hbac7b35c),
	.w5(32'hbcb962dd),
	.w6(32'hbc4da823),
	.w7(32'h395c7e77),
	.w8(32'hbc359af8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8aa5b),
	.w1(32'hbb5461b1),
	.w2(32'hba79c670),
	.w3(32'hba364288),
	.w4(32'hbb9636cd),
	.w5(32'hbbec6000),
	.w6(32'hba915b02),
	.w7(32'hbb0334df),
	.w8(32'hbae2c4a4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab55ca),
	.w1(32'h3bf0a603),
	.w2(32'hbb986680),
	.w3(32'hbc104c2e),
	.w4(32'hbb11ef5d),
	.w5(32'hbc00fd36),
	.w6(32'hbb63606a),
	.w7(32'h3c2b9cfd),
	.w8(32'hbbc8c741),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08808a),
	.w1(32'hbbab6b60),
	.w2(32'hbb68a497),
	.w3(32'h3a6f903a),
	.w4(32'hbbd5d3bf),
	.w5(32'hbb058153),
	.w6(32'hbb47ad88),
	.w7(32'h3a51d3ef),
	.w8(32'h3a88a434),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91aa77),
	.w1(32'h3bc37b5f),
	.w2(32'hbab21355),
	.w3(32'hba530c49),
	.w4(32'hbcad3e68),
	.w5(32'h3c40920b),
	.w6(32'hbbef4721),
	.w7(32'hbbb1519c),
	.w8(32'h3ae5e0e6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd033c63),
	.w1(32'hbce3b605),
	.w2(32'h3b2c0819),
	.w3(32'h3c07c279),
	.w4(32'h3bb6e0cd),
	.w5(32'hbcfee3fe),
	.w6(32'h3bc95867),
	.w7(32'h3c818c9a),
	.w8(32'hbc573776),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d9858),
	.w1(32'hbc154215),
	.w2(32'hbc481e3b),
	.w3(32'hbc6d6e5c),
	.w4(32'hbc23fbeb),
	.w5(32'hbc3936f9),
	.w6(32'hbaddc8ed),
	.w7(32'hbb666e6d),
	.w8(32'hbc117944),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58d026),
	.w1(32'hbb9eb453),
	.w2(32'h3c8c3dc8),
	.w3(32'hbbaaa935),
	.w4(32'hbc55ee32),
	.w5(32'hb9d0df3c),
	.w6(32'h3c01d100),
	.w7(32'h3c4eaa65),
	.w8(32'hbbda7e02),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba28dfb),
	.w1(32'h3b128f7d),
	.w2(32'hbcbb6973),
	.w3(32'h3c7c9a35),
	.w4(32'h3c827609),
	.w5(32'h3d0bee2b),
	.w6(32'hbcd5df23),
	.w7(32'hbc48f5fb),
	.w8(32'hbbad1d74),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3dc89),
	.w1(32'hba7f2d84),
	.w2(32'h3a27b065),
	.w3(32'hbafaaa1d),
	.w4(32'hbaa4fa93),
	.w5(32'h3a125b38),
	.w6(32'h3b0230c9),
	.w7(32'h3b8f2f07),
	.w8(32'h3b86fd84),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fae4df),
	.w1(32'hbb1bbd13),
	.w2(32'hbbdf2429),
	.w3(32'h39b697dc),
	.w4(32'h3c211a04),
	.w5(32'hbc3d6daf),
	.w6(32'h3bc838f8),
	.w7(32'h3b2ecedc),
	.w8(32'h3bf956a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc60654),
	.w1(32'hbc4b58b6),
	.w2(32'h3d48da1a),
	.w3(32'hbc43e581),
	.w4(32'h3c21907d),
	.w5(32'h3bf24fd3),
	.w6(32'h3c8ae06b),
	.w7(32'h3c3b2420),
	.w8(32'hbc431993),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e2bdd),
	.w1(32'h3c3c3066),
	.w2(32'hbc389434),
	.w3(32'h3c9eb9b9),
	.w4(32'h3c872f4c),
	.w5(32'h3c79421c),
	.w6(32'hba45a189),
	.w7(32'hbb794765),
	.w8(32'h3c13abcb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2a3e1),
	.w1(32'h3b77a8af),
	.w2(32'hbc4d484a),
	.w3(32'hbce54f7e),
	.w4(32'hbca499f5),
	.w5(32'h3ab34727),
	.w6(32'hbba133fa),
	.w7(32'hbbd8863d),
	.w8(32'h3afaddd0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc6a99),
	.w1(32'hbc407e15),
	.w2(32'hbc217440),
	.w3(32'h3b2ee09e),
	.w4(32'hbb3fd135),
	.w5(32'hbb4c5f26),
	.w6(32'hbbdedbf4),
	.w7(32'h3abc20a5),
	.w8(32'hbbb4f9f2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddef91),
	.w1(32'hbc08e7be),
	.w2(32'hbbb0918e),
	.w3(32'hbbae21d5),
	.w4(32'hbb4adc40),
	.w5(32'h3bb3e6e5),
	.w6(32'h3b85ec86),
	.w7(32'hbbb07c95),
	.w8(32'hbaae9deb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd210),
	.w1(32'hbc1b5784),
	.w2(32'hbb826ec5),
	.w3(32'hbb36a160),
	.w4(32'hbc97a035),
	.w5(32'hbc7946ed),
	.w6(32'hba72784e),
	.w7(32'hbc66c337),
	.w8(32'hbc9ca5e2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d8194),
	.w1(32'hbca46050),
	.w2(32'hbb9bad5f),
	.w3(32'hbbdd7fdc),
	.w4(32'hbcaf8ce6),
	.w5(32'h3b22ccb3),
	.w6(32'hbace5c82),
	.w7(32'hb9abca82),
	.w8(32'h3a4268cb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39a9d0),
	.w1(32'h3b91096b),
	.w2(32'h3c49df3a),
	.w3(32'hbc313a7f),
	.w4(32'hbcabe282),
	.w5(32'hbc0d9cb3),
	.w6(32'hbb435d5b),
	.w7(32'hbb800266),
	.w8(32'hbc77757d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523b61),
	.w1(32'h3b491b7f),
	.w2(32'h3b803584),
	.w3(32'h3b9fc5a2),
	.w4(32'hbb28e60a),
	.w5(32'h3baac1bf),
	.w6(32'h3aadde29),
	.w7(32'hbb2bddc4),
	.w8(32'hbaeaecc8),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe17159),
	.w1(32'hbb8333e3),
	.w2(32'hbc817d86),
	.w3(32'hbc043a1d),
	.w4(32'hbc41efed),
	.w5(32'h3b66d36a),
	.w6(32'hba9e709d),
	.w7(32'hbbe65b45),
	.w8(32'h3aa75705),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061012),
	.w1(32'hbc859077),
	.w2(32'hbbccef69),
	.w3(32'h3bf2c54a),
	.w4(32'hbc578c53),
	.w5(32'hbce0b65f),
	.w6(32'hbb91f123),
	.w7(32'hbbca2749),
	.w8(32'hbbaa463c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445b47),
	.w1(32'hba1a4215),
	.w2(32'hbc2cb423),
	.w3(32'hbc6c3c6c),
	.w4(32'h3c6e84b7),
	.w5(32'hbc8efc7e),
	.w6(32'hbbb1d8e0),
	.w7(32'hbaeaf30c),
	.w8(32'hbba60dfc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e8a43),
	.w1(32'hbbb3b27e),
	.w2(32'hbc2be9cc),
	.w3(32'hbc884090),
	.w4(32'hbba24925),
	.w5(32'hbc2a7fb9),
	.w6(32'hbb832ff1),
	.w7(32'hbb11fa70),
	.w8(32'h3c10866b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4c5d),
	.w1(32'hbb4c1e5d),
	.w2(32'hbb5411c8),
	.w3(32'hbb3be1f7),
	.w4(32'h3c06f64b),
	.w5(32'h3bfd9bf5),
	.w6(32'hb988671c),
	.w7(32'hbab9ec40),
	.w8(32'hbc0ff83b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc471922),
	.w1(32'hbb16c466),
	.w2(32'hbb1df7fa),
	.w3(32'hbb5098a2),
	.w4(32'h3b3a1efd),
	.w5(32'h3b8720ce),
	.w6(32'hbaa41524),
	.w7(32'hbb2675ea),
	.w8(32'h3b448a77),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2086af),
	.w1(32'h3b18fe9f),
	.w2(32'h3c81ad6d),
	.w3(32'hbc1429f4),
	.w4(32'hbc3a5ea3),
	.w5(32'h3b46e13d),
	.w6(32'h3c0d015d),
	.w7(32'h3bb487ec),
	.w8(32'h3ba6f301),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52049d),
	.w1(32'hbbf7b06c),
	.w2(32'hbc42810d),
	.w3(32'h3bc39a5b),
	.w4(32'h3be309fe),
	.w5(32'h3c04b9b0),
	.w6(32'hbc85ad97),
	.w7(32'hbc7ac088),
	.w8(32'hbc6b5c4d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67cabd),
	.w1(32'h3bf5f463),
	.w2(32'hbc8b287b),
	.w3(32'hbaa498b4),
	.w4(32'h3c38eb2b),
	.w5(32'h3cebf0a4),
	.w6(32'hbc505da9),
	.w7(32'hbbd0d7b6),
	.w8(32'hbbaa3248),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc944519),
	.w1(32'h3b992c0c),
	.w2(32'h395be25f),
	.w3(32'hbc8042be),
	.w4(32'h3b17fe61),
	.w5(32'hbbb6cdd9),
	.w6(32'h39884841),
	.w7(32'h3bb81e47),
	.w8(32'h3b6f0611),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17bf30),
	.w1(32'h3c8de4b4),
	.w2(32'h3ca843f1),
	.w3(32'hbb0f7c62),
	.w4(32'hbba068b0),
	.w5(32'hbba4023f),
	.w6(32'h3c2b7b70),
	.w7(32'h3c927c71),
	.w8(32'h3c80dfdc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2de808),
	.w1(32'h3a552e54),
	.w2(32'h3aae4c46),
	.w3(32'h3c69daa8),
	.w4(32'hbacf990a),
	.w5(32'hbb8afa30),
	.w6(32'h3bd54798),
	.w7(32'h3b89e855),
	.w8(32'h3b8254d1),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa3a4d),
	.w1(32'h399ae357),
	.w2(32'h39955608),
	.w3(32'h3b27e72a),
	.w4(32'h3a917b6c),
	.w5(32'h3b0b1326),
	.w6(32'h3bb6a665),
	.w7(32'h3bd953c2),
	.w8(32'h3b9298cb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107098),
	.w1(32'hbaeb9425),
	.w2(32'h3c80346a),
	.w3(32'hbb3308a9),
	.w4(32'hbc80cbfe),
	.w5(32'hbb8e1cee),
	.w6(32'h3c3eb778),
	.w7(32'h3c1d03ad),
	.w8(32'h3bcf200c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8844dc),
	.w1(32'hbbcb5445),
	.w2(32'h3b255abd),
	.w3(32'h3ca75045),
	.w4(32'hbc2c7952),
	.w5(32'hbc15585e),
	.w6(32'hbb988bef),
	.w7(32'hbc1f9252),
	.w8(32'hbc0b315d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1fb79),
	.w1(32'hbbc2cbec),
	.w2(32'hbc9e2ed9),
	.w3(32'hbc9cd28a),
	.w4(32'h3b107cfe),
	.w5(32'hbc42cdfc),
	.w6(32'hbc85f6ea),
	.w7(32'h3b91619a),
	.w8(32'hbc0fad13),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dce8c),
	.w1(32'h3abb19cb),
	.w2(32'hbbcbb5ab),
	.w3(32'hbb99d506),
	.w4(32'h3ab43fc4),
	.w5(32'h39b9f5ff),
	.w6(32'h3b04020a),
	.w7(32'h3b697bfc),
	.w8(32'hbac6deef),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fa94e),
	.w1(32'hbadfb001),
	.w2(32'hbb6e2b95),
	.w3(32'hbbebd62f),
	.w4(32'h3c16d39f),
	.w5(32'hbad815dd),
	.w6(32'hb97a9304),
	.w7(32'h3bdc4ddf),
	.w8(32'hb98a7774),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d3fa),
	.w1(32'hba421ed0),
	.w2(32'hbb908d28),
	.w3(32'hbbc16a20),
	.w4(32'hba6f9d3c),
	.w5(32'hba9ebbd0),
	.w6(32'h3b20a5b3),
	.w7(32'hbb80b557),
	.w8(32'h3a27d5ee),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc364282),
	.w1(32'hbc4ae1fb),
	.w2(32'hbc282230),
	.w3(32'hbc50e4a8),
	.w4(32'hbb46b5cf),
	.w5(32'hbb157adb),
	.w6(32'hbbec411f),
	.w7(32'h3be0461c),
	.w8(32'hbc2338b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e948),
	.w1(32'hbb9140ab),
	.w2(32'h3b1aee5c),
	.w3(32'hbb91a048),
	.w4(32'hbbe532ac),
	.w5(32'hbba59bb8),
	.w6(32'hbb44dc34),
	.w7(32'h3b3427a3),
	.w8(32'hbabfa8fe),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f49f90),
	.w1(32'hbbf2d8e4),
	.w2(32'hbc2445c2),
	.w3(32'hbbbde0ae),
	.w4(32'hbbeae715),
	.w5(32'hbbe651c2),
	.w6(32'h3909c604),
	.w7(32'hbaa377d1),
	.w8(32'hbbbb4223),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc484d95),
	.w1(32'h3b5cba19),
	.w2(32'h3b1b75a9),
	.w3(32'hbc3250a4),
	.w4(32'hbc851e23),
	.w5(32'hbcb23121),
	.w6(32'h3a8ae56d),
	.w7(32'h3aac89ec),
	.w8(32'h3a85c013),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1ec88),
	.w1(32'h3c5be289),
	.w2(32'h3b335276),
	.w3(32'h39620ebf),
	.w4(32'hbc010487),
	.w5(32'hbc996ac4),
	.w6(32'h3b8a1ddc),
	.w7(32'h3b344b04),
	.w8(32'h3aa5735c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f38096),
	.w1(32'h3b6094ff),
	.w2(32'h3a40f5c2),
	.w3(32'hbc2149fe),
	.w4(32'h3c20c89e),
	.w5(32'h3c26f871),
	.w6(32'hbc0956fc),
	.w7(32'h3b44fe8c),
	.w8(32'h3c0c2702),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124b3f),
	.w1(32'h3aa2f437),
	.w2(32'hbbf45872),
	.w3(32'h3c3045b9),
	.w4(32'h3b987b3e),
	.w5(32'hbbb62389),
	.w6(32'h3b71c995),
	.w7(32'hb96d6d5a),
	.w8(32'hbac264f7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb603ab),
	.w1(32'hbbaddbf6),
	.w2(32'hbbd0bf1f),
	.w3(32'hbca50388),
	.w4(32'hbc33e923),
	.w5(32'hbc18a6f8),
	.w6(32'hbc042bee),
	.w7(32'h3c5937a9),
	.w8(32'h3aef237b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ff88a),
	.w1(32'hbbc2e113),
	.w2(32'hbb328998),
	.w3(32'hbb0b68b6),
	.w4(32'hbb7ac382),
	.w5(32'hbaa6d43b),
	.w6(32'h3b071485),
	.w7(32'h3a165ee0),
	.w8(32'h39ff091f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5313d),
	.w1(32'h3c0acd7f),
	.w2(32'hbbe0652d),
	.w3(32'hba1e0398),
	.w4(32'h3b84b9a8),
	.w5(32'hbc6ba26e),
	.w6(32'h3ab07485),
	.w7(32'h39e4a6d7),
	.w8(32'h3a2f898b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd32f96),
	.w1(32'h3c435ad8),
	.w2(32'h3b87677e),
	.w3(32'hbc0c53fd),
	.w4(32'hbb8140d7),
	.w5(32'h3ca25a35),
	.w6(32'hbb286c70),
	.w7(32'hbc8e3596),
	.w8(32'h3a619494),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9853d6),
	.w1(32'hbb2299c2),
	.w2(32'hbcf61422),
	.w3(32'h3a98c2ce),
	.w4(32'h3b218ebd),
	.w5(32'h3c2f5a33),
	.w6(32'hbc253f92),
	.w7(32'hbc56e884),
	.w8(32'h3b531ab6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71ca71),
	.w1(32'h3bc52def),
	.w2(32'h3c0c942a),
	.w3(32'hbcc9631f),
	.w4(32'hbc37e01c),
	.w5(32'h3b92a22c),
	.w6(32'h3b1967fa),
	.w7(32'hbbdb8959),
	.w8(32'hbc4f9994),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc902f17),
	.w1(32'h3bd84e72),
	.w2(32'h3bd99f1d),
	.w3(32'hbc700e4e),
	.w4(32'h3aab34b6),
	.w5(32'h3b6ac026),
	.w6(32'h3b98b6d7),
	.w7(32'h3c2b1251),
	.w8(32'h3adc2097),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5c46),
	.w1(32'hbbbbda54),
	.w2(32'hbbcc71e4),
	.w3(32'hbba726b7),
	.w4(32'hbbef8c1d),
	.w5(32'hbc0db096),
	.w6(32'hbb1ae78c),
	.w7(32'hbbd3ff65),
	.w8(32'hbb414650),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc287a21),
	.w1(32'hbbfedd88),
	.w2(32'h3a54132a),
	.w3(32'hbc047455),
	.w4(32'hbc81e184),
	.w5(32'hbb1fef96),
	.w6(32'h3b327eee),
	.w7(32'hbb8d583e),
	.w8(32'hbc7dd06e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b82f63),
	.w1(32'hbba03bf2),
	.w2(32'hbaf44bf8),
	.w3(32'h3bbf2f74),
	.w4(32'hbc8736fd),
	.w5(32'hbbe1a619),
	.w6(32'hbc093f81),
	.w7(32'hbbeaf950),
	.w8(32'hbc0a3b38),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99d0be),
	.w1(32'hbb9a6240),
	.w2(32'h3b2f0587),
	.w3(32'hba2e6e33),
	.w4(32'hba5b295f),
	.w5(32'h3a96f9c0),
	.w6(32'h3b05feae),
	.w7(32'h3bd5ff79),
	.w8(32'h3c641655),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23e5c2),
	.w1(32'h3ad68770),
	.w2(32'hbbb8f09d),
	.w3(32'hbc485fae),
	.w4(32'h3ba628cf),
	.w5(32'hbb418941),
	.w6(32'h3ba2874a),
	.w7(32'h3c505c33),
	.w8(32'h3bf23448),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb79c9),
	.w1(32'hbbf96120),
	.w2(32'hbc63f3cc),
	.w3(32'hbb481f52),
	.w4(32'hbbfdda9e),
	.w5(32'hbc2ae2d5),
	.w6(32'hbbfe30db),
	.w7(32'hbc1baeb7),
	.w8(32'hbc1c56a4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a5e94),
	.w1(32'h3a74a6c4),
	.w2(32'h3a17e1db),
	.w3(32'hbc797536),
	.w4(32'hba97a3cd),
	.w5(32'hbb0d0a00),
	.w6(32'h3bdf2550),
	.w7(32'h3b87d446),
	.w8(32'h3b4a04f5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba04325),
	.w1(32'hbb186f17),
	.w2(32'hbb1cddbc),
	.w3(32'hbb046f35),
	.w4(32'hbc2d7af2),
	.w5(32'h3b3c1954),
	.w6(32'hbb68b00e),
	.w7(32'hbbba443c),
	.w8(32'hbbe94c1f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d106b),
	.w1(32'hbcb6aa31),
	.w2(32'hbd02e13b),
	.w3(32'hbb65c7ab),
	.w4(32'hbc05af5d),
	.w5(32'hbbb021b2),
	.w6(32'hbc56d076),
	.w7(32'hb9237ed5),
	.w8(32'h3c17ee2c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd93c04),
	.w1(32'hbc682ef8),
	.w2(32'hbc83277c),
	.w3(32'hbc6a88bb),
	.w4(32'hbc831b3c),
	.w5(32'hbc216c37),
	.w6(32'hbb9e9321),
	.w7(32'hbbe90c5e),
	.w8(32'hb9973221),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c7d4),
	.w1(32'h3d07e7e1),
	.w2(32'hbbfcea41),
	.w3(32'hbbc7bd4a),
	.w4(32'h3ce7921b),
	.w5(32'h3d5c528d),
	.w6(32'hbc556320),
	.w7(32'hbb06d976),
	.w8(32'h3c00e7d9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3b411),
	.w1(32'hbb3835c1),
	.w2(32'h3b6b14ae),
	.w3(32'hbc7d844c),
	.w4(32'hbc1058ab),
	.w5(32'hbc9030b4),
	.w6(32'hbc04bd5c),
	.w7(32'h3b8f097b),
	.w8(32'h3bb77653),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b65ebe),
	.w1(32'hbb82243e),
	.w2(32'h3b848c92),
	.w3(32'h3b8f7799),
	.w4(32'hbb83f34b),
	.w5(32'hbb8488c1),
	.w6(32'h39f8b2d0),
	.w7(32'h3b672419),
	.w8(32'hbc127eb1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0aa33),
	.w1(32'hbc09a59f),
	.w2(32'hbc441aca),
	.w3(32'hbbb35cb7),
	.w4(32'h3a141193),
	.w5(32'hbac14048),
	.w6(32'h398ce9d0),
	.w7(32'hbb0c1be3),
	.w8(32'h3b8a6b43),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89a681),
	.w1(32'hbbcadb05),
	.w2(32'h3bf649d1),
	.w3(32'h3b625a8d),
	.w4(32'hbc2d34ca),
	.w5(32'hbc05da74),
	.w6(32'h3cb588f6),
	.w7(32'h3bbb4c28),
	.w8(32'h3c172d30),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e638e),
	.w1(32'hbbd00351),
	.w2(32'h3c0ff94f),
	.w3(32'h3c08ba80),
	.w4(32'hbbe9b5bc),
	.w5(32'hbbe63bd2),
	.w6(32'hbb15ff5b),
	.w7(32'h3bc667f3),
	.w8(32'hba04ef28),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3dc6),
	.w1(32'hb9e3f059),
	.w2(32'h3bc25739),
	.w3(32'h392faaf2),
	.w4(32'hb95dc210),
	.w5(32'h3ba89890),
	.w6(32'h3a7c30bc),
	.w7(32'h3adb1960),
	.w8(32'h3b563eb5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68d274),
	.w1(32'h3b962188),
	.w2(32'h3c2dc91e),
	.w3(32'hbb6fab02),
	.w4(32'hba8442ea),
	.w5(32'h3b2dbff1),
	.w6(32'hbabbd525),
	.w7(32'h3b378964),
	.w8(32'h3c254ae5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77019),
	.w1(32'h3a4cb3a2),
	.w2(32'h3b8584e6),
	.w3(32'h3bd427d1),
	.w4(32'hbae7ebc3),
	.w5(32'hbabe9d66),
	.w6(32'hbb3fad91),
	.w7(32'h3a13644f),
	.w8(32'hbb182b91),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fcc16),
	.w1(32'h3a39e1b6),
	.w2(32'hbc3ab6cd),
	.w3(32'hbc4f00fa),
	.w4(32'h3b54beb4),
	.w5(32'hbbb2a42b),
	.w6(32'hbbd640a0),
	.w7(32'hba8a5d16),
	.w8(32'hbb7f5fc7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b4de),
	.w1(32'h3b48a0b5),
	.w2(32'hbc4647ca),
	.w3(32'hbb8df591),
	.w4(32'h3c22c007),
	.w5(32'h3b6362f4),
	.w6(32'hbc38d35e),
	.w7(32'h3b70399b),
	.w8(32'h3b92eaad),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4170b9),
	.w1(32'hbbcdbd89),
	.w2(32'hbcd0074d),
	.w3(32'hbc2e94c0),
	.w4(32'h3cdeeacd),
	.w5(32'hbc02499d),
	.w6(32'hbc8255e9),
	.w7(32'hbbc03a24),
	.w8(32'h3ba07d19),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd16335),
	.w1(32'hbb9fe312),
	.w2(32'hbc7bb1c3),
	.w3(32'hbcb94f1d),
	.w4(32'h3b547c47),
	.w5(32'h3bfebc80),
	.w6(32'hbc3bd9e3),
	.w7(32'hbbf178b0),
	.w8(32'hbb722666),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9300bc),
	.w1(32'h3cc86685),
	.w2(32'hbc9826fa),
	.w3(32'hbc20fe75),
	.w4(32'h3cdadef8),
	.w5(32'h3d2c42c0),
	.w6(32'hbccc96f1),
	.w7(32'hbb699e11),
	.w8(32'h3a22c387),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce86592),
	.w1(32'hba7fd6cb),
	.w2(32'hbc07df3d),
	.w3(32'hbc74384d),
	.w4(32'hbb94a933),
	.w5(32'hbbbf5d98),
	.w6(32'hbbf7b20f),
	.w7(32'h39b30313),
	.w8(32'hbc2c0dcd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc791d95),
	.w1(32'h3b939bce),
	.w2(32'hbc9ce7a6),
	.w3(32'hbc2a7e52),
	.w4(32'h3baa4812),
	.w5(32'hbcbe25f2),
	.w6(32'hbc9f997c),
	.w7(32'h3b13e156),
	.w8(32'hbc2fe2fe),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc847f3b),
	.w1(32'hbc27e214),
	.w2(32'hbcde434d),
	.w3(32'hbb9a9fbf),
	.w4(32'h3c526df2),
	.w5(32'h3cba36f2),
	.w6(32'hbcb17f59),
	.w7(32'hbab8d626),
	.w8(32'h3ba53cdb),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcc48b),
	.w1(32'hbc449c74),
	.w2(32'hbc0503bd),
	.w3(32'hbc94bd77),
	.w4(32'h3b80c6ee),
	.w5(32'hbb2f2eaf),
	.w6(32'hbc6dd924),
	.w7(32'hbb600611),
	.w8(32'hbb8234d2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16b57d),
	.w1(32'hbaccf6ce),
	.w2(32'hbb114ba0),
	.w3(32'hb9da19f3),
	.w4(32'hba89fc6d),
	.w5(32'h3a39da87),
	.w6(32'hb9ced8e7),
	.w7(32'hbaf74434),
	.w8(32'hbad997a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f386cb),
	.w1(32'hbb8981ca),
	.w2(32'hbb2c7aa9),
	.w3(32'hb9540249),
	.w4(32'hbb6fe43d),
	.w5(32'h3901e1ee),
	.w6(32'hbba36067),
	.w7(32'hbbba8767),
	.w8(32'hbb9ffe73),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1421a5),
	.w1(32'hbb13a455),
	.w2(32'h393f3be6),
	.w3(32'hbb245b80),
	.w4(32'hba8227b0),
	.w5(32'h3af1ae98),
	.w6(32'h3b64874c),
	.w7(32'hba60785d),
	.w8(32'hbb1ec9c6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9285955),
	.w1(32'hba2f3e3c),
	.w2(32'hbba88ed4),
	.w3(32'h3af04d25),
	.w4(32'hbc10d07b),
	.w5(32'hbc717eb4),
	.w6(32'h3c8905a5),
	.w7(32'hba3e979a),
	.w8(32'h3c0f9a3c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5c572),
	.w1(32'hbb7672b9),
	.w2(32'h3a005ea2),
	.w3(32'hbb250fc0),
	.w4(32'hbb98292e),
	.w5(32'hbc602ad5),
	.w6(32'h3c02403f),
	.w7(32'h3bfb6948),
	.w8(32'h3b9d5dcb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15eb34),
	.w1(32'hbc077857),
	.w2(32'hbc65f94b),
	.w3(32'hbad62164),
	.w4(32'h3c7b61e7),
	.w5(32'h3cdf1d0e),
	.w6(32'hbc5f3db3),
	.w7(32'hbc17e942),
	.w8(32'hbc2efdfb),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65b5be),
	.w1(32'h3ae5891d),
	.w2(32'hba5e5186),
	.w3(32'hbb8a3512),
	.w4(32'hb83baa90),
	.w5(32'hbb3c0593),
	.w6(32'hbbebd14d),
	.w7(32'hbb32211c),
	.w8(32'hbbf65a34),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda30ea),
	.w1(32'hbb27bf6e),
	.w2(32'hbb1c2ada),
	.w3(32'hbb6d2d59),
	.w4(32'hbabaf7a6),
	.w5(32'hbb635dda),
	.w6(32'hba92ab22),
	.w7(32'hba835b17),
	.w8(32'hbb5c915d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d6cb4),
	.w1(32'h3c800101),
	.w2(32'h3ab0e50a),
	.w3(32'h38e491eb),
	.w4(32'hb99c4f4e),
	.w5(32'hbb59ef5a),
	.w6(32'h3b6e4cd3),
	.w7(32'hbbddfbcc),
	.w8(32'h3c198205),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4276b7),
	.w1(32'h3b01f5f7),
	.w2(32'hba53f185),
	.w3(32'hbb6c7173),
	.w4(32'h3b188135),
	.w5(32'h3ab38801),
	.w6(32'h3a1074b0),
	.w7(32'hbb01f202),
	.w8(32'hba77a88a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7dccb9),
	.w1(32'hbc4fa4d9),
	.w2(32'h3b87e249),
	.w3(32'hbbed91fa),
	.w4(32'hbc6f79fc),
	.w5(32'hbc8801fe),
	.w6(32'h3c0729d3),
	.w7(32'h3c1a379f),
	.w8(32'hb96430a1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95d6cc),
	.w1(32'h3aa52882),
	.w2(32'h3beea9b3),
	.w3(32'h3c5f56a1),
	.w4(32'hbb682433),
	.w5(32'h3a22ad4a),
	.w6(32'h3c41b060),
	.w7(32'hbb0fd7ea),
	.w8(32'h3b25e047),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a93c5),
	.w1(32'hba4867f7),
	.w2(32'h3c2c6a0e),
	.w3(32'h3c8b8270),
	.w4(32'hbc1c439b),
	.w5(32'h3b74a636),
	.w6(32'h3c3a0726),
	.w7(32'h3c0e8b78),
	.w8(32'h3b8218c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57e98b),
	.w1(32'hbc89c583),
	.w2(32'hbcb5381e),
	.w3(32'h3c5b47d8),
	.w4(32'h3c83c7b0),
	.w5(32'hbca36b67),
	.w6(32'hbaecdd4d),
	.w7(32'hba9cbb47),
	.w8(32'hbb415875),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b913c56),
	.w1(32'h3c523097),
	.w2(32'hbbb57eb2),
	.w3(32'hbc6521df),
	.w4(32'h3ca7d69e),
	.w5(32'h3d1efd67),
	.w6(32'hbbb86d2a),
	.w7(32'h3a77909e),
	.w8(32'hbb3fea4b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5be96),
	.w1(32'hbbc813e3),
	.w2(32'h3c5939e0),
	.w3(32'hbb318607),
	.w4(32'hbafdf965),
	.w5(32'hbc5a2169),
	.w6(32'h3bc91495),
	.w7(32'hba5bf601),
	.w8(32'h3bdcdd5f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba411a55),
	.w1(32'hbba8000f),
	.w2(32'hbcb81fbd),
	.w3(32'h3a9295df),
	.w4(32'h3ca9c0b4),
	.w5(32'h3d28281b),
	.w6(32'hbc876b55),
	.w7(32'hbc5f6cb6),
	.w8(32'hbc0f863e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d1010),
	.w1(32'hbc24e4ca),
	.w2(32'h3aac68f4),
	.w3(32'hbc499909),
	.w4(32'hbb341528),
	.w5(32'hbb5a7bcc),
	.w6(32'h3c12d35b),
	.w7(32'h3cb98de8),
	.w8(32'h3c58f07b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4ef6b),
	.w1(32'h3c4e6215),
	.w2(32'h3c1285c5),
	.w3(32'hbb7ea586),
	.w4(32'h39add9b8),
	.w5(32'hbaa28090),
	.w6(32'h3bf2a9fd),
	.w7(32'h3b9cf0f8),
	.w8(32'h3c8057d3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f852e),
	.w1(32'hbc146f8b),
	.w2(32'hbb849f1c),
	.w3(32'hb880a24a),
	.w4(32'hbc536ef1),
	.w5(32'hbc0cd10d),
	.w6(32'hb9bd8e10),
	.w7(32'hba3fc699),
	.w8(32'h3a366d8a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dde07),
	.w1(32'hbb4ccd9f),
	.w2(32'h3c0cb65b),
	.w3(32'hbbce6680),
	.w4(32'hbb9aac6b),
	.w5(32'hbabce395),
	.w6(32'hb8c44787),
	.w7(32'hbb4de2db),
	.w8(32'h3af1d901),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf189fa),
	.w1(32'h3b9f2205),
	.w2(32'hbc2d3f44),
	.w3(32'hbb0b278d),
	.w4(32'h3c452d57),
	.w5(32'h3c90dc5c),
	.w6(32'hbbfd98e9),
	.w7(32'hbaeedadb),
	.w8(32'hbb1c0f64),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565b2b),
	.w1(32'h3b4d0c69),
	.w2(32'hbc2237c2),
	.w3(32'h3a7d103d),
	.w4(32'h3aa3d0a4),
	.w5(32'hbc1c8e67),
	.w6(32'h3a0c163c),
	.w7(32'h3b103701),
	.w8(32'h3c80b8f0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67b0d0),
	.w1(32'hbacc9ed8),
	.w2(32'hb9d56ad0),
	.w3(32'h3b8028bb),
	.w4(32'h3aa1c8a2),
	.w5(32'hbaf79293),
	.w6(32'h3b7da7c4),
	.w7(32'h3b0b31ba),
	.w8(32'h3af0ff5c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeffc1d),
	.w1(32'hbc9b678e),
	.w2(32'hbcb0dbc1),
	.w3(32'hbb8d7561),
	.w4(32'h3ce7d257),
	.w5(32'h3c2d3809),
	.w6(32'hbc629d3a),
	.w7(32'h3a066fe1),
	.w8(32'hbbc40c72),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf67a16),
	.w1(32'hb995e157),
	.w2(32'hbbcb667a),
	.w3(32'hbca6ec65),
	.w4(32'hbacddfc0),
	.w5(32'hbae224db),
	.w6(32'hbbb7232a),
	.w7(32'h3b0e0f4a),
	.w8(32'hbaca5985),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb328612),
	.w1(32'h3c11c9f9),
	.w2(32'h3b6bd35b),
	.w3(32'h3aac26c6),
	.w4(32'h3b607051),
	.w5(32'h3bdc7ca6),
	.w6(32'h398cd63f),
	.w7(32'hbb88c413),
	.w8(32'hb99c8681),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff4e8c),
	.w1(32'hbba22e7e),
	.w2(32'hbc8bd071),
	.w3(32'h3b8be95d),
	.w4(32'hbc0b2971),
	.w5(32'h3bba7f6a),
	.w6(32'h3c12705a),
	.w7(32'h3aab5d7b),
	.w8(32'h3c7b7fe4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257da0),
	.w1(32'hbb61c41c),
	.w2(32'hbbdfd806),
	.w3(32'h3bcb3997),
	.w4(32'hbba0b39e),
	.w5(32'hbc16d596),
	.w6(32'h3ab314b3),
	.w7(32'hb9de82af),
	.w8(32'hbace2d39),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f643),
	.w1(32'hbb501582),
	.w2(32'hbb5ab40a),
	.w3(32'hbbf6bfd0),
	.w4(32'hbb16ea6e),
	.w5(32'hbb8cea94),
	.w6(32'h38af17ef),
	.w7(32'hbabf88ef),
	.w8(32'hba91913a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddb2b8),
	.w1(32'h3aa1194b),
	.w2(32'h3b3a97c2),
	.w3(32'hbb89e29e),
	.w4(32'h3c2f6954),
	.w5(32'h3b9cdd75),
	.w6(32'hb92dd64a),
	.w7(32'h3aa9ccb3),
	.w8(32'h3b78bdb4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824bbf),
	.w1(32'hbbe1bc00),
	.w2(32'hbc1d875a),
	.w3(32'hba71aafa),
	.w4(32'h3a993833),
	.w5(32'h3aac9eca),
	.w6(32'hbc103eb2),
	.w7(32'h3b228a71),
	.w8(32'hbb7a7992),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059f31),
	.w1(32'h3ca4e2cf),
	.w2(32'hbadc2053),
	.w3(32'hbc0e3c5b),
	.w4(32'h3c122421),
	.w5(32'h3d3048f2),
	.w6(32'hbc316880),
	.w7(32'hbcae4510),
	.w8(32'hb9a2a7ab),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd445b),
	.w1(32'hbb0229a5),
	.w2(32'h3b59db52),
	.w3(32'h3bb6775b),
	.w4(32'hbbda6d21),
	.w5(32'h3b462029),
	.w6(32'hbb2010a0),
	.w7(32'hbbb064cc),
	.w8(32'hbacbe036),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabad7d4),
	.w1(32'h3c943c1d),
	.w2(32'hbc94a89a),
	.w3(32'h3a508b01),
	.w4(32'h3c9891ce),
	.w5(32'h3ce70e40),
	.w6(32'hbca3b270),
	.w7(32'hbc5857d8),
	.w8(32'h3b54ac6e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1dd6c),
	.w1(32'hbb92307c),
	.w2(32'hbc096899),
	.w3(32'hbc5ebeee),
	.w4(32'hb9918ec5),
	.w5(32'h3c28545a),
	.w6(32'hbb90b214),
	.w7(32'hbbc13705),
	.w8(32'hbaf761e1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b59b1),
	.w1(32'hbb1ac523),
	.w2(32'hbb2b7f3a),
	.w3(32'hbc2199c9),
	.w4(32'hbb860f37),
	.w5(32'hbb180d56),
	.w6(32'hb9fe5e75),
	.w7(32'hbb34cdfb),
	.w8(32'hba578897),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7681dc),
	.w1(32'hbbab7d21),
	.w2(32'h3b06a3f7),
	.w3(32'hbafb62db),
	.w4(32'hbad4c534),
	.w5(32'hbb24ef1c),
	.w6(32'hba3c901b),
	.w7(32'h3b754620),
	.w8(32'h3ba50b3d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287e23),
	.w1(32'h3d4a47c3),
	.w2(32'h3ce1aed7),
	.w3(32'h3bd25bc6),
	.w4(32'hbc655f65),
	.w5(32'h3d4b79c4),
	.w6(32'h3bdd9ee8),
	.w7(32'hbbde91fc),
	.w8(32'h3c5a7fa1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e467c),
	.w1(32'h3c16d954),
	.w2(32'h3c2842b5),
	.w3(32'h3d159268),
	.w4(32'hbc14799a),
	.w5(32'hbc928e02),
	.w6(32'h3aa9bd4d),
	.w7(32'h3aede4b8),
	.w8(32'hba44df90),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4f848),
	.w1(32'hbac8aafb),
	.w2(32'hba47c09c),
	.w3(32'h3af23e94),
	.w4(32'h3a621585),
	.w5(32'h391b1c43),
	.w6(32'hbabb6e1a),
	.w7(32'h3ae28173),
	.w8(32'hba65d073),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e35ec),
	.w1(32'hbc8cebb0),
	.w2(32'hbc1bb620),
	.w3(32'hbb711fa0),
	.w4(32'hbca85cf0),
	.w5(32'hbc366c9f),
	.w6(32'hbc995324),
	.w7(32'hbc55cac2),
	.w8(32'hbc4a8257),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule