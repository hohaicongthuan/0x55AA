module layer_8_featuremap_199(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b845dcb),
	.w1(32'h3a8a545c),
	.w2(32'h3c7d66d4),
	.w3(32'hbaae73cf),
	.w4(32'hba4f8d21),
	.w5(32'h3c92e3b6),
	.w6(32'h39a61d48),
	.w7(32'h3b795e8f),
	.w8(32'hbab466d2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99201a0),
	.w1(32'h3ab3b82a),
	.w2(32'h38f5b31f),
	.w3(32'h3b70c2b8),
	.w4(32'hbb54b487),
	.w5(32'hb9bc06b4),
	.w6(32'hba5d130f),
	.w7(32'h3a0b723f),
	.w8(32'hbb0a7946),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c7e6d),
	.w1(32'h3b457757),
	.w2(32'hbc2d1122),
	.w3(32'h3b21811a),
	.w4(32'h3c29b5cd),
	.w5(32'hba8713d7),
	.w6(32'h3bcf76cf),
	.w7(32'hbb8f0ff7),
	.w8(32'hbb9280d5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcec6db),
	.w1(32'h3b9749d3),
	.w2(32'h3af173d7),
	.w3(32'hbbb97cb9),
	.w4(32'hbaf39db5),
	.w5(32'hbc070fb6),
	.w6(32'h3c4a64d5),
	.w7(32'h3bb73c75),
	.w8(32'h3b1148f8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb02e5a),
	.w1(32'hbbc8cfea),
	.w2(32'hbb513b64),
	.w3(32'hba93c443),
	.w4(32'hbb17aa8c),
	.w5(32'hbb2b1ec3),
	.w6(32'hba14ee06),
	.w7(32'h3bbb9035),
	.w8(32'h38bcac56),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98f7aa),
	.w1(32'h3baefc73),
	.w2(32'h3ab31bea),
	.w3(32'h3a0f4d78),
	.w4(32'hba9dc7f8),
	.w5(32'hbc9e1b20),
	.w6(32'h3be8830f),
	.w7(32'h3c6f835a),
	.w8(32'hbbea8a3f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d907a),
	.w1(32'h3af0f5af),
	.w2(32'h3a0bb425),
	.w3(32'hbbe2d65f),
	.w4(32'hbab92fc7),
	.w5(32'hbb596d1d),
	.w6(32'hbb9690be),
	.w7(32'hbb42e2f2),
	.w8(32'hbb78adaf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef8e9),
	.w1(32'hbbb2d16b),
	.w2(32'h3b12ae49),
	.w3(32'hbb6e74b4),
	.w4(32'hbbefa44d),
	.w5(32'hbad20bfc),
	.w6(32'h3ba545f0),
	.w7(32'h3bfd3dfc),
	.w8(32'hbbc3108b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b885aef),
	.w1(32'h3b59e7ab),
	.w2(32'h3b773ffd),
	.w3(32'hbc4763b1),
	.w4(32'h3b69cd3b),
	.w5(32'h3b99a218),
	.w6(32'hbc17c480),
	.w7(32'hbb45a275),
	.w8(32'hbc0c698b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9bfff),
	.w1(32'h3b85511c),
	.w2(32'hbc022419),
	.w3(32'h3b1a832f),
	.w4(32'h3b9c6091),
	.w5(32'h3c6c4ae2),
	.w6(32'hbbcbdfad),
	.w7(32'hb8285224),
	.w8(32'h3b6adf88),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7000bd),
	.w1(32'h3b83feac),
	.w2(32'hbbdd7f68),
	.w3(32'h3bed8e6d),
	.w4(32'h3b4a6a4c),
	.w5(32'hbb971ab9),
	.w6(32'hbc5e3f9d),
	.w7(32'hbc4afd04),
	.w8(32'hbc29f07d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985c97),
	.w1(32'h3baa624a),
	.w2(32'h3c18450c),
	.w3(32'hbac44f66),
	.w4(32'h3b7a4ca8),
	.w5(32'h3b897d2a),
	.w6(32'h38bafdca),
	.w7(32'h3bc42ffc),
	.w8(32'hbb1f8a1a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072a0a),
	.w1(32'hbc043a68),
	.w2(32'hbc433b39),
	.w3(32'h3a875225),
	.w4(32'hbae7409b),
	.w5(32'h3b23ad8f),
	.w6(32'hbb865927),
	.w7(32'hbc0fe50f),
	.w8(32'hbae67ace),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1278c0),
	.w1(32'h3d1b4fc3),
	.w2(32'h3d22e141),
	.w3(32'hbaabd7ef),
	.w4(32'h3cbf06e9),
	.w5(32'h3d0190c4),
	.w6(32'h3d03ac1e),
	.w7(32'h3d2434be),
	.w8(32'h3cea6604),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff72c8),
	.w1(32'h3a75e2f5),
	.w2(32'hbb221874),
	.w3(32'h3cb38158),
	.w4(32'h3b3d4f6f),
	.w5(32'hbae50d8f),
	.w6(32'hbba6573e),
	.w7(32'hbc04075a),
	.w8(32'hbbb61e12),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ade27),
	.w1(32'h3b73c27b),
	.w2(32'h3c5e30e0),
	.w3(32'hbb382db7),
	.w4(32'hbaff3be5),
	.w5(32'h3bd7b370),
	.w6(32'hbc0def4e),
	.w7(32'hbbb67481),
	.w8(32'hbc2b52fb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba404bed),
	.w1(32'hbc496d6e),
	.w2(32'hba6fe9cb),
	.w3(32'hbb446ab9),
	.w4(32'hbc9a055a),
	.w5(32'h3b777b5d),
	.w6(32'hbbb895ba),
	.w7(32'hbbd4b869),
	.w8(32'hbba29207),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45c58a),
	.w1(32'hba8c297c),
	.w2(32'hbc18df29),
	.w3(32'h3aac22f5),
	.w4(32'hbb2c3d51),
	.w5(32'hb794f44d),
	.w6(32'hbc09d85d),
	.w7(32'hbc5ceaca),
	.w8(32'hbae25cae),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96bfec),
	.w1(32'h3a6ff04b),
	.w2(32'hbabed66f),
	.w3(32'h3abea8fc),
	.w4(32'hbba0833d),
	.w5(32'h3ba5be24),
	.w6(32'hbad26397),
	.w7(32'h3ac1fe73),
	.w8(32'h39bb2dc4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c78d),
	.w1(32'h3ba84a7d),
	.w2(32'h3ad57082),
	.w3(32'h3b220fb7),
	.w4(32'h3bb341fb),
	.w5(32'h3b771418),
	.w6(32'hbb2ccd26),
	.w7(32'hbbd4396b),
	.w8(32'hbb25068a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9b6b7),
	.w1(32'h39dd31ea),
	.w2(32'h3c2cd0fc),
	.w3(32'hba0a723f),
	.w4(32'hbb28f790),
	.w5(32'h3c01bb35),
	.w6(32'h3b449f93),
	.w7(32'h3c67d2dc),
	.w8(32'h3adb1e3c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29ea22),
	.w1(32'hbc1f1d62),
	.w2(32'hbd020a6c),
	.w3(32'hba459ac6),
	.w4(32'hbc3727f6),
	.w5(32'hbca8c3a5),
	.w6(32'hbb0483c4),
	.w7(32'hbc15d378),
	.w8(32'hbc23a1d7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85cdd5),
	.w1(32'hbc79f715),
	.w2(32'hbc2de3fa),
	.w3(32'h3b84048b),
	.w4(32'hbb7f854e),
	.w5(32'h3c26074a),
	.w6(32'hbc6000dd),
	.w7(32'hbc96144a),
	.w8(32'hbc141e10),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8b8b1),
	.w1(32'hbb94a10d),
	.w2(32'hbcea8a00),
	.w3(32'h3c402255),
	.w4(32'hbc8d8fd7),
	.w5(32'hbc8ff58a),
	.w6(32'h3b4eefd6),
	.w7(32'hbc4eb40a),
	.w8(32'hbc288387),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54f104),
	.w1(32'hbc1d184b),
	.w2(32'hbc0874a6),
	.w3(32'hb9b5aa48),
	.w4(32'hbc23724e),
	.w5(32'hbbd44eb3),
	.w6(32'h39be6b7d),
	.w7(32'hbbc485e9),
	.w8(32'hbb7c9ca6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3f14c),
	.w1(32'hbc06c7d8),
	.w2(32'hbc0691a0),
	.w3(32'h3c1595b7),
	.w4(32'hbbc48d7f),
	.w5(32'h3c0f5a9d),
	.w6(32'hba63b58d),
	.w7(32'h3ad3303b),
	.w8(32'hbbe264ff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87e3cb),
	.w1(32'h3b78e362),
	.w2(32'h3a1b97f1),
	.w3(32'h3a272bcd),
	.w4(32'hbb6f4fcf),
	.w5(32'hbc515b36),
	.w6(32'h3b9b373c),
	.w7(32'h3c90131e),
	.w8(32'hbb6efc13),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6be40),
	.w1(32'h3a9c18cd),
	.w2(32'hbc3e081a),
	.w3(32'hbbbbd70c),
	.w4(32'h3b10420d),
	.w5(32'hbb8e2e27),
	.w6(32'hbbe8ae99),
	.w7(32'hbc462a2b),
	.w8(32'hbbe22d42),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c30032),
	.w1(32'hbb88a54e),
	.w2(32'h3ba236a3),
	.w3(32'hbb7ebbe0),
	.w4(32'h3a6f9a1f),
	.w5(32'h3c09cdc7),
	.w6(32'hbc5d04fb),
	.w7(32'hbba40fbe),
	.w8(32'hbc161b7e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb3c34),
	.w1(32'h3acd8d6c),
	.w2(32'hbb46dbe3),
	.w3(32'h3a16e97f),
	.w4(32'hbaa1d414),
	.w5(32'h3b27f8e4),
	.w6(32'h3b359d88),
	.w7(32'h3b2cd984),
	.w8(32'hbb86e637),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff8f64),
	.w1(32'hbaec5aeb),
	.w2(32'hbbaa0aa1),
	.w3(32'h3bca2980),
	.w4(32'hbac63127),
	.w5(32'hbb44fd50),
	.w6(32'hbbd6859d),
	.w7(32'hbc0aabe5),
	.w8(32'hbc31aab9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1169e3),
	.w1(32'h3bb02125),
	.w2(32'hbad5c619),
	.w3(32'h3bebcf23),
	.w4(32'h3b5da018),
	.w5(32'h3bf4d661),
	.w6(32'hbb9ccbd6),
	.w7(32'h3a0e298d),
	.w8(32'hbc1efa1d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aade4c4),
	.w1(32'h3b737793),
	.w2(32'hbc8510ad),
	.w3(32'h3c05527a),
	.w4(32'h3b9f268e),
	.w5(32'hbb348b1a),
	.w6(32'hbbf8c5dd),
	.w7(32'hbb118daf),
	.w8(32'h3b10a344),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb295549),
	.w1(32'hbb8d40c3),
	.w2(32'h3c8b4efc),
	.w3(32'h3a802aed),
	.w4(32'h3ac676d1),
	.w5(32'h3c52c46b),
	.w6(32'hbc07c373),
	.w7(32'hbb05b42f),
	.w8(32'hbc00c065),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfded7f),
	.w1(32'h3c916890),
	.w2(32'h3c338dcb),
	.w3(32'h3c14bf5c),
	.w4(32'h3c555764),
	.w5(32'h3c4a7c7c),
	.w6(32'h3be3d28d),
	.w7(32'h3b2ccbf2),
	.w8(32'hbb4cad68),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e265b),
	.w1(32'hbcacde37),
	.w2(32'hbd5300b3),
	.w3(32'h3c31be52),
	.w4(32'hbcbe20b7),
	.w5(32'hbd3b2bbd),
	.w6(32'hbb884d83),
	.w7(32'hbc67c687),
	.w8(32'hbc31d834),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce25209),
	.w1(32'hbb2afb41),
	.w2(32'hbb6f9e98),
	.w3(32'hbd1a5582),
	.w4(32'hbaed499a),
	.w5(32'hbb1fa110),
	.w6(32'hba10d483),
	.w7(32'hbb37837d),
	.w8(32'hbb4bc3f8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03e4c),
	.w1(32'hbb4fb14b),
	.w2(32'hba80d58f),
	.w3(32'hbb831267),
	.w4(32'h3b680cd3),
	.w5(32'h3b93f9a1),
	.w6(32'hbbb9134f),
	.w7(32'hbbbeab60),
	.w8(32'hbba2b9c0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba15698),
	.w1(32'h3cd60b8a),
	.w2(32'h3d0b73be),
	.w3(32'h3b500451),
	.w4(32'h3c4a119f),
	.w5(32'h3d01c131),
	.w6(32'h3c9aa2c9),
	.w7(32'h3c9c834c),
	.w8(32'h3cb9b4aa),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf03f6c),
	.w1(32'hbd0e2f46),
	.w2(32'hbd8f3072),
	.w3(32'h3cb18cb6),
	.w4(32'hbce01d09),
	.w5(32'hbd4d1717),
	.w6(32'hbc86ddc7),
	.w7(32'hbd1d615c),
	.w8(32'hbcd819fd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2cccc7),
	.w1(32'h3bb56bbf),
	.w2(32'h3b6af133),
	.w3(32'hbcdffc16),
	.w4(32'h3ba2b849),
	.w5(32'h3b9c3ce3),
	.w6(32'h3bd3ce08),
	.w7(32'h3b88d33a),
	.w8(32'h3b885176),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b248339),
	.w1(32'h3c16414e),
	.w2(32'h3b6aab39),
	.w3(32'h3b4e33b9),
	.w4(32'h3c284d13),
	.w5(32'h3b4a7a5e),
	.w6(32'hbc3db329),
	.w7(32'hbc2e162b),
	.w8(32'hbc2a680b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9047a35),
	.w1(32'h3bc6fe3f),
	.w2(32'h3bc5e830),
	.w3(32'hbb353f44),
	.w4(32'h3afa27bd),
	.w5(32'hbb9e519d),
	.w6(32'h3b6c6c5b),
	.w7(32'h3b97debf),
	.w8(32'h3b3555b3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e5feb),
	.w1(32'h3b948302),
	.w2(32'h3c58adfb),
	.w3(32'hb921973c),
	.w4(32'hbbe73217),
	.w5(32'h3c5850c6),
	.w6(32'hbba912aa),
	.w7(32'hba3e5b67),
	.w8(32'hbb501189),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d6772),
	.w1(32'hbb849582),
	.w2(32'hbc86b6f2),
	.w3(32'h3c540a4b),
	.w4(32'hbb842c06),
	.w5(32'hbc46b5a4),
	.w6(32'h3b88b774),
	.w7(32'hbb48bc33),
	.w8(32'hbb32f799),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac56e7),
	.w1(32'h3bbb4efa),
	.w2(32'h39b14843),
	.w3(32'hbc6c2e6c),
	.w4(32'h3ab56bdb),
	.w5(32'hbaf5582a),
	.w6(32'h3abff684),
	.w7(32'hb9ff8eb2),
	.w8(32'h3a92c329),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951906),
	.w1(32'hb9aec5b5),
	.w2(32'hba85ff53),
	.w3(32'h3b184272),
	.w4(32'hbbbfb6d3),
	.w5(32'hbc214344),
	.w6(32'hb8c6c70e),
	.w7(32'hbad64e58),
	.w8(32'h3a7c108b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b65e),
	.w1(32'hbd232964),
	.w2(32'hbd7ff147),
	.w3(32'h3b4b4c84),
	.w4(32'hbcf7e909),
	.w5(32'hbd1a79cf),
	.w6(32'hbbe0674a),
	.w7(32'hbd03c6fd),
	.w8(32'hbd01486c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ecf80),
	.w1(32'hbcf8b3f9),
	.w2(32'hbd8e5edb),
	.w3(32'hbc5e2200),
	.w4(32'hbcb81bb1),
	.w5(32'hbce3b8c7),
	.w6(32'hbc6d075f),
	.w7(32'hbcffdac0),
	.w8(32'hbd1a65cb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1ae93c),
	.w1(32'hbb968afb),
	.w2(32'hbaa7a6ce),
	.w3(32'hbbc736c3),
	.w4(32'h39fa5ea5),
	.w5(32'hbb4f3f70),
	.w6(32'hbbb2a0e3),
	.w7(32'hba9f4454),
	.w8(32'h3603d9ac),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ff6ee),
	.w1(32'h3bb2352a),
	.w2(32'h3c0b2eff),
	.w3(32'h3abf25d4),
	.w4(32'hba73bd92),
	.w5(32'h3b9bb2a5),
	.w6(32'h3b413284),
	.w7(32'h3c26ce0a),
	.w8(32'hba0b1b15),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5eb2ce),
	.w1(32'hbb43efa9),
	.w2(32'hbac3c364),
	.w3(32'hbb25704d),
	.w4(32'hbbeec8cc),
	.w5(32'hbb3923c8),
	.w6(32'hbbd24e08),
	.w7(32'h3b112640),
	.w8(32'hbbb29dcb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba10ec9),
	.w1(32'h3ad23435),
	.w2(32'h36c57560),
	.w3(32'hbbd7eeb9),
	.w4(32'hbb29a562),
	.w5(32'hbac46e40),
	.w6(32'h3b1d3294),
	.w7(32'h3b263e36),
	.w8(32'h3b12cdd6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad201b),
	.w1(32'h3a8f5676),
	.w2(32'h3c90d4c7),
	.w3(32'h3af03f25),
	.w4(32'hbc0273ec),
	.w5(32'h3c652268),
	.w6(32'h3ab36dd1),
	.w7(32'h394bc3c7),
	.w8(32'hbb28c5b3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d4ae),
	.w1(32'hbc3506bf),
	.w2(32'hbc302499),
	.w3(32'hb91d8f81),
	.w4(32'h3a2d40b2),
	.w5(32'hbbaf9ba8),
	.w6(32'hbba42866),
	.w7(32'hbb8901df),
	.w8(32'h3a2bff14),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca765c),
	.w1(32'hbc929ffd),
	.w2(32'hbcdba974),
	.w3(32'h3b1af958),
	.w4(32'hbbdfc70d),
	.w5(32'hbbfe22e6),
	.w6(32'hbcb01958),
	.w7(32'hbcefa2f1),
	.w8(32'hbc95d4b8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8a5ff),
	.w1(32'h3c247939),
	.w2(32'h3c4fdfb6),
	.w3(32'hbc0bb1e1),
	.w4(32'h3b30a200),
	.w5(32'h3ca643fe),
	.w6(32'h3b3ded6e),
	.w7(32'hbbb005c5),
	.w8(32'hb9823561),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88cbd9),
	.w1(32'hbb6b7f3a),
	.w2(32'hbbeaadea),
	.w3(32'h3ca135ad),
	.w4(32'hb9bf635b),
	.w5(32'hbb7e931b),
	.w6(32'hbb41532a),
	.w7(32'hbbefb29b),
	.w8(32'hbb8748d5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50c623),
	.w1(32'h3b066651),
	.w2(32'hba496c16),
	.w3(32'h3b79fc63),
	.w4(32'hbb10a8e8),
	.w5(32'h3a052949),
	.w6(32'h3a3cbb33),
	.w7(32'hba40b295),
	.w8(32'hbaf83aba),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba831bb0),
	.w1(32'hbc07f8b6),
	.w2(32'hbccc1655),
	.w3(32'hbb044015),
	.w4(32'hbbeedc73),
	.w5(32'hbca97e93),
	.w6(32'hbb866831),
	.w7(32'hbc2f09ec),
	.w8(32'hbb1075b8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd80d08),
	.w1(32'h3bb2beee),
	.w2(32'hba969342),
	.w3(32'h3bae86f5),
	.w4(32'hba657099),
	.w5(32'hbaff545f),
	.w6(32'h3b0de8b3),
	.w7(32'h3b7b42c7),
	.w8(32'hbb24238b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe74734),
	.w1(32'h3b4f8322),
	.w2(32'h3b2af567),
	.w3(32'hbb293896),
	.w4(32'h3bac1a71),
	.w5(32'h3aebae77),
	.w6(32'hbb300526),
	.w7(32'hbbb2e3d4),
	.w8(32'h3afa066a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3be15b),
	.w1(32'h3bc798a6),
	.w2(32'h3c5ff902),
	.w3(32'h3c2219f0),
	.w4(32'h3c2968a8),
	.w5(32'h3c2c812f),
	.w6(32'hbc5ee5bb),
	.w7(32'hbb24b798),
	.w8(32'h392f7c4a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ffba1),
	.w1(32'h3a8c4e5b),
	.w2(32'hba2b9fce),
	.w3(32'h3ae4331a),
	.w4(32'hba0d3f73),
	.w5(32'hbb1d729b),
	.w6(32'h3aa6378f),
	.w7(32'h3b381337),
	.w8(32'hba823fc1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40b431),
	.w1(32'hba829556),
	.w2(32'h3b7e0a67),
	.w3(32'hbba3773d),
	.w4(32'hbac0c90b),
	.w5(32'h3ba9a44c),
	.w6(32'hbbb2b67c),
	.w7(32'hbb6e85da),
	.w8(32'h392aee15),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9498cd),
	.w1(32'hbcf24627),
	.w2(32'hbd7ca113),
	.w3(32'h3b3ebce1),
	.w4(32'hbcea3e09),
	.w5(32'hbd5b4978),
	.w6(32'hbc7a5f98),
	.w7(32'hbd0556cb),
	.w8(32'hbce71d32),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28cfe5),
	.w1(32'h3bf923bf),
	.w2(32'h3c075794),
	.w3(32'hbccccfb1),
	.w4(32'h3bd8a016),
	.w5(32'h3bc10410),
	.w6(32'h3c0e4875),
	.w7(32'h3bc036af),
	.w8(32'hbbac5dea),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0379b5),
	.w1(32'h3940012a),
	.w2(32'h3c57d0f8),
	.w3(32'h3bdbebb4),
	.w4(32'hba7172d8),
	.w5(32'h3bd48d23),
	.w6(32'h3c1e055e),
	.w7(32'h3bbe1c4b),
	.w8(32'h3b1f962c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e3038),
	.w1(32'hbb579a8b),
	.w2(32'hbb8a8bc2),
	.w3(32'h3b371c7e),
	.w4(32'hbb19e2c0),
	.w5(32'h3b9d829b),
	.w6(32'hbc5ae156),
	.w7(32'hbbb42d8e),
	.w8(32'h3a289885),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ac6d7),
	.w1(32'hbc530136),
	.w2(32'hbcc35eb7),
	.w3(32'h3b861102),
	.w4(32'hbbe68446),
	.w5(32'hbbd0fa44),
	.w6(32'hbb7d3b1c),
	.w7(32'hbc7d31a2),
	.w8(32'hbc966fe3),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc98a410),
	.w1(32'hbaa3b5c7),
	.w2(32'h3a17f2a9),
	.w3(32'h3982519a),
	.w4(32'hbb6a7cb5),
	.w5(32'hb8fe57e5),
	.w6(32'hbc091758),
	.w7(32'hbb9c2f4c),
	.w8(32'hba63b42b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4340b),
	.w1(32'h3c675ed7),
	.w2(32'hbaf960e7),
	.w3(32'h39ac766b),
	.w4(32'h3c60c770),
	.w5(32'h3b9e6ba8),
	.w6(32'h3bf70922),
	.w7(32'h3b945586),
	.w8(32'h38071869),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd00a04),
	.w1(32'hbcdab536),
	.w2(32'hbd2f211b),
	.w3(32'hbc053181),
	.w4(32'hbbb63f38),
	.w5(32'hbcb95d91),
	.w6(32'hbbf3f169),
	.w7(32'hbc88ecc1),
	.w8(32'hbbf17b04),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdd9b16),
	.w1(32'h3c00f64e),
	.w2(32'h3b830d4e),
	.w3(32'hbccd1a59),
	.w4(32'h3c187a4a),
	.w5(32'hbb04ed62),
	.w6(32'hbb8b6674),
	.w7(32'hba2d47b8),
	.w8(32'h3a6b458c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0acda8),
	.w1(32'hbc59de90),
	.w2(32'hbc1edfe8),
	.w3(32'h3c3b6726),
	.w4(32'hbc0d6b90),
	.w5(32'hbac96d61),
	.w6(32'hbae3d95c),
	.w7(32'hbb88641b),
	.w8(32'hbc0f5daa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6fcfa),
	.w1(32'h3c86ad8c),
	.w2(32'h3cb9710d),
	.w3(32'h39ee7c7b),
	.w4(32'h3b0412b4),
	.w5(32'h3c8c2c62),
	.w6(32'h3b4dd3e2),
	.w7(32'h3c3015b5),
	.w8(32'h3b3e80c2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b905085),
	.w1(32'hbc07ceaf),
	.w2(32'hbc3e4d3e),
	.w3(32'h3c10c4a0),
	.w4(32'hbb8ba8c5),
	.w5(32'hba49bc3b),
	.w6(32'hbbe21780),
	.w7(32'hbc094012),
	.w8(32'hbc0df20d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ff56),
	.w1(32'h3a8b0c91),
	.w2(32'h3ba1176b),
	.w3(32'h39d78ee8),
	.w4(32'h3b612a87),
	.w5(32'h3b9ce348),
	.w6(32'hbb967229),
	.w7(32'h3ad95ec2),
	.w8(32'hbafe5224),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b0f47),
	.w1(32'hbb31741a),
	.w2(32'hbbc4862f),
	.w3(32'h3b222e09),
	.w4(32'hbbcda04b),
	.w5(32'hbc131527),
	.w6(32'hbb212297),
	.w7(32'h3b85e204),
	.w8(32'hba5894bb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd5654),
	.w1(32'hbcc95157),
	.w2(32'hbc9143a5),
	.w3(32'hbbfaeb38),
	.w4(32'hbb5a1f83),
	.w5(32'hb9ed601f),
	.w6(32'hbcd195f4),
	.w7(32'hbcdcc2e1),
	.w8(32'hbc29b22a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86dce3),
	.w1(32'h3baa9601),
	.w2(32'h39e9f6db),
	.w3(32'hbc41c697),
	.w4(32'h3bc5d227),
	.w5(32'h3b6a763d),
	.w6(32'h3c14398f),
	.w7(32'h3bd39bdb),
	.w8(32'h3b57ffeb),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90f401),
	.w1(32'h3ccafc66),
	.w2(32'h3d289297),
	.w3(32'hbb90cf8e),
	.w4(32'h3ca1f5ca),
	.w5(32'h3cf8a948),
	.w6(32'h3c403af4),
	.w7(32'h3d13b1ca),
	.w8(32'h3ce21c38),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d151c09),
	.w1(32'h3c69f8ae),
	.w2(32'h3c264308),
	.w3(32'h3caa8495),
	.w4(32'h3988a3c4),
	.w5(32'h3c44c160),
	.w6(32'h3c151174),
	.w7(32'h3bb24bac),
	.w8(32'h3b7ad29d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd4e6),
	.w1(32'h3c6fa274),
	.w2(32'h3c3272fb),
	.w3(32'h3be6c0e7),
	.w4(32'hba16e8a0),
	.w5(32'hbbbd410a),
	.w6(32'h3c5101d1),
	.w7(32'h3c9644ee),
	.w8(32'hbbb4220c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16abf9),
	.w1(32'h3c1ba9e3),
	.w2(32'h3c1a9a6f),
	.w3(32'h3bc7e081),
	.w4(32'h3c4939de),
	.w5(32'h3c4cb25b),
	.w6(32'h3c83f35f),
	.w7(32'h3c96b140),
	.w8(32'h3c7a31ab),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65ff80),
	.w1(32'h3b9f06a0),
	.w2(32'hbc178989),
	.w3(32'h3c21bfdb),
	.w4(32'hbad970c7),
	.w5(32'hbc46b758),
	.w6(32'h3932caf4),
	.w7(32'h3bfab107),
	.w8(32'hbb22354a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854486),
	.w1(32'hbbe095af),
	.w2(32'hbb929ff2),
	.w3(32'hbc3113b1),
	.w4(32'hbb133620),
	.w5(32'hbb10ada4),
	.w6(32'hbbe901c2),
	.w7(32'hba85f88f),
	.w8(32'h3bad036a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5d16),
	.w1(32'h3bf8626a),
	.w2(32'h3b0fbfc3),
	.w3(32'hba89108f),
	.w4(32'h3bcd4f83),
	.w5(32'hb981c91e),
	.w6(32'hbb9fce3e),
	.w7(32'hbad8c24f),
	.w8(32'hbb16fe4a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16dfdc),
	.w1(32'hbb512c22),
	.w2(32'hbb305877),
	.w3(32'hbb9e03d6),
	.w4(32'h39871fc2),
	.w5(32'h39fa8784),
	.w6(32'h3bc54fce),
	.w7(32'h3bcb0d1d),
	.w8(32'h3b0004b7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23aebe),
	.w1(32'hbc4d91aa),
	.w2(32'hbcbc8ff9),
	.w3(32'h3ae06b85),
	.w4(32'hbba1c70a),
	.w5(32'hbc27491a),
	.w6(32'hbb6dd330),
	.w7(32'hbc7ed447),
	.w8(32'hbc7e707d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63f4e0),
	.w1(32'hbc51333f),
	.w2(32'hbd021929),
	.w3(32'hbbae41db),
	.w4(32'hb9fbcc0e),
	.w5(32'hbcd66338),
	.w6(32'hbbd42684),
	.w7(32'hbc077c66),
	.w8(32'h3ac7d31e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e96b5),
	.w1(32'h3c6afa64),
	.w2(32'h3d2c28f6),
	.w3(32'hbce12501),
	.w4(32'h3c2441e3),
	.w5(32'h3cd11446),
	.w6(32'h3aeaa741),
	.w7(32'h3c81612f),
	.w8(32'h3be866d5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1d4c33),
	.w1(32'hbab50987),
	.w2(32'hb9bd98bd),
	.w3(32'h3c858180),
	.w4(32'hba33ef6d),
	.w5(32'hba2f4249),
	.w6(32'hbb80485d),
	.w7(32'hba946eef),
	.w8(32'hba867550),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba9802),
	.w1(32'h3a7031f2),
	.w2(32'h39f2b534),
	.w3(32'hb925fad5),
	.w4(32'hbb2228e4),
	.w5(32'hbb63db7b),
	.w6(32'hbb9ddc8b),
	.w7(32'hbb411135),
	.w8(32'hbb79815f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0525bb),
	.w1(32'h3b4f1c5c),
	.w2(32'hbb4b65f0),
	.w3(32'h3b3631b0),
	.w4(32'hbc0f2db0),
	.w5(32'hbb931422),
	.w6(32'hbb06c590),
	.w7(32'hbc14c61d),
	.w8(32'hbc3ab232),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73d77),
	.w1(32'h3b8b3cf6),
	.w2(32'h3bfd825b),
	.w3(32'h3b6436a1),
	.w4(32'h3ba77bfb),
	.w5(32'h3bc65961),
	.w6(32'hbb6cbc1a),
	.w7(32'hbac0c78a),
	.w8(32'hbb353ec4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6dca),
	.w1(32'h3bacbaa7),
	.w2(32'h3cc2aa7a),
	.w3(32'h3af87182),
	.w4(32'h3ade1357),
	.w5(32'h3c5ca2a5),
	.w6(32'h3c163dc7),
	.w7(32'h3bb315cf),
	.w8(32'hbbad0479),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be10f7c),
	.w1(32'h3cb55132),
	.w2(32'h3d27527a),
	.w3(32'h3c7551ef),
	.w4(32'h3c89812f),
	.w5(32'h3d0126b3),
	.w6(32'h3c83526f),
	.w7(32'h3ce1f6bd),
	.w8(32'h3c756e60),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03ec4c),
	.w1(32'h3d0ad36d),
	.w2(32'h3d7273ff),
	.w3(32'h3ccd5a2a),
	.w4(32'h3c76e79a),
	.w5(32'h3d28a24c),
	.w6(32'h3cb35db2),
	.w7(32'h3d1d1509),
	.w8(32'h3c887ca1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c9a27),
	.w1(32'hbb01a621),
	.w2(32'hbc1e048c),
	.w3(32'h3cf24e63),
	.w4(32'h3b9139b9),
	.w5(32'hbae95cf2),
	.w6(32'hbc0324de),
	.w7(32'hbbc317aa),
	.w8(32'hbb23ac84),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18bb89),
	.w1(32'hbc8631af),
	.w2(32'hbbaa3dde),
	.w3(32'h3a85f88b),
	.w4(32'hbc53acf5),
	.w5(32'hbbe2ac91),
	.w6(32'hbb4ead74),
	.w7(32'hbbbbb0b2),
	.w8(32'hbbb2a9e4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb4b2c),
	.w1(32'h3a85433b),
	.w2(32'hbb3d32d2),
	.w3(32'hbbf530a4),
	.w4(32'h3a4af98c),
	.w5(32'hbc136708),
	.w6(32'hbb316038),
	.w7(32'h3b755856),
	.w8(32'h3bbf536a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944443),
	.w1(32'h3d1325ef),
	.w2(32'h3d99f437),
	.w3(32'hbba6e0ba),
	.w4(32'h3ca5e201),
	.w5(32'h3d424c6c),
	.w6(32'h3d05fa08),
	.w7(32'h3d1a60a4),
	.w8(32'h3cad3188),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d244327),
	.w1(32'hbd301966),
	.w2(32'hbd56e1ec),
	.w3(32'h3cfa4bfa),
	.w4(32'hbcd40902),
	.w5(32'hbbe65c97),
	.w6(32'hbccbcd38),
	.w7(32'hbd2facd0),
	.w8(32'hbcc36323),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc72383),
	.w1(32'h3cde0a35),
	.w2(32'h3cac2903),
	.w3(32'hbb99c1aa),
	.w4(32'h3c9356ab),
	.w5(32'h3cb29ccb),
	.w6(32'h3c48e702),
	.w7(32'h3bf3b41f),
	.w8(32'h3c0ad5f0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bb6a4),
	.w1(32'h3b44c125),
	.w2(32'hbb201ad6),
	.w3(32'h3c516c86),
	.w4(32'hb9086a66),
	.w5(32'hbb934b47),
	.w6(32'hbb9c7dbc),
	.w7(32'hbbe7714e),
	.w8(32'hbbd53bec),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cd75f),
	.w1(32'hbb1a4a2b),
	.w2(32'hbc2eced4),
	.w3(32'hbabc63a6),
	.w4(32'hbb8a55be),
	.w5(32'hbbf20885),
	.w6(32'hb9dd3509),
	.w7(32'hba0f166d),
	.w8(32'hbbbb77ce),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd44ba),
	.w1(32'hb9ffd2b0),
	.w2(32'hbb9cf00d),
	.w3(32'h3ae551e0),
	.w4(32'h3acfc650),
	.w5(32'hbc09c15e),
	.w6(32'h3b0bf67e),
	.w7(32'hbbba466b),
	.w8(32'hbb0a8344),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d8e1),
	.w1(32'h3c3742b7),
	.w2(32'h3ccadd54),
	.w3(32'h3a9d9723),
	.w4(32'h3c1afd24),
	.w5(32'h3c1d8ca2),
	.w6(32'h3c2bd9b0),
	.w7(32'h3c7c64e3),
	.w8(32'h3c6a6f9c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e33f2),
	.w1(32'hbac10c95),
	.w2(32'hb9dc7d0b),
	.w3(32'h3c2ae95d),
	.w4(32'hbab5a823),
	.w5(32'h3ab359ce),
	.w6(32'hb9d5f8ff),
	.w7(32'hbaf5e939),
	.w8(32'hb9f692cf),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61cfac),
	.w1(32'h3d156324),
	.w2(32'h3d6fd82f),
	.w3(32'h3b4c7e9b),
	.w4(32'h3ca1a2b0),
	.w5(32'h3d23713e),
	.w6(32'h3ce18cf8),
	.w7(32'h3ce7b5bc),
	.w8(32'h3c82a3ea),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3e83f6),
	.w1(32'h3b1b6137),
	.w2(32'h3bdf34ca),
	.w3(32'h3ccd35ea),
	.w4(32'h3b4f92df),
	.w5(32'h3b804590),
	.w6(32'hbb83c6ba),
	.w7(32'h3a3abac1),
	.w8(32'hb98ace0b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9f229),
	.w1(32'h3996cf4b),
	.w2(32'hbc055415),
	.w3(32'h3b6741dc),
	.w4(32'h38340d08),
	.w5(32'hbc1a1d17),
	.w6(32'h3a85040e),
	.w7(32'hbbd9e8b7),
	.w8(32'hbc25aa45),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69ceee),
	.w1(32'hbc72fb91),
	.w2(32'hbcc00c4f),
	.w3(32'h3b5d8a9a),
	.w4(32'hbb5689b1),
	.w5(32'h3b90efa9),
	.w6(32'hbbcf62a8),
	.w7(32'hbcb88624),
	.w8(32'hbc3e9000),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2aa5c),
	.w1(32'hbb971506),
	.w2(32'hbb184d78),
	.w3(32'h3bf0f7f4),
	.w4(32'h3a7fec96),
	.w5(32'hbb412aa3),
	.w6(32'hbb5adfc5),
	.w7(32'h3b57340c),
	.w8(32'h3af24e38),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7add332),
	.w1(32'hb998eec8),
	.w2(32'h3b0ed18b),
	.w3(32'hba9b9518),
	.w4(32'hb9d05046),
	.w5(32'h3b83099a),
	.w6(32'hba5d31ff),
	.w7(32'h3a515f20),
	.w8(32'h3ac8009b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8ba9),
	.w1(32'h3be3838a),
	.w2(32'h3c034085),
	.w3(32'h3b247a88),
	.w4(32'h3bf9c052),
	.w5(32'h3bc6a348),
	.w6(32'h3c5ba6b4),
	.w7(32'h3c7cf510),
	.w8(32'h3c36d497),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e2b98),
	.w1(32'h38e6ef35),
	.w2(32'h3b1fc9da),
	.w3(32'h3bc78040),
	.w4(32'h3c14086c),
	.w5(32'h3bad9045),
	.w6(32'hbb6862db),
	.w7(32'hb99a37b3),
	.w8(32'h3b62a7e9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d8e79),
	.w1(32'hbbb94241),
	.w2(32'hbb973158),
	.w3(32'hbb43b393),
	.w4(32'h3c153f28),
	.w5(32'h3bb952c1),
	.w6(32'hb97a54e8),
	.w7(32'hbbc5ca96),
	.w8(32'hba9323b9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb580c7d),
	.w1(32'hbbb9d580),
	.w2(32'hbb80e5fd),
	.w3(32'hba37740b),
	.w4(32'hbbc96ee7),
	.w5(32'hba8d26cd),
	.w6(32'hb9469688),
	.w7(32'hbbcfad69),
	.w8(32'hbb6175b1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20889d),
	.w1(32'hbc2721de),
	.w2(32'hbc8de56f),
	.w3(32'h3b4a9265),
	.w4(32'h3be3426e),
	.w5(32'hbb1628f4),
	.w6(32'hbc29a8bb),
	.w7(32'hbca94636),
	.w8(32'hbb7a5423),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefba70),
	.w1(32'hb9f3dc06),
	.w2(32'h3981d1ea),
	.w3(32'h3a40e6c5),
	.w4(32'h3b13cd44),
	.w5(32'h3ae678d0),
	.w6(32'h3b9980bf),
	.w7(32'h3ac40bbd),
	.w8(32'h3aee232d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c001742),
	.w1(32'h3b83a9d6),
	.w2(32'h3ba16ffc),
	.w3(32'hba64c3b8),
	.w4(32'h3a5afbe5),
	.w5(32'h3b879ad6),
	.w6(32'h39be1adc),
	.w7(32'h3b5ae940),
	.w8(32'hbb11a90f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8450e4),
	.w1(32'hbb68d2f8),
	.w2(32'hbcb2da25),
	.w3(32'h39037a5c),
	.w4(32'hbabefaf3),
	.w5(32'hbc760edf),
	.w6(32'hbb6cc2b1),
	.w7(32'hbba724ef),
	.w8(32'hbaac709c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15707b),
	.w1(32'h3c08c23b),
	.w2(32'h3c17e9af),
	.w3(32'h3a8ca83f),
	.w4(32'h3c580af8),
	.w5(32'h3c2d4710),
	.w6(32'h3c0ee09b),
	.w7(32'h3c825ea5),
	.w8(32'h3c3e8838),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b865391),
	.w1(32'hbcd7ec08),
	.w2(32'hbd5b65b6),
	.w3(32'h3cb7ed4c),
	.w4(32'hbca968e8),
	.w5(32'hbceedb5a),
	.w6(32'hbb44d432),
	.w7(32'hbcdd7b5b),
	.w8(32'hbd11e503),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd029b46),
	.w1(32'hbaa021ff),
	.w2(32'h3b20e6b6),
	.w3(32'h3a0e6adb),
	.w4(32'hba83ee3a),
	.w5(32'h3a6a63e5),
	.w6(32'hba942457),
	.w7(32'hb9d67b96),
	.w8(32'h36f4aa76),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3b5d4),
	.w1(32'hbcd564dd),
	.w2(32'hbbf39f90),
	.w3(32'hba50d074),
	.w4(32'hbc83df6a),
	.w5(32'hbade7d8f),
	.w6(32'hbc7c3bf5),
	.w7(32'hbc5d74b0),
	.w8(32'h3b441292),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule