module layer_10_featuremap_351(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8945b8),
	.w1(32'h3b497194),
	.w2(32'h38f9e683),
	.w3(32'h3b50ba56),
	.w4(32'hbb147eb8),
	.w5(32'h3acaae05),
	.w6(32'h3b857cdb),
	.w7(32'hbb2ac0bf),
	.w8(32'h3c138097),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b777fe9),
	.w1(32'h3bf0ba71),
	.w2(32'h3b109105),
	.w3(32'h3bf18403),
	.w4(32'h3b630b33),
	.w5(32'h3880e15f),
	.w6(32'h3c79450d),
	.w7(32'h3ba3cc61),
	.w8(32'hb89d3879),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac76667),
	.w1(32'h3ad8f296),
	.w2(32'h3931b54b),
	.w3(32'hbb754b03),
	.w4(32'hba885d48),
	.w5(32'hbb05f1d0),
	.w6(32'hb9a3e3eb),
	.w7(32'h3b8f209d),
	.w8(32'h392c6939),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9c31),
	.w1(32'h3ae99505),
	.w2(32'hb9bf1524),
	.w3(32'hba73185d),
	.w4(32'hbaa34a47),
	.w5(32'hba945756),
	.w6(32'hba9b8967),
	.w7(32'hba4470bf),
	.w8(32'hbb4384b8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8b061),
	.w1(32'h3b32cce3),
	.w2(32'h3aa6ada0),
	.w3(32'hba67e410),
	.w4(32'hb90650c5),
	.w5(32'h3a0104ab),
	.w6(32'hbbe54046),
	.w7(32'hbb586308),
	.w8(32'h3ab1ab11),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1000ae),
	.w1(32'h3b06533c),
	.w2(32'hb8d8f4f3),
	.w3(32'h3ae581a6),
	.w4(32'h3acfe1cd),
	.w5(32'hba7a0f3a),
	.w6(32'h3b061eea),
	.w7(32'h3a989392),
	.w8(32'h3a524c22),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9a9df),
	.w1(32'h3c0b9c07),
	.w2(32'h3b20aa4b),
	.w3(32'h3b8d5d5b),
	.w4(32'h3b0f49a9),
	.w5(32'h3b61e22d),
	.w6(32'h3b19ed70),
	.w7(32'h38355b59),
	.w8(32'h3a15436a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb435f62),
	.w1(32'hbb265650),
	.w2(32'hbade5895),
	.w3(32'hbb800989),
	.w4(32'hbb0c7fcd),
	.w5(32'hbb4890c4),
	.w6(32'hbbc0365d),
	.w7(32'h3b611451),
	.w8(32'h3a3bff40),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b903),
	.w1(32'h3b36b438),
	.w2(32'h3b21fb9a),
	.w3(32'h3b1e419f),
	.w4(32'h3ba90e21),
	.w5(32'hbaf588bd),
	.w6(32'h3b287922),
	.w7(32'h3b1bfcfc),
	.w8(32'hbaec01fa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919a4e0),
	.w1(32'hb920d36f),
	.w2(32'hb89120ef),
	.w3(32'hba5f016f),
	.w4(32'hba97171a),
	.w5(32'h3b71b647),
	.w6(32'hbb3e32df),
	.w7(32'hbb393dea),
	.w8(32'h3b6cea3d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fa0ca),
	.w1(32'h3b9943a0),
	.w2(32'h3b1d5e01),
	.w3(32'h3b570606),
	.w4(32'h3b309174),
	.w5(32'hbace328c),
	.w6(32'h3b28c0ef),
	.w7(32'h3a80b157),
	.w8(32'hbb569fee),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f838),
	.w1(32'h3aa2b927),
	.w2(32'hba868548),
	.w3(32'h3b0ca10d),
	.w4(32'h3b62dbbf),
	.w5(32'hbb14ef19),
	.w6(32'hbb3c9ff0),
	.w7(32'h3b8f1a2b),
	.w8(32'hbbccbb30),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb487a3e),
	.w1(32'hbba76868),
	.w2(32'hbb2e9b18),
	.w3(32'hbb48f1e2),
	.w4(32'hbaac019c),
	.w5(32'hba2c6c16),
	.w6(32'hbbb07e64),
	.w7(32'hbaf176c4),
	.w8(32'hbb01b3ab),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52363f),
	.w1(32'hbb7849c7),
	.w2(32'hbab099a1),
	.w3(32'hbb3f5831),
	.w4(32'hbb30ea54),
	.w5(32'hbb1fd3d6),
	.w6(32'hbb517c38),
	.w7(32'hbb210aab),
	.w8(32'hbb8bef3c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d3c25),
	.w1(32'h3983018b),
	.w2(32'hb9e89cf2),
	.w3(32'h396c69e0),
	.w4(32'hb99c8111),
	.w5(32'hba011731),
	.w6(32'hbb3c9e8e),
	.w7(32'hbb3555ac),
	.w8(32'hbb4927af),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c564),
	.w1(32'hbb6c88d3),
	.w2(32'hbb840f55),
	.w3(32'hbba9cdc0),
	.w4(32'hbbd37363),
	.w5(32'h3b373a34),
	.w6(32'hbb9408de),
	.w7(32'hbc10665e),
	.w8(32'hbb2bb6e4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5df56),
	.w1(32'hbae587c6),
	.w2(32'hbab51967),
	.w3(32'h39a681d7),
	.w4(32'h39dc2878),
	.w5(32'h3ab1644a),
	.w6(32'hb92b43dc),
	.w7(32'h3b345737),
	.w8(32'h3b99de89),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb366914),
	.w1(32'hbc13db6d),
	.w2(32'hbc2571e9),
	.w3(32'hbc06a9fb),
	.w4(32'hbc16fe97),
	.w5(32'hbc4daadb),
	.w6(32'hbb7fd648),
	.w7(32'hbc00a4fd),
	.w8(32'hbba3fc3c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a179),
	.w1(32'hbc139e69),
	.w2(32'hbc14e0a1),
	.w3(32'hbbe3d69f),
	.w4(32'hbbc7e05e),
	.w5(32'hbbef558a),
	.w6(32'h3b26718a),
	.w7(32'h39ee2ef4),
	.w8(32'hbbd25ff0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44d804),
	.w1(32'hb997aa63),
	.w2(32'hbb458240),
	.w3(32'hbb2ec359),
	.w4(32'hba6a3b13),
	.w5(32'hbb41aebe),
	.w6(32'hbbb18cb6),
	.w7(32'hbb2944d7),
	.w8(32'hb9efbb2c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52cf9f),
	.w1(32'hbb35f7c0),
	.w2(32'hbb61fd62),
	.w3(32'hbb6c10b2),
	.w4(32'hbb88f9e0),
	.w5(32'hb8d9ceed),
	.w6(32'hbb196923),
	.w7(32'hbb664136),
	.w8(32'hbb2e4634),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a835fd6),
	.w1(32'h3a9c3385),
	.w2(32'h39f9ab78),
	.w3(32'h3acc2dd7),
	.w4(32'h3a6f95aa),
	.w5(32'hbabd1108),
	.w6(32'hbafca5ae),
	.w7(32'hba687f1f),
	.w8(32'hb9a01100),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6566c4),
	.w1(32'hbc231fba),
	.w2(32'hbc5133dc),
	.w3(32'hbbfbb01a),
	.w4(32'hbc09f1cb),
	.w5(32'hbc3264fc),
	.w6(32'hbc01e5fa),
	.w7(32'hbbfbb83f),
	.w8(32'hbc24b9a6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bced5),
	.w1(32'h3b41421d),
	.w2(32'h3baee053),
	.w3(32'h3ad62e7a),
	.w4(32'hba5b2d65),
	.w5(32'h3b4e49ac),
	.w6(32'h3bc00adb),
	.w7(32'h3b8793b4),
	.w8(32'hbabf1d1f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4117fd),
	.w1(32'h3b4a7cad),
	.w2(32'h3bbd6f0b),
	.w3(32'h3bd602f6),
	.w4(32'h3bd5b732),
	.w5(32'h3bd8fd17),
	.w6(32'h3b757225),
	.w7(32'h3b046370),
	.w8(32'h3a5d5380),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab70434),
	.w1(32'h3b489d98),
	.w2(32'h3afbb80c),
	.w3(32'h3b1f9157),
	.w4(32'hb94d19d4),
	.w5(32'hb8d381b8),
	.w6(32'hbb1c6f36),
	.w7(32'hbaad202e),
	.w8(32'h3b1149c5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d36762),
	.w1(32'h39384407),
	.w2(32'h3aa2d4db),
	.w3(32'hbb2b3e73),
	.w4(32'hbb1b72ff),
	.w5(32'hbaea16a9),
	.w6(32'h3a294459),
	.w7(32'h3a6cf9d7),
	.w8(32'hbaed2459),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ccd1a),
	.w1(32'h39859bf4),
	.w2(32'h3ae5cdb1),
	.w3(32'h3ba4de3b),
	.w4(32'h3b92cd07),
	.w5(32'h3b618f92),
	.w6(32'h3ada7e38),
	.w7(32'hbb32a89d),
	.w8(32'hbb3ba8d7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19fbf6),
	.w1(32'hb9f0592c),
	.w2(32'hbb028bd7),
	.w3(32'h3b376ec1),
	.w4(32'h3ad2d780),
	.w5(32'hbaa098cb),
	.w6(32'hbafadfbb),
	.w7(32'h3ab425fc),
	.w8(32'hbab72099),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84312f),
	.w1(32'hb94619e8),
	.w2(32'hba8d99db),
	.w3(32'h3b1a0022),
	.w4(32'hbaa93291),
	.w5(32'hbafcefe6),
	.w6(32'h3a984b71),
	.w7(32'hb91273ee),
	.w8(32'h3ad4caab),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396922c6),
	.w1(32'h3a7d9e13),
	.w2(32'h3b21159c),
	.w3(32'hbc0dc958),
	.w4(32'hbaa0a513),
	.w5(32'hba2d2fb0),
	.w6(32'hbbc981cb),
	.w7(32'hbb9e72a9),
	.w8(32'hba7c94b1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4045),
	.w1(32'h3aa91b6f),
	.w2(32'h39f71f1e),
	.w3(32'hbaf9a993),
	.w4(32'hb98eda33),
	.w5(32'hbbe0e16d),
	.w6(32'hbb4508df),
	.w7(32'hb9e5460c),
	.w8(32'hbb3734e7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0f541),
	.w1(32'hbb03db75),
	.w2(32'hbbb17aba),
	.w3(32'hbb769d25),
	.w4(32'hbb18b381),
	.w5(32'h3aa0ec36),
	.w6(32'hbbc9ef01),
	.w7(32'hbb86def4),
	.w8(32'h3ab64cb1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa81852),
	.w1(32'hbad649bc),
	.w2(32'h3a04cfcf),
	.w3(32'h38843d34),
	.w4(32'h3b327698),
	.w5(32'h3b5d18d0),
	.w6(32'h3ace4e1f),
	.w7(32'h3b03c656),
	.w8(32'h3a158bd7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0462c4),
	.w1(32'hba18a68a),
	.w2(32'h3ade5cd6),
	.w3(32'h3b2a3c8a),
	.w4(32'hba9d6ebf),
	.w5(32'h3a9f67bd),
	.w6(32'h3a874478),
	.w7(32'hba1ed903),
	.w8(32'h39e12623),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace1400),
	.w1(32'h3b14da10),
	.w2(32'h3b88d02b),
	.w3(32'hbb1a8bed),
	.w4(32'h3b0f8da2),
	.w5(32'h39b48c38),
	.w6(32'h3b0aa453),
	.w7(32'h3b7af14a),
	.w8(32'hbbf60393),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ae143),
	.w1(32'hba708f75),
	.w2(32'hbbd02062),
	.w3(32'h39ea5aa5),
	.w4(32'hbae89760),
	.w5(32'h3c600c3d),
	.w6(32'hbbce1b4d),
	.w7(32'h3b8ee1dc),
	.w8(32'h3c895d4a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c832d82),
	.w1(32'h3c980ee5),
	.w2(32'h3c8b6c9e),
	.w3(32'h3c9673db),
	.w4(32'h3c681fe3),
	.w5(32'h3c0d2ede),
	.w6(32'h3cc59b38),
	.w7(32'h3c86efda),
	.w8(32'h3c0688a3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dd2c4),
	.w1(32'h3c5e1584),
	.w2(32'h3c1f7ea1),
	.w3(32'h3c5c114c),
	.w4(32'h3c295413),
	.w5(32'h3bc0708e),
	.w6(32'h3c56da80),
	.w7(32'h3bd8799b),
	.w8(32'hb802210f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5585c8),
	.w1(32'h39190424),
	.w2(32'hb987c658),
	.w3(32'h3ae78f72),
	.w4(32'hb91c4ce3),
	.w5(32'h3af3986d),
	.w6(32'hbae374bb),
	.w7(32'hbae47c40),
	.w8(32'h39a54bb4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e328),
	.w1(32'hbb69a850),
	.w2(32'h39bab3cf),
	.w3(32'hba111a48),
	.w4(32'hbaba1bde),
	.w5(32'hba66c4ad),
	.w6(32'hba27d77e),
	.w7(32'hb97610f4),
	.w8(32'hbb8d7c71),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b391b6e),
	.w1(32'h3bada373),
	.w2(32'h3b0fd30a),
	.w3(32'h3b4b2fdf),
	.w4(32'hb90efc20),
	.w5(32'h3bd79ce8),
	.w6(32'hbbbda24c),
	.w7(32'hbb363123),
	.w8(32'h3c3ebe9b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc33384),
	.w1(32'h3b749628),
	.w2(32'h3b4c4a55),
	.w3(32'h3bb9bb47),
	.w4(32'h3c02fb03),
	.w5(32'hbb3f0253),
	.w6(32'h3bea53a8),
	.w7(32'h3b147d6a),
	.w8(32'h3b1756b8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0817bb),
	.w1(32'hbc348010),
	.w2(32'hbb84d896),
	.w3(32'hbc45c600),
	.w4(32'hbbcaee9a),
	.w5(32'hbb10bc4c),
	.w6(32'hbb077217),
	.w7(32'hbbcb7753),
	.w8(32'hbbb0dbf5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0eec3),
	.w1(32'h3afabcd9),
	.w2(32'hba331d4a),
	.w3(32'h3a6349a6),
	.w4(32'hb899303f),
	.w5(32'hbaa71b3b),
	.w6(32'hbbad2503),
	.w7(32'hbaeba5dc),
	.w8(32'hbb5cdd1a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9ac21),
	.w1(32'hbb5bebb0),
	.w2(32'h3b8c5d7f),
	.w3(32'hbb221fb0),
	.w4(32'hbaaeb390),
	.w5(32'h3a9ee053),
	.w6(32'hbb0a03ae),
	.w7(32'hbb027630),
	.w8(32'h3ab7ad7d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2df31e),
	.w1(32'hbb3c21cb),
	.w2(32'hbac3b31b),
	.w3(32'hbac3f7cb),
	.w4(32'hbaa43436),
	.w5(32'h3b7b42a9),
	.w6(32'hbb86a2c4),
	.w7(32'hbb2d5c18),
	.w8(32'h39a5d66c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab1536),
	.w1(32'hbbc250f3),
	.w2(32'hbc0dc0a0),
	.w3(32'hbbc344db),
	.w4(32'hbbfbe3a1),
	.w5(32'hbc292fec),
	.w6(32'hbc211e17),
	.w7(32'hbc1686fa),
	.w8(32'hbc11fc9f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38500302),
	.w1(32'hbb15bc31),
	.w2(32'hba9cf204),
	.w3(32'hba6ba0de),
	.w4(32'h3aeb3210),
	.w5(32'h3a982e69),
	.w6(32'hbaddc8f2),
	.w7(32'hbabe5539),
	.w8(32'hbafdab95),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b179202),
	.w1(32'h3b3693fe),
	.w2(32'hba2e5901),
	.w3(32'h3a97037c),
	.w4(32'hba7e77bd),
	.w5(32'hbb9c8085),
	.w6(32'hbb5996f5),
	.w7(32'hbb35796d),
	.w8(32'hbb49da8a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af300e2),
	.w1(32'h3b01190e),
	.w2(32'h392e3918),
	.w3(32'hba4c615e),
	.w4(32'h3a7ad609),
	.w5(32'h3ba99bf9),
	.w6(32'hb9396d22),
	.w7(32'h3a143ce4),
	.w8(32'h3c9347d3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e52c),
	.w1(32'h3a7c05ba),
	.w2(32'h3b83b327),
	.w3(32'h3b05f4be),
	.w4(32'h39a5916e),
	.w5(32'hbae5648e),
	.w6(32'h3c956012),
	.w7(32'h3c14d873),
	.w8(32'hbb15f9f9),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023780),
	.w1(32'hbaa7106a),
	.w2(32'h3aa53519),
	.w3(32'hb9dcc338),
	.w4(32'hbaa9022f),
	.w5(32'hbb217ef3),
	.w6(32'hba2c55aa),
	.w7(32'h3b0b8c32),
	.w8(32'hbb7f8684),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9dc67),
	.w1(32'hbbc642fa),
	.w2(32'hbc2530f0),
	.w3(32'hbbfaba38),
	.w4(32'hbc3571c7),
	.w5(32'hbb4723c0),
	.w6(32'hbbd3fb1e),
	.w7(32'hbc300485),
	.w8(32'hbb7c9664),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb145d56),
	.w1(32'hb931634e),
	.w2(32'hbb4bd198),
	.w3(32'hba427f8d),
	.w4(32'hb9735cac),
	.w5(32'h3acbf6a3),
	.w6(32'hba0893e9),
	.w7(32'h3a32853d),
	.w8(32'hbac1a429),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a690638),
	.w1(32'h3b1616c0),
	.w2(32'h3afafc29),
	.w3(32'h3b22c0c5),
	.w4(32'h3abe584a),
	.w5(32'h3b56ac55),
	.w6(32'hbaf42ea1),
	.w7(32'hbb2f0deb),
	.w8(32'hbaa75105),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ff379),
	.w1(32'hba94a402),
	.w2(32'h3af0b6c7),
	.w3(32'h3a909ed0),
	.w4(32'h3a8f6101),
	.w5(32'hbafd898c),
	.w6(32'hbaca8d9e),
	.w7(32'hb99c3a92),
	.w8(32'hbac8b739),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394915bd),
	.w1(32'hba6fc9d9),
	.w2(32'hbb637963),
	.w3(32'hbb0958e0),
	.w4(32'hba98abbb),
	.w5(32'h3aad2b91),
	.w6(32'hbb7e39dd),
	.w7(32'hbb816673),
	.w8(32'hba47d4fe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eb0ae),
	.w1(32'h3bbd8c69),
	.w2(32'h3b3da7a4),
	.w3(32'h3b5fd01d),
	.w4(32'h3a83bccc),
	.w5(32'h3bbc3f54),
	.w6(32'hb7e2deb7),
	.w7(32'h389150b3),
	.w8(32'h3abda02f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaf326),
	.w1(32'h3afd38a3),
	.w2(32'h3c047fbb),
	.w3(32'h3b20d2c9),
	.w4(32'h3b380cfb),
	.w5(32'hbb1be0d4),
	.w6(32'h3ba20d01),
	.w7(32'h3bc6234f),
	.w8(32'hbb8b48a5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41f95a),
	.w1(32'hbb975793),
	.w2(32'hbbcd235d),
	.w3(32'hbb9b1135),
	.w4(32'hbb376da9),
	.w5(32'hbbd2a64a),
	.w6(32'hbbea443a),
	.w7(32'hbbd3aec9),
	.w8(32'hbc37de11),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff833c),
	.w1(32'hba44faf4),
	.w2(32'hbb4821d7),
	.w3(32'hbbaf55ac),
	.w4(32'hbbbcaf31),
	.w5(32'hbb5180bd),
	.w6(32'hbbf949f9),
	.w7(32'hbbf68861),
	.w8(32'hbb1f5ac5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb603310),
	.w1(32'hbb5fedaa),
	.w2(32'hbae7146e),
	.w3(32'h3a6c575d),
	.w4(32'hb9b9083e),
	.w5(32'h3a88f08d),
	.w6(32'h3b7807a1),
	.w7(32'h3b2d9a4e),
	.w8(32'hbaaf0271),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd6ef4),
	.w1(32'hbaae4cf0),
	.w2(32'hb73828da),
	.w3(32'hbaa96e06),
	.w4(32'hbb2651c6),
	.w5(32'hb9bf991c),
	.w6(32'hbabde352),
	.w7(32'hbaacb6d5),
	.w8(32'hb9b8c821),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27effe),
	.w1(32'h3a1be971),
	.w2(32'hbae54f9e),
	.w3(32'hba36831b),
	.w4(32'hbb3eadc8),
	.w5(32'hba9c35ea),
	.w6(32'hba75df7d),
	.w7(32'hbaae0dda),
	.w8(32'h3b2c1c0f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba344a91),
	.w1(32'hbb10ef3b),
	.w2(32'hbb1c24ea),
	.w3(32'hb8480364),
	.w4(32'hba92352f),
	.w5(32'h3b80eadd),
	.w6(32'h3b7905f8),
	.w7(32'h3b6559b3),
	.w8(32'h39897c62),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c47c),
	.w1(32'hbac6274c),
	.w2(32'h3a908b62),
	.w3(32'h3b6a6616),
	.w4(32'h3ba01770),
	.w5(32'h3b047820),
	.w6(32'hbb00e3ca),
	.w7(32'hbb42a913),
	.w8(32'hbbda9993),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dd513),
	.w1(32'h39bed12b),
	.w2(32'h3ba258ff),
	.w3(32'hba71868c),
	.w4(32'h3b3a25ef),
	.w5(32'hbbae2381),
	.w6(32'hbb572313),
	.w7(32'hba4579b1),
	.w8(32'h395a4bba),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977e01),
	.w1(32'hbb981813),
	.w2(32'hbbdfcdda),
	.w3(32'hbbb1df28),
	.w4(32'hbbb89cd4),
	.w5(32'hbbc8535d),
	.w6(32'hbbc17831),
	.w7(32'hbc0e2052),
	.w8(32'hbc14c989),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770b01),
	.w1(32'h3bc1fa65),
	.w2(32'h3c20e5e3),
	.w3(32'h3b9bd7e5),
	.w4(32'h3c3b5a45),
	.w5(32'h3c548237),
	.w6(32'h3b5bd42b),
	.w7(32'h3bad793b),
	.w8(32'h3c30de2c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b879403),
	.w1(32'h3a53f3ac),
	.w2(32'h3a8a79f7),
	.w3(32'h3b61e629),
	.w4(32'h3b1116d7),
	.w5(32'hb9937900),
	.w6(32'h3a105732),
	.w7(32'h3b52a7b6),
	.w8(32'hbb070091),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac88fb8),
	.w1(32'hbaba80ba),
	.w2(32'h39434bc7),
	.w3(32'hbadbc486),
	.w4(32'hbb2a8ed5),
	.w5(32'h3bfec024),
	.w6(32'hbb12faeb),
	.w7(32'h3a906f87),
	.w8(32'h3c06fc2a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a4fba),
	.w1(32'h3c3de80b),
	.w2(32'h3c1ad37c),
	.w3(32'h3b682e2e),
	.w4(32'h3a3c0831),
	.w5(32'hba7e6a4b),
	.w6(32'h3c3552fb),
	.w7(32'h3c021a2b),
	.w8(32'hbb08f9bc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e4ec),
	.w1(32'hbb21fb3f),
	.w2(32'hbb82c832),
	.w3(32'h39687cc5),
	.w4(32'hba42ded0),
	.w5(32'h3ba0852e),
	.w6(32'h396c87bb),
	.w7(32'hbb5125b0),
	.w8(32'h3b17116a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb49e40),
	.w1(32'h3b0051ae),
	.w2(32'h3a3ccf25),
	.w3(32'h3b7f38aa),
	.w4(32'h3b466f67),
	.w5(32'h3b28c086),
	.w6(32'h3b8ba3fd),
	.w7(32'hb9781d73),
	.w8(32'h3b93e16f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0def79),
	.w1(32'hbbc939ac),
	.w2(32'hbb3e8d5b),
	.w3(32'hbb229b6f),
	.w4(32'hbb4ee713),
	.w5(32'hbb9d1544),
	.w6(32'hbb132912),
	.w7(32'hbac62aa0),
	.w8(32'hbbb3090e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9f0df),
	.w1(32'hbbc9f28d),
	.w2(32'hbc24ac76),
	.w3(32'hbbcf0ae3),
	.w4(32'hbc4d410a),
	.w5(32'hbbe69eff),
	.w6(32'hbbf02ef0),
	.w7(32'hbbcce5c8),
	.w8(32'hbbacb3ec),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a838ba4),
	.w1(32'h3b3d7dde),
	.w2(32'h3b9f86cb),
	.w3(32'h3b536ac6),
	.w4(32'h3b51ee8f),
	.w5(32'h3920478e),
	.w6(32'h3b239f09),
	.w7(32'h3b7af725),
	.w8(32'h397d7b75),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44c233),
	.w1(32'hbb90f602),
	.w2(32'hbae25faa),
	.w3(32'hbb72b7cc),
	.w4(32'hbb64e010),
	.w5(32'hbb6fd263),
	.w6(32'hbb51b354),
	.w7(32'hbb92328d),
	.w8(32'hbbfa709f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5996ac),
	.w1(32'hbb879b89),
	.w2(32'hbb293452),
	.w3(32'hbb215dd7),
	.w4(32'hb8e7f8ce),
	.w5(32'hbad4eaa0),
	.w6(32'hbbbc3011),
	.w7(32'hbb6fcd73),
	.w8(32'hbbe1b2a4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb5fc5),
	.w1(32'hbc161783),
	.w2(32'hbbe6ef96),
	.w3(32'hbbc2791a),
	.w4(32'hbb2ef51b),
	.w5(32'h3aebf1e9),
	.w6(32'hbc10c27a),
	.w7(32'hbb89db07),
	.w8(32'h3aebe5f7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa9f41),
	.w1(32'hbb901c2b),
	.w2(32'hbb950f07),
	.w3(32'hbb52406b),
	.w4(32'hbb198282),
	.w5(32'hbb5fe3f5),
	.w6(32'hbb8b0340),
	.w7(32'hbb940b20),
	.w8(32'hbb5ac99f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a9c18),
	.w1(32'h38977798),
	.w2(32'hbb4509f0),
	.w3(32'hba9f0350),
	.w4(32'hbb23d333),
	.w5(32'hb7b8d3e0),
	.w6(32'h3a5240ce),
	.w7(32'hbac10dd4),
	.w8(32'hbb346acc),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925aca),
	.w1(32'hbb7e90c5),
	.w2(32'hbb034d86),
	.w3(32'hbb09fd3c),
	.w4(32'hbb605db3),
	.w5(32'hb99063eb),
	.w6(32'hbb139d3c),
	.w7(32'hbb1e1f5c),
	.w8(32'hba724ae9),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07b6a3),
	.w1(32'hbb190d5b),
	.w2(32'hbb86d03b),
	.w3(32'hba978f70),
	.w4(32'hba9e6832),
	.w5(32'hbb3b19ba),
	.w6(32'h3988822a),
	.w7(32'hba163944),
	.w8(32'hb8312481),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac64c65),
	.w1(32'hbabc1df6),
	.w2(32'h3b9047b9),
	.w3(32'hb944ef8d),
	.w4(32'h3a931180),
	.w5(32'h3924ebe2),
	.w6(32'h3a8ab44d),
	.w7(32'h3b35df09),
	.w8(32'hbb0e6ff9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ce07),
	.w1(32'h3c041e9e),
	.w2(32'h3ba61f53),
	.w3(32'h3b853ba4),
	.w4(32'h3b4ed5cc),
	.w5(32'h3af2bc56),
	.w6(32'hbb15a69f),
	.w7(32'h3a42aef9),
	.w8(32'h3be64410),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afed96b),
	.w1(32'hb99a4c87),
	.w2(32'hbaaf66ec),
	.w3(32'hbae2448d),
	.w4(32'hbabb197c),
	.w5(32'hb8f646f7),
	.w6(32'h3b7f650c),
	.w7(32'h3b17660c),
	.w8(32'hbb29ee0f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31913a),
	.w1(32'h3954d689),
	.w2(32'hbaeec26c),
	.w3(32'h3a7ec43a),
	.w4(32'h3ab293c5),
	.w5(32'hbadc11ad),
	.w6(32'hb8de3a41),
	.w7(32'h3a70f62a),
	.w8(32'h3aa7f832),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f04c5),
	.w1(32'hbc28b7a2),
	.w2(32'hbbf830de),
	.w3(32'hbbfadd8f),
	.w4(32'hbc6b8d7e),
	.w5(32'hbc49adbd),
	.w6(32'hbc471e17),
	.w7(32'hbc3cc3dd),
	.w8(32'hbc2e04de),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375d0b70),
	.w1(32'h3b957bac),
	.w2(32'h3b51073a),
	.w3(32'h3b9b3aa9),
	.w4(32'h3b1c70d8),
	.w5(32'h3a029118),
	.w6(32'h3b07a05e),
	.w7(32'hb9ebfd33),
	.w8(32'h3998ef5a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985fac9),
	.w1(32'hbb45e03f),
	.w2(32'hbb98e965),
	.w3(32'hbaaab041),
	.w4(32'hb99dc672),
	.w5(32'h3ad00072),
	.w6(32'hbb7c89a0),
	.w7(32'hbb4d1671),
	.w8(32'hba95c17e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01020f),
	.w1(32'h3bcbc2d3),
	.w2(32'h3b197568),
	.w3(32'h3b502eb4),
	.w4(32'h3aa2bebe),
	.w5(32'h38cfb00c),
	.w6(32'hbb866d91),
	.w7(32'hbab27971),
	.w8(32'h3c22c5fa),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae265f),
	.w1(32'hbbe61e5f),
	.w2(32'hbba1e16c),
	.w3(32'hbb832a4f),
	.w4(32'hbba91fb9),
	.w5(32'h3aff01bf),
	.w6(32'h3bedc6bc),
	.w7(32'h3abee9a0),
	.w8(32'h3b2f04a6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb94f02),
	.w1(32'h3b8b2aff),
	.w2(32'h3ba82e96),
	.w3(32'h3c1c791c),
	.w4(32'h3b712f6f),
	.w5(32'h3c2e79ca),
	.w6(32'h3bba83af),
	.w7(32'h39f08f6e),
	.w8(32'h3c4a86c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9fec5),
	.w1(32'h3bbfca9c),
	.w2(32'h3c024db1),
	.w3(32'h3c0cc3a0),
	.w4(32'h3c351c02),
	.w5(32'hb964e1f1),
	.w6(32'h3c72e7eb),
	.w7(32'h3c430e47),
	.w8(32'hba9310a9),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41cc42),
	.w1(32'hbb14db27),
	.w2(32'hbb05262d),
	.w3(32'hbb872770),
	.w4(32'hbb91692c),
	.w5(32'h3baf23c6),
	.w6(32'hbae1693b),
	.w7(32'hbb86d0f4),
	.w8(32'h3bb47cce),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3671eb),
	.w1(32'hbaef9fca),
	.w2(32'hba8ae55f),
	.w3(32'h3c03a0dd),
	.w4(32'h3b9a2ee2),
	.w5(32'hbaafa4ec),
	.w6(32'h3bbdfb97),
	.w7(32'h3ba765dd),
	.w8(32'hbb3374ef),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a33dd8),
	.w1(32'hbac66f14),
	.w2(32'h3a5fcc2d),
	.w3(32'h38fdfc90),
	.w4(32'h3b343aef),
	.w5(32'h3b3608f1),
	.w6(32'hb727cac8),
	.w7(32'hb93a8877),
	.w8(32'hbb87e50e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab15a42),
	.w1(32'hbbf2beb2),
	.w2(32'hbc2486dc),
	.w3(32'hbbf39133),
	.w4(32'hbbce2e6d),
	.w5(32'hbbc12a4d),
	.w6(32'hbc01d61c),
	.w7(32'hbb9661b2),
	.w8(32'hbb97dc08),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990229f),
	.w1(32'h3bcf199b),
	.w2(32'h3bc533c3),
	.w3(32'h3bd92e23),
	.w4(32'h3c0d2f7a),
	.w5(32'h3c12b2bd),
	.w6(32'h3b6ce79c),
	.w7(32'h3ba8b920),
	.w8(32'h3b973dd6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa8cf),
	.w1(32'h3b1707f6),
	.w2(32'h3b6f7b14),
	.w3(32'h3b9dc6dc),
	.w4(32'h3b8e8791),
	.w5(32'h3bbb0c88),
	.w6(32'h3b8d0829),
	.w7(32'h3b420e4f),
	.w8(32'h3ba21651),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c93d8f),
	.w1(32'hbb832f74),
	.w2(32'hbb834947),
	.w3(32'hbb1e39de),
	.w4(32'h3ae0a44f),
	.w5(32'hbb09de9e),
	.w6(32'hbb3af913),
	.w7(32'h3933e4c6),
	.w8(32'hbbd4237e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb592717),
	.w1(32'hbb13889f),
	.w2(32'hba59f2d7),
	.w3(32'hbb1e47a2),
	.w4(32'hb8feec72),
	.w5(32'h3afbad3b),
	.w6(32'hbba9bef2),
	.w7(32'hbb1c14e5),
	.w8(32'h3a6612f7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5b30),
	.w1(32'hbc4098fb),
	.w2(32'hbc8c99d8),
	.w3(32'hbc38714f),
	.w4(32'hbc321c9e),
	.w5(32'hbc394c36),
	.w6(32'hbc3a38d8),
	.w7(32'hbba9c27f),
	.w8(32'hbc0e0528),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60fc14),
	.w1(32'h38ed9011),
	.w2(32'hba73c396),
	.w3(32'hba9f873a),
	.w4(32'h3a88f199),
	.w5(32'hba04b738),
	.w6(32'hba9d50f9),
	.w7(32'h3b1d056f),
	.w8(32'h3989f4db),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5710bf),
	.w1(32'hba1029a3),
	.w2(32'hba8027b0),
	.w3(32'hba077396),
	.w4(32'hba1dc459),
	.w5(32'h38c86cfa),
	.w6(32'hbb10316c),
	.w7(32'hba9cc3b6),
	.w8(32'h38de31fc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd7fee),
	.w1(32'h3a101982),
	.w2(32'h39aa3ec8),
	.w3(32'h38a0bfc0),
	.w4(32'h3a7c1ecc),
	.w5(32'h39d7a3a7),
	.w6(32'hb984fe4b),
	.w7(32'hba15ad45),
	.w8(32'hb88d6545),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ce22e),
	.w1(32'h3aa6f09d),
	.w2(32'h3b5c467f),
	.w3(32'h3a93fc4d),
	.w4(32'h3b403b79),
	.w5(32'h3b231731),
	.w6(32'h3a2bf532),
	.w7(32'h3ae6c857),
	.w8(32'h3a998ab0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd2ec7),
	.w1(32'h3afe17f8),
	.w2(32'h3b90affd),
	.w3(32'h3b668cd2),
	.w4(32'h3b6d5379),
	.w5(32'h3ba1fcb8),
	.w6(32'h3bb3691b),
	.w7(32'h3b897f55),
	.w8(32'h3b93cb5e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebba96),
	.w1(32'h39ad4ff5),
	.w2(32'h39b4896d),
	.w3(32'h3b361a86),
	.w4(32'h39b9403e),
	.w5(32'h39789e18),
	.w6(32'h3b17ef18),
	.w7(32'hbacdc03d),
	.w8(32'hba12c25b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821af1),
	.w1(32'hb4342880),
	.w2(32'hba509cd6),
	.w3(32'h39cecbee),
	.w4(32'hba3aeb7d),
	.w5(32'h3a1173d7),
	.w6(32'hb941ecdc),
	.w7(32'hbaf081df),
	.w8(32'hb9e1852a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac283fa),
	.w1(32'h39d1039d),
	.w2(32'h3b103fe5),
	.w3(32'hbb077fe1),
	.w4(32'h3a2e2df5),
	.w5(32'hba06b713),
	.w6(32'h3a6bdf08),
	.w7(32'h3bb6c6e3),
	.w8(32'h3b9da520),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06a17),
	.w1(32'hbb3b04bd),
	.w2(32'hbb11d621),
	.w3(32'hbb5cffbd),
	.w4(32'hbb228a8d),
	.w5(32'hbb587de5),
	.w6(32'hbb52125b),
	.w7(32'hbba42b4e),
	.w8(32'hbb3b0275),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77325f),
	.w1(32'h3a42d3d9),
	.w2(32'h3b59a79d),
	.w3(32'h39994e06),
	.w4(32'h3b0afac5),
	.w5(32'h3b1e9ebf),
	.w6(32'h3b335fac),
	.w7(32'h3b6dfff3),
	.w8(32'h3ab0cc5d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b9906),
	.w1(32'hbad17797),
	.w2(32'hba7a4c5c),
	.w3(32'hb9e0550d),
	.w4(32'hba89098e),
	.w5(32'h3ab982a7),
	.w6(32'hbb16d038),
	.w7(32'hbac0c195),
	.w8(32'h3a839e8d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab451fc),
	.w1(32'h3a9db140),
	.w2(32'h3a032f64),
	.w3(32'h3aa7b8be),
	.w4(32'h3abf918d),
	.w5(32'h38e39f0d),
	.w6(32'h3a31a527),
	.w7(32'h3a2bb9c4),
	.w8(32'hb88d130b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e759af),
	.w1(32'hbaa4ac04),
	.w2(32'hbaaec4d6),
	.w3(32'hbac432a0),
	.w4(32'hb8838549),
	.w5(32'h3707e92c),
	.w6(32'h39d69c37),
	.w7(32'h3a10468b),
	.w8(32'hb8fea397),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a6feb),
	.w1(32'hbad2fc20),
	.w2(32'hba384c9e),
	.w3(32'hbaa83306),
	.w4(32'hb9d3c5af),
	.w5(32'hbb0951fe),
	.w6(32'hbaefe725),
	.w7(32'hb91328f1),
	.w8(32'hbb4bf1c8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dbd7d),
	.w1(32'hba808c35),
	.w2(32'h3b1cc6e0),
	.w3(32'hbaae0253),
	.w4(32'hba340dce),
	.w5(32'h3b775050),
	.w6(32'h39bfd65a),
	.w7(32'hba0579c7),
	.w8(32'h3b943792),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b5ae9),
	.w1(32'hba16967b),
	.w2(32'hba7a5e22),
	.w3(32'h39f046fe),
	.w4(32'hba786f06),
	.w5(32'hba1ea3cd),
	.w6(32'hb984dc0b),
	.w7(32'hb97fb296),
	.w8(32'hba2e31b3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae125f0),
	.w1(32'hbb6506d1),
	.w2(32'hbb2c3335),
	.w3(32'hbb1eef00),
	.w4(32'hbb148813),
	.w5(32'hbaaea541),
	.w6(32'hbb0b3fa3),
	.w7(32'hbb1e0619),
	.w8(32'hbb12c46a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf7a9f),
	.w1(32'h3b7501e1),
	.w2(32'h3ba58dba),
	.w3(32'h3b7f4ca7),
	.w4(32'h3b3c6542),
	.w5(32'h3b1ca48b),
	.w6(32'h3b869147),
	.w7(32'h39ff0ff3),
	.w8(32'hb99e5ace),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb927027d),
	.w1(32'h39f0c9c2),
	.w2(32'hbace193b),
	.w3(32'hba20916f),
	.w4(32'hba922507),
	.w5(32'h3a51112b),
	.w6(32'hba0f0a6c),
	.w7(32'hbb041031),
	.w8(32'h39cf157c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38380f81),
	.w1(32'h3a675836),
	.w2(32'h3aa8d2e9),
	.w3(32'h3a77b0e9),
	.w4(32'h3a1cce4c),
	.w5(32'hb91fecee),
	.w6(32'h3aa1b02c),
	.w7(32'h394ed637),
	.w8(32'h38eef326),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf47e5),
	.w1(32'h398ecc45),
	.w2(32'hba05c7ae),
	.w3(32'hb8ff9fa9),
	.w4(32'hb95a75da),
	.w5(32'hb9e31817),
	.w6(32'hb9262dce),
	.w7(32'hba825b0b),
	.w8(32'hba35147d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df3f6c),
	.w1(32'h3a43b5a8),
	.w2(32'h3b007f19),
	.w3(32'h3a4bc736),
	.w4(32'h3abb60cd),
	.w5(32'h399a46b9),
	.w6(32'h3a6b5a83),
	.w7(32'h3ac72e93),
	.w8(32'h3a947e67),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4b936),
	.w1(32'hb73ccfa7),
	.w2(32'h39d030d4),
	.w3(32'hba0279b0),
	.w4(32'hbb218105),
	.w5(32'hbb9f5580),
	.w6(32'h3ad4b571),
	.w7(32'h38aef7be),
	.w8(32'h3a24c9c4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0263a),
	.w1(32'hba9e8c0c),
	.w2(32'h39a9e646),
	.w3(32'hbb3997a9),
	.w4(32'hbb13ed78),
	.w5(32'h3a327b0f),
	.w6(32'hba3f78f2),
	.w7(32'hbafe1d10),
	.w8(32'hb9f11b31),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bad0cf),
	.w1(32'hba52cf13),
	.w2(32'h3972543c),
	.w3(32'hba3be28d),
	.w4(32'hba8337dd),
	.w5(32'hba1414c7),
	.w6(32'hb9945a77),
	.w7(32'hb964329c),
	.w8(32'hbaa6ae21),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37077e),
	.w1(32'hbab9555f),
	.w2(32'hba0b9b90),
	.w3(32'hba011ba5),
	.w4(32'hbb00419f),
	.w5(32'h393f3677),
	.w6(32'hbaf1aaaa),
	.w7(32'hbaace818),
	.w8(32'h3a466329),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99baf0),
	.w1(32'h3aa955b2),
	.w2(32'h3b108780),
	.w3(32'h3ab76d77),
	.w4(32'h3ae20161),
	.w5(32'h39afdbb7),
	.w6(32'h3b1190e5),
	.w7(32'h3adc54a3),
	.w8(32'hb8cea808),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a09a6a),
	.w1(32'h3a2e9e0c),
	.w2(32'h3aad3be3),
	.w3(32'h3a3dda96),
	.w4(32'h3ad7a944),
	.w5(32'hb99a193a),
	.w6(32'hb8787a01),
	.w7(32'h39d92d32),
	.w8(32'h3851e5e2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9398e4),
	.w1(32'h39220823),
	.w2(32'h3b113113),
	.w3(32'h39fc2e9c),
	.w4(32'h3b267d38),
	.w5(32'h3b1201ab),
	.w6(32'h3ad0a571),
	.w7(32'h3a32df88),
	.w8(32'h3a193e24),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8e6cb),
	.w1(32'hbbd50fa4),
	.w2(32'hbba2a7e0),
	.w3(32'hbbacb7cb),
	.w4(32'hbb55e8ae),
	.w5(32'hbb2defad),
	.w6(32'hbbb27e0e),
	.w7(32'hbbc5709c),
	.w8(32'hbbd12f9f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a381da1),
	.w1(32'h38633979),
	.w2(32'h392df817),
	.w3(32'h3b0880fa),
	.w4(32'h3b1eed5b),
	.w5(32'h3b518b3e),
	.w6(32'h3a6993b4),
	.w7(32'hb8d50fcc),
	.w8(32'h3b5d827e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e15970),
	.w1(32'hba731134),
	.w2(32'hb9d15a1d),
	.w3(32'hba0de794),
	.w4(32'h3a8582c3),
	.w5(32'hb9fc9ed3),
	.w6(32'hb97af1a7),
	.w7(32'hba0f5a95),
	.w8(32'hbabab3f8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166e20),
	.w1(32'hbb9a3b69),
	.w2(32'hbb4a824d),
	.w3(32'hbb869570),
	.w4(32'hbb5fe1f1),
	.w5(32'hbadc614e),
	.w6(32'hbb0dfcab),
	.w7(32'hbb073cc2),
	.w8(32'hbb6a09b3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabc768),
	.w1(32'h390cef0d),
	.w2(32'h3a9ad42d),
	.w3(32'hb9e1f50c),
	.w4(32'h38a95d4a),
	.w5(32'h3aa89cfe),
	.w6(32'hb9c2f7db),
	.w7(32'h3956b139),
	.w8(32'h3b59973c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398340bd),
	.w1(32'hba808426),
	.w2(32'h394d579b),
	.w3(32'hba53bcbd),
	.w4(32'hba4c2d69),
	.w5(32'hbaeb396a),
	.w6(32'hba8f520b),
	.w7(32'hbab51f76),
	.w8(32'hbb708ff8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb363f9d),
	.w1(32'hbb1ca023),
	.w2(32'hbb574f40),
	.w3(32'hbb10c2a4),
	.w4(32'hbb30f3d0),
	.w5(32'hb9526dce),
	.w6(32'hbb149b6d),
	.w7(32'hbb8100d1),
	.w8(32'hbad16080),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7db0f1),
	.w1(32'h3ab5720e),
	.w2(32'h3b60d085),
	.w3(32'h3bce3fbc),
	.w4(32'h3b832ad9),
	.w5(32'h3b8c8171),
	.w6(32'h3bae6d4c),
	.w7(32'h3b3a9e01),
	.w8(32'h3b6caaca),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1ea29),
	.w1(32'hba1a045b),
	.w2(32'hba84be24),
	.w3(32'hb914a06f),
	.w4(32'hb9f6cbff),
	.w5(32'h39f37210),
	.w6(32'hba2482a2),
	.w7(32'hba9b224f),
	.w8(32'hba144cdb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a71a3),
	.w1(32'h3a82a935),
	.w2(32'h3b1cf381),
	.w3(32'h3abe864b),
	.w4(32'h3af5f85e),
	.w5(32'h3aaacd11),
	.w6(32'h3b1f00f5),
	.w7(32'h3b08a764),
	.w8(32'h3af6358d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4122ac),
	.w1(32'h3acb52b8),
	.w2(32'h3ad16900),
	.w3(32'h3a70dab7),
	.w4(32'h3ab0491a),
	.w5(32'hbb1a0010),
	.w6(32'h3acf1bed),
	.w7(32'h3ac2dac0),
	.w8(32'hbabcdbd5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb242e),
	.w1(32'hba256c1e),
	.w2(32'hb9c2ea7f),
	.w3(32'hbad9fc11),
	.w4(32'hba333474),
	.w5(32'hb894773c),
	.w6(32'hba4e8684),
	.w7(32'hb9e65374),
	.w8(32'hba4ba2bc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39897d8d),
	.w1(32'h39170740),
	.w2(32'hb9399e7f),
	.w3(32'h3b2d1237),
	.w4(32'h3acb3219),
	.w5(32'h3a419c1f),
	.w6(32'h3a1f2668),
	.w7(32'h3a05390e),
	.w8(32'h3a4e084f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989a20d),
	.w1(32'h3a41232d),
	.w2(32'h3a0cad33),
	.w3(32'hbaa40a91),
	.w4(32'h38d51be5),
	.w5(32'h3ac7331c),
	.w6(32'h3ac70cb1),
	.w7(32'hb8d20877),
	.w8(32'h3a1f22e8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b7aed),
	.w1(32'h3a282a3b),
	.w2(32'h3ad1e3aa),
	.w3(32'h3af29886),
	.w4(32'h3ad8530c),
	.w5(32'h3b1ffda6),
	.w6(32'h3b06caea),
	.w7(32'h3b10a272),
	.w8(32'h3b1305cd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4656f4),
	.w1(32'h3b015dbe),
	.w2(32'h3b49710f),
	.w3(32'h3b382b0c),
	.w4(32'h3b4e8ca1),
	.w5(32'h3afbeaa7),
	.w6(32'h3a9bbbde),
	.w7(32'h3ad4da85),
	.w8(32'hb76b83c9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accea9c),
	.w1(32'h39abfe1d),
	.w2(32'h3a7cd666),
	.w3(32'h3af3c354),
	.w4(32'h3a47369a),
	.w5(32'h3ad9d4f1),
	.w6(32'h3ac4b545),
	.w7(32'h38bfaef5),
	.w8(32'h3a13b647),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d94af),
	.w1(32'hbb15ce55),
	.w2(32'hbbbf408b),
	.w3(32'hbb0bf899),
	.w4(32'hbb0059ab),
	.w5(32'hbb458b1c),
	.w6(32'hba3be551),
	.w7(32'hbaffa185),
	.w8(32'hbbd55357),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad168d7),
	.w1(32'h3abedb28),
	.w2(32'h3a84a113),
	.w3(32'h3b9c57e7),
	.w4(32'h3b2f753f),
	.w5(32'h3b8d8e15),
	.w6(32'h3b898209),
	.w7(32'hba7c0a72),
	.w8(32'h3b453a4b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b286bb5),
	.w1(32'h3b325fa0),
	.w2(32'h3b23a6f4),
	.w3(32'h3b5df8dc),
	.w4(32'h3b503e2f),
	.w5(32'h3afc6015),
	.w6(32'h3b8167dd),
	.w7(32'h3aeef5d5),
	.w8(32'h3a8c5d07),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6eb81),
	.w1(32'h3a31af60),
	.w2(32'h3ac621b7),
	.w3(32'h3b2af1eb),
	.w4(32'h3b3bc17a),
	.w5(32'h3b6c12ce),
	.w6(32'h3b0c3434),
	.w7(32'h3b0e0be0),
	.w8(32'h3b18febd),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ea6ee),
	.w1(32'hba1ef3c5),
	.w2(32'h39965033),
	.w3(32'hba446484),
	.w4(32'hb9565959),
	.w5(32'hbaaa8252),
	.w6(32'h3a08f1e2),
	.w7(32'h3a895f17),
	.w8(32'hbaf385ce),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9a116),
	.w1(32'h394b2119),
	.w2(32'h3aac0b50),
	.w3(32'h3ad7b7a6),
	.w4(32'h3b03d958),
	.w5(32'h3b1d9849),
	.w6(32'h3af9f012),
	.w7(32'hbac1a8b9),
	.w8(32'h3a2b3cd7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fc47a),
	.w1(32'h3abc1594),
	.w2(32'h3ac93811),
	.w3(32'h3a645314),
	.w4(32'h3a7b5853),
	.w5(32'h39879a86),
	.w6(32'h3ad9324a),
	.w7(32'h3a018ea0),
	.w8(32'h39b6963a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e8dd31),
	.w1(32'hbb561ff7),
	.w2(32'hbb5c2d64),
	.w3(32'hbb3bd9d7),
	.w4(32'hbac9cfbc),
	.w5(32'h38d31c6e),
	.w6(32'hbb20e52d),
	.w7(32'hb89acd7b),
	.w8(32'hba37a0c3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b8cbdb),
	.w1(32'h3aec44eb),
	.w2(32'h3a8057b0),
	.w3(32'h3ac25706),
	.w4(32'h3aa1740e),
	.w5(32'hb92286f8),
	.w6(32'h3a490355),
	.w7(32'h3a21ee94),
	.w8(32'h391bd65f),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb824de38),
	.w1(32'hbab6a783),
	.w2(32'hba2af44a),
	.w3(32'hbaa5ce60),
	.w4(32'hbabef12d),
	.w5(32'hbb04f6e4),
	.w6(32'hb8cfe678),
	.w7(32'hba85711d),
	.w8(32'hbb1c9403),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba543647),
	.w1(32'hb9b7080e),
	.w2(32'hba8285c8),
	.w3(32'hbaeafb4e),
	.w4(32'hbac89f4b),
	.w5(32'h39461abe),
	.w6(32'h38b7276d),
	.w7(32'hbaec41db),
	.w8(32'hbac47efb),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0f02),
	.w1(32'hba5c8f44),
	.w2(32'h3a501fbe),
	.w3(32'h3975cabe),
	.w4(32'h3a8c3edf),
	.w5(32'h3ad13a1e),
	.w6(32'h3a48fac4),
	.w7(32'h3a547d10),
	.w8(32'h3aaffb81),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24ab7e),
	.w1(32'hb821be0d),
	.w2(32'hbafa33a4),
	.w3(32'hba3f4dd5),
	.w4(32'hba8f195a),
	.w5(32'hb9df583d),
	.w6(32'hba9aa89d),
	.w7(32'hba298718),
	.w8(32'h37a7b6e4),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b946944),
	.w1(32'h3a8a10a1),
	.w2(32'h3a0db04a),
	.w3(32'h3b6f9d1e),
	.w4(32'h3a5c9196),
	.w5(32'hba918895),
	.w6(32'h3b650284),
	.w7(32'hb8cc7c2a),
	.w8(32'hbadb7c89),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd4bcc),
	.w1(32'h38b99a26),
	.w2(32'h368af6cb),
	.w3(32'h3a408926),
	.w4(32'h3a61ac40),
	.w5(32'hba3ff096),
	.w6(32'h3a11147e),
	.w7(32'h3a81eae7),
	.w8(32'hba088241),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa004a),
	.w1(32'h3a7350ed),
	.w2(32'hba87197c),
	.w3(32'hb99df787),
	.w4(32'hba972bfe),
	.w5(32'h3988c3e2),
	.w6(32'hb99552ac),
	.w7(32'hbaa4f083),
	.w8(32'h390f24eb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a56ae4),
	.w1(32'h3a2d78cc),
	.w2(32'h3aeeee4a),
	.w3(32'h3b68a1ba),
	.w4(32'h3b8096c3),
	.w5(32'h3b05c9ef),
	.w6(32'h3b431710),
	.w7(32'h3b6ecb85),
	.w8(32'h3aa67fa8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997bc6a),
	.w1(32'hbb1d388f),
	.w2(32'hbb3b5e2b),
	.w3(32'hbb846608),
	.w4(32'hbb9a55e4),
	.w5(32'hbb808543),
	.w6(32'hbbd9a924),
	.w7(32'hbb9e8c5a),
	.w8(32'hbb13c7f3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae310),
	.w1(32'h3ad451a4),
	.w2(32'h3ac72b83),
	.w3(32'h3ae981d2),
	.w4(32'h3adfb0f4),
	.w5(32'hb9c3f7d1),
	.w6(32'h3ad8f668),
	.w7(32'h3ad667fe),
	.w8(32'h3a46e8a3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954ead),
	.w1(32'h3b35b176),
	.w2(32'h3b47da52),
	.w3(32'h3b2aef49),
	.w4(32'h3b3f9f30),
	.w5(32'hb899ae0f),
	.w6(32'h3bc32d1c),
	.w7(32'h3b837b54),
	.w8(32'h3a80d75f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba815c3c),
	.w1(32'hbabe7f88),
	.w2(32'hbaf5e7c4),
	.w3(32'hbaf7f4ef),
	.w4(32'hbade9578),
	.w5(32'hbb2c268f),
	.w6(32'hbac0f73e),
	.w7(32'hbab80459),
	.w8(32'hbb58fc6b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7a4d3),
	.w1(32'hbb16e28d),
	.w2(32'hba879643),
	.w3(32'hbb1444c7),
	.w4(32'hba5a373e),
	.w5(32'hb98c8aa8),
	.w6(32'hba89f449),
	.w7(32'hbb0f4e74),
	.w8(32'hb92c7f79),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47849d),
	.w1(32'hbb1d25f0),
	.w2(32'hba8ae4ec),
	.w3(32'hba8d49e3),
	.w4(32'hba6fdcaf),
	.w5(32'hba8cff67),
	.w6(32'hbacbaa35),
	.w7(32'hba3e262e),
	.w8(32'hbb10772b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb8632),
	.w1(32'hbb744d75),
	.w2(32'hbb2af1e1),
	.w3(32'hbb8349a3),
	.w4(32'hbb73da4f),
	.w5(32'h3a99d469),
	.w6(32'hbb8a10df),
	.w7(32'hbb9f3037),
	.w8(32'h397ab075),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6def94),
	.w1(32'h3b3405a0),
	.w2(32'h3b223ab1),
	.w3(32'h3b47e21b),
	.w4(32'h3b648f2a),
	.w5(32'hbabfe167),
	.w6(32'h3b2e141a),
	.w7(32'h3b615487),
	.w8(32'hba6161b2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68ba43),
	.w1(32'hbb8cda47),
	.w2(32'hbb71c307),
	.w3(32'hbb36dd7f),
	.w4(32'hbb194e5d),
	.w5(32'h3b4fdfe9),
	.w6(32'hbabe5344),
	.w7(32'hbb315747),
	.w8(32'h3b00f90b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b440585),
	.w1(32'h3af3a766),
	.w2(32'h3b220b71),
	.w3(32'h3b3fc9d6),
	.w4(32'h3b54cc5f),
	.w5(32'h3a220ed1),
	.w6(32'h3ae3f115),
	.w7(32'h3b1d2f85),
	.w8(32'h391c23c7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d26a0),
	.w1(32'hb97bfa95),
	.w2(32'hb95955d3),
	.w3(32'h39861c3d),
	.w4(32'hb8d0019f),
	.w5(32'hb7e15449),
	.w6(32'hb97c3802),
	.w7(32'hba1ee75c),
	.w8(32'h3a92e443),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3893b4e7),
	.w1(32'hba53b551),
	.w2(32'h3a5c862e),
	.w3(32'hba31a85e),
	.w4(32'h3a8e925f),
	.w5(32'h387aab52),
	.w6(32'hb8240785),
	.w7(32'h3ae9422c),
	.w8(32'hb9486637),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219175),
	.w1(32'hbaee331e),
	.w2(32'hba0e0c0b),
	.w3(32'hba6a874f),
	.w4(32'hbab03e63),
	.w5(32'hba8cd741),
	.w6(32'hbab2dddd),
	.w7(32'hbb3d6731),
	.w8(32'hba724f27),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a30c8c),
	.w1(32'hba245757),
	.w2(32'h3ab07e40),
	.w3(32'h3a4fc629),
	.w4(32'hb9681cf9),
	.w5(32'hba80d91a),
	.w6(32'h3b34fb2c),
	.w7(32'h386014cd),
	.w8(32'hba3d9cbc),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391e3b19),
	.w1(32'hb826b894),
	.w2(32'hba3a0445),
	.w3(32'hb94c34a5),
	.w4(32'h37b7e2ee),
	.w5(32'hb9881168),
	.w6(32'h3986a284),
	.w7(32'h39af4446),
	.w8(32'hba9873c5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9199a5),
	.w1(32'hb9ad70aa),
	.w2(32'h3a7fb1ea),
	.w3(32'h3a40bcd7),
	.w4(32'h39b3e45a),
	.w5(32'h3ab2ece7),
	.w6(32'h3973fa6b),
	.w7(32'hba9afbda),
	.w8(32'h3a76d7ee),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125286),
	.w1(32'hba60aefd),
	.w2(32'h3a46e381),
	.w3(32'h3b69c34a),
	.w4(32'h3aea5995),
	.w5(32'h3a98fe39),
	.w6(32'h3b94527d),
	.w7(32'hba7628bc),
	.w8(32'hba234c55),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e79f80),
	.w1(32'hb86b2830),
	.w2(32'hba3ab446),
	.w3(32'hbb0a97d0),
	.w4(32'h3b0e97de),
	.w5(32'h3b78cd35),
	.w6(32'hbb30a62a),
	.w7(32'h3b0b55c0),
	.w8(32'h3b254b24),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9dea5),
	.w1(32'h3926b051),
	.w2(32'h3a32e0eb),
	.w3(32'h3a1d4ce3),
	.w4(32'h3ab82bbe),
	.w5(32'hba72a42a),
	.w6(32'h3a6c2998),
	.w7(32'h39c3af6c),
	.w8(32'hb819ce1a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5020b6),
	.w1(32'hbbb1b3a2),
	.w2(32'hbb3f0d62),
	.w3(32'hbb80f83f),
	.w4(32'hbb07c9af),
	.w5(32'hbb80b4c1),
	.w6(32'hbb797e54),
	.w7(32'hbb16477b),
	.w8(32'hbb39755d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe74e5),
	.w1(32'h3ac9f85a),
	.w2(32'h3b86b95b),
	.w3(32'h3ba6d244),
	.w4(32'h3bbb3df0),
	.w5(32'h3bdd8b6e),
	.w6(32'h3ba79ad3),
	.w7(32'h3a34fbac),
	.w8(32'h3a8911fb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7c966),
	.w1(32'h39a1cabc),
	.w2(32'hb7a54084),
	.w3(32'hb7945116),
	.w4(32'h392ce3d0),
	.w5(32'hba1d363d),
	.w6(32'h39e96e4f),
	.w7(32'h3a859555),
	.w8(32'hbb301374),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1023d),
	.w1(32'hbab5e609),
	.w2(32'hbab45d68),
	.w3(32'hb90a5cc2),
	.w4(32'hb9fd3220),
	.w5(32'hba09e133),
	.w6(32'hbac85fb6),
	.w7(32'hbae9533f),
	.w8(32'hbaec05cc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3ebcc),
	.w1(32'hbac57020),
	.w2(32'hba8d1ca9),
	.w3(32'hba41e0b4),
	.w4(32'hba4d31e8),
	.w5(32'h3891472a),
	.w6(32'h397df09c),
	.w7(32'hbab45674),
	.w8(32'hbab6b61a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93384d),
	.w1(32'hba731f0b),
	.w2(32'hbab5b970),
	.w3(32'h3980ad01),
	.w4(32'hba7f1b5a),
	.w5(32'hba1c2bf4),
	.w6(32'hb90d5dfc),
	.w7(32'hba8bc6e6),
	.w8(32'hb97b41f0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b293c37),
	.w1(32'h3ac1a094),
	.w2(32'h3a1d87a1),
	.w3(32'h39c9bff8),
	.w4(32'h3a9ada9a),
	.w5(32'h39b5ecf1),
	.w6(32'hb9ead342),
	.w7(32'h399275f0),
	.w8(32'hba87e228),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f9ba0),
	.w1(32'hba99d604),
	.w2(32'hba9c6baf),
	.w3(32'h3aa43aeb),
	.w4(32'h39bec066),
	.w5(32'hbb7f433f),
	.w6(32'hb8e9b6ee),
	.w7(32'hbb1b72ff),
	.w8(32'hbb9efc5f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13e40b),
	.w1(32'hb9a884e0),
	.w2(32'h3a71bfcd),
	.w3(32'hba011433),
	.w4(32'h3adec6e4),
	.w5(32'h3b7dfdfb),
	.w6(32'h3a932cde),
	.w7(32'h3ac86f19),
	.w8(32'h3b639b62),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a6c08),
	.w1(32'hb9cca536),
	.w2(32'h39b05a3f),
	.w3(32'h39ae9988),
	.w4(32'hba97ff6f),
	.w5(32'hbb09bbc7),
	.w6(32'h38cd98b1),
	.w7(32'hba2000c4),
	.w8(32'hbac8306a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87a60a),
	.w1(32'hba360e8a),
	.w2(32'hb92d994d),
	.w3(32'hbaf05f74),
	.w4(32'h39344649),
	.w5(32'hba15a3b5),
	.w6(32'hb9cf5908),
	.w7(32'h39c687ef),
	.w8(32'hba875ab3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f621b6),
	.w1(32'h37ce262d),
	.w2(32'h3a2a2cbf),
	.w3(32'h3a766992),
	.w4(32'h3a8ca1fd),
	.w5(32'h39ae8ca3),
	.w6(32'h3a0dc3b6),
	.w7(32'h3b336e36),
	.w8(32'h3a143ca2),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebbed5),
	.w1(32'hba8d749e),
	.w2(32'hba992913),
	.w3(32'hbaa7b093),
	.w4(32'hba526ced),
	.w5(32'hb997d51d),
	.w6(32'hbadf5d2f),
	.w7(32'h3958ab52),
	.w8(32'hba4a406d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae254e2),
	.w1(32'hbacd233c),
	.w2(32'hbab86506),
	.w3(32'hbb21f162),
	.w4(32'hbb0e705e),
	.w5(32'hbb3f353d),
	.w6(32'hbb0af4c0),
	.w7(32'h3a6d734f),
	.w8(32'hbb15f4a3),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd171d),
	.w1(32'hbab30b11),
	.w2(32'hbaeea901),
	.w3(32'hbb351527),
	.w4(32'hbb70da26),
	.w5(32'hb8a3d50a),
	.w6(32'hba6819bb),
	.w7(32'hbb1ce986),
	.w8(32'h39da793d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80ed29),
	.w1(32'hb848fa59),
	.w2(32'h3a3c262e),
	.w3(32'hb95902be),
	.w4(32'h39f6833f),
	.w5(32'hbb873c7b),
	.w6(32'h3a84c39e),
	.w7(32'h39900098),
	.w8(32'hbb9cb64e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39e4a),
	.w1(32'hb990ccfe),
	.w2(32'hb98218c2),
	.w3(32'h3a742199),
	.w4(32'hb95d6782),
	.w5(32'h3b857d0f),
	.w6(32'h3850ec9d),
	.w7(32'hbb0aaf45),
	.w8(32'h3b228b76),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27a7a4),
	.w1(32'h3a16631a),
	.w2(32'h3aec888b),
	.w3(32'h3adbdd95),
	.w4(32'h3aa99612),
	.w5(32'h3905472b),
	.w6(32'h3acbb70d),
	.w7(32'h3a6b4793),
	.w8(32'h3a6a3fdc),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c1fca),
	.w1(32'hba25afe0),
	.w2(32'hb9c92f3c),
	.w3(32'hbab23e85),
	.w4(32'h390fb1dc),
	.w5(32'hba2f94b9),
	.w6(32'hba7cf93c),
	.w7(32'h37b3a987),
	.w8(32'hba32f0cc),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a0413),
	.w1(32'h39eeef6e),
	.w2(32'h3b28fe4f),
	.w3(32'h3b396b8b),
	.w4(32'h3b5392a6),
	.w5(32'h3b6a9dfc),
	.w6(32'h3b03ee8d),
	.w7(32'h3ae9b9f3),
	.w8(32'h3b9685ce),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87d8a4),
	.w1(32'hbaba4529),
	.w2(32'h39e9d047),
	.w3(32'hbb0104b2),
	.w4(32'hba927472),
	.w5(32'hb9c040f8),
	.w6(32'hba2cd58f),
	.w7(32'hb8b4e799),
	.w8(32'hba77a708),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b7a97),
	.w1(32'h390fff8b),
	.w2(32'h3b084124),
	.w3(32'hbaebb287),
	.w4(32'h38043e3a),
	.w5(32'hba6b9f17),
	.w6(32'hbacafbfd),
	.w7(32'hb9d8a05e),
	.w8(32'hba0fce2b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae90ce7),
	.w1(32'hbaee368f),
	.w2(32'hbb0f8efc),
	.w3(32'hbb1ab7d1),
	.w4(32'hbaf060cb),
	.w5(32'h393626db),
	.w6(32'hba898151),
	.w7(32'hbace9039),
	.w8(32'hba162a60),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba110d24),
	.w1(32'hba5feb70),
	.w2(32'hbabf12ac),
	.w3(32'hb9d455e4),
	.w4(32'hba705e02),
	.w5(32'hba8c7088),
	.w6(32'hba9add69),
	.w7(32'hbac6c208),
	.w8(32'hbae43970),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9220e57),
	.w1(32'h3acb0c76),
	.w2(32'h3b6adf44),
	.w3(32'h3b0ff805),
	.w4(32'h3b075d7d),
	.w5(32'hb9d4e5bc),
	.w6(32'h3a8c2315),
	.w7(32'h3b31118f),
	.w8(32'h3b1f1ea6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7d0c6),
	.w1(32'hbb8dd0e7),
	.w2(32'hbb7e5056),
	.w3(32'hbb0f6a5d),
	.w4(32'hbb252abb),
	.w5(32'hbb389f77),
	.w6(32'hbbbe69a9),
	.w7(32'hbb99bee2),
	.w8(32'hbb28841d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21a98a),
	.w1(32'h3a253273),
	.w2(32'h3b5cebe2),
	.w3(32'h3aa516d6),
	.w4(32'h3b073806),
	.w5(32'h3b4c113a),
	.w6(32'h3ade4c08),
	.w7(32'h3b0c3c92),
	.w8(32'h3b4265cc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c0010),
	.w1(32'hbabe87cf),
	.w2(32'hb9e7f09d),
	.w3(32'h3a78f444),
	.w4(32'h3ba2c280),
	.w5(32'h3b6cc96b),
	.w6(32'h3a68b707),
	.w7(32'h3a928e6b),
	.w8(32'hbb275779),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8701d4),
	.w1(32'h3905960d),
	.w2(32'h39c756b1),
	.w3(32'hb996cd0a),
	.w4(32'h392373db),
	.w5(32'h3a09c1e3),
	.w6(32'hb94dc4b7),
	.w7(32'hb9c25956),
	.w8(32'h39c73739),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c212ff),
	.w1(32'hba6308af),
	.w2(32'hb8fb41d5),
	.w3(32'hb9e2dbd9),
	.w4(32'h399d9d7f),
	.w5(32'h3ac9c638),
	.w6(32'h38ce5867),
	.w7(32'hb952f393),
	.w8(32'h3a2e9d30),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe1771),
	.w1(32'h3b36dec4),
	.w2(32'hbb1e9e8b),
	.w3(32'hba853247),
	.w4(32'h3ab6b260),
	.w5(32'hbb01491e),
	.w6(32'hbb0b7c24),
	.w7(32'h3aa43821),
	.w8(32'hb985b0f6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e9f09),
	.w1(32'hbb6effc9),
	.w2(32'hbb16ea4a),
	.w3(32'hbb82871b),
	.w4(32'hbba1c2fb),
	.w5(32'hbb86562e),
	.w6(32'hba689d58),
	.w7(32'hbb44808d),
	.w8(32'hbb979917),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d448f),
	.w1(32'hbb0a3e75),
	.w2(32'hbb82e059),
	.w3(32'hbb33cb96),
	.w4(32'hbb111351),
	.w5(32'hbb4e90cd),
	.w6(32'hbbc722c2),
	.w7(32'hbb2374f3),
	.w8(32'hbb86b768),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae219e),
	.w1(32'h3b26e1ce),
	.w2(32'h3b32df42),
	.w3(32'h3acc2ad9),
	.w4(32'h3b24d35d),
	.w5(32'h3b930fc1),
	.w6(32'h3b6c1dbe),
	.w7(32'h3aca1af5),
	.w8(32'h3b80651e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906e589),
	.w1(32'h3ae777b3),
	.w2(32'h3b3d5f2a),
	.w3(32'h3b3cc67c),
	.w4(32'h3b48d6de),
	.w5(32'h3b59db59),
	.w6(32'h3b342cd6),
	.w7(32'h3ae6caff),
	.w8(32'h3abc6ba5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ee2bd),
	.w1(32'hba01c580),
	.w2(32'hb90b9a5d),
	.w3(32'hb8659de6),
	.w4(32'hba24d192),
	.w5(32'h3a39a50d),
	.w6(32'hb949787f),
	.w7(32'hb9027104),
	.w8(32'h3b02ec8d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4136a7),
	.w1(32'h3b0107bf),
	.w2(32'h3ae6d622),
	.w3(32'h3a642025),
	.w4(32'h3ae37f25),
	.w5(32'hb9a210f0),
	.w6(32'h3a84acba),
	.w7(32'h3ad811f7),
	.w8(32'hba69a5dd),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5da778),
	.w1(32'hb9ee9424),
	.w2(32'h3a91e4ce),
	.w3(32'hb98fbe4f),
	.w4(32'h3a60d019),
	.w5(32'h3b06bd0a),
	.w6(32'hbb07370b),
	.w7(32'hb9f18a05),
	.w8(32'h3b0753f3),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff5fc1),
	.w1(32'h3a523c61),
	.w2(32'hba0af52e),
	.w3(32'h3a8ab60f),
	.w4(32'hba2457e5),
	.w5(32'h3b208cdd),
	.w6(32'h3b0f8f1f),
	.w7(32'hb9a2563e),
	.w8(32'h3af6def9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287335),
	.w1(32'h3c0844c6),
	.w2(32'h3aeb49cf),
	.w3(32'h3bf4326b),
	.w4(32'h3aa44549),
	.w5(32'hbbcdf4d3),
	.w6(32'h3bd5825b),
	.w7(32'h3b6127c1),
	.w8(32'hbbefb3dc),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd110e),
	.w1(32'hbb8e0f97),
	.w2(32'hbb66ebcd),
	.w3(32'hbb032dbe),
	.w4(32'hb98e8f39),
	.w5(32'hbc2aed5c),
	.w6(32'hbafc5533),
	.w7(32'hbbb04c09),
	.w8(32'hbbf0e9ea),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f15b1),
	.w1(32'hbb339bd8),
	.w2(32'hbb8df57e),
	.w3(32'hbb3c395b),
	.w4(32'hbb59de66),
	.w5(32'h3b13a23b),
	.w6(32'hba81edb6),
	.w7(32'hba9a129c),
	.w8(32'h3b806b99),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17abcb),
	.w1(32'hbbaeca72),
	.w2(32'hbb7bfa68),
	.w3(32'hbaf73031),
	.w4(32'hbb484205),
	.w5(32'h3b0514f8),
	.w6(32'hbb83b0b4),
	.w7(32'hbbb9a238),
	.w8(32'h3acd53eb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b112871),
	.w1(32'hba6dbb9b),
	.w2(32'hbbccc520),
	.w3(32'hbb988c3c),
	.w4(32'hbb74f2ac),
	.w5(32'hbc0ac9e3),
	.w6(32'hbb8691a0),
	.w7(32'hbba6f769),
	.w8(32'hbc15a1ea),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75a04e),
	.w1(32'hbbdcdb96),
	.w2(32'hbb4a94d2),
	.w3(32'hbc0fda32),
	.w4(32'hbb9a1992),
	.w5(32'hbb7761e9),
	.w6(32'hbbb8cc4c),
	.w7(32'hbb350e6f),
	.w8(32'hba5c3d1c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87dcf47),
	.w1(32'hba00c785),
	.w2(32'h395afbab),
	.w3(32'hbb42915d),
	.w4(32'h39ea22c4),
	.w5(32'hb95714b4),
	.w6(32'h3aeb7bfe),
	.w7(32'h3adb756c),
	.w8(32'hbab6e0d4),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01679b),
	.w1(32'hbb9a03b7),
	.w2(32'hbb68ec1c),
	.w3(32'hbba692ed),
	.w4(32'hbb8b13be),
	.w5(32'h3a45d0e4),
	.w6(32'hbbaab384),
	.w7(32'hbb921e61),
	.w8(32'h3b48fff0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9b3d),
	.w1(32'hbbb6ff76),
	.w2(32'hbab3eae9),
	.w3(32'hbb9f1ef5),
	.w4(32'h3b089f09),
	.w5(32'h3b679fa2),
	.w6(32'hbb2f29dd),
	.w7(32'h39e908de),
	.w8(32'h3bdf714a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a877242),
	.w1(32'h3c182c47),
	.w2(32'h3b990372),
	.w3(32'h3c095770),
	.w4(32'h3bb2f8ef),
	.w5(32'h3ba535ba),
	.w6(32'h3c5fc168),
	.w7(32'h3bcf2aa4),
	.w8(32'h3b62f3f6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b944249),
	.w1(32'h3b86bdf1),
	.w2(32'h3ad46e9f),
	.w3(32'h3b0cf9dd),
	.w4(32'hbafbfbfd),
	.w5(32'h3bea6b2f),
	.w6(32'h39412447),
	.w7(32'h3a2ebd21),
	.w8(32'h3bce6908),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29611),
	.w1(32'h3c883a22),
	.w2(32'h3c513ff3),
	.w3(32'h3c96697c),
	.w4(32'h3c5b30ed),
	.w5(32'hbbf076b0),
	.w6(32'h3cae6202),
	.w7(32'h3c6ace07),
	.w8(32'hbb61399c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a445b),
	.w1(32'hb88aa61b),
	.w2(32'hbb0c72cf),
	.w3(32'hb893a93d),
	.w4(32'hbb65cb75),
	.w5(32'h3b90d81c),
	.w6(32'h3c0bfe98),
	.w7(32'hbace4d19),
	.w8(32'h3b821d37),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f69db),
	.w1(32'hbb101854),
	.w2(32'hbaecb538),
	.w3(32'h3af413a5),
	.w4(32'hb959fd93),
	.w5(32'h3b12f1db),
	.w6(32'hb8d82c45),
	.w7(32'hbb839d67),
	.w8(32'hb7eeb10e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fa4e0),
	.w1(32'h3b2a2e9f),
	.w2(32'hba94d878),
	.w3(32'h3b5814bf),
	.w4(32'hbaaa918f),
	.w5(32'hbb04420b),
	.w6(32'h3b6abd73),
	.w7(32'hbadbc1af),
	.w8(32'hbac7bc73),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf42c70),
	.w1(32'hbb4d3931),
	.w2(32'hbb0dd245),
	.w3(32'hbb606d7c),
	.w4(32'hbb2a53ba),
	.w5(32'h3a924305),
	.w6(32'hbb34d6ea),
	.w7(32'hbba9fbc1),
	.w8(32'h3b29078a),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa39c4),
	.w1(32'h3b804025),
	.w2(32'hbb262cdc),
	.w3(32'hbb406ddb),
	.w4(32'hbb0bd366),
	.w5(32'hba84995a),
	.w6(32'h3948d1a5),
	.w7(32'hbb5e1a12),
	.w8(32'hbaa26cff),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf82c2),
	.w1(32'h3aeee54a),
	.w2(32'hbb606663),
	.w3(32'h39f48424),
	.w4(32'hbae8f92f),
	.w5(32'h3914a346),
	.w6(32'h398f3bc7),
	.w7(32'hbb994e17),
	.w8(32'hbab2536b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbe6dd),
	.w1(32'h3bb27d11),
	.w2(32'h3c10e620),
	.w3(32'hbabb4373),
	.w4(32'h3ba76a39),
	.w5(32'hbb43dcfc),
	.w6(32'hb8cf9f98),
	.w7(32'h3bd1cc92),
	.w8(32'hba4274d3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85299c),
	.w1(32'hbb227df3),
	.w2(32'hbb6e793f),
	.w3(32'hbb36af00),
	.w4(32'hbb82d04c),
	.w5(32'hbbf921a1),
	.w6(32'hb9baa0cc),
	.w7(32'h39ffce05),
	.w8(32'hbb3f23bf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd378cd),
	.w1(32'hbade90c6),
	.w2(32'hbbc93f76),
	.w3(32'hbb7f10bf),
	.w4(32'hbc11bc95),
	.w5(32'h3afc8a6b),
	.w6(32'hba85a584),
	.w7(32'hbb704256),
	.w8(32'h3be15591),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc4760),
	.w1(32'h3c76c571),
	.w2(32'h3c0af156),
	.w3(32'h3c3f8444),
	.w4(32'h3bb613d0),
	.w5(32'hbb370198),
	.w6(32'h3c995957),
	.w7(32'h3c47bd07),
	.w8(32'hbb9a619b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e7788),
	.w1(32'hbb2084e0),
	.w2(32'hb947fc39),
	.w3(32'hbb64e6f2),
	.w4(32'h3b7b9e9a),
	.w5(32'hbb82fd00),
	.w6(32'hbbc35cc0),
	.w7(32'h3ac75b6b),
	.w8(32'hbbabbad7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa6ec8),
	.w1(32'hbbb763be),
	.w2(32'hba5646ae),
	.w3(32'hb9c97647),
	.w4(32'hbb24041f),
	.w5(32'h3c0a16c0),
	.w6(32'hbb4f5c2b),
	.w7(32'h3aea98fe),
	.w8(32'h3c63a353),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b352c5b),
	.w1(32'hbbf0d592),
	.w2(32'hbb8825cf),
	.w3(32'h3a81c0c1),
	.w4(32'hbb74de2d),
	.w5(32'hba2ae248),
	.w6(32'h3b3719b3),
	.w7(32'hbc0ab8f5),
	.w8(32'hbbf35865),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea1da1),
	.w1(32'hbb9b3808),
	.w2(32'hbb8e9377),
	.w3(32'hba1b3d5d),
	.w4(32'h3ac7a168),
	.w5(32'h3b027350),
	.w6(32'hbb3a8501),
	.w7(32'hbb33b895),
	.w8(32'h3c31641b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae13fcf),
	.w1(32'hbb755126),
	.w2(32'hbbe24589),
	.w3(32'hbb573cf7),
	.w4(32'hbb8e2768),
	.w5(32'hba8db695),
	.w6(32'hb95c9e46),
	.w7(32'hbc38720e),
	.w8(32'hb98c444a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91f4a0),
	.w1(32'hbb9a6e64),
	.w2(32'hbae5c70f),
	.w3(32'hbb4ba458),
	.w4(32'hbb875db3),
	.w5(32'hbb81fbda),
	.w6(32'hba892b2e),
	.w7(32'hbbcca7ae),
	.w8(32'hbae0acba),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8df83),
	.w1(32'hb93ea22e),
	.w2(32'hba80db45),
	.w3(32'h3a7c983e),
	.w4(32'h3a8c19ea),
	.w5(32'h3b558e4d),
	.w6(32'h3bf19716),
	.w7(32'h3a8568ef),
	.w8(32'h3bcf31db),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1586a4),
	.w1(32'hbbdf8a80),
	.w2(32'hba6240f8),
	.w3(32'hbbb79016),
	.w4(32'hbbbdc5b4),
	.w5(32'hbb9d4d2c),
	.w6(32'hbbd1e839),
	.w7(32'hb97e175b),
	.w8(32'hbb85b7e6),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule