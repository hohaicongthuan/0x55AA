module layer_8_featuremap_103(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3f4a2),
	.w1(32'h3b9c9a86),
	.w2(32'h3bc13dea),
	.w3(32'hb905f8b5),
	.w4(32'h3c4d455e),
	.w5(32'hbbfb7d91),
	.w6(32'h3ad33d5b),
	.w7(32'h3c1499a1),
	.w8(32'hbc3101be),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acff6),
	.w1(32'h3c547274),
	.w2(32'h3be382e7),
	.w3(32'h3b6a2d2a),
	.w4(32'hbaf5596e),
	.w5(32'h3941a30f),
	.w6(32'h3c35a44b),
	.w7(32'h3be4ea8b),
	.w8(32'h3d019fe7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c910037),
	.w1(32'hbc7af5ef),
	.w2(32'h3c79b661),
	.w3(32'hb9953519),
	.w4(32'hbcdbc6d0),
	.w5(32'h3c523848),
	.w6(32'h39fdc753),
	.w7(32'h3c133358),
	.w8(32'h3d41e84a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafddbf),
	.w1(32'hbc06a260),
	.w2(32'hb9950a1f),
	.w3(32'hbc9b9d52),
	.w4(32'h3be112fc),
	.w5(32'h3b085928),
	.w6(32'hbd0058b7),
	.w7(32'h3b1f3e3e),
	.w8(32'h3c02f22c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb8aad),
	.w1(32'hbc11fc9e),
	.w2(32'hbbb2fc1e),
	.w3(32'hbc8447a7),
	.w4(32'hbc00cd27),
	.w5(32'h392a1961),
	.w6(32'hbc0a1cf8),
	.w7(32'hb9dac2ea),
	.w8(32'hbcd6652d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f7b4),
	.w1(32'h3a170374),
	.w2(32'h3c7e6a97),
	.w3(32'hbad31911),
	.w4(32'h3993fc42),
	.w5(32'hbb2e3889),
	.w6(32'h3b90b21a),
	.w7(32'h3b1b6914),
	.w8(32'hbca20b40),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02f8cd),
	.w1(32'hbb8323d2),
	.w2(32'h3c384975),
	.w3(32'h3c8c1f50),
	.w4(32'hbb9027ee),
	.w5(32'h3c83b33e),
	.w6(32'h3a9aff92),
	.w7(32'h3c2c7456),
	.w8(32'hbc4de11a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4313dd),
	.w1(32'hbc17468f),
	.w2(32'hbc010173),
	.w3(32'h3ca40ddf),
	.w4(32'hbca15b2d),
	.w5(32'h3c10d76c),
	.w6(32'h3c780b4c),
	.w7(32'hbcc8ed68),
	.w8(32'h3a77a20f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b9c7f),
	.w1(32'h3c4bc1bb),
	.w2(32'h3ac12b46),
	.w3(32'h3c0781bf),
	.w4(32'h3bbc2823),
	.w5(32'hbc81271e),
	.w6(32'h3c8362b5),
	.w7(32'h3c6e24cd),
	.w8(32'hbc30e449),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d8809),
	.w1(32'h3c00b610),
	.w2(32'h3cc8e456),
	.w3(32'h3b863e3e),
	.w4(32'h3c5362f4),
	.w5(32'hbd5ac0fe),
	.w6(32'h3c80cb30),
	.w7(32'h3d3d12f4),
	.w8(32'hbd97d448),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd028ed),
	.w1(32'hbbc5a296),
	.w2(32'h3c4a5c93),
	.w3(32'h3cdca166),
	.w4(32'hbbc30cf6),
	.w5(32'h3bfb617b),
	.w6(32'h3be855b5),
	.w7(32'hbbf4e455),
	.w8(32'h3cafd98f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00aa28),
	.w1(32'hbc8510ad),
	.w2(32'hbc12589d),
	.w3(32'hbc92d590),
	.w4(32'hbc39cbe9),
	.w5(32'hbae311e1),
	.w6(32'hbc7de3ab),
	.w7(32'hbcbae618),
	.w8(32'hbc861dae),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f31d2),
	.w1(32'h3a59b735),
	.w2(32'h3c03f026),
	.w3(32'hbba9acb9),
	.w4(32'h3b5f2470),
	.w5(32'hbbe59113),
	.w6(32'h3b0e7d1c),
	.w7(32'h3c7ced0a),
	.w8(32'hbbf038a4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb422fd),
	.w1(32'hbada4580),
	.w2(32'hbb2ef282),
	.w3(32'hbb70a4c3),
	.w4(32'hba81565f),
	.w5(32'hba8395ee),
	.w6(32'hbb19eeb8),
	.w7(32'hba9717ab),
	.w8(32'hba1d41d2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ff1ef),
	.w1(32'hbb4c5b6e),
	.w2(32'hbb9c4544),
	.w3(32'h3a2d1930),
	.w4(32'hbb8fb35d),
	.w5(32'h3a12f587),
	.w6(32'hbb9aa42a),
	.w7(32'hbbb283e8),
	.w8(32'h3a7e32fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad69252),
	.w1(32'h39efb524),
	.w2(32'hbc9f7c8c),
	.w3(32'h3b062b24),
	.w4(32'h3b1a752e),
	.w5(32'hbc927894),
	.w6(32'hba5ee7b0),
	.w7(32'h3b289b13),
	.w8(32'hbc3d18be),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f2bf3),
	.w1(32'hbb029ffb),
	.w2(32'h3afe1c31),
	.w3(32'hbc845fbc),
	.w4(32'hbc1f4c47),
	.w5(32'hbd0ac7e5),
	.w6(32'hbc1cc9ac),
	.w7(32'h3cb3968b),
	.w8(32'hbcdc9baa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc333bf8),
	.w1(32'hbc0874c7),
	.w2(32'h3a892c5d),
	.w3(32'hba8ff90c),
	.w4(32'h3c185912),
	.w5(32'h3c9239fb),
	.w6(32'h3ab4a314),
	.w7(32'h3a445de4),
	.w8(32'h3b581152),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd22e5),
	.w1(32'h3a87e83d),
	.w2(32'hbb0be1c3),
	.w3(32'hbc13aec3),
	.w4(32'h3c554fe8),
	.w5(32'h3bc5157b),
	.w6(32'h3b697ed4),
	.w7(32'h3cae690d),
	.w8(32'hbc48510e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc47151),
	.w1(32'h3bc17873),
	.w2(32'hbc30ffec),
	.w3(32'h3bf422ed),
	.w4(32'h39ae14a6),
	.w5(32'hbbbfe1f0),
	.w6(32'h3c2f5845),
	.w7(32'h3bc108ce),
	.w8(32'hbba29d43),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba411d77),
	.w1(32'h3b609d0e),
	.w2(32'hbca7766f),
	.w3(32'hbbd15630),
	.w4(32'h3ac0f46e),
	.w5(32'hbbca8806),
	.w6(32'hbbcd6435),
	.w7(32'hbba9a270),
	.w8(32'h3bfea3ed),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0768a0),
	.w1(32'h3cccc94b),
	.w2(32'h3c852a75),
	.w3(32'h3c508bae),
	.w4(32'hbb9b4d15),
	.w5(32'h3c3666cf),
	.w6(32'h3cd11b07),
	.w7(32'h3c9498a6),
	.w8(32'h3cd362f2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceba84c),
	.w1(32'hbc51b5ef),
	.w2(32'hbca72464),
	.w3(32'hbd038988),
	.w4(32'hbc967ae6),
	.w5(32'hbce6f086),
	.w6(32'hbb68077f),
	.w7(32'hbd509e0e),
	.w8(32'hbcce3819),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc663316),
	.w1(32'hbc0deaa2),
	.w2(32'hba8e04d0),
	.w3(32'hbb8c252c),
	.w4(32'hbb18211a),
	.w5(32'hbc5aa64b),
	.w6(32'h3a8ab139),
	.w7(32'hbbb3a65f),
	.w8(32'hbbcab0fd),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce2c665),
	.w1(32'hbc95a650),
	.w2(32'hbcbb91c6),
	.w3(32'hbcc4b58a),
	.w4(32'hbbd3896c),
	.w5(32'hbc567081),
	.w6(32'hbc9abdf3),
	.w7(32'hbcca9ae0),
	.w8(32'hbc8b47c7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d5d6),
	.w1(32'hba19945a),
	.w2(32'hbb8d5b84),
	.w3(32'h3ac2fc02),
	.w4(32'h3c0693e3),
	.w5(32'hbb90ac3e),
	.w6(32'h3b9bb9db),
	.w7(32'h3c34a7dd),
	.w8(32'h3c22f83e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0397d5),
	.w1(32'hbb9ed9ae),
	.w2(32'h3c30a60d),
	.w3(32'hbb419360),
	.w4(32'h3c5a9d2d),
	.w5(32'hbae1d5dc),
	.w6(32'h3bb0c29c),
	.w7(32'h3b885d46),
	.w8(32'hbb2b8012),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1694),
	.w1(32'hbc39a50a),
	.w2(32'h3ca99195),
	.w3(32'hbcbc2de1),
	.w4(32'h3a431e52),
	.w5(32'hbcc7c7f9),
	.w6(32'hbc82dcf2),
	.w7(32'hbc27772f),
	.w8(32'hbce764ca),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46b040),
	.w1(32'h3a86f413),
	.w2(32'hbb34f0a3),
	.w3(32'h3bca584e),
	.w4(32'hbc261aba),
	.w5(32'hbc2a3380),
	.w6(32'h3c38c482),
	.w7(32'h3bd973f1),
	.w8(32'hbc431492),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4474a),
	.w1(32'hbc0690ac),
	.w2(32'hbb9bcb96),
	.w3(32'h3b39224c),
	.w4(32'hba9a5529),
	.w5(32'h398f3b98),
	.w6(32'hbb7f29c5),
	.w7(32'hbc14e93b),
	.w8(32'h3c817469),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198c58),
	.w1(32'h3bb13b01),
	.w2(32'h3c0dd5c0),
	.w3(32'h3c6043e7),
	.w4(32'h3c0ac220),
	.w5(32'h3c6b0b2f),
	.w6(32'h3bf46e82),
	.w7(32'h3c119acf),
	.w8(32'h3c5e16e2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c5c4b),
	.w1(32'h3b729652),
	.w2(32'h3a6c4a2d),
	.w3(32'h3b32c5a2),
	.w4(32'h3c04cbc4),
	.w5(32'hbcb989cc),
	.w6(32'hb9a9d9c6),
	.w7(32'h3c6f89df),
	.w8(32'hbcb8955d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a238c),
	.w1(32'hbc0134a6),
	.w2(32'hbbb17d6e),
	.w3(32'hbca8f81a),
	.w4(32'h3b6641c7),
	.w5(32'h3c332af2),
	.w6(32'hbc38ebd4),
	.w7(32'hbc88df6f),
	.w8(32'h37c59995),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9cdd1),
	.w1(32'hbc3d07f4),
	.w2(32'h3c4057a9),
	.w3(32'hba478ac2),
	.w4(32'h3c0ffa70),
	.w5(32'hbaeaf770),
	.w6(32'hbbd7141d),
	.w7(32'h3cb0ab14),
	.w8(32'h3cb9c534),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49f124),
	.w1(32'hbc771f50),
	.w2(32'hbb80d52d),
	.w3(32'hbc4ce1fb),
	.w4(32'h3b98d867),
	.w5(32'h3c57a756),
	.w6(32'h3ba648b1),
	.w7(32'hbb4c43cb),
	.w8(32'h3c887f04),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc296a2),
	.w1(32'h3c28e454),
	.w2(32'hbce7c981),
	.w3(32'h3c25b9ca),
	.w4(32'hbc9ddda8),
	.w5(32'h3abd19b9),
	.w6(32'h3c156023),
	.w7(32'hbd9c1d8b),
	.w8(32'hbc5b1e48),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27efe4),
	.w1(32'h3ce59191),
	.w2(32'h3c44c76f),
	.w3(32'h3cb8205a),
	.w4(32'h3b5e2768),
	.w5(32'hbbad3ca4),
	.w6(32'h3cec5e79),
	.w7(32'h3b80d578),
	.w8(32'hbcaca1c8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb524436),
	.w1(32'h3bf163dc),
	.w2(32'h3bf58bfc),
	.w3(32'hbbf3a1b9),
	.w4(32'h3ae0ed6d),
	.w5(32'h3ac0fd1f),
	.w6(32'hbb25d7d5),
	.w7(32'h3bc1d731),
	.w8(32'hbc5d0a05),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a5f9c),
	.w1(32'hbc100a40),
	.w2(32'h3c181bcc),
	.w3(32'h3ace5de1),
	.w4(32'h3c8b9b11),
	.w5(32'hbcbc3093),
	.w6(32'hbbad160a),
	.w7(32'h3d01ce92),
	.w8(32'hbc74d935),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88e349),
	.w1(32'hbcb2bd6f),
	.w2(32'h3c2e44ef),
	.w3(32'hbc71f932),
	.w4(32'hbb5fb5a3),
	.w5(32'hba0598b0),
	.w6(32'hbcb1229a),
	.w7(32'hbb4aada3),
	.w8(32'h3b534ea2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fb1df),
	.w1(32'h3c063f88),
	.w2(32'hbc0fc52b),
	.w3(32'hbb05b359),
	.w4(32'hbaec44d6),
	.w5(32'hbc34fbea),
	.w6(32'h3c48ea43),
	.w7(32'h3c10bf88),
	.w8(32'hbb88248e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace97d6),
	.w1(32'hbbac7bcc),
	.w2(32'hbc9f525e),
	.w3(32'hbad00abb),
	.w4(32'hbad3b8f8),
	.w5(32'h3c843e5c),
	.w6(32'h3b87837d),
	.w7(32'hbd3cf653),
	.w8(32'h3c664dc5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4418),
	.w1(32'h3c6a542e),
	.w2(32'h3c728483),
	.w3(32'h3c8582c6),
	.w4(32'h3ad566db),
	.w5(32'hbbc0e098),
	.w6(32'h3c4d0dd9),
	.w7(32'hbb9c2975),
	.w8(32'hbc1382dc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b6e1),
	.w1(32'hbc922460),
	.w2(32'h3bc1fad5),
	.w3(32'h3b912d58),
	.w4(32'hbaf80bee),
	.w5(32'hbc4b88bc),
	.w6(32'hbbeaf359),
	.w7(32'h3c1b4e37),
	.w8(32'hbc68c53c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8658a),
	.w1(32'h3be35e2a),
	.w2(32'h3bc4d2e5),
	.w3(32'h3bc73b7f),
	.w4(32'h3b8bb5c5),
	.w5(32'hbbf31c23),
	.w6(32'h3bf71325),
	.w7(32'h3ce5093e),
	.w8(32'h3aa549e8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c224488),
	.w1(32'hbb65f80e),
	.w2(32'h3c933343),
	.w3(32'h3c153a32),
	.w4(32'h3babc9c8),
	.w5(32'h3bdccf22),
	.w6(32'h3ba1a145),
	.w7(32'hbc5b6d70),
	.w8(32'h3bf7b304),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c835040),
	.w1(32'h3baa1fb8),
	.w2(32'h3c083279),
	.w3(32'hbb0528d4),
	.w4(32'hbc3f99d2),
	.w5(32'hba42cf3e),
	.w6(32'h3bae1666),
	.w7(32'hbb9c0e63),
	.w8(32'h3c440295),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e226),
	.w1(32'h3c6511f0),
	.w2(32'hbc0e3212),
	.w3(32'hbbfbfa25),
	.w4(32'hbb31e3d2),
	.w5(32'hbcf45b36),
	.w6(32'h3be59590),
	.w7(32'h3c4e7109),
	.w8(32'hbc6c755c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c476e37),
	.w1(32'h39a0da3a),
	.w2(32'h3d1e8426),
	.w3(32'hbcaba7bd),
	.w4(32'h3b163224),
	.w5(32'h3a53b430),
	.w6(32'hbbccf627),
	.w7(32'h3cbfd315),
	.w8(32'hbc8158db),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9de1f),
	.w1(32'hbc53b587),
	.w2(32'h3d3e45ce),
	.w3(32'hbc9b1ffb),
	.w4(32'h3d03c976),
	.w5(32'hbcae9a60),
	.w6(32'hbc92bc68),
	.w7(32'h3d8a738d),
	.w8(32'hbc8cb379),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba738d7),
	.w1(32'hbd0d7ea8),
	.w2(32'hbbd9c3a6),
	.w3(32'hbd1c4828),
	.w4(32'h3c3b6fc1),
	.w5(32'h399092e4),
	.w6(32'hbcea98b6),
	.w7(32'hba35738b),
	.w8(32'h3cc65965),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c311da2),
	.w1(32'h3c622c64),
	.w2(32'h3c1384bc),
	.w3(32'hbc1e7f3e),
	.w4(32'hb9e007dd),
	.w5(32'h3cb88424),
	.w6(32'hbbcb1071),
	.w7(32'h3d3fa94d),
	.w8(32'h3db7d4c4),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c327ab2),
	.w1(32'hbc914bc1),
	.w2(32'h39a07ae2),
	.w3(32'hbb8fccca),
	.w4(32'h3ace948a),
	.w5(32'hbc9bc620),
	.w6(32'h3c0cf496),
	.w7(32'h39b2acb6),
	.w8(32'hbd1ba792),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a2816),
	.w1(32'hbad31e25),
	.w2(32'h3b069f68),
	.w3(32'hbb612fb8),
	.w4(32'h3b3c705a),
	.w5(32'hbc04cd44),
	.w6(32'hbb969003),
	.w7(32'h3bd21df1),
	.w8(32'hbc086f01),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fd51e),
	.w1(32'hbb82aef0),
	.w2(32'h3c201a5a),
	.w3(32'hbb2a7322),
	.w4(32'hbc261ee9),
	.w5(32'hbbdb4afb),
	.w6(32'hbb939c97),
	.w7(32'hbb1064a8),
	.w8(32'h3bf145c4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca4f94a),
	.w1(32'hbbbd085e),
	.w2(32'h3cd7df21),
	.w3(32'hbc1c4693),
	.w4(32'h3c228090),
	.w5(32'hbc8ecce8),
	.w6(32'h3b0dd0b0),
	.w7(32'h3d27a967),
	.w8(32'hbcd65aff),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee50ea),
	.w1(32'hbc750e7b),
	.w2(32'hb9f01f90),
	.w3(32'hbc561a9b),
	.w4(32'hbba19272),
	.w5(32'hbbb15f4d),
	.w6(32'hbc9df3b3),
	.w7(32'hbcade66c),
	.w8(32'hbc2c6157),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64e4d1),
	.w1(32'h3a2173bb),
	.w2(32'hbc05a850),
	.w3(32'hbbe7b0c5),
	.w4(32'hbb9d281a),
	.w5(32'hbc5e2031),
	.w6(32'hbc014c5f),
	.w7(32'hbca04d0f),
	.w8(32'hbb392012),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c993b15),
	.w1(32'h3c0c5f5e),
	.w2(32'h3bc24c7c),
	.w3(32'hbc0c84bd),
	.w4(32'h3a155301),
	.w5(32'hbbf51911),
	.w6(32'hbafd19c3),
	.w7(32'h3c1303df),
	.w8(32'hbc12d20a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8c59d),
	.w1(32'hbbb9ca2a),
	.w2(32'h3bb4476e),
	.w3(32'hbbd965ca),
	.w4(32'h3b668f53),
	.w5(32'h3b8d29cb),
	.w6(32'hbc035fe0),
	.w7(32'h3bc35ce3),
	.w8(32'hbd165708),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91a34d),
	.w1(32'hbc2507a9),
	.w2(32'hbc813229),
	.w3(32'hbbc82d84),
	.w4(32'h3b248632),
	.w5(32'h3becf3ef),
	.w6(32'hbc2ccf00),
	.w7(32'hbc90dcc9),
	.w8(32'h3b8d3d77),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeae1e),
	.w1(32'h3b4c9f1b),
	.w2(32'hbb599419),
	.w3(32'h3cb64254),
	.w4(32'hbad17a7f),
	.w5(32'hbaf31b8e),
	.w6(32'h3c740689),
	.w7(32'hbbdc35f0),
	.w8(32'hbbcc861e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc560621),
	.w1(32'h3a99d9c5),
	.w2(32'h3c8f7143),
	.w3(32'hbb9dc1ff),
	.w4(32'hbbd9f458),
	.w5(32'h3b8be0af),
	.w6(32'hba2db1d4),
	.w7(32'h3c4dfc61),
	.w8(32'hbc63e2a5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e1b83),
	.w1(32'h3c22f5df),
	.w2(32'h3b87d5c8),
	.w3(32'h3bed252e),
	.w4(32'h3a88e40b),
	.w5(32'hbc1c3424),
	.w6(32'h3bf93c68),
	.w7(32'h3c4423ed),
	.w8(32'hbc46b875),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c33ac),
	.w1(32'hbc635536),
	.w2(32'hbb4593d0),
	.w3(32'hbc03b1bd),
	.w4(32'hbad87d2e),
	.w5(32'h3c0afcff),
	.w6(32'hbc928595),
	.w7(32'hbcb3a042),
	.w8(32'h3c144ddb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb98d8d),
	.w1(32'h3bede908),
	.w2(32'hbc64be25),
	.w3(32'h3b94b130),
	.w4(32'hbc4e0f32),
	.w5(32'hbc43266c),
	.w6(32'h3c8193eb),
	.w7(32'hbca756f5),
	.w8(32'hbbe77619),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bd659),
	.w1(32'hbc21d10b),
	.w2(32'h3c1d143f),
	.w3(32'hbbd361de),
	.w4(32'hba92b23e),
	.w5(32'h3b0162e6),
	.w6(32'h3afd996b),
	.w7(32'hbb92f751),
	.w8(32'h3ce092f0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbdc6fb),
	.w1(32'hbc9ef544),
	.w2(32'hbcd8046e),
	.w3(32'hbbbb2489),
	.w4(32'h3bf0ac17),
	.w5(32'h3c14c50c),
	.w6(32'hbcf84103),
	.w7(32'h3a848c43),
	.w8(32'h3d0d4ff8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73e9bd),
	.w1(32'h3bd1ad79),
	.w2(32'h3c1d8e6c),
	.w3(32'hbaac2d66),
	.w4(32'hbbbc51f7),
	.w5(32'hbc9c5bd0),
	.w6(32'h3c46c0d6),
	.w7(32'h3c7deba9),
	.w8(32'hbc8969c3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc1098),
	.w1(32'hbb093001),
	.w2(32'hb9bef18a),
	.w3(32'hbc8e1879),
	.w4(32'hbbeb9eef),
	.w5(32'hbc33316f),
	.w6(32'hbc811478),
	.w7(32'h3c0bc0aa),
	.w8(32'hbceb320a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc935f8f),
	.w1(32'h3b9a8fad),
	.w2(32'hbc36bcd2),
	.w3(32'hbbd887a9),
	.w4(32'h3c278054),
	.w5(32'h3c662952),
	.w6(32'h3b8c82eb),
	.w7(32'hbc6b9b02),
	.w8(32'h3a4dfaf7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a431843),
	.w1(32'h3befae3c),
	.w2(32'h3c6a457d),
	.w3(32'h3c345b76),
	.w4(32'h3bd3fc1b),
	.w5(32'hbb6c9372),
	.w6(32'h3c33c6fc),
	.w7(32'h3c80272d),
	.w8(32'hbc468b89),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83d0d9),
	.w1(32'hbc48384d),
	.w2(32'hbb0e176f),
	.w3(32'hbc8b897c),
	.w4(32'h3c41056a),
	.w5(32'hba1600c1),
	.w6(32'hbcbc9100),
	.w7(32'hbba015cb),
	.w8(32'h3a922c1e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ec653),
	.w1(32'h3b3ea2f5),
	.w2(32'hb8d7b00e),
	.w3(32'hbc949e99),
	.w4(32'hbcdcddbb),
	.w5(32'hbcb70433),
	.w6(32'h3aa6f311),
	.w7(32'hbcc9707a),
	.w8(32'hbcfd47ba),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e6ae),
	.w1(32'h397c51ad),
	.w2(32'h3cda879b),
	.w3(32'hba0ff690),
	.w4(32'h3b352552),
	.w5(32'hbb06a782),
	.w6(32'h3a8a1d35),
	.w7(32'hb7f4663f),
	.w8(32'hbce66672),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc852452),
	.w1(32'hbbd9208d),
	.w2(32'h3c0f27fa),
	.w3(32'hbc82dbd2),
	.w4(32'hbb388d24),
	.w5(32'hbca2e8c3),
	.w6(32'hbbb75d49),
	.w7(32'h3c4ce8a9),
	.w8(32'hbcba3c06),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65ce36),
	.w1(32'hbc290df7),
	.w2(32'h38a49d0c),
	.w3(32'hbb63fc01),
	.w4(32'hb99db314),
	.w5(32'hba082048),
	.w6(32'hbc1bb6b5),
	.w7(32'hb7b2af78),
	.w8(32'hba220f10),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a26194),
	.w1(32'h3853a523),
	.w2(32'hba21e09b),
	.w3(32'hb88cf147),
	.w4(32'hb9fb8198),
	.w5(32'hba337a38),
	.w6(32'hb89121a2),
	.w7(32'hba10ab1a),
	.w8(32'hba1ee53a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2718c),
	.w1(32'h390791de),
	.w2(32'hbad3d0f1),
	.w3(32'hbb786c70),
	.w4(32'hbb909c29),
	.w5(32'hbb33ae72),
	.w6(32'hbb6468ab),
	.w7(32'hbbe9587f),
	.w8(32'hbbc89614),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd3c8f),
	.w1(32'hbbaff769),
	.w2(32'hbbd0a57f),
	.w3(32'hbb3ad8f7),
	.w4(32'hbba2bf05),
	.w5(32'hbb95e8ef),
	.w6(32'hbba020fd),
	.w7(32'hbb336cfe),
	.w8(32'hbb6180c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fad7bf),
	.w1(32'h380bfe96),
	.w2(32'h38814b77),
	.w3(32'h38a79574),
	.w4(32'h3889533e),
	.w5(32'h3938e433),
	.w6(32'hb8e909f6),
	.w7(32'hb79fb276),
	.w8(32'h38b86472),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f8a92),
	.w1(32'h3ae173b8),
	.w2(32'h3a99a137),
	.w3(32'h3a8ed9b1),
	.w4(32'h39b1f0be),
	.w5(32'h38ad4c52),
	.w6(32'h3addc2f8),
	.w7(32'h3a862992),
	.w8(32'h3a13b353),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb584f4),
	.w1(32'h3bc0688a),
	.w2(32'h3b2a07b9),
	.w3(32'h3bec3ed5),
	.w4(32'h3bbccc62),
	.w5(32'h3b9d80a5),
	.w6(32'h3c2a826a),
	.w7(32'h3c1a2b67),
	.w8(32'h3bd2df16),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a034),
	.w1(32'h3b038b3c),
	.w2(32'h3a8cd1aa),
	.w3(32'h3a913ad8),
	.w4(32'h39b9c786),
	.w5(32'hb9ac02ae),
	.w6(32'h3b4f1c27),
	.w7(32'h3b202825),
	.w8(32'h3b0fd02a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7d25),
	.w1(32'hbb939dce),
	.w2(32'hbc05168e),
	.w3(32'hbc2b07e7),
	.w4(32'hbc39c57b),
	.w5(32'hbc28e52f),
	.w6(32'hbc4bb922),
	.w7(32'hbc8adc3c),
	.w8(32'hbc8f2c1c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e307),
	.w1(32'hbad281f9),
	.w2(32'hba32c16e),
	.w3(32'hbb2cd854),
	.w4(32'hbb57dcd5),
	.w5(32'hbb3150db),
	.w6(32'hbb89cea9),
	.w7(32'hbb9cd313),
	.w8(32'hbb2a8560),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b50dfd),
	.w1(32'h39e90c76),
	.w2(32'h3a0c2cff),
	.w3(32'h3a040937),
	.w4(32'h3a2bbc6a),
	.w5(32'h3a368e7b),
	.w6(32'h3a34896e),
	.w7(32'h3a4883f1),
	.w8(32'h3a24d8fd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8205dc0),
	.w1(32'hb7463d45),
	.w2(32'hb6f40d35),
	.w3(32'h3759ed7c),
	.w4(32'hb7e94b35),
	.w5(32'hb79794d8),
	.w6(32'hb8612ded),
	.w7(32'hb8a3c192),
	.w8(32'hb8cb435b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85dcd7),
	.w1(32'h3a495775),
	.w2(32'h3a0ce516),
	.w3(32'h3a887f01),
	.w4(32'h3a475137),
	.w5(32'h395dfb8b),
	.w6(32'h3a48e93f),
	.w7(32'h39699ba7),
	.w8(32'h3964f2ce),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964ce91),
	.w1(32'hb90629f2),
	.w2(32'hb8b672f6),
	.w3(32'hb9683416),
	.w4(32'h38aafd8e),
	.w5(32'hba028610),
	.w6(32'hb9e8bcbb),
	.w7(32'hb9dca277),
	.w8(32'hb997663c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27892d),
	.w1(32'h3a111a67),
	.w2(32'h3a117462),
	.w3(32'h3a73488e),
	.w4(32'h3a692d40),
	.w5(32'h39febeff),
	.w6(32'h3abff465),
	.w7(32'h3aab4ef2),
	.w8(32'h3aab19d9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67f816),
	.w1(32'hbb5313a4),
	.w2(32'hba4f2240),
	.w3(32'hbbadcf9b),
	.w4(32'hbb3c9f99),
	.w5(32'hbaf8f036),
	.w6(32'hbb31b4e4),
	.w7(32'hbb2c89e4),
	.w8(32'h3a19220b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbe214),
	.w1(32'h398b03a3),
	.w2(32'h3987b4c2),
	.w3(32'h3aed5ea6),
	.w4(32'h3b236905),
	.w5(32'h3ad7a73c),
	.w6(32'h3b52de17),
	.w7(32'h3b562d65),
	.w8(32'h3b70783d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c829330),
	.w1(32'h3c732f49),
	.w2(32'h3c54e411),
	.w3(32'h3c70e432),
	.w4(32'h3c4f44cc),
	.w5(32'h3c331a10),
	.w6(32'h3c809883),
	.w7(32'h3c5b13eb),
	.w8(32'h3c31dcb1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b4772),
	.w1(32'h3c8944f9),
	.w2(32'h3c431154),
	.w3(32'h3c958345),
	.w4(32'h3c8613c4),
	.w5(32'h3c3ba7ef),
	.w6(32'h3c8a09fd),
	.w7(32'h3c828913),
	.w8(32'h3c5acec4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaf739),
	.w1(32'hbba90275),
	.w2(32'hbb0b7903),
	.w3(32'hbbb3a18f),
	.w4(32'hbb8bbaaf),
	.w5(32'hbad8c90a),
	.w6(32'hba96ede3),
	.w7(32'h3a53290d),
	.w8(32'h3b0cc969),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e2c2ff),
	.w1(32'h39392775),
	.w2(32'hb9b119e1),
	.w3(32'h391b1e06),
	.w4(32'hb7cc83ed),
	.w5(32'hb91d7994),
	.w6(32'h38d7841e),
	.w7(32'h390f2b60),
	.w8(32'hb8a46f90),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8532bc5),
	.w1(32'hb8e3bef3),
	.w2(32'hb8c0c638),
	.w3(32'hb909401b),
	.w4(32'h3814e926),
	.w5(32'h36d48b1b),
	.w6(32'hb90f9e33),
	.w7(32'hb8ce9ce6),
	.w8(32'hb7b21235),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8990689),
	.w1(32'hb8d0b561),
	.w2(32'hb8f2a338),
	.w3(32'hb83a825f),
	.w4(32'hb92b33cf),
	.w5(32'hb951495d),
	.w6(32'hb97c0090),
	.w7(32'hb9bb3494),
	.w8(32'hb9d84eed),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818275c),
	.w1(32'hb89ac5c7),
	.w2(32'hb7bb0ad5),
	.w3(32'hb80539d6),
	.w4(32'hb89130b4),
	.w5(32'h37114c0d),
	.w6(32'hb94f1bf1),
	.w7(32'hb93506a8),
	.w8(32'hb90b1bc2),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cbd4f),
	.w1(32'hba00c64c),
	.w2(32'hb7f069ee),
	.w3(32'hbad8704a),
	.w4(32'hba172d37),
	.w5(32'hb99f0d28),
	.w6(32'hb982d816),
	.w7(32'h3990541d),
	.w8(32'h3a275be4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8dd5),
	.w1(32'h3bcfde53),
	.w2(32'h3b93333c),
	.w3(32'h3c030275),
	.w4(32'h3bc6ea9e),
	.w5(32'h3bfa2f23),
	.w6(32'h3c1ad794),
	.w7(32'h3c3c76c9),
	.w8(32'h3bf323da),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48b131),
	.w1(32'hbc6c708e),
	.w2(32'hbc652018),
	.w3(32'hbc8ae216),
	.w4(32'hbc862a49),
	.w5(32'hbc7bbc09),
	.w6(32'hbcb434ba),
	.w7(32'hbcbccc65),
	.w8(32'hbca194fb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcf1ba),
	.w1(32'hbb5f9ce2),
	.w2(32'hbb73af7f),
	.w3(32'hbb2e48c7),
	.w4(32'hbb87904c),
	.w5(32'hbb8f80ae),
	.w6(32'hbb66e332),
	.w7(32'hbbbb5d3b),
	.w8(32'hbba21770),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae35573),
	.w1(32'h3b0801ba),
	.w2(32'h3afcd741),
	.w3(32'h3a606a0e),
	.w4(32'h3afce2e9),
	.w5(32'h3a84dcfd),
	.w6(32'h3b07b0cc),
	.w7(32'h3b1249ae),
	.w8(32'h3b08ef1a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03c1f6),
	.w1(32'hbc2b69d6),
	.w2(32'hbc6936d3),
	.w3(32'hbc8e73d2),
	.w4(32'hbca703f7),
	.w5(32'hbcbe4a7a),
	.w6(32'hbcaeefc7),
	.w7(32'hbcb47ba8),
	.w8(32'hbcd732dd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf52601),
	.w1(32'h3c1b81b4),
	.w2(32'h3bdb18f6),
	.w3(32'h3c38622f),
	.w4(32'h3c3a9ca4),
	.w5(32'h3c2fe152),
	.w6(32'h3c50eb4b),
	.w7(32'h3c6e446c),
	.w8(32'h3c4a9d14),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af595a0),
	.w1(32'h3ac8c400),
	.w2(32'h3af2ba26),
	.w3(32'h3b64cbfd),
	.w4(32'h3b0d8c58),
	.w5(32'h3b91667a),
	.w6(32'h3bbfffd8),
	.w7(32'h3be8ae8c),
	.w8(32'h3bc467bb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becb3c3),
	.w1(32'h3c0e737d),
	.w2(32'h3c109b82),
	.w3(32'h3bc05db2),
	.w4(32'h3c042d44),
	.w5(32'h3bf370d7),
	.w6(32'h3bed78c1),
	.w7(32'h3c092493),
	.w8(32'h3c026388),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c57c),
	.w1(32'h3b582c32),
	.w2(32'h3a25c7aa),
	.w3(32'h3b988af2),
	.w4(32'h3b1e372d),
	.w5(32'h3ad27b01),
	.w6(32'h3b92fad0),
	.w7(32'h3b3954df),
	.w8(32'h39ba1ccc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87326e),
	.w1(32'hb9d836ee),
	.w2(32'hbadb56c8),
	.w3(32'h3acdf4c4),
	.w4(32'hb9b90b58),
	.w5(32'h3aa70371),
	.w6(32'h3ba051ae),
	.w7(32'h3ba8e20f),
	.w8(32'h3b59360e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988ae96),
	.w1(32'h3990ca75),
	.w2(32'h39b23d43),
	.w3(32'h3a92bd70),
	.w4(32'h3ab42bba),
	.w5(32'h3ae0d670),
	.w6(32'h3b315d19),
	.w7(32'h3b6303f1),
	.w8(32'h3b53f570),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7bb29),
	.w1(32'h3a1112ee),
	.w2(32'h3b1cc2d5),
	.w3(32'h3b5c0a7a),
	.w4(32'hb9cbd391),
	.w5(32'h3a81b789),
	.w6(32'h3afd8ce4),
	.w7(32'hbb15b47a),
	.w8(32'hb95655b8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fdd46a),
	.w1(32'hb97234b2),
	.w2(32'hb912d9e5),
	.w3(32'hb9a3d8a7),
	.w4(32'hb93e6059),
	.w5(32'hb98e2f4e),
	.w6(32'hba1524d9),
	.w7(32'hba6d83c7),
	.w8(32'hba59e724),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de440a),
	.w1(32'h398beb7a),
	.w2(32'h36b6ae80),
	.w3(32'h392d9a9d),
	.w4(32'h398d0907),
	.w5(32'hb8b971b4),
	.w6(32'hb92088df),
	.w7(32'hb9bfd4e5),
	.w8(32'hb9aa0dd6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6eb8),
	.w1(32'hbb8f103b),
	.w2(32'hbbb83207),
	.w3(32'hbbe8739a),
	.w4(32'hbbed61a4),
	.w5(32'hbbe710ad),
	.w6(32'hbbd64d8d),
	.w7(32'hbc004140),
	.w8(32'hbbec257e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ac257),
	.w1(32'h385f9d64),
	.w2(32'h39e3b304),
	.w3(32'hbadc7721),
	.w4(32'hba23f581),
	.w5(32'hba8c5ce9),
	.w6(32'h3a6ea1d2),
	.w7(32'h3aec4c17),
	.w8(32'h3abde06b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb9d48),
	.w1(32'hb9a2b472),
	.w2(32'hb9d364c8),
	.w3(32'hb9a0b926),
	.w4(32'hb9c4a4b3),
	.w5(32'hb9723ea5),
	.w6(32'h3a36e994),
	.w7(32'h3a501031),
	.w8(32'h3a2f1da5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84d9101),
	.w1(32'hb86f0faf),
	.w2(32'hb80b701e),
	.w3(32'hb8374070),
	.w4(32'hb8d358a0),
	.w5(32'h38884793),
	.w6(32'hb8c10cb8),
	.w7(32'hb8a5b25e),
	.w8(32'hb8fcb3dd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb600366f),
	.w1(32'hb99f8f6d),
	.w2(32'hb9afa187),
	.w3(32'h35a9a582),
	.w4(32'hb9a2d423),
	.w5(32'hba331a5e),
	.w6(32'hb7b196d2),
	.w7(32'hb952065f),
	.w8(32'hb9f98284),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4974a),
	.w1(32'hbb011c1e),
	.w2(32'hbb30b3d2),
	.w3(32'hbae673f7),
	.w4(32'hbb0f5fbb),
	.w5(32'hbb26b5f9),
	.w6(32'hbab99203),
	.w7(32'hbb1fa2cc),
	.w8(32'hbb1317b2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88a2c3),
	.w1(32'hb8a9352f),
	.w2(32'hba9cc576),
	.w3(32'hba962c40),
	.w4(32'hbac44c37),
	.w5(32'hbb2a5922),
	.w6(32'h39cc922e),
	.w7(32'hb9a47481),
	.w8(32'hbb010bba),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8f003),
	.w1(32'h39cc7b8e),
	.w2(32'h3a8ccbab),
	.w3(32'h39bcf56e),
	.w4(32'h3972b6a1),
	.w5(32'h3a278eae),
	.w6(32'hb89c6893),
	.w7(32'h39cbb3e6),
	.w8(32'h3a09543a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae26763),
	.w1(32'hbb0fcf4f),
	.w2(32'hbae87d0d),
	.w3(32'hbaaa2d29),
	.w4(32'hba70b5ed),
	.w5(32'hba23bb85),
	.w6(32'hbaea28df),
	.w7(32'hbaeb6d73),
	.w8(32'hb8c24124),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9782c),
	.w1(32'h3af0c8d3),
	.w2(32'h3af62e13),
	.w3(32'h3ade442c),
	.w4(32'h3b22265c),
	.w5(32'h3b3dcae2),
	.w6(32'h3b8a6783),
	.w7(32'h3bc0ce95),
	.w8(32'h3b7a5f61),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41c682),
	.w1(32'h3afca890),
	.w2(32'h3ad6c8e7),
	.w3(32'h3b83ad73),
	.w4(32'h3ac750c0),
	.w5(32'h3b4a6911),
	.w6(32'h3bc19344),
	.w7(32'h3b8db9e1),
	.w8(32'h3b865a06),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3cc22),
	.w1(32'hbbe409ed),
	.w2(32'hbc1231fc),
	.w3(32'hbbdcff02),
	.w4(32'hbc013713),
	.w5(32'hbbcd568f),
	.w6(32'hbb90bd82),
	.w7(32'hbc264337),
	.w8(32'hbbfb8899),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71b213),
	.w1(32'hbb5a41a4),
	.w2(32'hbb35d6b6),
	.w3(32'hbb284074),
	.w4(32'hbac5fae8),
	.w5(32'hbaaf9702),
	.w6(32'hba902ebb),
	.w7(32'hba117d70),
	.w8(32'h39dbbdfe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule