module layer_8_featuremap_124(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161b9a),
	.w1(32'hba95bb8f),
	.w2(32'h3be45a3e),
	.w3(32'hbb4729c4),
	.w4(32'h3c02e468),
	.w5(32'h3c25f702),
	.w6(32'h3aecaf02),
	.w7(32'h3ca77d43),
	.w8(32'hbc9d6e65),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe399),
	.w1(32'h3b8c9476),
	.w2(32'hbc7627b4),
	.w3(32'hbc31b959),
	.w4(32'h3c15a628),
	.w5(32'hbc82ff3f),
	.w6(32'hbb864a50),
	.w7(32'h3a92ddf7),
	.w8(32'h398c7c76),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfce82),
	.w1(32'h3b82ef41),
	.w2(32'hbafd2cd5),
	.w3(32'hbc448c9d),
	.w4(32'h3bd6d583),
	.w5(32'hbc0155a8),
	.w6(32'h3bae44d1),
	.w7(32'h3b4c7ea5),
	.w8(32'hbc85eacc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ba9c4),
	.w1(32'hbb9673ea),
	.w2(32'h3be0ffc8),
	.w3(32'hbb0bee63),
	.w4(32'hbb665dc1),
	.w5(32'hbc8c1f19),
	.w6(32'hbcb927ba),
	.w7(32'h39a9c820),
	.w8(32'h3b719048),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2d79e),
	.w1(32'hbbf9421e),
	.w2(32'hbc2ca889),
	.w3(32'h3c9fb6f9),
	.w4(32'hbc48d473),
	.w5(32'hbc5b4752),
	.w6(32'hbb1f087b),
	.w7(32'hbbf8059b),
	.w8(32'hbc206e2f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad80121),
	.w1(32'hbc241123),
	.w2(32'h3c84054b),
	.w3(32'hb8cab39b),
	.w4(32'h39130bf2),
	.w5(32'hbbdffd35),
	.w6(32'hbc2a7845),
	.w7(32'hbc9adbef),
	.w8(32'h3d6760d6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd615f),
	.w1(32'hbd293809),
	.w2(32'hbc8de48a),
	.w3(32'h3c5cc4be),
	.w4(32'h3bac360c),
	.w5(32'hbcea4120),
	.w6(32'h3b2c6a47),
	.w7(32'hbcaaf944),
	.w8(32'h3ca9b16d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc015e4),
	.w1(32'hbb2e696e),
	.w2(32'hbcbbcb15),
	.w3(32'hbc43e9ad),
	.w4(32'h3c9ffd44),
	.w5(32'hbc13929e),
	.w6(32'hbc3ebe78),
	.w7(32'hbbd3d20a),
	.w8(32'h3bddbe23),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b947f02),
	.w1(32'h3b8b9879),
	.w2(32'h3c6ad7e6),
	.w3(32'h3ac26c80),
	.w4(32'hbbaaa780),
	.w5(32'h3bb6b50b),
	.w6(32'h3c91272e),
	.w7(32'hbbee1dc5),
	.w8(32'h3c06192a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836436),
	.w1(32'hbbcac452),
	.w2(32'hbbbac932),
	.w3(32'h3b59751b),
	.w4(32'hbc51783e),
	.w5(32'hbca79f13),
	.w6(32'hbb9776f9),
	.w7(32'hbc9023ac),
	.w8(32'h3d30844f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e620c),
	.w1(32'hb9bb5212),
	.w2(32'h38b72309),
	.w3(32'h3bf8044b),
	.w4(32'hbc2dd97c),
	.w5(32'h3c30c091),
	.w6(32'hbb0ac007),
	.w7(32'h3c9f6341),
	.w8(32'hbcafa68b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a8185),
	.w1(32'hba199fee),
	.w2(32'hbbe93817),
	.w3(32'h3a2259e7),
	.w4(32'hba38045a),
	.w5(32'hbb02b24e),
	.w6(32'h3a2f4d53),
	.w7(32'hbd0d2cd3),
	.w8(32'h3cab2f7c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15e61),
	.w1(32'h3c349ebd),
	.w2(32'h3a7c786d),
	.w3(32'h3c0a6e8c),
	.w4(32'hba554cfd),
	.w5(32'hba198903),
	.w6(32'h3c5d29f7),
	.w7(32'hbba0410a),
	.w8(32'hbbececd5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad953eb),
	.w1(32'hba4ae514),
	.w2(32'h398d344d),
	.w3(32'hba8d966f),
	.w4(32'hbb409e51),
	.w5(32'hba6b9f55),
	.w6(32'hbc0b3ccb),
	.w7(32'hb97b350d),
	.w8(32'h3b699098),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30a499),
	.w1(32'h3b661ad9),
	.w2(32'hba6c91bf),
	.w3(32'h39aeaffe),
	.w4(32'hba885326),
	.w5(32'hba20723e),
	.w6(32'h3ba9c39c),
	.w7(32'hbaa4c50e),
	.w8(32'hba924586),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac946),
	.w1(32'h38f05f08),
	.w2(32'hbbf3e84f),
	.w3(32'h3abdbea2),
	.w4(32'h3b2a6cf4),
	.w5(32'hbabc270c),
	.w6(32'h3ad43905),
	.w7(32'h3c180344),
	.w8(32'h3c8f207c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20911b),
	.w1(32'hbc4e961a),
	.w2(32'hb98c40fd),
	.w3(32'h3b377f12),
	.w4(32'h3b87ed22),
	.w5(32'h3bcfaa95),
	.w6(32'h3c1aec0f),
	.w7(32'hbaa884fd),
	.w8(32'hba91fdc7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa0225),
	.w1(32'hbbefb366),
	.w2(32'h3ac9b69f),
	.w3(32'hba28c0d3),
	.w4(32'h3bb79f73),
	.w5(32'hba5c5e07),
	.w6(32'hbba56f22),
	.w7(32'hbb1d31d8),
	.w8(32'hbbe36e75),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b527e0d),
	.w1(32'hb89ec967),
	.w2(32'hbb896324),
	.w3(32'hbc28c621),
	.w4(32'h3b807cbc),
	.w5(32'hbbe662ca),
	.w6(32'h3799fd29),
	.w7(32'hbb140c19),
	.w8(32'h3b83d1ce),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b0dc),
	.w1(32'hbc822619),
	.w2(32'hbbe0897a),
	.w3(32'hbba67091),
	.w4(32'h3b9eb712),
	.w5(32'hbb98819f),
	.w6(32'hbbba9563),
	.w7(32'h3cd81d66),
	.w8(32'h3d2c5f42),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcecd7),
	.w1(32'hbc0ce2ea),
	.w2(32'hba82f1ee),
	.w3(32'h3bfe24c6),
	.w4(32'h3b2d8437),
	.w5(32'h3c48f215),
	.w6(32'h3ca429cb),
	.w7(32'hbc4f4eb8),
	.w8(32'hbc75448b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10eaa3),
	.w1(32'hbba28041),
	.w2(32'h3a4362f1),
	.w3(32'h3b723b4c),
	.w4(32'h3aab7357),
	.w5(32'h3c515fa3),
	.w6(32'hba047b57),
	.w7(32'hbb22fa44),
	.w8(32'hbb8be966),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bbc06),
	.w1(32'h3a4ef2b9),
	.w2(32'h3b175888),
	.w3(32'h3bff57be),
	.w4(32'h3b1c21d9),
	.w5(32'h3b20911c),
	.w6(32'hba8e9f55),
	.w7(32'hba2a128f),
	.w8(32'hbb9dd599),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5626f5),
	.w1(32'hbc090b5d),
	.w2(32'hbb4c312a),
	.w3(32'hbb4d4373),
	.w4(32'h39deadcf),
	.w5(32'hbb9ebdfb),
	.w6(32'hba480c3c),
	.w7(32'h398f172a),
	.w8(32'hbb9fcc24),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc2848),
	.w1(32'h3ba602c9),
	.w2(32'hbb8d053c),
	.w3(32'h3bf62641),
	.w4(32'h3b8aadcd),
	.w5(32'h3a7149e4),
	.w6(32'h3ba8fc16),
	.w7(32'h38cada22),
	.w8(32'hbbac7e9f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb940a3),
	.w1(32'hbaa068e0),
	.w2(32'h3c2f44aa),
	.w3(32'hbb2b95ac),
	.w4(32'h3bb4b34e),
	.w5(32'h3cad66ce),
	.w6(32'hbb0735a2),
	.w7(32'hbc43a11f),
	.w8(32'hbd1a50af),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadf091),
	.w1(32'h3c1cf673),
	.w2(32'hbc2425b4),
	.w3(32'hbb1f2238),
	.w4(32'h3a8c2e52),
	.w5(32'hbbb9e036),
	.w6(32'hbbbf3043),
	.w7(32'hbbfec534),
	.w8(32'hbc0af7a5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31162e),
	.w1(32'hbc376cfc),
	.w2(32'hba261488),
	.w3(32'hbbf2c41a),
	.w4(32'h3c399c26),
	.w5(32'h3ce26f4f),
	.w6(32'hbc28d392),
	.w7(32'h3b666795),
	.w8(32'h3c77eab2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81bc4a),
	.w1(32'hbb155d50),
	.w2(32'h3b21b658),
	.w3(32'h3bce1a4a),
	.w4(32'hbade49b1),
	.w5(32'hba2bb590),
	.w6(32'h3b80a96a),
	.w7(32'h3b3c05ab),
	.w8(32'h3cbfd002),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6c68c),
	.w1(32'h3c62cef3),
	.w2(32'h3c1a8de8),
	.w3(32'h3c2efb56),
	.w4(32'hbb030e43),
	.w5(32'h3c1a12cc),
	.w6(32'h3ba91d0f),
	.w7(32'hba4ad204),
	.w8(32'hbc0ce82b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32ae5b),
	.w1(32'h3c526f79),
	.w2(32'hba6e8fbd),
	.w3(32'h3bc2baab),
	.w4(32'hbafca330),
	.w5(32'h3a71298b),
	.w6(32'h3b56aa65),
	.w7(32'hbaefc56a),
	.w8(32'h39867d16),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ded41),
	.w1(32'hb8fb51f1),
	.w2(32'hbc06d16f),
	.w3(32'hb952467b),
	.w4(32'hbbc6ecb8),
	.w5(32'hbd016726),
	.w6(32'hba47833f),
	.w7(32'h3b5e10a1),
	.w8(32'h3c550ff2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf0a041),
	.w1(32'hbc76f5ce),
	.w2(32'h3bcc723c),
	.w3(32'hbc2d93dc),
	.w4(32'hbc012c8e),
	.w5(32'h3b76b8da),
	.w6(32'h3ba12932),
	.w7(32'h3b1e36cc),
	.w8(32'hbc27e056),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95d478),
	.w1(32'h3baafd04),
	.w2(32'hba59f2ab),
	.w3(32'h3c364864),
	.w4(32'h3bb1dd81),
	.w5(32'h3b9545a4),
	.w6(32'hbc07b6d8),
	.w7(32'h39880e31),
	.w8(32'hbbcb158e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c3f36),
	.w1(32'hbba001e6),
	.w2(32'h3bfb40f4),
	.w3(32'hbb2591b6),
	.w4(32'h3bc2a58b),
	.w5(32'hbb5cb494),
	.w6(32'h3a626ac6),
	.w7(32'h3b6755be),
	.w8(32'hbc32a91d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eadd8),
	.w1(32'h3b8f0ba8),
	.w2(32'h3be43e42),
	.w3(32'hbb040d6f),
	.w4(32'hbc911b60),
	.w5(32'hbbf33c4b),
	.w6(32'hbb506748),
	.w7(32'hba7652e5),
	.w8(32'hbbf2f5f2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69a4c7),
	.w1(32'h3b5391ec),
	.w2(32'h3b6ad5f0),
	.w3(32'h3ae3c514),
	.w4(32'hbaa7da5d),
	.w5(32'hbc19c9de),
	.w6(32'hbaaddde5),
	.w7(32'h3c1788e2),
	.w8(32'h3c029787),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dbb38),
	.w1(32'hbb7a0864),
	.w2(32'hbba66891),
	.w3(32'hbb972511),
	.w4(32'h3b93d7e4),
	.w5(32'h3c41c60d),
	.w6(32'hbb63180f),
	.w7(32'h39337f3e),
	.w8(32'h3b2da488),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d338a),
	.w1(32'h3b2cd862),
	.w2(32'h3b41f541),
	.w3(32'h3bd9e6d1),
	.w4(32'hbb2b3310),
	.w5(32'hbc83f4fb),
	.w6(32'h3c16fafb),
	.w7(32'h38cb5540),
	.w8(32'h3c4f1220),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc684add),
	.w1(32'hbb6c36eb),
	.w2(32'hbbf5a717),
	.w3(32'h3866c5ef),
	.w4(32'hbc1e0fd2),
	.w5(32'hbc266078),
	.w6(32'hbadf83bf),
	.w7(32'hbc512682),
	.w8(32'hbbf36fdb),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc337433),
	.w1(32'hbbd20a03),
	.w2(32'hbb58ed54),
	.w3(32'hbc20562a),
	.w4(32'hbb40a0a7),
	.w5(32'hbc28b2fc),
	.w6(32'hbc39a1d7),
	.w7(32'h3cc9a4f5),
	.w8(32'h3d26c5d3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb0700),
	.w1(32'hbb8339be),
	.w2(32'h3b8dc2cf),
	.w3(32'h3b0dc778),
	.w4(32'h3bb94df3),
	.w5(32'h3c0470be),
	.w6(32'h3c2298ea),
	.w7(32'hbb94bcda),
	.w8(32'hbcb738ef),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2cb00),
	.w1(32'hbc0b38dc),
	.w2(32'h3c187700),
	.w3(32'hbc8285af),
	.w4(32'h3ba69cf5),
	.w5(32'h3afd2779),
	.w6(32'hbc3fca91),
	.w7(32'hbc134df2),
	.w8(32'h3c18540b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad184e3),
	.w1(32'h3c510948),
	.w2(32'h3addc26c),
	.w3(32'h3c12c3b7),
	.w4(32'hbab6f0ba),
	.w5(32'h3a3992f3),
	.w6(32'hbb4d13c8),
	.w7(32'hbb9acbbd),
	.w8(32'hbbbed20e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a4616),
	.w1(32'h39b02711),
	.w2(32'h3c28531b),
	.w3(32'hb9e4645b),
	.w4(32'h3abdfdfe),
	.w5(32'h3bf45c87),
	.w6(32'hbbe8d058),
	.w7(32'h3b4e2694),
	.w8(32'h3c29f2b3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dd90a),
	.w1(32'h3c3c5cb3),
	.w2(32'hbb25a582),
	.w3(32'h3b817e93),
	.w4(32'h3ae209ac),
	.w5(32'h3b21b9a0),
	.w6(32'hbb49bc8d),
	.w7(32'hbb18de7f),
	.w8(32'h3bd756dd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04aee4),
	.w1(32'h3bfae519),
	.w2(32'hbb4334f0),
	.w3(32'hba69895e),
	.w4(32'hbb7782ab),
	.w5(32'h3ada9bc4),
	.w6(32'hbbcc3de9),
	.w7(32'hbc120352),
	.w8(32'hba6bdc2e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab268d2),
	.w1(32'h3a5b464e),
	.w2(32'hbbc0b931),
	.w3(32'h3c05d3ca),
	.w4(32'hbc000c88),
	.w5(32'h3b9c076b),
	.w6(32'hbb8cb7bd),
	.w7(32'hbc2b7312),
	.w8(32'hbc7812c1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaee202),
	.w1(32'h39ee9104),
	.w2(32'hbba55d1b),
	.w3(32'h3ba9dbb9),
	.w4(32'h393c2117),
	.w5(32'h3a65031d),
	.w6(32'hbc0261dc),
	.w7(32'h3a2e8ecb),
	.w8(32'hbca5baca),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5217cc),
	.w1(32'hbc9a7447),
	.w2(32'hbcb5ff9c),
	.w3(32'h3b04de8a),
	.w4(32'hbba6169b),
	.w5(32'hbbc66f27),
	.w6(32'hbbd21768),
	.w7(32'hbbe1540f),
	.w8(32'h3c2d0c98),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb2132f),
	.w1(32'hbc67482a),
	.w2(32'h3b44a7d1),
	.w3(32'h3b81463d),
	.w4(32'h3c2171db),
	.w5(32'h3ceaff3a),
	.w6(32'h3b0ea3fa),
	.w7(32'hbc233b7c),
	.w8(32'hbd4acb59),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8571cc),
	.w1(32'h39d24b09),
	.w2(32'hb8b3cc4b),
	.w3(32'h3b8bf288),
	.w4(32'h3bcb224c),
	.w5(32'h3c6ca8a1),
	.w6(32'hbc16d939),
	.w7(32'hbb8eca07),
	.w8(32'h3a7b1150),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130dea),
	.w1(32'hba9e7e73),
	.w2(32'h3a988db1),
	.w3(32'hbbacc78a),
	.w4(32'h3bac15f0),
	.w5(32'hbb43f5b5),
	.w6(32'hbbfe4c44),
	.w7(32'hbb68ec61),
	.w8(32'h3cc52ada),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a20f9),
	.w1(32'h3a190e97),
	.w2(32'h3ad33dc2),
	.w3(32'h3bc7913c),
	.w4(32'hbad2fce6),
	.w5(32'h3a1da50e),
	.w6(32'h3cc80d58),
	.w7(32'hbb0dee6f),
	.w8(32'hba978311),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2472a),
	.w1(32'h3a9b8246),
	.w2(32'h3ba8faa6),
	.w3(32'hba244a98),
	.w4(32'hbb9ec39c),
	.w5(32'h3bb2b99c),
	.w6(32'hbaf339fd),
	.w7(32'hbc669018),
	.w8(32'hbc0e419d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb56a82),
	.w1(32'h3a5b628e),
	.w2(32'hbc71ef79),
	.w3(32'h3bbdd987),
	.w4(32'hb9c75a5f),
	.w5(32'hbb004890),
	.w6(32'hbb447695),
	.w7(32'hbbf3a2d6),
	.w8(32'hbb183b23),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b421f),
	.w1(32'hbc051ab2),
	.w2(32'hbbfe950c),
	.w3(32'hb9e0c02b),
	.w4(32'hbbe9393e),
	.w5(32'hbbf37bbf),
	.w6(32'hbc020350),
	.w7(32'hbb96d95b),
	.w8(32'hba9efecf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4f5c),
	.w1(32'hbb2113c1),
	.w2(32'h3c016531),
	.w3(32'hbaed9745),
	.w4(32'h3c87b412),
	.w5(32'h3d02d951),
	.w6(32'h3a9bf1f7),
	.w7(32'h3c8248cc),
	.w8(32'h3d0dd5f0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c803030),
	.w1(32'hbb292fee),
	.w2(32'h3ae86675),
	.w3(32'h3ba9149c),
	.w4(32'hba9ff57e),
	.w5(32'h3ac0ba43),
	.w6(32'h3ba58d44),
	.w7(32'hbb39294e),
	.w8(32'hbb149a20),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a931a27),
	.w1(32'h3ad12186),
	.w2(32'h3b93ae6d),
	.w3(32'h39ea543d),
	.w4(32'h3c827133),
	.w5(32'hbb235638),
	.w6(32'hbb7ef3b0),
	.w7(32'hbb8580d1),
	.w8(32'h39546ae2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52cbac),
	.w1(32'h3a342a8b),
	.w2(32'h3c3cc8a4),
	.w3(32'h399a3b92),
	.w4(32'h3b82ece0),
	.w5(32'h39d726bd),
	.w6(32'hb930ecb6),
	.w7(32'hb8a3f8ac),
	.w8(32'h39a88978),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa71330),
	.w1(32'h3b53b6b2),
	.w2(32'hbb3fd2f2),
	.w3(32'hbc6a88f8),
	.w4(32'hb9942410),
	.w5(32'h3b2a6fea),
	.w6(32'hbc2386ef),
	.w7(32'hbb42c424),
	.w8(32'hbb236323),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8718fcb),
	.w1(32'h3a2f8358),
	.w2(32'h3b2b620b),
	.w3(32'h3bb50250),
	.w4(32'hbc476ba6),
	.w5(32'hbbfb07a5),
	.w6(32'hb97fa97d),
	.w7(32'hbbff63c0),
	.w8(32'hbc1bee8c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb608c23),
	.w1(32'hbc27fae2),
	.w2(32'h3bde39ca),
	.w3(32'hbb9239bb),
	.w4(32'hbb6250b1),
	.w5(32'hbc14d90c),
	.w6(32'hbc8c366b),
	.w7(32'h3b977b67),
	.w8(32'h3c04ec70),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bf93d),
	.w1(32'h3bc26b2e),
	.w2(32'hbbc7f15a),
	.w3(32'hbb1461fa),
	.w4(32'hbad9faac),
	.w5(32'h3b0dbdac),
	.w6(32'h3ac74d3a),
	.w7(32'hbbaff957),
	.w8(32'h39f4a947),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f569b),
	.w1(32'hbac76387),
	.w2(32'h3bb5fb4c),
	.w3(32'h39471fc5),
	.w4(32'hbb2893b1),
	.w5(32'h3bdf6b00),
	.w6(32'h3b989ff0),
	.w7(32'h3a71d87c),
	.w8(32'h3aeea37d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cf746),
	.w1(32'h3c067e1a),
	.w2(32'h3ba1f586),
	.w3(32'hba70d8cc),
	.w4(32'h3b7d71ad),
	.w5(32'h3a5ff52c),
	.w6(32'h3c205d87),
	.w7(32'h3bb14a77),
	.w8(32'h3bf4b568),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38caad),
	.w1(32'h3ba9c4a6),
	.w2(32'hbb333c73),
	.w3(32'hbc70e33b),
	.w4(32'h3ba82a50),
	.w5(32'hbb535710),
	.w6(32'h3a8923a8),
	.w7(32'hbb59dfd5),
	.w8(32'h3aec85ee),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b46d3),
	.w1(32'hbb8a6741),
	.w2(32'hbbc0fb74),
	.w3(32'h3b862525),
	.w4(32'h3ba7a4d9),
	.w5(32'h39127542),
	.w6(32'h395cf5e6),
	.w7(32'h3c71d49b),
	.w8(32'h3d0fd6f9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74ac3c),
	.w1(32'hb9d91262),
	.w2(32'hbbc77e56),
	.w3(32'h3ba623a0),
	.w4(32'h3b22a4d9),
	.w5(32'h38185415),
	.w6(32'h3c5749d8),
	.w7(32'hbc3a5e0c),
	.w8(32'hbb2a2952),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b1cd),
	.w1(32'h3ab174ba),
	.w2(32'hbb120665),
	.w3(32'h3b04ce57),
	.w4(32'h3ba8dd93),
	.w5(32'h3b0e8a24),
	.w6(32'h3a35ac95),
	.w7(32'h37fe321c),
	.w8(32'h3bca4998),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbbe84),
	.w1(32'hbb981567),
	.w2(32'hbc5cd4d5),
	.w3(32'hbbce46ec),
	.w4(32'h3bbe5f9c),
	.w5(32'hbc4cd94b),
	.w6(32'hbb2e7714),
	.w7(32'hbc19d4be),
	.w8(32'hbc81baf6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65ea29),
	.w1(32'hbbcaeef8),
	.w2(32'hbb5b8742),
	.w3(32'hbc1bf77b),
	.w4(32'h3b5264ff),
	.w5(32'h3b9b720c),
	.w6(32'hbc89830c),
	.w7(32'h3c51f7c3),
	.w8(32'h3cae444c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90753d5),
	.w1(32'hbb468055),
	.w2(32'hb8e01df2),
	.w3(32'h3bc7ae85),
	.w4(32'hb96b4814),
	.w5(32'h3ac40bb7),
	.w6(32'h3c8f890a),
	.w7(32'hbc31871a),
	.w8(32'hbc1ed3ed),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37df91),
	.w1(32'hb979e47b),
	.w2(32'hbbce7572),
	.w3(32'h3c5d0940),
	.w4(32'h3bb4b4a4),
	.w5(32'h3acf1358),
	.w6(32'hbb2d1c71),
	.w7(32'hbc13f788),
	.w8(32'hbc52b1e0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc998962),
	.w1(32'hbc5a3d62),
	.w2(32'hbc2512ae),
	.w3(32'h3bc5c180),
	.w4(32'hbb588a7b),
	.w5(32'hbc445b8d),
	.w6(32'hbc0aab5a),
	.w7(32'hbc13881c),
	.w8(32'hbb4c5192),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17540c),
	.w1(32'hbbea6495),
	.w2(32'h3a2591ed),
	.w3(32'hbc467518),
	.w4(32'h3a96eed4),
	.w5(32'h3badeb0f),
	.w6(32'hbc4e17c9),
	.w7(32'hb9b82bce),
	.w8(32'hba0e9548),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba327f60),
	.w1(32'hb996d2d3),
	.w2(32'h3a340812),
	.w3(32'h3ab7cc85),
	.w4(32'h3a9cc606),
	.w5(32'h3a90b3b4),
	.w6(32'hbaed6234),
	.w7(32'h3a5d01f5),
	.w8(32'hbad7893a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c948a),
	.w1(32'hbab38db6),
	.w2(32'h3b2ab380),
	.w3(32'hb8d9015e),
	.w4(32'h3b324c99),
	.w5(32'h3b1074e3),
	.w6(32'hbb1c4091),
	.w7(32'h3b1651b9),
	.w8(32'h39a74dda),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9543d5),
	.w1(32'hba16c1b6),
	.w2(32'hbba6ebbf),
	.w3(32'h3a80c639),
	.w4(32'hbb4459ee),
	.w5(32'hbbc9db45),
	.w6(32'hba3dd378),
	.w7(32'hbba0fa05),
	.w8(32'hbba67f6a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9516f2),
	.w1(32'hbb8d616f),
	.w2(32'h3b7945f4),
	.w3(32'hbb5cacd9),
	.w4(32'hb9188aae),
	.w5(32'h3bad17a5),
	.w6(32'hbb9b0e56),
	.w7(32'h3b78dec6),
	.w8(32'h3a03ba98),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb6ac),
	.w1(32'hba67b777),
	.w2(32'h3a82386a),
	.w3(32'h3bfcdfeb),
	.w4(32'h3a5ebd11),
	.w5(32'hbb840cbb),
	.w6(32'h3bb2a2b3),
	.w7(32'h39fa03c3),
	.w8(32'hbb896457),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88d19a),
	.w1(32'hbbad8220),
	.w2(32'h3b45f3f8),
	.w3(32'hbb7571d6),
	.w4(32'h3a7ec424),
	.w5(32'hbb4eaeab),
	.w6(32'hbb92a1e7),
	.w7(32'hbb138047),
	.w8(32'hba37dce0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fc3d3),
	.w1(32'hbbe53f13),
	.w2(32'hbb108492),
	.w3(32'hbbdbf555),
	.w4(32'hba23d44c),
	.w5(32'h3a2858ae),
	.w6(32'hbbd1d3b7),
	.w7(32'hbbfc7c20),
	.w8(32'hbc17e98d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8ae2f),
	.w1(32'hbc191e28),
	.w2(32'hbb8c9674),
	.w3(32'hbbc43df7),
	.w4(32'hbb9c0f7a),
	.w5(32'h3ad1f87b),
	.w6(32'hbc6b17bd),
	.w7(32'hbba9d78c),
	.w8(32'h3af3d8a2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6cb01),
	.w1(32'h3bbe6c8c),
	.w2(32'hbbf6c021),
	.w3(32'hbb6114ac),
	.w4(32'hbc012f4c),
	.w5(32'hba822baa),
	.w6(32'h3bd14acf),
	.w7(32'hbc23bab6),
	.w8(32'hbc09d84d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeddea8),
	.w1(32'hbb4e9cdf),
	.w2(32'h3bccbedd),
	.w3(32'hb9426020),
	.w4(32'h3b7a312e),
	.w5(32'h3bb56cb6),
	.w6(32'hba9bc253),
	.w7(32'h3bb7c603),
	.w8(32'h3b47769f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854c9c),
	.w1(32'h3a50cfe3),
	.w2(32'h3beef43d),
	.w3(32'h389edfa8),
	.w4(32'h3a8b213a),
	.w5(32'hba5323c2),
	.w6(32'hbaa0906a),
	.w7(32'h3b18036d),
	.w8(32'h3974f41e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3eb5f4),
	.w1(32'hba9e0e0c),
	.w2(32'hbaf21c9a),
	.w3(32'h3bd7fc9d),
	.w4(32'h3b2d2c0b),
	.w5(32'hbc0523d2),
	.w6(32'h3b01d9b9),
	.w7(32'h3a87cc94),
	.w8(32'hbbe88969),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e29a),
	.w1(32'hbaa4a532),
	.w2(32'hbbc72b17),
	.w3(32'hbb4f1e95),
	.w4(32'hb7746b22),
	.w5(32'h3842287e),
	.w6(32'hba9573bd),
	.w7(32'hbab2bdf5),
	.w8(32'hbb61cc52),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ce346),
	.w1(32'hba4bd64c),
	.w2(32'h3b17ee95),
	.w3(32'hbbb30fc6),
	.w4(32'h3babad74),
	.w5(32'h3bf4acf9),
	.w6(32'h3a3d93cf),
	.w7(32'h3b2457f3),
	.w8(32'h3adca7a9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bc454),
	.w1(32'hbb28dbf2),
	.w2(32'hbc21e2f6),
	.w3(32'h3baf0517),
	.w4(32'h3aa36bc6),
	.w5(32'h3cba554f),
	.w6(32'hbadbbd55),
	.w7(32'hbc4e902b),
	.w8(32'h3c4b3b08),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ff28b),
	.w1(32'h3bddf7be),
	.w2(32'hbbec6274),
	.w3(32'h3b8b0e29),
	.w4(32'hbbdc777b),
	.w5(32'hbb1c41e8),
	.w6(32'hbb8d2094),
	.w7(32'hbc115b60),
	.w8(32'hbbe71e7b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ea7eb),
	.w1(32'hbc374023),
	.w2(32'hbc29aed9),
	.w3(32'hbb7e865d),
	.w4(32'hbafd375c),
	.w5(32'h3babb22f),
	.w6(32'hbbd44950),
	.w7(32'hbba637f1),
	.w8(32'hbb842cc7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f295),
	.w1(32'hbc76ffb9),
	.w2(32'hba0848ef),
	.w3(32'h3c06609e),
	.w4(32'hba043fb8),
	.w5(32'h3a99589b),
	.w6(32'hbb3cd24e),
	.w7(32'hb9391338),
	.w8(32'h38b8b2e9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4e39a),
	.w1(32'hba9795e6),
	.w2(32'hbaec320f),
	.w3(32'hba71ac61),
	.w4(32'h3b7f562c),
	.w5(32'hbad4ac85),
	.w6(32'hba66bbf5),
	.w7(32'h3b9bfc80),
	.w8(32'h3b33e7c8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2273a),
	.w1(32'hbb8a636a),
	.w2(32'hbc98798d),
	.w3(32'hbb0a1ec0),
	.w4(32'hbcc50444),
	.w5(32'hbcd61f83),
	.w6(32'h3a1c75cb),
	.w7(32'hbc306380),
	.w8(32'hbc711f0f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc964e55),
	.w1(32'hbc44522f),
	.w2(32'h3b55c308),
	.w3(32'hbc6be93f),
	.w4(32'hbb01f757),
	.w5(32'hbb369402),
	.w6(32'hbbbb2434),
	.w7(32'h3afd3f82),
	.w8(32'hbab319d3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab83a00),
	.w1(32'h3c1f36a0),
	.w2(32'h3b4c0212),
	.w3(32'hbb6dcfc6),
	.w4(32'h3b766396),
	.w5(32'h39d5408e),
	.w6(32'h3bc19893),
	.w7(32'h3bc496e3),
	.w8(32'h3abddec1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d4a2d),
	.w1(32'hba0c709a),
	.w2(32'hbba1ceda),
	.w3(32'h3a8eef86),
	.w4(32'hbc517a3f),
	.w5(32'hbc117803),
	.w6(32'h3a9fac3b),
	.w7(32'hbb12cd72),
	.w8(32'hbb9a2dab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f72af),
	.w1(32'hbb2cfc34),
	.w2(32'hbbbf483b),
	.w3(32'hbc02fa9a),
	.w4(32'hbb8e24e7),
	.w5(32'hbc0cdfe2),
	.w6(32'hbb4acc65),
	.w7(32'h3b4def70),
	.w8(32'hbba109f2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc265635),
	.w1(32'hbb947a98),
	.w2(32'hbb0cc350),
	.w3(32'hbb4ca42f),
	.w4(32'h3b182e50),
	.w5(32'hbc153fc6),
	.w6(32'h3b574936),
	.w7(32'hbb095cfb),
	.w8(32'hbc42dab0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc201801),
	.w1(32'h3af3c5af),
	.w2(32'h3b802d5f),
	.w3(32'hbbbe4676),
	.w4(32'h3aec0a4f),
	.w5(32'h390e09ce),
	.w6(32'hbb0530f2),
	.w7(32'hba100ce0),
	.w8(32'hbb221af8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38e34a),
	.w1(32'hbb8da402),
	.w2(32'hbb481732),
	.w3(32'hbb2773b2),
	.w4(32'hbb833cb5),
	.w5(32'hbbdc11d0),
	.w6(32'hbaed28e3),
	.w7(32'hbc102abd),
	.w8(32'hbc3826b0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51e9b),
	.w1(32'hbbe7f4a7),
	.w2(32'hbbda88d9),
	.w3(32'hbc0646d7),
	.w4(32'hbbd8f426),
	.w5(32'hbbc2ef41),
	.w6(32'hbc634ccf),
	.w7(32'hbc0c0472),
	.w8(32'hbbdd4b80),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89758b),
	.w1(32'hbb6424dc),
	.w2(32'hbc372bad),
	.w3(32'hbb9dba4c),
	.w4(32'hbc2504a8),
	.w5(32'hbb95ce6a),
	.w6(32'hbbe666c0),
	.w7(32'hbc41ceaf),
	.w8(32'hbc05a3cc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c528c),
	.w1(32'hbc8d6cbb),
	.w2(32'h3ba903a0),
	.w3(32'hbc3c18c0),
	.w4(32'hbbebf292),
	.w5(32'hbbc339c5),
	.w6(32'hbc6158a1),
	.w7(32'h3b355110),
	.w8(32'hbbaad787),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6665d3),
	.w1(32'h3b09c0c5),
	.w2(32'h3a48eaf1),
	.w3(32'h3b7c322d),
	.w4(32'h3ae8ea14),
	.w5(32'h3bfc82a7),
	.w6(32'h3bd66267),
	.w7(32'h3728ab5f),
	.w8(32'h39a89238),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba991cf5),
	.w1(32'hba39099b),
	.w2(32'hb98f9abd),
	.w3(32'h3b6aeb00),
	.w4(32'h3b8f4e96),
	.w5(32'h3c4d0967),
	.w6(32'hb981b659),
	.w7(32'h3b2d9db7),
	.w8(32'h3bf22ee9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98473b),
	.w1(32'h3b741bd0),
	.w2(32'hbbaad8fa),
	.w3(32'h3c2a7be7),
	.w4(32'hbb977779),
	.w5(32'h3b319e23),
	.w6(32'h3c1085b9),
	.w7(32'hbbe248da),
	.w8(32'hbbbca6c5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8680a),
	.w1(32'hbc0bd7f1),
	.w2(32'hbb8ead6b),
	.w3(32'h3b554eba),
	.w4(32'hb78a77c1),
	.w5(32'h3b3aee49),
	.w6(32'hbbb212b8),
	.w7(32'hbb910f3c),
	.w8(32'hbb53d138),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955bb6),
	.w1(32'hbc13bba4),
	.w2(32'h3b9814e6),
	.w3(32'h3ab30c8f),
	.w4(32'h3b9b5eb8),
	.w5(32'h3bedd50c),
	.w6(32'hbba852f4),
	.w7(32'h3c00b100),
	.w8(32'h3ae3cc30),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bea15),
	.w1(32'h3b7db5a2),
	.w2(32'hbb6f2ff4),
	.w3(32'h3c2ced55),
	.w4(32'hb9a5a5b3),
	.w5(32'h3932bbad),
	.w6(32'h3b96cc9f),
	.w7(32'hbb1c872d),
	.w8(32'h3ad31543),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70ac39),
	.w1(32'hbc4b6778),
	.w2(32'hbba7244d),
	.w3(32'h3ac6689b),
	.w4(32'hbb1b0d71),
	.w5(32'hbba02eac),
	.w6(32'hbbb09104),
	.w7(32'hbbdbd645),
	.w8(32'hbc2d4b8b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c7a8d),
	.w1(32'hbc5b9fd2),
	.w2(32'hbb203767),
	.w3(32'h3b13a559),
	.w4(32'hbb503211),
	.w5(32'hbb487e92),
	.w6(32'hbbd1559d),
	.w7(32'hbb987888),
	.w8(32'hbb3b9039),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf4506),
	.w1(32'h3a85f35d),
	.w2(32'hbbb7bc78),
	.w3(32'hbb86a7bc),
	.w4(32'h3a1fce7f),
	.w5(32'h3b84681f),
	.w6(32'hbb63133f),
	.w7(32'hbb454cf9),
	.w8(32'h3ba38258),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d86f4),
	.w1(32'h3c0d7890),
	.w2(32'h3ac83570),
	.w3(32'h3b40c728),
	.w4(32'hbb801a17),
	.w5(32'hbb97fa99),
	.w6(32'h3bb42bfb),
	.w7(32'hbb3735b3),
	.w8(32'hb9b33c87),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28ce79),
	.w1(32'hbaf9e1f7),
	.w2(32'h3aa6e49b),
	.w3(32'hbba5aec9),
	.w4(32'h3af3bcb1),
	.w5(32'h3b963e5a),
	.w6(32'hb9dc255d),
	.w7(32'h3a785725),
	.w8(32'h38330a2d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41ba80),
	.w1(32'hb919d809),
	.w2(32'hbb34650c),
	.w3(32'h3b01e21e),
	.w4(32'hb9d5cb8a),
	.w5(32'hba9cea6d),
	.w6(32'hba2ce0af),
	.w7(32'h3b13693c),
	.w8(32'h3a708ff6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a1090),
	.w1(32'hb8835b97),
	.w2(32'hbbc4c7a7),
	.w3(32'hbb217308),
	.w4(32'hba6b01c0),
	.w5(32'h39b125af),
	.w6(32'hbb52a3f8),
	.w7(32'hbb866cbd),
	.w8(32'h3a80f0a8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba769551),
	.w1(32'hbb5f7757),
	.w2(32'hbbecad6c),
	.w3(32'h39121c57),
	.w4(32'hbc19eda4),
	.w5(32'hbc11bf53),
	.w6(32'hbb2802aa),
	.w7(32'hbc3a5f5e),
	.w8(32'hbc583a5b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130675),
	.w1(32'hbb9b487d),
	.w2(32'hba456ce9),
	.w3(32'hbb9dabaa),
	.w4(32'h3c87b37a),
	.w5(32'h3d07ec10),
	.w6(32'hbbfe9777),
	.w7(32'hbb004a20),
	.w8(32'h3c731a32),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92b636),
	.w1(32'h3b8bb291),
	.w2(32'h3a8b2714),
	.w3(32'h3c1eb42f),
	.w4(32'h3aeeaa06),
	.w5(32'h3bd2d39e),
	.w6(32'hbaecbb9e),
	.w7(32'h3a055bad),
	.w8(32'h3a1f1723),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bccb5),
	.w1(32'hb9ad60c5),
	.w2(32'hb702466e),
	.w3(32'h3b4df41c),
	.w4(32'hbc0ccf67),
	.w5(32'hbc5a50c3),
	.w6(32'hb977732d),
	.w7(32'hbbfc57d7),
	.w8(32'hbbc01e5c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b0c86),
	.w1(32'hbb2a3635),
	.w2(32'h3acce060),
	.w3(32'hbc33f8ef),
	.w4(32'hbbd4d3ff),
	.w5(32'h3a39fc54),
	.w6(32'hbc0dc779),
	.w7(32'hbb76fa65),
	.w8(32'hbbd22174),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb501ea3),
	.w1(32'h3b5e5703),
	.w2(32'h3ad4efd6),
	.w3(32'hbbf627a8),
	.w4(32'hbb0b53ce),
	.w5(32'hb98926f3),
	.w6(32'hbb98418e),
	.w7(32'h397e6768),
	.w8(32'hbb07be7f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22c1ed),
	.w1(32'hba6de63f),
	.w2(32'h39da4cdb),
	.w3(32'h3bca39c0),
	.w4(32'hbb47aeb2),
	.w5(32'hbb0c8b06),
	.w6(32'h3b401c68),
	.w7(32'hb924bff5),
	.w8(32'hba181b81),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ff14f),
	.w1(32'h3a62c24c),
	.w2(32'h3ac1f6cd),
	.w3(32'hbbe81f09),
	.w4(32'hba108ed1),
	.w5(32'hba3e825a),
	.w6(32'hbbd28043),
	.w7(32'hbb57881e),
	.w8(32'hba46afbd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule