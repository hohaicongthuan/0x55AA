module layer_8_featuremap_98(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3883d),
	.w1(32'hbb79a370),
	.w2(32'hbc552de5),
	.w3(32'hbb8aec30),
	.w4(32'hbc1a1c8b),
	.w5(32'hbb7e493e),
	.w6(32'hbbc77ce7),
	.w7(32'hbd47dc0e),
	.w8(32'hbc1316f8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28fde),
	.w1(32'hbb212414),
	.w2(32'h3d2a2e12),
	.w3(32'h3c8f4184),
	.w4(32'hbc92e7e2),
	.w5(32'hbd1e9dfb),
	.w6(32'h3d48db3a),
	.w7(32'h3bcdbf7e),
	.w8(32'h3c053151),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d975512),
	.w1(32'h3c14da0c),
	.w2(32'h3c5904f1),
	.w3(32'hbd15a1b4),
	.w4(32'hbc4b1394),
	.w5(32'hbcd3262d),
	.w6(32'hbc522752),
	.w7(32'hbba94849),
	.w8(32'hbc190ec0),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d34f278),
	.w1(32'h3c4e3fae),
	.w2(32'hbd380149),
	.w3(32'hbcac70fb),
	.w4(32'h3ab63471),
	.w5(32'h3cda66b3),
	.w6(32'hbc5e67f9),
	.w7(32'h3c0627c6),
	.w8(32'h3a1d2c61),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4de70),
	.w1(32'hbbdb0b06),
	.w2(32'hbc82078e),
	.w3(32'h3c71e8c1),
	.w4(32'hbca7bf21),
	.w5(32'hbc9c6006),
	.w6(32'hbc81ca26),
	.w7(32'hbc462a59),
	.w8(32'hbac4a577),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e6c6),
	.w1(32'h3c97a946),
	.w2(32'h3d2c83fa),
	.w3(32'hbb9b5377),
	.w4(32'h3cadd4b8),
	.w5(32'h3d1b1d55),
	.w6(32'h3c98cb2f),
	.w7(32'h3d1b4a6f),
	.w8(32'h3c4f8c81),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f5fa4),
	.w1(32'hbb3cfe38),
	.w2(32'hbc244b7d),
	.w3(32'hbc0bdf88),
	.w4(32'h3c15803d),
	.w5(32'h3cab7fb2),
	.w6(32'hbcd0e93a),
	.w7(32'hba9b6f6d),
	.w8(32'h3c01f6fd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f9388),
	.w1(32'hbc808ba3),
	.w2(32'hbb14bc63),
	.w3(32'h3ca3c264),
	.w4(32'hbbbab482),
	.w5(32'hbca9d9c4),
	.w6(32'hbc50922b),
	.w7(32'hbaad54f6),
	.w8(32'hb8b34cda),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061e47),
	.w1(32'hbb6a0d3e),
	.w2(32'hbc96fc5d),
	.w3(32'hbd032d43),
	.w4(32'hbc6aaf5d),
	.w5(32'h3cb45ba6),
	.w6(32'hbc8c0ca5),
	.w7(32'hbcd1cfd4),
	.w8(32'hbc43121a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32a092),
	.w1(32'h3c9886d7),
	.w2(32'hbb652f20),
	.w3(32'h3d1263aa),
	.w4(32'hbbea03eb),
	.w5(32'h3c320c66),
	.w6(32'h3c23aef5),
	.w7(32'h3c6f1170),
	.w8(32'hbc3be485),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f95a),
	.w1(32'h3b46ba03),
	.w2(32'hbcc40c8c),
	.w3(32'h3be75693),
	.w4(32'hbc31b372),
	.w5(32'hbc7298a9),
	.w6(32'hbcd64028),
	.w7(32'hbd06e27d),
	.w8(32'hbb89d7b8),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3069),
	.w1(32'h3d118a88),
	.w2(32'h3c4837c5),
	.w3(32'h36ff9468),
	.w4(32'hbc55c046),
	.w5(32'hbc8d6111),
	.w6(32'h3cb504f9),
	.w7(32'hbbed7d5f),
	.w8(32'hbc5baaad),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed7b32),
	.w1(32'hbc0a65e7),
	.w2(32'hba3403f6),
	.w3(32'hbb363777),
	.w4(32'hbb89f603),
	.w5(32'h39d24fe4),
	.w6(32'h3b8b37bc),
	.w7(32'h3bb17d56),
	.w8(32'h3bb94234),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a941d6c),
	.w1(32'h39a9006b),
	.w2(32'h39254660),
	.w3(32'h3a9de019),
	.w4(32'h39f5790b),
	.w5(32'h3a360327),
	.w6(32'h3ab6366e),
	.w7(32'h3a0bfeb6),
	.w8(32'h39f610df),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997755b),
	.w1(32'h391f44d7),
	.w2(32'h3882e35a),
	.w3(32'h392655c3),
	.w4(32'h389ba1ba),
	.w5(32'h386c24b2),
	.w6(32'hb75bac5b),
	.w7(32'hb9161dfc),
	.w8(32'hb780c3ad),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39655096),
	.w1(32'h35bffe90),
	.w2(32'hb981d253),
	.w3(32'hba67c930),
	.w4(32'hba949177),
	.w5(32'hba2888e1),
	.w6(32'hba2f5228),
	.w7(32'hb98b535d),
	.w8(32'h37939543),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b5ad5f),
	.w1(32'h3b90046c),
	.w2(32'h3b821bd9),
	.w3(32'h3a218bd5),
	.w4(32'h3b89f064),
	.w5(32'h3b478802),
	.w6(32'hb9b43faa),
	.w7(32'h38cc3a3e),
	.w8(32'hbac20c65),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40222e),
	.w1(32'h3b9f16de),
	.w2(32'hbb877c44),
	.w3(32'hbae75549),
	.w4(32'hbbd28913),
	.w5(32'hbbb9dc52),
	.w6(32'hbb32638d),
	.w7(32'hbc0fc558),
	.w8(32'hbba81ae8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6655ab),
	.w1(32'h3d2c8caa),
	.w2(32'h3c47dd16),
	.w3(32'hbbe7a397),
	.w4(32'hba35af9a),
	.w5(32'h3c0b78f8),
	.w6(32'hbc69bfb8),
	.w7(32'hbcdf19a2),
	.w8(32'h3c9f9668),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdc3a9),
	.w1(32'hbb8ce5a1),
	.w2(32'hbbe020b1),
	.w3(32'h3749c57b),
	.w4(32'hbbd1984b),
	.w5(32'hb8f7ff1f),
	.w6(32'h3b9e1de3),
	.w7(32'h3a9efea9),
	.w8(32'h3bd24754),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad1718),
	.w1(32'h3bc76654),
	.w2(32'h3c0359cb),
	.w3(32'hbbb5be29),
	.w4(32'h3c2fac7e),
	.w5(32'h3c770f48),
	.w6(32'h3c8869f4),
	.w7(32'h3c37dc79),
	.w8(32'h3bd33dd4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be211ba),
	.w1(32'hbb10300d),
	.w2(32'hba678f7f),
	.w3(32'h3c45c369),
	.w4(32'h3bb7d496),
	.w5(32'h3b5d11d6),
	.w6(32'h3c88df94),
	.w7(32'h3c137f67),
	.w8(32'h3b9608ae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4f6f8),
	.w1(32'hbb904d87),
	.w2(32'hbd0619e1),
	.w3(32'hbc984025),
	.w4(32'hbd0f9954),
	.w5(32'hbd129ccd),
	.w6(32'hbc88dcd5),
	.w7(32'hbd3eb525),
	.w8(32'hbce4ed84),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eaa4c),
	.w1(32'hbb42127b),
	.w2(32'hbb065c1a),
	.w3(32'h39020b10),
	.w4(32'h3977d827),
	.w5(32'h3a819266),
	.w6(32'hb94714eb),
	.w7(32'h3a942e13),
	.w8(32'h3b423278),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b302b),
	.w1(32'h3b221cb8),
	.w2(32'h3c08846f),
	.w3(32'h3b746af8),
	.w4(32'h3a78d436),
	.w5(32'h3bdd0f05),
	.w6(32'h3b9532e6),
	.w7(32'h3a4e1663),
	.w8(32'h3b55bcce),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf3aaf),
	.w1(32'h3c0b2e0e),
	.w2(32'hbb91606b),
	.w3(32'hbbd745f8),
	.w4(32'hbc0f05c8),
	.w5(32'hbc22f03c),
	.w6(32'hbc3b5443),
	.w7(32'hbcabace1),
	.w8(32'hbc1390db),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c84e7),
	.w1(32'h3a06be59),
	.w2(32'h3a810e98),
	.w3(32'hba977cc0),
	.w4(32'h382be701),
	.w5(32'h3a5633f2),
	.w6(32'hbabc6c17),
	.w7(32'hb9edb13f),
	.w8(32'h3a0a5b3b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f36d0),
	.w1(32'h3dae55b9),
	.w2(32'h3cb224ac),
	.w3(32'hba34697c),
	.w4(32'h3db0a7c1),
	.w5(32'h3d8ad203),
	.w6(32'h3bdeddda),
	.w7(32'hbcec5716),
	.w8(32'h3c4a126c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a4f84),
	.w1(32'h3ba1490d),
	.w2(32'hba4e7569),
	.w3(32'hbb4736a5),
	.w4(32'hbc09dde5),
	.w5(32'hbbc7e66d),
	.w6(32'hbbb00011),
	.w7(32'hbc24063f),
	.w8(32'hbb7d6a29),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010faa),
	.w1(32'hba3dac0b),
	.w2(32'hbaac4c90),
	.w3(32'h39d0942f),
	.w4(32'hbae217cd),
	.w5(32'hbaeed77f),
	.w6(32'h3a3d4d99),
	.w7(32'hbac099cc),
	.w8(32'hba992af4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485931),
	.w1(32'h3b12ba83),
	.w2(32'h3b55ba45),
	.w3(32'hb9ddf3dd),
	.w4(32'h3b88f860),
	.w5(32'h3b8becac),
	.w6(32'h3ae70ded),
	.w7(32'h3b9c68cd),
	.w8(32'h3b8bb8b2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057b58),
	.w1(32'hba96b5cc),
	.w2(32'hbb7c7d03),
	.w3(32'hb9a55cbf),
	.w4(32'h3af2d7f6),
	.w5(32'h3ac3b18d),
	.w6(32'h3b92bb01),
	.w7(32'h3b3d98b4),
	.w8(32'h3b16c561),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392100f6),
	.w1(32'h38c23981),
	.w2(32'hb896a245),
	.w3(32'h3993d23b),
	.w4(32'h3919c2fa),
	.w5(32'h38773ead),
	.w6(32'h38be8d60),
	.w7(32'h3933a5b8),
	.w8(32'hb8091fc6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aae7b7),
	.w1(32'hb69f5344),
	.w2(32'hb944700a),
	.w3(32'h38929d11),
	.w4(32'h39110112),
	.w5(32'hb9010baa),
	.w6(32'h38915e9d),
	.w7(32'h38272ab4),
	.w8(32'hb891c1f7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c1b3a),
	.w1(32'hbb102207),
	.w2(32'h3b2528c5),
	.w3(32'h3b32063f),
	.w4(32'h3b94344c),
	.w5(32'h3c06c567),
	.w6(32'h3c8c839a),
	.w7(32'h3c892fee),
	.w8(32'h3c44a73e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9a388),
	.w1(32'h3c6c0a8e),
	.w2(32'h3c19dc8a),
	.w3(32'h39811bd1),
	.w4(32'h39ae368b),
	.w5(32'h3ba99da0),
	.w6(32'hb8f4ffc5),
	.w7(32'hbbac51a1),
	.w8(32'h3b6cb562),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c23c40),
	.w1(32'h391bc743),
	.w2(32'h39854226),
	.w3(32'hba00a179),
	.w4(32'hb9f46d8d),
	.w5(32'h3903e2bf),
	.w6(32'hba49e3c1),
	.w7(32'hba53e74f),
	.w8(32'hb8f0038c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1d13),
	.w1(32'hbadc671b),
	.w2(32'hbbb5abef),
	.w3(32'h3ab84242),
	.w4(32'hbb776c8e),
	.w5(32'hbbbb43a5),
	.w6(32'h3b156d41),
	.w7(32'hbaee932f),
	.w8(32'hbb5f5635),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392222eb),
	.w1(32'hb90d991c),
	.w2(32'hb9cb158d),
	.w3(32'h39d38e33),
	.w4(32'hb869fc9e),
	.w5(32'hba11bc3d),
	.w6(32'h38bc715b),
	.w7(32'hb9382f35),
	.w8(32'hb9feb947),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957d165),
	.w1(32'h38e6a5cc),
	.w2(32'h3903015d),
	.w3(32'h3aa21792),
	.w4(32'h3aa25352),
	.w5(32'h39ed5217),
	.w6(32'h3a3e1ab4),
	.w7(32'h3935b19f),
	.w8(32'hba185def),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c726077),
	.w1(32'h3b01584c),
	.w2(32'hbc88b17b),
	.w3(32'hbc4b4a79),
	.w4(32'hbcd7877e),
	.w5(32'hbcc5e42f),
	.w6(32'hbc85f68c),
	.w7(32'hbcb57c7d),
	.w8(32'hbc1d6c23),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe6816),
	.w1(32'h3b81406f),
	.w2(32'h3b482bc2),
	.w3(32'hbab656c7),
	.w4(32'h3b3d97bd),
	.w5(32'h3b419c86),
	.w6(32'hba85c82c),
	.w7(32'h3999a56c),
	.w8(32'h3b3538c0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3795a2ce),
	.w1(32'h3a94361c),
	.w2(32'h3ade475e),
	.w3(32'h3a2916a8),
	.w4(32'h3a98714d),
	.w5(32'h3b025c26),
	.w6(32'h3af96ef7),
	.w7(32'h3b110c28),
	.w8(32'h3ada776b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a57bc6),
	.w1(32'h3b265876),
	.w2(32'hbb530c83),
	.w3(32'hbab5a645),
	.w4(32'hb9f71fc3),
	.w5(32'hbb0868b4),
	.w6(32'hbb72e72b),
	.w7(32'hbc07459c),
	.w8(32'hbb4aed84),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e99f1),
	.w1(32'h3c23696b),
	.w2(32'hbbce6b45),
	.w3(32'hb9f5098b),
	.w4(32'h38936522),
	.w5(32'hbb0ecfb5),
	.w6(32'hbbc86cf9),
	.w7(32'hbc6ad9c7),
	.w8(32'hbb668f53),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe8441),
	.w1(32'h3bddd067),
	.w2(32'h3ad69de5),
	.w3(32'hba363e98),
	.w4(32'hb964393d),
	.w5(32'hb9f93764),
	.w6(32'h3a018a65),
	.w7(32'h3afcec5f),
	.w8(32'h3ba9df51),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377f6038),
	.w1(32'h3833a3e6),
	.w2(32'hb878a26b),
	.w3(32'hb8734a0d),
	.w4(32'hb80767d0),
	.w5(32'hb8e1b164),
	.w6(32'hb858c1a7),
	.w7(32'hb8e259a9),
	.w8(32'hb8b78592),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28631e),
	.w1(32'h3c011b86),
	.w2(32'hbbc7a81c),
	.w3(32'h3b635b88),
	.w4(32'hbb3cd170),
	.w5(32'hbbdd8c04),
	.w6(32'h3ac94c54),
	.w7(32'hbc6c6a8f),
	.w8(32'hbbcb6110),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ce329),
	.w1(32'hbb5122e7),
	.w2(32'hbaddfa2c),
	.w3(32'hbb0442ae),
	.w4(32'hbb83280c),
	.w5(32'hbaf02235),
	.w6(32'hb9afc7d0),
	.w7(32'hbb1c0d06),
	.w8(32'hb8ea263f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1feb09),
	.w1(32'h3b31daf7),
	.w2(32'hbc02c4e6),
	.w3(32'h3907268f),
	.w4(32'hbbd158ef),
	.w5(32'hbbfcc624),
	.w6(32'hbc3fbf19),
	.w7(32'hbc5f3f84),
	.w8(32'hbbeefa5c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cfd22),
	.w1(32'hbbb92e2a),
	.w2(32'hbba7721e),
	.w3(32'h3b2f1c46),
	.w4(32'hbb883e17),
	.w5(32'hbb1039c4),
	.w6(32'h3c5e43d6),
	.w7(32'h3c0e947f),
	.w8(32'h3b9c5445),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d110f8d),
	.w1(32'h3cdacbb3),
	.w2(32'h3c0029c3),
	.w3(32'h3cd38f8b),
	.w4(32'h3ca3bf4e),
	.w5(32'h3c118d0c),
	.w6(32'hbc88d0f2),
	.w7(32'hbc9f5e12),
	.w8(32'h3c3c8c65),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9bfa),
	.w1(32'hbb56b2d8),
	.w2(32'hbb536bf4),
	.w3(32'hb9eed70e),
	.w4(32'hbbcaf9dc),
	.w5(32'hbb43f7b5),
	.w6(32'hbc037119),
	.w7(32'hbc1008f0),
	.w8(32'hba400625),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1567a9),
	.w1(32'h3b31e0ea),
	.w2(32'hbbcd3eb7),
	.w3(32'hbb122fa0),
	.w4(32'hbc861515),
	.w5(32'hbc8abdbe),
	.w6(32'h3a4324e4),
	.w7(32'hbbd9cccd),
	.w8(32'hbba4df69),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39031537),
	.w1(32'h3801e53c),
	.w2(32'hb7806498),
	.w3(32'h38817b81),
	.w4(32'hb83022c4),
	.w5(32'hb777bee0),
	.w6(32'hb881b79a),
	.w7(32'hb8dc1ee2),
	.w8(32'hb9536040),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66e025),
	.w1(32'h3cafd2dd),
	.w2(32'h3b38629e),
	.w3(32'hbc0d282a),
	.w4(32'hbc405e4b),
	.w5(32'hbc53fb47),
	.w6(32'h3c868556),
	.w7(32'hbbbd5f72),
	.w8(32'hb9f7e9e9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c1e7c),
	.w1(32'hbb7ce518),
	.w2(32'hb9f4d648),
	.w3(32'hb7596e5e),
	.w4(32'h39f573f9),
	.w5(32'h3b58a041),
	.w6(32'h3b87d593),
	.w7(32'h3b300661),
	.w8(32'hb9254c55),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c4b4a),
	.w1(32'h3c292050),
	.w2(32'h3b88874c),
	.w3(32'h3bb515f3),
	.w4(32'h3b6c1fae),
	.w5(32'h3accdcf8),
	.w6(32'hbb8a1e3f),
	.w7(32'hbb9a6b69),
	.w8(32'h3b59d5eb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a857a21),
	.w1(32'h3ba45d54),
	.w2(32'hbaea86fa),
	.w3(32'h3b9bab14),
	.w4(32'h3b9a4d73),
	.w5(32'hbac6cbf9),
	.w6(32'h3b145129),
	.w7(32'hbbbc1eab),
	.w8(32'hbbce63fd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19fbb5),
	.w1(32'h3a0877bd),
	.w2(32'hbc0e74b3),
	.w3(32'h3bee3cf4),
	.w4(32'hb881d4dd),
	.w5(32'hbba325ce),
	.w6(32'h3baa47e5),
	.w7(32'hb9b912e1),
	.w8(32'hbbb39991),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24cfc7),
	.w1(32'h39dc96e3),
	.w2(32'h3ab4be66),
	.w3(32'hb9341257),
	.w4(32'hb96abf75),
	.w5(32'h3a25f24f),
	.w6(32'hba04641d),
	.w7(32'hb9286b91),
	.w8(32'h3a5f48ae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df09b3),
	.w1(32'h37f34bf1),
	.w2(32'hba552634),
	.w3(32'h3a153827),
	.w4(32'hb90f1344),
	.w5(32'hbad8e5fc),
	.w6(32'h39625c68),
	.w7(32'hba8575f6),
	.w8(32'hbb016ae3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc8b30c),
	.w1(32'h3c738d72),
	.w2(32'h3b583313),
	.w3(32'hbb9840fb),
	.w4(32'hbc866ac6),
	.w5(32'hbc2427b1),
	.w6(32'hbbb38082),
	.w7(32'hbc22cb56),
	.w8(32'hb838d884),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa77b67),
	.w1(32'hba574d82),
	.w2(32'h3b7049a7),
	.w3(32'h3b1ec343),
	.w4(32'h3a92b29a),
	.w5(32'h3b317c78),
	.w6(32'hbae5934c),
	.w7(32'hbac053f0),
	.w8(32'h3b711c1c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15e51c),
	.w1(32'hbb03cb31),
	.w2(32'hba84bddf),
	.w3(32'hbb3e6080),
	.w4(32'hbb24fa5d),
	.w5(32'hbadbea0c),
	.w6(32'hbb3c8ee6),
	.w7(32'hbb077a8e),
	.w8(32'hba9dd828),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabf0cd),
	.w1(32'h3b3f221a),
	.w2(32'hb969788f),
	.w3(32'hbacf795f),
	.w4(32'hbb1947d3),
	.w5(32'h37311d51),
	.w6(32'hbb7558bb),
	.w7(32'hbc01a29d),
	.w8(32'hbb120eeb),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295a31),
	.w1(32'h3a95e98d),
	.w2(32'hbaa2579f),
	.w3(32'h3ba56a33),
	.w4(32'hb9673e13),
	.w5(32'hbaebe3ca),
	.w6(32'h3b7251a5),
	.w7(32'h39004352),
	.w8(32'h3a89681f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62aeec),
	.w1(32'h3bf50b22),
	.w2(32'h3bc70c29),
	.w3(32'hbbdd1a52),
	.w4(32'hbb91b27f),
	.w5(32'h3b2ebf86),
	.w6(32'h3abadb83),
	.w7(32'hbb200e1f),
	.w8(32'h3bd1a223),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d2cfd),
	.w1(32'h38db05c7),
	.w2(32'h37634cad),
	.w3(32'hbb085954),
	.w4(32'hba9f7ce8),
	.w5(32'hba136f20),
	.w6(32'hbb425bc9),
	.w7(32'hbafbc6e8),
	.w8(32'hba789a8d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af94f6e),
	.w1(32'h3ca1a061),
	.w2(32'hbc76498e),
	.w3(32'h3c44e438),
	.w4(32'h3c85f57e),
	.w5(32'hbb5d6520),
	.w6(32'h3c1c962b),
	.w7(32'hbca23a85),
	.w8(32'hbcb5984b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89815d),
	.w1(32'hb9cfb45a),
	.w2(32'hb9750639),
	.w3(32'hba20113e),
	.w4(32'hb99e12d2),
	.w5(32'hb81c6065),
	.w6(32'hba4ba09c),
	.w7(32'hb97ebe63),
	.w8(32'hb9b5a261),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cf39),
	.w1(32'hbb695004),
	.w2(32'hbbeb8337),
	.w3(32'h3ac9c870),
	.w4(32'hbb85a0e4),
	.w5(32'hbb84845d),
	.w6(32'h3a57fee2),
	.w7(32'hbb9bc445),
	.w8(32'hbb62e1e1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba134927),
	.w1(32'hba73516c),
	.w2(32'hba9b8183),
	.w3(32'hbae5a9c4),
	.w4(32'hbaee7693),
	.w5(32'hbad176f1),
	.w6(32'hbb2563d2),
	.w7(32'hbb18150b),
	.w8(32'hbab88f43),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58fb43),
	.w1(32'h3be7fc4b),
	.w2(32'hbbc813bb),
	.w3(32'hbbe63b61),
	.w4(32'hbc5c273a),
	.w5(32'hbc298c7b),
	.w6(32'h3b733351),
	.w7(32'hbba87055),
	.w8(32'hbb4c8003),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb716b21d),
	.w1(32'hb8e37154),
	.w2(32'h38b7ecb2),
	.w3(32'hb8abc5e8),
	.w4(32'hb85adfbc),
	.w5(32'hb7ad7abc),
	.w6(32'hb709d020),
	.w7(32'hb8e63e6d),
	.w8(32'h384a1fbb),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79d8074),
	.w1(32'h3a50ef39),
	.w2(32'h3b869904),
	.w3(32'hbb77bd30),
	.w4(32'hbb208a81),
	.w5(32'h3ab31edd),
	.w6(32'hbb654bd6),
	.w7(32'hbb3e058f),
	.w8(32'h399fa693),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387ec687),
	.w1(32'h39798d18),
	.w2(32'h3bda8397),
	.w3(32'hb8c771ee),
	.w4(32'h3a8ed3cb),
	.w5(32'hbbc2a378),
	.w6(32'hb98e2561),
	.w7(32'h378797e1),
	.w8(32'hbb620ba6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce024be),
	.w1(32'h3b86e7d9),
	.w2(32'hba02c7ed),
	.w3(32'hbba50afe),
	.w4(32'hbc1741e1),
	.w5(32'hbc0849d3),
	.w6(32'hbc2d2bab),
	.w7(32'hbc912b95),
	.w8(32'hbb5b12b0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8403ba),
	.w1(32'h3be0a62c),
	.w2(32'hbb2ff12c),
	.w3(32'hba9682ad),
	.w4(32'hbba62119),
	.w5(32'hbc44f965),
	.w6(32'h3bfee44c),
	.w7(32'hba40b9ed),
	.w8(32'h3a8044c3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ca3b5),
	.w1(32'hbb5c0e70),
	.w2(32'h3b6f1926),
	.w3(32'hba38c920),
	.w4(32'hbbfb6263),
	.w5(32'hbc24f8c9),
	.w6(32'hba39f566),
	.w7(32'hbad59976),
	.w8(32'hbb5052db),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa431ff),
	.w1(32'hbb8fc288),
	.w2(32'hbb4b1541),
	.w3(32'hbbbbc6f6),
	.w4(32'h3b298029),
	.w5(32'hbc09c2fe),
	.w6(32'hbbdb508b),
	.w7(32'hbb925eff),
	.w8(32'hbc2d8375),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9969e),
	.w1(32'h3c089391),
	.w2(32'hbcc0092d),
	.w3(32'hbb3f0cc1),
	.w4(32'h3bff87c9),
	.w5(32'hbb425af8),
	.w6(32'hbaff854a),
	.w7(32'h3c222e5d),
	.w8(32'hbbb78237),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e5c93),
	.w1(32'h3a905d31),
	.w2(32'hbbb00eb4),
	.w3(32'hbc013963),
	.w4(32'hbb707395),
	.w5(32'hbc4c5a53),
	.w6(32'hbcce3d96),
	.w7(32'hbc3a01e9),
	.w8(32'hbc6fbc60),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4eaa20),
	.w1(32'h3ce07b37),
	.w2(32'hbc172966),
	.w3(32'hbb12608d),
	.w4(32'hbd17f82f),
	.w5(32'hbd110085),
	.w6(32'hbc6f7a25),
	.w7(32'hbb23cb86),
	.w8(32'hbc93f91e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d207969),
	.w1(32'h3cce340e),
	.w2(32'hbc863e36),
	.w3(32'hbc3179e0),
	.w4(32'hbcc21b36),
	.w5(32'hbc393c18),
	.w6(32'hbd076c78),
	.w7(32'hbd80ef1f),
	.w8(32'hbc951f71),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d7d9c),
	.w1(32'h3b13c9f5),
	.w2(32'hbb697c7e),
	.w3(32'h3b07ef43),
	.w4(32'hbc25c69a),
	.w5(32'hbceb6e72),
	.w6(32'h3a9e0e3c),
	.w7(32'hbc900e6f),
	.w8(32'hbbe16a28),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95e5b3),
	.w1(32'hbc9093f6),
	.w2(32'hbc30d84e),
	.w3(32'hbc8a36c0),
	.w4(32'hbbbbb399),
	.w5(32'hba84dce6),
	.w6(32'h3af17261),
	.w7(32'hbc0f1e1c),
	.w8(32'hbbcb76bb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdfc664),
	.w1(32'hbc988550),
	.w2(32'hbc18a3d7),
	.w3(32'hbc3ddf08),
	.w4(32'h3bf068e5),
	.w5(32'h3abe1264),
	.w6(32'hbc0fc70b),
	.w7(32'h3ba0b10d),
	.w8(32'hb9f87705),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b02bb),
	.w1(32'hbb0a13c6),
	.w2(32'hb7fa80f1),
	.w3(32'hbbcbc5cc),
	.w4(32'hbad271af),
	.w5(32'hba3a6f99),
	.w6(32'hbb19db72),
	.w7(32'hb9842b02),
	.w8(32'h3b6ebdd5),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf525f9),
	.w1(32'hbc1f98f2),
	.w2(32'h3bff8a82),
	.w3(32'h3b903135),
	.w4(32'h3b3d0693),
	.w5(32'hbbf1cf0d),
	.w6(32'h3a6b913c),
	.w7(32'hbb923d21),
	.w8(32'h3b6ea960),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3ca6f),
	.w1(32'h3bb8e551),
	.w2(32'h3bd6b1cc),
	.w3(32'hbaae69e4),
	.w4(32'h3ace9b83),
	.w5(32'hbb1e3f57),
	.w6(32'h3c46e0f7),
	.w7(32'h3c6bf061),
	.w8(32'hbc2ec6f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e1d05),
	.w1(32'h3c065d0e),
	.w2(32'hbc3a2d49),
	.w3(32'hbbadfe1b),
	.w4(32'hbc72d3ce),
	.w5(32'hba1e4fd3),
	.w6(32'hbbe497cd),
	.w7(32'hbc2ba91c),
	.w8(32'hbc711c6a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0ac1c7),
	.w1(32'hbbf8a4f4),
	.w2(32'hbc9a9a91),
	.w3(32'h3bbbb49a),
	.w4(32'hbc455813),
	.w5(32'h3c00d7ec),
	.w6(32'h3c887a40),
	.w7(32'hbc1f4038),
	.w8(32'hbc33732b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc61b4),
	.w1(32'h3c58e6d3),
	.w2(32'hbb0b1845),
	.w3(32'h3c281000),
	.w4(32'hbbebf50a),
	.w5(32'hbb8edcc1),
	.w6(32'hbbcf372a),
	.w7(32'hbc5ea138),
	.w8(32'h3b5ef828),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a015e7d),
	.w1(32'h3aaf38af),
	.w2(32'hbb83696e),
	.w3(32'hbb05c7ff),
	.w4(32'hbbab4a63),
	.w5(32'h3a38ecb1),
	.w6(32'h3c273fa8),
	.w7(32'h3b7af8fc),
	.w8(32'h3bcd73b1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c242a29),
	.w1(32'h3c5e3d91),
	.w2(32'h3ce4e85b),
	.w3(32'h3c1a72b6),
	.w4(32'hbc4ac9d2),
	.w5(32'hbc690d9d),
	.w6(32'h3c3db639),
	.w7(32'hbcf23173),
	.w8(32'hbd2827c1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4da61e),
	.w1(32'hbb1515a4),
	.w2(32'h3cb86afd),
	.w3(32'hbcb8c8a2),
	.w4(32'hbd0d1da1),
	.w5(32'hbc88886d),
	.w6(32'hbd116f09),
	.w7(32'hbc5ce097),
	.w8(32'h3d62f211),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7895d1),
	.w1(32'h3bbe9574),
	.w2(32'hbc2bd51d),
	.w3(32'hbc89e5bd),
	.w4(32'h3b8254cd),
	.w5(32'hbbed9f35),
	.w6(32'hbb03d7a1),
	.w7(32'h3b05c812),
	.w8(32'h3c38e787),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5f87c),
	.w1(32'hba44bcf0),
	.w2(32'h3955c4dd),
	.w3(32'hbc0d78ee),
	.w4(32'h3c83309b),
	.w5(32'h3c16c1dc),
	.w6(32'h3b1e86a0),
	.w7(32'h3c68500d),
	.w8(32'h3b8af0be),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb67dd),
	.w1(32'hbc171b75),
	.w2(32'h3c796a89),
	.w3(32'hbac5ec98),
	.w4(32'h3c2e033e),
	.w5(32'h3be8c580),
	.w6(32'h3af85faf),
	.w7(32'h3cfac1c9),
	.w8(32'h3c06fb7e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb907),
	.w1(32'hbcb9938f),
	.w2(32'hba7925d1),
	.w3(32'hbb8c2261),
	.w4(32'hb9676d0d),
	.w5(32'h3b9d8469),
	.w6(32'hbc2b7bea),
	.w7(32'hbcbe92e4),
	.w8(32'hbb88be6f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c923121),
	.w1(32'hbcd50309),
	.w2(32'hbc3560a3),
	.w3(32'h3b33ffc6),
	.w4(32'hbc0fd6b3),
	.w5(32'hbaee3a12),
	.w6(32'hbc500eb8),
	.w7(32'hbbdda22b),
	.w8(32'h3b8ca39c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc465706),
	.w1(32'hbaa8e75b),
	.w2(32'h3c5ebd94),
	.w3(32'hbad390b3),
	.w4(32'hbca31e80),
	.w5(32'hbcc4a699),
	.w6(32'h3b9dc081),
	.w7(32'hbb58f101),
	.w8(32'hbd19e408),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b8e75),
	.w1(32'h3c68efb3),
	.w2(32'hbc89219a),
	.w3(32'hbb5c4723),
	.w4(32'hbbb16b51),
	.w5(32'hbc494d2a),
	.w6(32'hbcc67f94),
	.w7(32'h3c1264ed),
	.w8(32'h3a843feb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cbfa7),
	.w1(32'hbbcea0fc),
	.w2(32'h3c111a56),
	.w3(32'hbc204ebf),
	.w4(32'hbba978b4),
	.w5(32'hbc337c49),
	.w6(32'h3b66ce6f),
	.w7(32'h3bab8572),
	.w8(32'hbc6aff70),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96e01f),
	.w1(32'h3c9b6bd4),
	.w2(32'hb87cb3a1),
	.w3(32'hbbc22444),
	.w4(32'h3b956962),
	.w5(32'h3b54e0d2),
	.w6(32'hbbf7f146),
	.w7(32'hbcc2ea59),
	.w8(32'h3aef69ee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf155e),
	.w1(32'h3b843371),
	.w2(32'hbbdb0f44),
	.w3(32'hbaada2ad),
	.w4(32'hbc4e572a),
	.w5(32'h3a0c8edc),
	.w6(32'hbc360313),
	.w7(32'h3a2b697e),
	.w8(32'hbbe6b401),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b0c7e),
	.w1(32'hbc0c3f59),
	.w2(32'h3b9126e6),
	.w3(32'hbaca25b8),
	.w4(32'hba20549e),
	.w5(32'hbbf49e56),
	.w6(32'h3b8f8155),
	.w7(32'h3b177724),
	.w8(32'h3807c7cb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83b628),
	.w1(32'hbc10bd3a),
	.w2(32'h3bce9563),
	.w3(32'hbb668c6c),
	.w4(32'hbc464b4d),
	.w5(32'hbabc1037),
	.w6(32'hbb3ee18f),
	.w7(32'h3b98836b),
	.w8(32'hbc14f646),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc29b2),
	.w1(32'hbbf668dd),
	.w2(32'hbae82148),
	.w3(32'h3c0bb407),
	.w4(32'hba477154),
	.w5(32'hb9b08526),
	.w6(32'hbb53185c),
	.w7(32'h3b1129b2),
	.w8(32'hbc388dac),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac498a5),
	.w1(32'hbb7b1e38),
	.w2(32'h3c25ca22),
	.w3(32'hbbc30486),
	.w4(32'hbcb30bab),
	.w5(32'hbc036441),
	.w6(32'hbbf50e44),
	.w7(32'h3bb52233),
	.w8(32'h3b0f023c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabf2d5),
	.w1(32'hbb269275),
	.w2(32'h3af217f7),
	.w3(32'hbbfe3a77),
	.w4(32'h3c190d24),
	.w5(32'h3c8e2f63),
	.w6(32'hbc6fb6b8),
	.w7(32'h3b2e84da),
	.w8(32'h3c876dbd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2941a7),
	.w1(32'hbce72324),
	.w2(32'hbaa8a1e9),
	.w3(32'hbc2778e2),
	.w4(32'hbc55563e),
	.w5(32'hbc717618),
	.w6(32'hba92b6b6),
	.w7(32'hbbd831d5),
	.w8(32'hbc558549),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32d284),
	.w1(32'hb95f7d73),
	.w2(32'h3cdd0d20),
	.w3(32'hbc2cef9f),
	.w4(32'hbd0aa0de),
	.w5(32'hbd003d7f),
	.w6(32'hbc386def),
	.w7(32'hbcaa79ca),
	.w8(32'hbcd9f042),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57739c),
	.w1(32'h3c6b3eee),
	.w2(32'hbcbe67e6),
	.w3(32'hbce840eb),
	.w4(32'h3aa42cff),
	.w5(32'h3c5c8ec2),
	.w6(32'hbce883f1),
	.w7(32'h3c2fc50e),
	.w8(32'h3d49cdf7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ee638),
	.w1(32'h3bac0897),
	.w2(32'h3b98d60b),
	.w3(32'h3c6c8a6f),
	.w4(32'hbbcd690a),
	.w5(32'hbbc085b3),
	.w6(32'h3cb35b0f),
	.w7(32'hbc2ceadc),
	.w8(32'h3c291ec4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c41345),
	.w1(32'h3ca3a061),
	.w2(32'h3be11faf),
	.w3(32'hbabcdc3f),
	.w4(32'h3bb8df54),
	.w5(32'h38dae263),
	.w6(32'h3cb516c6),
	.w7(32'hbc1781a2),
	.w8(32'hbc2fae03),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c431021),
	.w1(32'h3c87fd4a),
	.w2(32'h3c207b30),
	.w3(32'hbbd9b318),
	.w4(32'hb8f011c7),
	.w5(32'hbb873e3e),
	.w6(32'hbb8e8552),
	.w7(32'hbb9f022c),
	.w8(32'hbb57f83d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68a88c),
	.w1(32'hbb9bf650),
	.w2(32'h3c0df693),
	.w3(32'hbaf46370),
	.w4(32'hbc32840f),
	.w5(32'hbc53a4ee),
	.w6(32'hbb34feea),
	.w7(32'hb9f18460),
	.w8(32'hbbc7474c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99a8a6),
	.w1(32'h3be88927),
	.w2(32'h3cac4006),
	.w3(32'hbc80e1f4),
	.w4(32'hbc8211be),
	.w5(32'hbbf0a888),
	.w6(32'hbb0fc7f9),
	.w7(32'hbc4f04dd),
	.w8(32'hbc95fd8a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc22cea),
	.w1(32'hbacaa90d),
	.w2(32'hbc691f99),
	.w3(32'hbb1ac88f),
	.w4(32'h3a7ecbfa),
	.w5(32'hbbd29f14),
	.w6(32'h3bd7a066),
	.w7(32'h3c8c6b39),
	.w8(32'h3a975a88),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc173a5f),
	.w1(32'hbaa17375),
	.w2(32'hbd48d529),
	.w3(32'hbbd42f01),
	.w4(32'h3c9cc8db),
	.w5(32'h3d19ca4d),
	.w6(32'h3b5fb30a),
	.w7(32'h3a9fa1f0),
	.w8(32'h3c9ada6c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda6975f),
	.w1(32'hbca7429b),
	.w2(32'h3bbaaa6f),
	.w3(32'h3d1477c4),
	.w4(32'h3a9873ec),
	.w5(32'hbbbeebbb),
	.w6(32'h3d0ca1c2),
	.w7(32'h3b5dc7e6),
	.w8(32'hba9de882),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36841d),
	.w1(32'hbbe9e812),
	.w2(32'hbadde3e6),
	.w3(32'hbbb329f2),
	.w4(32'h3adb7c19),
	.w5(32'h3b83aee2),
	.w6(32'hbbaa06f5),
	.w7(32'hba04afdd),
	.w8(32'hbb49dd65),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22bee),
	.w1(32'hb99ea22b),
	.w2(32'hbcb9cc46),
	.w3(32'h3b9426c6),
	.w4(32'hbbe4be14),
	.w5(32'hba880a62),
	.w6(32'h3bbc651c),
	.w7(32'hbc861426),
	.w8(32'h3b84280f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64265f),
	.w1(32'h3cadf479),
	.w2(32'hbc954014),
	.w3(32'h3b4d53bf),
	.w4(32'h3c2a5896),
	.w5(32'h3b56e096),
	.w6(32'h3cd8171d),
	.w7(32'hbb044e10),
	.w8(32'hbb87d9c6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab772d),
	.w1(32'hbca03270),
	.w2(32'hbae3cd0f),
	.w3(32'hbac93327),
	.w4(32'hbc064745),
	.w5(32'h37d831c4),
	.w6(32'hbb0392b8),
	.w7(32'hbc48ab10),
	.w8(32'hba83e111),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7631a3),
	.w1(32'hbba7ad33),
	.w2(32'h3cbc0fa5),
	.w3(32'hbb458958),
	.w4(32'h3c076c24),
	.w5(32'h3b04395c),
	.w6(32'h3c251dec),
	.w7(32'h3c4303b3),
	.w8(32'hbc1c69aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule