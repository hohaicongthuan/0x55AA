module layer_10_featuremap_11(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc261b3e),
	.w1(32'hbbac2fce),
	.w2(32'hbb07273d),
	.w3(32'hbc121b8b),
	.w4(32'hbbe3fb71),
	.w5(32'hba023818),
	.w6(32'h38adc8ee),
	.w7(32'h3b0d40ca),
	.w8(32'hbae0cf23),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7de327),
	.w1(32'hbb4a0945),
	.w2(32'h3bc815d7),
	.w3(32'hbae8f4e7),
	.w4(32'hbc1d5750),
	.w5(32'h3be31b14),
	.w6(32'h3ba6d71f),
	.w7(32'hbad5e314),
	.w8(32'h3c00cb39),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb906b),
	.w1(32'hbbf0fb20),
	.w2(32'h3bad9a0d),
	.w3(32'hba0b493d),
	.w4(32'hb9c44bc6),
	.w5(32'hbb463a5b),
	.w6(32'h3c0a2463),
	.w7(32'h3b60c5af),
	.w8(32'h396fd00b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26fd8c),
	.w1(32'hbbaaff54),
	.w2(32'hbbcf4684),
	.w3(32'hbab13c77),
	.w4(32'h3afd648a),
	.w5(32'hbc14db52),
	.w6(32'h3b7f663e),
	.w7(32'h3ba85973),
	.w8(32'h3ba4e6ee),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa1a06),
	.w1(32'h3aa0fcf4),
	.w2(32'h3bc9b61c),
	.w3(32'hbbaf6f64),
	.w4(32'h3b3f54dc),
	.w5(32'h3bf49935),
	.w6(32'h3c7768a7),
	.w7(32'h3c44fc66),
	.w8(32'h3bb19d8e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f7880),
	.w1(32'hbb9d57a5),
	.w2(32'hbd2e5585),
	.w3(32'h39d97788),
	.w4(32'hbbf5d9a1),
	.w5(32'hbc89d5f6),
	.w6(32'h3ad96f35),
	.w7(32'hbb8330e3),
	.w8(32'h3cea2392),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8f2702),
	.w1(32'hbd1d83b1),
	.w2(32'hbc1fd80d),
	.w3(32'h3c265d7c),
	.w4(32'h3c35908a),
	.w5(32'hbc9d63c2),
	.w6(32'h3da90009),
	.w7(32'h3d660584),
	.w8(32'h3b81d219),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92ab76),
	.w1(32'hbc2662d9),
	.w2(32'hbb9b50bf),
	.w3(32'hbce3fc43),
	.w4(32'hbc465804),
	.w5(32'hbb34a5d0),
	.w6(32'h3af873fe),
	.w7(32'h3c415829),
	.w8(32'hba49dfec),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb3f29),
	.w1(32'h3b830a6c),
	.w2(32'h3c045ca8),
	.w3(32'h3b614a12),
	.w4(32'h3b7ebd9e),
	.w5(32'h3b49f32c),
	.w6(32'h3c70102d),
	.w7(32'h3c2e94ab),
	.w8(32'hbc009a43),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10731f),
	.w1(32'h3c00d603),
	.w2(32'h3d2e554c),
	.w3(32'h3b9dc894),
	.w4(32'h3ae87ac7),
	.w5(32'h3cbf5bc9),
	.w6(32'hbc693c7a),
	.w7(32'hbc173f7e),
	.w8(32'hbc3acdb4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d802e60),
	.w1(32'h3d0bb360),
	.w2(32'hbaef14fc),
	.w3(32'h3b7d23e3),
	.w4(32'hbc2e0b04),
	.w5(32'hbb3212b5),
	.w6(32'hbd71ad9f),
	.w7(32'hbd3fdd15),
	.w8(32'hba2a0cbf),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23cf5c),
	.w1(32'h3b22e930),
	.w2(32'hbbf51083),
	.w3(32'h39199272),
	.w4(32'hbb560c08),
	.w5(32'hbb9e1223),
	.w6(32'hbb270972),
	.w7(32'hbb073e1b),
	.w8(32'h3bb4503b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc878615),
	.w1(32'hbc2c6883),
	.w2(32'hbb907873),
	.w3(32'hbaf1ff98),
	.w4(32'hba5f2d01),
	.w5(32'hbb3ed271),
	.w6(32'h3ca278eb),
	.w7(32'h3c7ff917),
	.w8(32'hbba7abad),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49fb48),
	.w1(32'hbbccb515),
	.w2(32'hba2b62c9),
	.w3(32'hbba43cfc),
	.w4(32'hbb74caa4),
	.w5(32'h3bc0e2d0),
	.w6(32'h3ab372e9),
	.w7(32'hbb5e0d59),
	.w8(32'h3b46aed2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dd947),
	.w1(32'h3a2792c7),
	.w2(32'hb9a93fb7),
	.w3(32'h3bc68bb9),
	.w4(32'h3b7295b5),
	.w5(32'hbafa2e56),
	.w6(32'hba42dbdf),
	.w7(32'h3a946a6c),
	.w8(32'hbb45a3e1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6095fe),
	.w1(32'h3ba99a9b),
	.w2(32'h3cc8437b),
	.w3(32'hbc596edd),
	.w4(32'hbc096476),
	.w5(32'h3c58561c),
	.w6(32'hbc2cfd17),
	.w7(32'hbc0f1b2d),
	.w8(32'hbc10b3bc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f6049),
	.w1(32'h3c8412a9),
	.w2(32'hbc2e8612),
	.w3(32'hba9a9667),
	.w4(32'hbc5a1cf4),
	.w5(32'hbc319e0f),
	.w6(32'hbd2353df),
	.w7(32'hbd0f8917),
	.w8(32'h3b19395c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfd78b),
	.w1(32'hbc52dd66),
	.w2(32'h39410b2c),
	.w3(32'hbb91a374),
	.w4(32'hbc0198fe),
	.w5(32'hbb6bc1a4),
	.w6(32'h3bf328fa),
	.w7(32'h3b81e706),
	.w8(32'hbbac4799),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a241fba),
	.w1(32'hbb0c66c8),
	.w2(32'hbaaf88d2),
	.w3(32'h3a3dfbc1),
	.w4(32'hbb57783b),
	.w5(32'h3b7af570),
	.w6(32'hbbf1d65b),
	.w7(32'hbb4fa489),
	.w8(32'h3c02641a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a39e5),
	.w1(32'h3b754c3e),
	.w2(32'h3ba91fde),
	.w3(32'h3c7d885e),
	.w4(32'h3c84da55),
	.w5(32'h3aa1388c),
	.w6(32'h3bebd18b),
	.w7(32'h3bcf37f0),
	.w8(32'h3bdce37e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a894e39),
	.w1(32'h3b7be0f8),
	.w2(32'hbbe72956),
	.w3(32'h3bd8c321),
	.w4(32'h3b8f0ca7),
	.w5(32'hbbe054bd),
	.w6(32'h3c7c5feb),
	.w7(32'h3bf6ad97),
	.w8(32'hbabea690),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025998),
	.w1(32'hbb7c247e),
	.w2(32'hbb9a65be),
	.w3(32'hbb6872a7),
	.w4(32'hba04d4b6),
	.w5(32'hba69bb7e),
	.w6(32'h3a4dd224),
	.w7(32'h3bd7edf5),
	.w8(32'h384412ff),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d4cc2),
	.w1(32'hbad9050e),
	.w2(32'h3d0b0ebf),
	.w3(32'hbbb0e109),
	.w4(32'hbb7d544a),
	.w5(32'h3c7ea62f),
	.w6(32'hbb10816c),
	.w7(32'hbbc1236c),
	.w8(32'hbcad1a40),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7f6b6f),
	.w1(32'h3d0311c9),
	.w2(32'hbb6aefcf),
	.w3(32'h3b612534),
	.w4(32'hbb94280d),
	.w5(32'hbc031123),
	.w6(32'hbd6d0e45),
	.w7(32'hbd31f9be),
	.w8(32'hbc05edb7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bc2d8),
	.w1(32'hbb0d3c3a),
	.w2(32'hbbe67b9e),
	.w3(32'hba257128),
	.w4(32'hbb3eb276),
	.w5(32'h3b6d009a),
	.w6(32'hbbd0ec31),
	.w7(32'h3aa2206f),
	.w8(32'h3b0c3d3c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7c12),
	.w1(32'h3ab692b5),
	.w2(32'hbb6a784a),
	.w3(32'h3c4095c1),
	.w4(32'h3c2e9b39),
	.w5(32'h3b91841e),
	.w6(32'h3c433443),
	.w7(32'h3c2cb1f8),
	.w8(32'h3be23c47),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fea0cf),
	.w1(32'hbb924f58),
	.w2(32'hb89905fa),
	.w3(32'h3af36e1e),
	.w4(32'h3b177780),
	.w5(32'h3943a345),
	.w6(32'h3b16e4fd),
	.w7(32'hbb3cf406),
	.w8(32'hb822e7bf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944aac4),
	.w1(32'hb8973249),
	.w2(32'hb97066a6),
	.w3(32'hb995736d),
	.w4(32'h390fd007),
	.w5(32'h3900a98a),
	.w6(32'hb9cdb8ae),
	.w7(32'hb8936f68),
	.w8(32'h3a43c5f5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09c3a3),
	.w1(32'hba740639),
	.w2(32'hba6dc693),
	.w3(32'hb9de8b40),
	.w4(32'hba71ba13),
	.w5(32'hbaeef16e),
	.w6(32'h39bccdc8),
	.w7(32'hba5cca58),
	.w8(32'hba0651b8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb125193),
	.w1(32'hba2c9293),
	.w2(32'hba7c11c1),
	.w3(32'hbb4fedb3),
	.w4(32'hbac7b0e7),
	.w5(32'hba72582e),
	.w6(32'hbad3733a),
	.w7(32'hbacb0af4),
	.w8(32'hba6e172e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa3c3d),
	.w1(32'hbaa89d0a),
	.w2(32'hbaa3897a),
	.w3(32'hba6cd830),
	.w4(32'hba870acb),
	.w5(32'h39edb5a3),
	.w6(32'hba8c5699),
	.w7(32'hba964ee3),
	.w8(32'hba19cbaf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043ab6),
	.w1(32'hba962724),
	.w2(32'hb966a2da),
	.w3(32'hb9f40e81),
	.w4(32'h3a2bf6ef),
	.w5(32'h39bdb209),
	.w6(32'hba7c7108),
	.w7(32'hba9f48be),
	.w8(32'h3a682cb3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fb50c0),
	.w1(32'h39e889d8),
	.w2(32'hb968de4f),
	.w3(32'hbaf99963),
	.w4(32'hba5a8b2c),
	.w5(32'hb93c9006),
	.w6(32'h3a837806),
	.w7(32'h3a579dee),
	.w8(32'h373e8251),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b89b7),
	.w1(32'h38bf22b4),
	.w2(32'hba153c78),
	.w3(32'hb998f6ef),
	.w4(32'hb7001534),
	.w5(32'hba1ae24c),
	.w6(32'hb9c6f487),
	.w7(32'hb98abd2d),
	.w8(32'h3a02cfd6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85a32a),
	.w1(32'hba25ea7e),
	.w2(32'h3aa414ec),
	.w3(32'hb9c2428f),
	.w4(32'hba483f91),
	.w5(32'h3ab5b325),
	.w6(32'hba02e5ff),
	.w7(32'h3955a8a1),
	.w8(32'h3a9d7a79),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa650b6),
	.w1(32'h3aaae759),
	.w2(32'hbac07bae),
	.w3(32'h3a7c5533),
	.w4(32'h3a9643f2),
	.w5(32'h3a33eae6),
	.w6(32'h3a9e893c),
	.w7(32'h3a8cdaee),
	.w8(32'h3ab13ab2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41cd76),
	.w1(32'h3a63f563),
	.w2(32'h3a95331c),
	.w3(32'h3911d384),
	.w4(32'h3b124821),
	.w5(32'h3ac70244),
	.w6(32'h39a25764),
	.w7(32'h3a9f4a80),
	.w8(32'h3b069468),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969eae4),
	.w1(32'h399320df),
	.w2(32'hb9118783),
	.w3(32'hbab28c48),
	.w4(32'hba0b4272),
	.w5(32'hbacc35ca),
	.w6(32'hba8651f0),
	.w7(32'hba84b65e),
	.w8(32'h3a3aa7b6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2143a9),
	.w1(32'hbac540ab),
	.w2(32'h3b011a3d),
	.w3(32'hbb5d1d93),
	.w4(32'hbb60ea10),
	.w5(32'h3b1eeb23),
	.w6(32'hb9578116),
	.w7(32'hbad1beba),
	.w8(32'h3aaf7078),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c934a),
	.w1(32'hb9c4b3d6),
	.w2(32'h38cf739c),
	.w3(32'h3a9ebb8e),
	.w4(32'hb911c2fa),
	.w5(32'hb9e60a41),
	.w6(32'h3a51114f),
	.w7(32'h39756106),
	.w8(32'hb9c181d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986663a),
	.w1(32'hba1fca82),
	.w2(32'hb9996e9f),
	.w3(32'hba435eea),
	.w4(32'hba8d9a19),
	.w5(32'hba9dc851),
	.w6(32'hba7e55a9),
	.w7(32'hbac752af),
	.w8(32'h3a2b3bda),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da24bd),
	.w1(32'hb882300c),
	.w2(32'h3a9696d3),
	.w3(32'hb987ee54),
	.w4(32'hba7542d3),
	.w5(32'h3ad2ff5d),
	.w6(32'h3a6020f3),
	.w7(32'hb9040141),
	.w8(32'h3a7e2ff0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972cd0e),
	.w1(32'hb816ff41),
	.w2(32'h3ac4ab33),
	.w3(32'h39d076b8),
	.w4(32'h37b3e261),
	.w5(32'h3abd0504),
	.w6(32'h3a063635),
	.w7(32'hba16f0e5),
	.w8(32'h3a9ea623),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec0772),
	.w1(32'h3b023981),
	.w2(32'h3a3aca74),
	.w3(32'h3a70b627),
	.w4(32'h3ac62b3f),
	.w5(32'hb94e7a0d),
	.w6(32'h3a178b19),
	.w7(32'h3a9d02ec),
	.w8(32'hba16c7d3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba237d6d),
	.w1(32'hba8b9395),
	.w2(32'h3ae32c3b),
	.w3(32'hbabd77c7),
	.w4(32'hbaefce99),
	.w5(32'h3ae41fad),
	.w6(32'hba662ae1),
	.w7(32'hbad6b80d),
	.w8(32'h3b2e5c13),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec5289),
	.w1(32'h3ae47cf4),
	.w2(32'h3b0f66ae),
	.w3(32'h3ae7603e),
	.w4(32'h3af13bec),
	.w5(32'h39ae9dce),
	.w6(32'h3b1f9487),
	.w7(32'h3a814c1e),
	.w8(32'h3adbee07),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08f71b),
	.w1(32'h3b54f0d0),
	.w2(32'hba2bf8f5),
	.w3(32'h3a7d099a),
	.w4(32'h3b31adf1),
	.w5(32'hbae7b1cf),
	.w6(32'h3a81930e),
	.w7(32'h3b3e4580),
	.w8(32'h393455c6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75129b3),
	.w1(32'hb9ff01b8),
	.w2(32'h3ac96514),
	.w3(32'hbac76f20),
	.w4(32'hba81f82c),
	.w5(32'h3ab3d1e0),
	.w6(32'hba561520),
	.w7(32'h38ef2b25),
	.w8(32'h3a8f6b9e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e6ecf),
	.w1(32'h3a9656f9),
	.w2(32'hb98fea5d),
	.w3(32'h3ab66849),
	.w4(32'h3a92e63f),
	.w5(32'h3937a0dd),
	.w6(32'h3a69ad87),
	.w7(32'h3a6a4e39),
	.w8(32'h39ef8307),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a624b5c),
	.w1(32'hb787cb94),
	.w2(32'h3ab6f9ec),
	.w3(32'hba454afb),
	.w4(32'h3a0939be),
	.w5(32'h3b1df810),
	.w6(32'hb74ca353),
	.w7(32'hba431d35),
	.w8(32'h3aebd299),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04b685),
	.w1(32'h3a43baf4),
	.w2(32'hb95a550b),
	.w3(32'hb8838208),
	.w4(32'h3a3f4464),
	.w5(32'hba67b6eb),
	.w6(32'hb9d5baf4),
	.w7(32'hb82cd8ca),
	.w8(32'hba26c869),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d35524),
	.w1(32'hb9def908),
	.w2(32'h3a86123d),
	.w3(32'h3aa8a013),
	.w4(32'hb9c65831),
	.w5(32'h3ad35a27),
	.w6(32'h39ad3c37),
	.w7(32'hba51f641),
	.w8(32'h3b0b6afb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac72e31),
	.w1(32'h3a936e1e),
	.w2(32'hb9c40bb2),
	.w3(32'h3a5f3b0a),
	.w4(32'h399285f6),
	.w5(32'h3a92c973),
	.w6(32'h39878f32),
	.w7(32'h37107177),
	.w8(32'h39dde211),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f6884c),
	.w1(32'h3a830cdd),
	.w2(32'h3a654e9c),
	.w3(32'h3b00c679),
	.w4(32'h3b0b36f0),
	.w5(32'h3a2528e3),
	.w6(32'h39c78a14),
	.w7(32'h3a37a60a),
	.w8(32'h3a8818b9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b56a8),
	.w1(32'h3902b106),
	.w2(32'hbb273fe8),
	.w3(32'hba8557dc),
	.w4(32'h38004aa9),
	.w5(32'hba99d4c1),
	.w6(32'hb9b82731),
	.w7(32'h39f49215),
	.w8(32'hba009d31),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb689c08),
	.w1(32'hbb24416b),
	.w2(32'h3acc4c4e),
	.w3(32'hba92cabf),
	.w4(32'hba6fde2f),
	.w5(32'h3abcd9ad),
	.w6(32'hb98d271c),
	.w7(32'hba334ef5),
	.w8(32'h3aa62f65),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3043d),
	.w1(32'h3aac0300),
	.w2(32'h39780615),
	.w3(32'h3abb9b62),
	.w4(32'h3acb65ed),
	.w5(32'h39d13081),
	.w6(32'h3abcbce6),
	.w7(32'h3ada1f5e),
	.w8(32'h3a3a55cc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9095e2c),
	.w1(32'hb9b6f27e),
	.w2(32'h39bc6522),
	.w3(32'hb902a20d),
	.w4(32'hb9f3dc00),
	.w5(32'h390d016e),
	.w6(32'h39617b52),
	.w7(32'hb93fffbc),
	.w8(32'hba65d719),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888da49),
	.w1(32'hbaab3b84),
	.w2(32'h392d41ce),
	.w3(32'hb9bbe85e),
	.w4(32'hbaed3eed),
	.w5(32'h39e4a574),
	.w6(32'hbab353ae),
	.w7(32'hbb587e2f),
	.w8(32'h3a510288),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a58a5d),
	.w1(32'h3a5e2340),
	.w2(32'h3a82a1f3),
	.w3(32'h3a32f933),
	.w4(32'h39bcd3b2),
	.w5(32'h39bc8c7c),
	.w6(32'h3a9b279b),
	.w7(32'h3a588e01),
	.w8(32'h3a3334a7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5619f),
	.w1(32'h39dd79c8),
	.w2(32'hb7193094),
	.w3(32'hb91460f0),
	.w4(32'hb9008565),
	.w5(32'hb9abded5),
	.w6(32'hb900cb22),
	.w7(32'hb8c65734),
	.w8(32'hba779336),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1769a4),
	.w1(32'hb9a3f807),
	.w2(32'hbae40cf7),
	.w3(32'hba5237ea),
	.w4(32'hba6ebf5b),
	.w5(32'hbae68431),
	.w6(32'hba90b882),
	.w7(32'hba82ddd3),
	.w8(32'hba96ff39),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba878c68),
	.w1(32'hbb0087fe),
	.w2(32'hba172fcc),
	.w3(32'hbaaf65a7),
	.w4(32'hbb243b2a),
	.w5(32'hba00b26f),
	.w6(32'hbac6e432),
	.w7(32'hbac680ff),
	.w8(32'hb91ddee0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c0e72),
	.w1(32'hb95b740d),
	.w2(32'hb916a816),
	.w3(32'hb8d323dc),
	.w4(32'hb7633e94),
	.w5(32'h3a4b26a0),
	.w6(32'hb8829865),
	.w7(32'hb983aa84),
	.w8(32'h3a9bfc3b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e1a7),
	.w1(32'h38d156c7),
	.w2(32'hb82abaa8),
	.w3(32'h3a8ae94f),
	.w4(32'h3a3694b7),
	.w5(32'h38817c7b),
	.w6(32'hb93d2c32),
	.w7(32'h39587d48),
	.w8(32'hb9c4561c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97575d8),
	.w1(32'hb9abd2ea),
	.w2(32'h3a27d699),
	.w3(32'h393912db),
	.w4(32'hb80b6ee1),
	.w5(32'h3a48f511),
	.w6(32'hb9a43b05),
	.w7(32'hb9679f16),
	.w8(32'h3a906981),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391858cd),
	.w1(32'h3a0d249f),
	.w2(32'hb9757d38),
	.w3(32'hb9cbb063),
	.w4(32'h3899f725),
	.w5(32'hba95e0de),
	.w6(32'h3940c070),
	.w7(32'h39bc5671),
	.w8(32'hb980b0ff),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80dde6),
	.w1(32'hba16c8df),
	.w2(32'h398f32d4),
	.w3(32'hbb197997),
	.w4(32'hbaa7008c),
	.w5(32'h3ace0d2e),
	.w6(32'hbb07c6a5),
	.w7(32'hbadbb041),
	.w8(32'h3a16a0ba),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd73c0),
	.w1(32'h39ea2049),
	.w2(32'h39d8367c),
	.w3(32'h39a5efa5),
	.w4(32'h3a100300),
	.w5(32'h392f6866),
	.w6(32'hb8d02843),
	.w7(32'hb9984800),
	.w8(32'hb80b8b60),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382f5f96),
	.w1(32'h39bd3499),
	.w2(32'h3ad90b87),
	.w3(32'hba29c4ea),
	.w4(32'hb97eb8a9),
	.w5(32'h3a84bbbe),
	.w6(32'hba8dce98),
	.w7(32'hba534db8),
	.w8(32'h3a6e921e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39952d91),
	.w1(32'hb8aaea5b),
	.w2(32'hb8f0a7b4),
	.w3(32'h3a3560ef),
	.w4(32'hb87b4fa6),
	.w5(32'h39907b1c),
	.w6(32'h3a2676a0),
	.w7(32'h38a5123f),
	.w8(32'h380ca6b4),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901f60f),
	.w1(32'hba51bae8),
	.w2(32'hb9e17cb4),
	.w3(32'h3acb151c),
	.w4(32'h38ddcf75),
	.w5(32'hba8e79d5),
	.w6(32'h3a81a387),
	.w7(32'hb95b5743),
	.w8(32'h39932aa6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c51eb6),
	.w1(32'h39ae088d),
	.w2(32'h381f1073),
	.w3(32'hbab47bee),
	.w4(32'h39c765e7),
	.w5(32'h3901a250),
	.w6(32'hb873b3aa),
	.w7(32'h398dde43),
	.w8(32'hba9ee994),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f06bd),
	.w1(32'hba5122aa),
	.w2(32'hbaa48734),
	.w3(32'hba4fa0ff),
	.w4(32'hb9da3c9f),
	.w5(32'hba88cdd0),
	.w6(32'hbab9524e),
	.w7(32'hba7cb858),
	.w8(32'hba97db94),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba54b0),
	.w1(32'hbab430be),
	.w2(32'h3a9129c3),
	.w3(32'hba90550d),
	.w4(32'hba918851),
	.w5(32'h3a7570e6),
	.w6(32'hbab2574c),
	.w7(32'hba9e505a),
	.w8(32'h3a39b804),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9afca6),
	.w1(32'h3a9aa08a),
	.w2(32'hba4f28dd),
	.w3(32'h3aaf78ce),
	.w4(32'h3aad08fe),
	.w5(32'h3a4907f6),
	.w6(32'h3a44a27b),
	.w7(32'h3a79ba2d),
	.w8(32'hb99e0719),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ac679),
	.w1(32'h3a86a5bb),
	.w2(32'h3ab97fc0),
	.w3(32'h3a76b6e9),
	.w4(32'h3a7a187a),
	.w5(32'h3a96d5a4),
	.w6(32'hb998e14f),
	.w7(32'h3a8f9a3d),
	.w8(32'hba0ec523),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36414c),
	.w1(32'h3ac11394),
	.w2(32'h3a20ea8e),
	.w3(32'hb96d73e6),
	.w4(32'h3aaa5bac),
	.w5(32'hba309102),
	.w6(32'hb9ebc258),
	.w7(32'hb8a2e794),
	.w8(32'h3a0f3d2e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89c892),
	.w1(32'h3a3f7655),
	.w2(32'h39daf784),
	.w3(32'h38c8ea89),
	.w4(32'h3a238b03),
	.w5(32'h3a4a3378),
	.w6(32'h39df4d99),
	.w7(32'h3a80fb0b),
	.w8(32'h3a37ee73),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e0e793),
	.w1(32'h390f6f32),
	.w2(32'h39ddd903),
	.w3(32'hb9d32a4e),
	.w4(32'h3932a492),
	.w5(32'h3969c6bf),
	.w6(32'hb8fde11e),
	.w7(32'h392ab536),
	.w8(32'h3a709634),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddb014),
	.w1(32'h39925811),
	.w2(32'hba5aeeef),
	.w3(32'h38ddac64),
	.w4(32'h3940a2cd),
	.w5(32'hba0adfec),
	.w6(32'h3a35de48),
	.w7(32'h3a5ccb93),
	.w8(32'hba11cb10),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8939d9),
	.w1(32'hba58d302),
	.w2(32'hba92d918),
	.w3(32'hba669996),
	.w4(32'hba188f64),
	.w5(32'hba94a53c),
	.w6(32'hba689c06),
	.w7(32'hba1d69fb),
	.w8(32'hb9e6fe8c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba679dc2),
	.w1(32'h3a54df8b),
	.w2(32'h3a1a79cf),
	.w3(32'hbae33779),
	.w4(32'h38f06eef),
	.w5(32'hb9327f2a),
	.w6(32'hba8bbed3),
	.w7(32'hba11e10d),
	.w8(32'h3aa6ad51),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e896b),
	.w1(32'h3a64a7af),
	.w2(32'hb9ca7ae5),
	.w3(32'h3740c823),
	.w4(32'h39b04e37),
	.w5(32'hba78120a),
	.w6(32'h3989c12a),
	.w7(32'h3afa974f),
	.w8(32'h392c2c5c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac95fb),
	.w1(32'h395bb855),
	.w2(32'hb9f7a6ed),
	.w3(32'hb7d869c6),
	.w4(32'hba1fc1c8),
	.w5(32'hbaa819cd),
	.w6(32'h3937fbe3),
	.w7(32'h3a472172),
	.w8(32'hba142183),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08064b),
	.w1(32'hba92bd6a),
	.w2(32'hb9138e0a),
	.w3(32'hbb0d151c),
	.w4(32'hbb193751),
	.w5(32'hb95e381e),
	.w6(32'hbb01a58a),
	.w7(32'hbb47a438),
	.w8(32'h3913420f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdaffc),
	.w1(32'hba47939e),
	.w2(32'hb98fb15d),
	.w3(32'h393a31ac),
	.w4(32'hba010416),
	.w5(32'hb983f36d),
	.w6(32'h39149d3b),
	.w7(32'hb9afcfe6),
	.w8(32'hb9528353),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c79aa),
	.w1(32'hb91d1f9a),
	.w2(32'h3a9428ef),
	.w3(32'hb908629b),
	.w4(32'hb9020f05),
	.w5(32'h3b7e9c4f),
	.w6(32'hb94d6a73),
	.w7(32'hb9bbdac8),
	.w8(32'h3a74edd4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a902ab7),
	.w1(32'h3a8fc075),
	.w2(32'h3997e658),
	.w3(32'h39edf2b2),
	.w4(32'h3b585d41),
	.w5(32'h3ae92357),
	.w6(32'h3adfe7b6),
	.w7(32'h3969ef4f),
	.w8(32'h3a9e3d02),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e1a2),
	.w1(32'h390cc8d8),
	.w2(32'h3abb7597),
	.w3(32'h3a56cd35),
	.w4(32'h3b114721),
	.w5(32'h3ad156a1),
	.w6(32'h3a4f8808),
	.w7(32'h39a5686c),
	.w8(32'h3a76f304),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3e4a6),
	.w1(32'h38cab281),
	.w2(32'h39b6f235),
	.w3(32'hb99924a7),
	.w4(32'hba0a94a6),
	.w5(32'h38e23c27),
	.w6(32'hba34de98),
	.w7(32'hba59206f),
	.w8(32'h3971cc69),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90fda0a),
	.w1(32'h39e0894a),
	.w2(32'h39b8b14d),
	.w3(32'hba88e8e8),
	.w4(32'hbaace82a),
	.w5(32'hb93691d1),
	.w6(32'hba87f231),
	.w7(32'hba80e213),
	.w8(32'hbabd292f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc39b),
	.w1(32'hbaafe389),
	.w2(32'h3a2afc31),
	.w3(32'hbacab8c9),
	.w4(32'hbae644d7),
	.w5(32'h36838052),
	.w6(32'hbaed8c28),
	.w7(32'hbb162e64),
	.w8(32'hb92b4e46),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37595d),
	.w1(32'h39e35054),
	.w2(32'h3a857979),
	.w3(32'h3906ae92),
	.w4(32'h36fb81a4),
	.w5(32'h3af34f1d),
	.w6(32'hba2e5555),
	.w7(32'hba215a3e),
	.w8(32'h3a99d774),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998a196),
	.w1(32'h379046d9),
	.w2(32'hb9fd859d),
	.w3(32'hb9bf8c02),
	.w4(32'h39cad467),
	.w5(32'hbaadd164),
	.w6(32'hb9eef291),
	.w7(32'h3953cb1f),
	.w8(32'hba2ca451),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0843b7),
	.w1(32'hba2f81f7),
	.w2(32'h3afe7801),
	.w3(32'hbaf88a35),
	.w4(32'hbaaca6aa),
	.w5(32'h3b090164),
	.w6(32'hbab950c4),
	.w7(32'hba0e2549),
	.w8(32'h3ad5c7a2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ce7e6),
	.w1(32'h3a631553),
	.w2(32'h3b5d6c23),
	.w3(32'h3a7ac652),
	.w4(32'h3b031b05),
	.w5(32'h3af97196),
	.w6(32'h3a02edb2),
	.w7(32'h3a2b9ef9),
	.w8(32'h3af9312a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b37d),
	.w1(32'h3af1bf58),
	.w2(32'h3aa537c1),
	.w3(32'h3b0d9813),
	.w4(32'h3a11c8d9),
	.w5(32'h3b09573f),
	.w6(32'h3967b5e3),
	.w7(32'h3aa0952f),
	.w8(32'h3ad7a2c8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d12d7),
	.w1(32'h3a27e519),
	.w2(32'h3a84f1ea),
	.w3(32'hba136989),
	.w4(32'h3ab24abf),
	.w5(32'h3a6ac223),
	.w6(32'h3a6a0374),
	.w7(32'h3adfa6d7),
	.w8(32'h3af3abbb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef75b7),
	.w1(32'h39c6a766),
	.w2(32'hba02807b),
	.w3(32'h398402d0),
	.w4(32'h39652093),
	.w5(32'h38b5d87a),
	.w6(32'h3911ee60),
	.w7(32'h39d5df18),
	.w8(32'h391a03c8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a416ef0),
	.w1(32'h3ab36aa9),
	.w2(32'h3a08d6c3),
	.w3(32'h39f7cfda),
	.w4(32'hb9e64045),
	.w5(32'h3a6e6e80),
	.w6(32'hbab8bb64),
	.w7(32'hbb0a2c9d),
	.w8(32'hba5df2f3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf717f2),
	.w1(32'hbabfb7c5),
	.w2(32'h3aad6904),
	.w3(32'hbabd7e03),
	.w4(32'h39745d59),
	.w5(32'h3aec1b90),
	.w6(32'hbb1f6e36),
	.w7(32'hbb1647fd),
	.w8(32'h3aa7968c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae4ce7),
	.w1(32'h3a2006b6),
	.w2(32'h39f541c6),
	.w3(32'h3a5759e4),
	.w4(32'h3ad61fc6),
	.w5(32'h3aa7407c),
	.w6(32'h3a0e866c),
	.w7(32'h39bf3e24),
	.w8(32'h3a121293),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c4b68),
	.w1(32'h39fce484),
	.w2(32'h3949fb22),
	.w3(32'h3ab4adad),
	.w4(32'h3aa877ae),
	.w5(32'hba90d2e3),
	.w6(32'h3a57730b),
	.w7(32'h3a1da660),
	.w8(32'h38b811db),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd27d4),
	.w1(32'hba1310bf),
	.w2(32'hb868a71a),
	.w3(32'hbaf6b155),
	.w4(32'hb963aa16),
	.w5(32'h3a606b75),
	.w6(32'hbaaaf565),
	.w7(32'hb90e714a),
	.w8(32'h3a350029),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43eb5b),
	.w1(32'hb946ec14),
	.w2(32'hba0133fa),
	.w3(32'h3a6621a7),
	.w4(32'h392b7d26),
	.w5(32'hb9ccd23e),
	.w6(32'h3a7e5dd5),
	.w7(32'hb862f16a),
	.w8(32'hb99d8c6c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a03fee),
	.w1(32'hba6629bf),
	.w2(32'h39383c62),
	.w3(32'hb9032a65),
	.w4(32'hb99f9a75),
	.w5(32'h398adff3),
	.w6(32'hb7d7ac75),
	.w7(32'hb9e13d60),
	.w8(32'h3a2f595a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7318f),
	.w1(32'hb94b7e00),
	.w2(32'h3a737346),
	.w3(32'h3a62dbae),
	.w4(32'h3a1093e3),
	.w5(32'h3a4350ee),
	.w6(32'h3a2ca702),
	.w7(32'h3aa283e9),
	.w8(32'hb895456b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3edc3),
	.w1(32'h3a376d13),
	.w2(32'hba5a0a6d),
	.w3(32'h3951d5a1),
	.w4(32'h39489e4f),
	.w5(32'h3926657b),
	.w6(32'h397c6fa2),
	.w7(32'hb74af625),
	.w8(32'hbad5ce14),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92e603),
	.w1(32'hba8c218c),
	.w2(32'h3ae1ea3e),
	.w3(32'hba887d3d),
	.w4(32'hb9eb2e33),
	.w5(32'h3a98a0c0),
	.w6(32'hbb2bd71f),
	.w7(32'hbb136f23),
	.w8(32'h3abc9cb2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961dcfa),
	.w1(32'h39c641cf),
	.w2(32'hb8e707d9),
	.w3(32'h39d5b73b),
	.w4(32'hb9f02e31),
	.w5(32'hbb066162),
	.w6(32'hba38b309),
	.w7(32'h39380ba6),
	.w8(32'hba105941),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7ee8a),
	.w1(32'hba4d1b07),
	.w2(32'h39752dee),
	.w3(32'hba763457),
	.w4(32'hba16241a),
	.w5(32'h3a880cc3),
	.w6(32'hba29e501),
	.w7(32'hb9753e97),
	.w8(32'h3b11078b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a702f7f),
	.w1(32'h3a8126e9),
	.w2(32'h3ab9ac7b),
	.w3(32'h39ad71f9),
	.w4(32'h3afa7d34),
	.w5(32'h3ac033ad),
	.w6(32'h3a87ea65),
	.w7(32'h3aafdee1),
	.w8(32'h3a8a04cf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48db7f),
	.w1(32'h3a9f3155),
	.w2(32'hba7dc326),
	.w3(32'h3a88a914),
	.w4(32'h3aaf6411),
	.w5(32'h39ec3412),
	.w6(32'h39e68d1b),
	.w7(32'h39fff9ff),
	.w8(32'h3aa21407),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c52b5),
	.w1(32'h3958cd6d),
	.w2(32'hba1f5a47),
	.w3(32'h3b1a671a),
	.w4(32'h3af95ec6),
	.w5(32'hb956ab99),
	.w6(32'h3ab8133f),
	.w7(32'h3ad15b0e),
	.w8(32'h3a16119e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c185c1),
	.w1(32'hba278aed),
	.w2(32'h3a05c6f4),
	.w3(32'h391ef423),
	.w4(32'hb91603c6),
	.w5(32'h3a9f5a00),
	.w6(32'h39f06dca),
	.w7(32'h39a46813),
	.w8(32'hb8aec3c1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a2947),
	.w1(32'hba182f7a),
	.w2(32'hba2c940a),
	.w3(32'h39defe08),
	.w4(32'h38561831),
	.w5(32'h399c8c5f),
	.w6(32'hba134061),
	.w7(32'hba0ffa82),
	.w8(32'h39d4c16a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba258697),
	.w1(32'hb9887b5b),
	.w2(32'hbaccaf8c),
	.w3(32'h39c2be6e),
	.w4(32'h39cf9c97),
	.w5(32'hba2103c4),
	.w6(32'h39bbd235),
	.w7(32'h389fb2a5),
	.w8(32'hba82155c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8984ed),
	.w1(32'hb9a72101),
	.w2(32'hb9a3936e),
	.w3(32'hba821350),
	.w4(32'h38a90232),
	.w5(32'h3986acbc),
	.w6(32'hba997795),
	.w7(32'hb9cc2057),
	.w8(32'hba037515),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba133d23),
	.w1(32'h3971b12c),
	.w2(32'h3aa59902),
	.w3(32'hba6633c1),
	.w4(32'hba468b80),
	.w5(32'h39c5a80a),
	.w6(32'hbaab6e21),
	.w7(32'hba893316),
	.w8(32'hba515a07),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c7e7f),
	.w1(32'hb98af0b1),
	.w2(32'hba2324ba),
	.w3(32'hb9a587ed),
	.w4(32'hb9c87ccb),
	.w5(32'hba0bc2e4),
	.w6(32'hba883113),
	.w7(32'hba865e87),
	.w8(32'hba644329),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba289298),
	.w1(32'hba24bdda),
	.w2(32'hb90c9bf9),
	.w3(32'hba2ec5c5),
	.w4(32'hba0556ed),
	.w5(32'hb9497600),
	.w6(32'hba69afdf),
	.w7(32'hba5a2802),
	.w8(32'hb991b4f1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26a148),
	.w1(32'hba326939),
	.w2(32'hb924596d),
	.w3(32'hb9cb0bcb),
	.w4(32'hba1018cf),
	.w5(32'h39abe842),
	.w6(32'hba1d880f),
	.w7(32'hba748990),
	.w8(32'h3aa918bf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58f179),
	.w1(32'h3972d5ca),
	.w2(32'hba588199),
	.w3(32'h3ac9625d),
	.w4(32'h3a6224bb),
	.w5(32'hba3b9549),
	.w6(32'h3b35120f),
	.w7(32'h3a8655f8),
	.w8(32'h38fbdccf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70cc02),
	.w1(32'hba425ac7),
	.w2(32'h38dc333f),
	.w3(32'hba51d98d),
	.w4(32'hba30ab6b),
	.w5(32'h3a694d05),
	.w6(32'hb81c5977),
	.w7(32'hb8bc88a1),
	.w8(32'h3ab49dff),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06dff1),
	.w1(32'h3a7a5852),
	.w2(32'hbb12e198),
	.w3(32'h39ccc2bd),
	.w4(32'h3a08fd44),
	.w5(32'hbaf0d418),
	.w6(32'h39c017de),
	.w7(32'h3a9d7de8),
	.w8(32'hba916427),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb181d1d),
	.w1(32'hbaa8637f),
	.w2(32'hbaba1a9f),
	.w3(32'hbb5541cc),
	.w4(32'hbaa0c72c),
	.w5(32'hbb10e473),
	.w6(32'hbb320621),
	.w7(32'hbb0a1754),
	.w8(32'hbab44135),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7364f),
	.w1(32'hba4a2caa),
	.w2(32'hbaad6204),
	.w3(32'hbae024ad),
	.w4(32'hba4b64b1),
	.w5(32'hba48e594),
	.w6(32'hbae7a863),
	.w7(32'hbab5cdd7),
	.w8(32'hba38e95f),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4aff1),
	.w1(32'hb9e8d954),
	.w2(32'h3916c6a4),
	.w3(32'hb82a82bb),
	.w4(32'h3a1e3984),
	.w5(32'h38fb0ac2),
	.w6(32'hb9f641df),
	.w7(32'h3943b446),
	.w8(32'h391fc1ae),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37fd7e),
	.w1(32'h3815dbf9),
	.w2(32'hbaf88b4b),
	.w3(32'h39dc8e13),
	.w4(32'hb9246aaa),
	.w5(32'hbb379e0b),
	.w6(32'hba5143ef),
	.w7(32'hb902c98c),
	.w8(32'hba70fd44),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb210a19),
	.w1(32'hbb0ab4b0),
	.w2(32'h3a78bba5),
	.w3(32'hbb514232),
	.w4(32'hbb0c5f3b),
	.w5(32'hb76e0ef4),
	.w6(32'hbaeb5636),
	.w7(32'hba8c6125),
	.w8(32'h3a7f5987),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958f508),
	.w1(32'h385fba15),
	.w2(32'h3b185803),
	.w3(32'h38dc7c43),
	.w4(32'hb90a7283),
	.w5(32'h3a902dda),
	.w6(32'h3947d764),
	.w7(32'hbad3846d),
	.w8(32'h3b0a93c4),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e06b6),
	.w1(32'h3b0c4907),
	.w2(32'hba71bd8c),
	.w3(32'h3ac3e76b),
	.w4(32'h3b022b4e),
	.w5(32'hbb1c801b),
	.w6(32'h3adc46d0),
	.w7(32'h3ab99e99),
	.w8(32'hbabcfabe),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945b573),
	.w1(32'hba1966e8),
	.w2(32'hb9a3edd0),
	.w3(32'h39897ef1),
	.w4(32'hbac6484a),
	.w5(32'hb9480832),
	.w6(32'h3b28415a),
	.w7(32'hba39bf43),
	.w8(32'hb98bdd4b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50049f),
	.w1(32'h381eef7a),
	.w2(32'hb93b9f68),
	.w3(32'hba41de47),
	.w4(32'hb9bfd542),
	.w5(32'h3a748dbf),
	.w6(32'hba563f03),
	.w7(32'hb9563113),
	.w8(32'h3a7158a0),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98094f0),
	.w1(32'h3a023974),
	.w2(32'h393279d8),
	.w3(32'h3a8e0c7a),
	.w4(32'h3abc5504),
	.w5(32'h3707f589),
	.w6(32'h3aabf5ad),
	.w7(32'h3a80f676),
	.w8(32'hb852a934),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a5181),
	.w1(32'hb7c0e880),
	.w2(32'h3ae6d927),
	.w3(32'h3aee327e),
	.w4(32'h3a5c509f),
	.w5(32'h3afed1f1),
	.w6(32'h399d4789),
	.w7(32'h3a7f073c),
	.w8(32'h3b0a5e80),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20b9b3),
	.w1(32'h3a89a4a6),
	.w2(32'hba2a22a8),
	.w3(32'h399b5c47),
	.w4(32'h3a4441c1),
	.w5(32'hba3cf259),
	.w6(32'h3a2aab9f),
	.w7(32'h3a691169),
	.w8(32'hba572b85),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99af42),
	.w1(32'hba7b3831),
	.w2(32'h39783bcc),
	.w3(32'hba61e40f),
	.w4(32'hba696871),
	.w5(32'h3a88d715),
	.w6(32'hba7d0886),
	.w7(32'hba59d64a),
	.w8(32'h3ab61416),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a274a18),
	.w1(32'h3a30cb13),
	.w2(32'hb9d78fac),
	.w3(32'h3ac79af2),
	.w4(32'h3a18dcea),
	.w5(32'hba35dd4f),
	.w6(32'h39477bb2),
	.w7(32'hb9656d15),
	.w8(32'hba7a2726),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa49250),
	.w1(32'hbab3a04e),
	.w2(32'h39edaed4),
	.w3(32'hbaa931ae),
	.w4(32'hbaafb936),
	.w5(32'h3a747251),
	.w6(32'hbaa845c0),
	.w7(32'hbaa72dd1),
	.w8(32'h3972ca27),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fd5fdd),
	.w1(32'h3a781ca6),
	.w2(32'h38fd090f),
	.w3(32'hb93b0441),
	.w4(32'h3aebe324),
	.w5(32'hbb165d72),
	.w6(32'hb84a8c03),
	.w7(32'h3a4524d7),
	.w8(32'hb8827397),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6fe5),
	.w1(32'hba12e0a6),
	.w2(32'h3923788a),
	.w3(32'hbb4d1a14),
	.w4(32'hbadb0c92),
	.w5(32'h380e8c37),
	.w6(32'hbaa2a6f1),
	.w7(32'hbaa2b38e),
	.w8(32'h3996dd83),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cb016),
	.w1(32'hb8a2bc2a),
	.w2(32'hba4ad582),
	.w3(32'h39182ca2),
	.w4(32'hb95a3158),
	.w5(32'hba6d31c7),
	.w6(32'h39f91a62),
	.w7(32'h3a250348),
	.w8(32'hba7500dc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88189e),
	.w1(32'hba83f3a6),
	.w2(32'hba1851bc),
	.w3(32'hba860d0f),
	.w4(32'hba93d48b),
	.w5(32'hb994277e),
	.w6(32'hba726aba),
	.w7(32'hba70153f),
	.w8(32'hba8edc04),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba859a7b),
	.w1(32'hba5bd545),
	.w2(32'hba58e410),
	.w3(32'hba2bc802),
	.w4(32'hba1016a3),
	.w5(32'hba326705),
	.w6(32'hbab4ed5c),
	.w7(32'hba367ef7),
	.w8(32'h395594b9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a2cf3),
	.w1(32'h3995003f),
	.w2(32'h3a98af2f),
	.w3(32'hb9f3497b),
	.w4(32'h39b05e96),
	.w5(32'hba1cd050),
	.w6(32'hba4f9898),
	.w7(32'h39bd343a),
	.w8(32'h3a0af2fb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa39210),
	.w1(32'hba5ce6e3),
	.w2(32'h37916263),
	.w3(32'h398f64a0),
	.w4(32'hbb04d61a),
	.w5(32'h39d9d294),
	.w6(32'hbb070802),
	.w7(32'hba8d883c),
	.w8(32'h39a44fba),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce05be),
	.w1(32'h393b2960),
	.w2(32'h3a616a4e),
	.w3(32'h394ab5c8),
	.w4(32'h39e67fe2),
	.w5(32'hba546063),
	.w6(32'h39c3ba92),
	.w7(32'h3a44a5cb),
	.w8(32'hb8bf4243),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391323fa),
	.w1(32'hb9c256ef),
	.w2(32'h3a5527a5),
	.w3(32'hba0a4b6c),
	.w4(32'hb9b5627e),
	.w5(32'hb883a669),
	.w6(32'hba8189ca),
	.w7(32'hb99e5d68),
	.w8(32'hb9083ce5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395725d9),
	.w1(32'h38843b8a),
	.w2(32'hb9a2b407),
	.w3(32'hb9e21c16),
	.w4(32'hba1d6356),
	.w5(32'hb8c42a79),
	.w6(32'hba32d678),
	.w7(32'hba18ce75),
	.w8(32'h39f52d15),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc611a),
	.w1(32'hba32e3c6),
	.w2(32'hb7d245d9),
	.w3(32'hb8a181b2),
	.w4(32'hb9c0a0b5),
	.w5(32'h38a6f496),
	.w6(32'hba1493c5),
	.w7(32'hba233e8b),
	.w8(32'h3ac46705),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbad88),
	.w1(32'h3a29b813),
	.w2(32'h3aeb7e9e),
	.w3(32'hbaadcb34),
	.w4(32'h3a123b8c),
	.w5(32'h3a6af762),
	.w6(32'hb93fe1c7),
	.w7(32'h3a364524),
	.w8(32'h3a4ac0ca),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f76e),
	.w1(32'h3a4d8029),
	.w2(32'h3a62f7ce),
	.w3(32'h3a483a78),
	.w4(32'hb9db0a8e),
	.w5(32'h3b28d2db),
	.w6(32'h39e85341),
	.w7(32'h3882125c),
	.w8(32'h37cc6ee2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa365cd),
	.w1(32'h3a96b291),
	.w2(32'hb9f79372),
	.w3(32'h3a745c23),
	.w4(32'h3b2b8510),
	.w5(32'hbae49761),
	.w6(32'h3aab3e59),
	.w7(32'h3aa91a2c),
	.w8(32'hba925da8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bb05e),
	.w1(32'hba0ee0fa),
	.w2(32'h3aff642d),
	.w3(32'hbb5ca435),
	.w4(32'hba599c8f),
	.w5(32'h3bde6616),
	.w6(32'hbb652698),
	.w7(32'hba3a5364),
	.w8(32'h3ab2b0fe),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b344973),
	.w1(32'h3bcaf8ce),
	.w2(32'hbcc569f8),
	.w3(32'h3bfdb41f),
	.w4(32'h3b8e1a26),
	.w5(32'hbcaf8365),
	.w6(32'h3b4cec7a),
	.w7(32'h3b197175),
	.w8(32'hbc003b5f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc75394),
	.w1(32'hbc799217),
	.w2(32'h39f4c9c0),
	.w3(32'hbd070c4b),
	.w4(32'hbc84e505),
	.w5(32'h3b8b51fc),
	.w6(32'hbcbcc49e),
	.w7(32'hbc57d1ed),
	.w8(32'h3b00353f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b864366),
	.w1(32'hba30d9e1),
	.w2(32'h3c166dcc),
	.w3(32'h3c0fb208),
	.w4(32'h3b4a31c0),
	.w5(32'h3c3cda14),
	.w6(32'h3b887d87),
	.w7(32'h3b86edb2),
	.w8(32'h3bbf5263),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ad9a5),
	.w1(32'h3b905d68),
	.w2(32'hbb5349f9),
	.w3(32'h3c650c13),
	.w4(32'h3cc1d762),
	.w5(32'hbc88c774),
	.w6(32'h3c1e4556),
	.w7(32'h3cd32567),
	.w8(32'hbc88e830),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf8be),
	.w1(32'h3c121280),
	.w2(32'hbbd44f6f),
	.w3(32'hbbe81958),
	.w4(32'h3c513c9f),
	.w5(32'h3b0e8a5e),
	.w6(32'hbc5a28a8),
	.w7(32'h3b6229f9),
	.w8(32'hbbdbaa27),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87dcb4),
	.w1(32'hbbff8a6f),
	.w2(32'h3bb982cf),
	.w3(32'h3ba1a2a3),
	.w4(32'hbb0ee816),
	.w5(32'hbba7f261),
	.w6(32'hbaa88309),
	.w7(32'hbc05966a),
	.w8(32'hbc273921),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37c8ec),
	.w1(32'hbc9ca505),
	.w2(32'hbb94d455),
	.w3(32'hbd09c2d3),
	.w4(32'hbd095057),
	.w5(32'hbb87d2be),
	.w6(32'hbd1cffe9),
	.w7(32'hbc909310),
	.w8(32'hbbc2a34a),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdf3ec),
	.w1(32'hbacf10e9),
	.w2(32'h3bc96f9c),
	.w3(32'hbbac1492),
	.w4(32'hbb98a0a2),
	.w5(32'h3cabf8b1),
	.w6(32'hbb7086d9),
	.w7(32'hbbc0bd60),
	.w8(32'h3c24b1c3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc418a9),
	.w1(32'hbbebd905),
	.w2(32'h3b3bcc1d),
	.w3(32'h3b965c78),
	.w4(32'h3b85ae92),
	.w5(32'h3c8ea813),
	.w6(32'h3c13b5a2),
	.w7(32'h3b4f8de9),
	.w8(32'h3bb2dd8b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfff8ac),
	.w1(32'hbbcd20de),
	.w2(32'hbbac4a7f),
	.w3(32'h3c82434c),
	.w4(32'hbb56f452),
	.w5(32'hbb99ff14),
	.w6(32'h3bd899e6),
	.w7(32'hbbc89718),
	.w8(32'h3bd355f5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f102),
	.w1(32'hbbb18ccb),
	.w2(32'hbc01c790),
	.w3(32'hbbd0352a),
	.w4(32'h3a395149),
	.w5(32'hbc9b2144),
	.w6(32'h3c338a54),
	.w7(32'h3bf0f71b),
	.w8(32'hbc199f18),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e97a7),
	.w1(32'hb95a0a2c),
	.w2(32'hbbaa06f1),
	.w3(32'hba9d09a9),
	.w4(32'h3bcb1171),
	.w5(32'hbc2d66ca),
	.w6(32'hbb700745),
	.w7(32'h3b8a7636),
	.w8(32'hbc27a6a4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceb38d),
	.w1(32'h3b9275ed),
	.w2(32'hbc2285f8),
	.w3(32'hbc4b86cb),
	.w4(32'hba52b4d9),
	.w5(32'hbc3428ea),
	.w6(32'hbbaec9c3),
	.w7(32'h3bdd6f60),
	.w8(32'hbbfa5b46),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02b8bb),
	.w1(32'h3bb07ef1),
	.w2(32'h3b1263ee),
	.w3(32'hbc6a3aef),
	.w4(32'h3a2f9fd3),
	.w5(32'hbb962366),
	.w6(32'hbc266ab8),
	.w7(32'hbb19d19f),
	.w8(32'h3bf910ba),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90258e),
	.w1(32'h3c17bb90),
	.w2(32'hbbbe8d82),
	.w3(32'h3bdad737),
	.w4(32'h3c42d015),
	.w5(32'hbc0491c2),
	.w6(32'h3c01d369),
	.w7(32'h3c71892f),
	.w8(32'hbb8d1294),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3718436e),
	.w1(32'h3b2817b7),
	.w2(32'hbc43fc2a),
	.w3(32'hbb1ea932),
	.w4(32'h3af8f263),
	.w5(32'hbcdde57c),
	.w6(32'h3aca0df8),
	.w7(32'h3b5fcb57),
	.w8(32'hbc90a5af),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd12b7ee),
	.w1(32'hbc66076f),
	.w2(32'hbb7d0f96),
	.w3(32'hbd21b8fa),
	.w4(32'hbcb42430),
	.w5(32'hbc13bf17),
	.w6(32'hbd1affc0),
	.w7(32'hbc5473bc),
	.w8(32'hbc5f0383),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2a437),
	.w1(32'hbbcd48e3),
	.w2(32'hbb42a401),
	.w3(32'hbbe3947c),
	.w4(32'hbb2e441b),
	.w5(32'hbadb4f18),
	.w6(32'hbbc1179b),
	.w7(32'h3bee9827),
	.w8(32'h3c0c03e8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39dced),
	.w1(32'hba61bc85),
	.w2(32'hba6ce582),
	.w3(32'hbb7d97f2),
	.w4(32'hbc18cf42),
	.w5(32'h3ba96c36),
	.w6(32'h3a7cb91e),
	.w7(32'h3bae8ea6),
	.w8(32'h3c642586),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f416a),
	.w1(32'hbc146236),
	.w2(32'h3aecec83),
	.w3(32'hbcc61765),
	.w4(32'hbc97bd9b),
	.w5(32'hbb4c3cc7),
	.w6(32'hbc69b9ae),
	.w7(32'hbc8189bf),
	.w8(32'hb9b409c2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82097ca),
	.w1(32'h3b337cb6),
	.w2(32'hbbe3d9f1),
	.w3(32'hbb68023d),
	.w4(32'hbaa7d7a3),
	.w5(32'hbba62142),
	.w6(32'hba326199),
	.w7(32'h3aef013c),
	.w8(32'hbb0470ef),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b0487),
	.w1(32'h3bbd65b6),
	.w2(32'h3c253e96),
	.w3(32'hbc83d1e2),
	.w4(32'hbc1b020d),
	.w5(32'h3a8356a6),
	.w6(32'hbc8e5f39),
	.w7(32'h3bafad6e),
	.w8(32'hbc409b6f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39945619),
	.w1(32'hbbe7bea5),
	.w2(32'hbc3ba750),
	.w3(32'hbb8fe8d6),
	.w4(32'hbb9429f0),
	.w5(32'hbc9eaa73),
	.w6(32'h3ba0c8ab),
	.w7(32'h3b2944f2),
	.w8(32'hbc96be31),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79a181),
	.w1(32'h39bec402),
	.w2(32'h3c4430f9),
	.w3(32'hbc8a52df),
	.w4(32'h3c4c2a35),
	.w5(32'h3b4595bf),
	.w6(32'hbb8cb941),
	.w7(32'h3cafb487),
	.w8(32'h3aa1c2d0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0740d0),
	.w1(32'h3b1748ae),
	.w2(32'h3b963ded),
	.w3(32'h3b278855),
	.w4(32'h3be8cbbb),
	.w5(32'hbb9d748c),
	.w6(32'h3c1bb4a5),
	.w7(32'h3c4566ba),
	.w8(32'h3bbfc0c3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b8216),
	.w1(32'h3c15fc4b),
	.w2(32'hbcc63d0f),
	.w3(32'hbbef1e16),
	.w4(32'h3bf65dc7),
	.w5(32'hbc538ff9),
	.w6(32'h3c5f77cd),
	.w7(32'h3c66e20c),
	.w8(32'h3ba3cbcd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8468e4),
	.w1(32'hbbe04084),
	.w2(32'hbbf10cf5),
	.w3(32'hbc92e446),
	.w4(32'hbbb576d7),
	.w5(32'hbcac45b9),
	.w6(32'h3c161c88),
	.w7(32'h3bfbdf50),
	.w8(32'hbcb85e19),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bee5e),
	.w1(32'hbc07d633),
	.w2(32'hbca445ec),
	.w3(32'hbcbbb70d),
	.w4(32'hbce52ae4),
	.w5(32'hbca5e347),
	.w6(32'hbd057927),
	.w7(32'hbc4b9364),
	.w8(32'hbc58915b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7f877),
	.w1(32'h3c30bc39),
	.w2(32'hba087ee7),
	.w3(32'hbc868fec),
	.w4(32'h3c103932),
	.w5(32'hbb5e2b9b),
	.w6(32'hbc792efa),
	.w7(32'hba50ea7b),
	.w8(32'h3ac1b21e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f2ada),
	.w1(32'hbb1477c3),
	.w2(32'hbaa98829),
	.w3(32'hbc2a16c9),
	.w4(32'hbc3c8950),
	.w5(32'h3a0ea3ff),
	.w6(32'hbbd99522),
	.w7(32'hbc44605b),
	.w8(32'h3b0abb4e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ce12),
	.w1(32'h3baf685c),
	.w2(32'h3a5bbabe),
	.w3(32'h3bd7b434),
	.w4(32'h3c578cc7),
	.w5(32'hbb5338e6),
	.w6(32'h3bb5e300),
	.w7(32'h3c2197af),
	.w8(32'hbb33ee81),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3fe70),
	.w1(32'h3be6117b),
	.w2(32'h3b1f22f5),
	.w3(32'h3a364d16),
	.w4(32'h3c2a4d59),
	.w5(32'h3bab4ea2),
	.w6(32'h3ac090c4),
	.w7(32'h3b5c8acd),
	.w8(32'h3b8d42e8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182adc),
	.w1(32'hbb269b59),
	.w2(32'hbc107ee2),
	.w3(32'h3c5fa5e0),
	.w4(32'h3ba7c860),
	.w5(32'h3b96b16e),
	.w6(32'h3bceff85),
	.w7(32'h3bf7f398),
	.w8(32'h3b9be94f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55aa5e),
	.w1(32'h3c0fdf58),
	.w2(32'hbbfd97be),
	.w3(32'h3aeb328a),
	.w4(32'h3bd6e40c),
	.w5(32'h3acd782d),
	.w6(32'h3b8712ce),
	.w7(32'h3b335d6d),
	.w8(32'h3b623f54),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc308539),
	.w1(32'hbbca7eca),
	.w2(32'h3c0661fa),
	.w3(32'hbc0553d4),
	.w4(32'hba040d30),
	.w5(32'h3c155126),
	.w6(32'h3a6d0f32),
	.w7(32'hbb2c75e9),
	.w8(32'h3b0d058a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77eed),
	.w1(32'h3c082983),
	.w2(32'h3b1c551f),
	.w3(32'h3c5f27e9),
	.w4(32'h3c5e89a7),
	.w5(32'hbb83d2ec),
	.w6(32'h3bc68ee3),
	.w7(32'h3c28efdc),
	.w8(32'hbbd2e44b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3907b8d6),
	.w1(32'h3a5d5038),
	.w2(32'h3ab9a4a3),
	.w3(32'h3b2556c9),
	.w4(32'h3bb37de6),
	.w5(32'h3a8967d7),
	.w6(32'h3bb3e920),
	.w7(32'h3bf4ddf3),
	.w8(32'hba9d5fb1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9f3ac),
	.w1(32'h3bede408),
	.w2(32'hbc002afd),
	.w3(32'h3be59637),
	.w4(32'h3bdbce97),
	.w5(32'hba28b773),
	.w6(32'hba8601a4),
	.w7(32'h3ab4a226),
	.w8(32'hbbb9966f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06fdfb),
	.w1(32'hbb7f2122),
	.w2(32'h3bd7c730),
	.w3(32'h3c102dd2),
	.w4(32'h3b7a7901),
	.w5(32'hba9342d2),
	.w6(32'h3b735b2e),
	.w7(32'hbaab1e5e),
	.w8(32'h39e68765),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb81be2),
	.w1(32'h3a883afc),
	.w2(32'hbb0254c9),
	.w3(32'h3c1736ab),
	.w4(32'h3b81c410),
	.w5(32'h3982ab0c),
	.w6(32'h3c2683f2),
	.w7(32'h3c29da55),
	.w8(32'h3a09a521),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35f5df),
	.w1(32'h3b8f0a10),
	.w2(32'h3c041aa9),
	.w3(32'h3c5cca55),
	.w4(32'h3b70be65),
	.w5(32'h3c29d311),
	.w6(32'h3ac25b15),
	.w7(32'h3b8c103c),
	.w8(32'h3bbd0fbc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b050bd5),
	.w1(32'hb9e3a664),
	.w2(32'h3ab3d35a),
	.w3(32'h3bac70d5),
	.w4(32'h3b1f4c76),
	.w5(32'hbb443fa6),
	.w6(32'hb927de94),
	.w7(32'hbae6f70f),
	.w8(32'hbb8d880a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a168950),
	.w1(32'h3c19bce1),
	.w2(32'hba87d039),
	.w3(32'hbc3a27a7),
	.w4(32'h3b13f9a0),
	.w5(32'h3b7380f0),
	.w6(32'hbbb21de7),
	.w7(32'h3bd1010a),
	.w8(32'h3bff1ed5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23fe1d),
	.w1(32'h3c399412),
	.w2(32'hbbe72bc8),
	.w3(32'hbaba1491),
	.w4(32'h3c4d5cf3),
	.w5(32'hbbdb930f),
	.w6(32'h3b38361f),
	.w7(32'h3b96e03f),
	.w8(32'h3bd9ba86),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb456def),
	.w1(32'h3c0c0c80),
	.w2(32'hbc4f0755),
	.w3(32'h3af371ad),
	.w4(32'hbb8d91ae),
	.w5(32'hbc953ca2),
	.w6(32'h3bc43dea),
	.w7(32'hb9fed11d),
	.w8(32'hbcdf838f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae7ebb),
	.w1(32'h3c6579d4),
	.w2(32'h3b5f47ff),
	.w3(32'hbc13dc17),
	.w4(32'h3c601f48),
	.w5(32'h3ba37b96),
	.w6(32'hbca5f082),
	.w7(32'h395df3fd),
	.w8(32'h3baaaa9b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad072),
	.w1(32'h3b3a5aee),
	.w2(32'hbcaca84c),
	.w3(32'h3b83f9bb),
	.w4(32'h3a8899f2),
	.w5(32'hbce62358),
	.w6(32'h3b92b9dd),
	.w7(32'h3bab2992),
	.w8(32'hbc7d1d44),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84ac7f),
	.w1(32'hbb9da8bc),
	.w2(32'h3bc34ac9),
	.w3(32'hbcb9c68e),
	.w4(32'hbbcf3023),
	.w5(32'h3af24983),
	.w6(32'hbc48df8a),
	.w7(32'h3b4c1b8d),
	.w8(32'h3b133be8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ea17d),
	.w1(32'h3c1be90e),
	.w2(32'h3bd9596d),
	.w3(32'h3adaa3bf),
	.w4(32'h3b810369),
	.w5(32'h3a723687),
	.w6(32'hbb7cc29e),
	.w7(32'h3bf54d6e),
	.w8(32'hbc01d69e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf57840),
	.w1(32'h3bde3e8a),
	.w2(32'hbb5ca492),
	.w3(32'hbaef4e7a),
	.w4(32'h37c4c3e3),
	.w5(32'h3b8ec199),
	.w6(32'h3b988422),
	.w7(32'h3c0e6fed),
	.w8(32'h3bfc543c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52ebd4),
	.w1(32'h3b0df25d),
	.w2(32'hbaf888b4),
	.w3(32'hbc4f733d),
	.w4(32'hbc149c8b),
	.w5(32'hba9a4591),
	.w6(32'hbc1f4feb),
	.w7(32'hb9d6cfd7),
	.w8(32'hbabcf9c1),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd77195),
	.w1(32'h39a90e4f),
	.w2(32'h3c520ac1),
	.w3(32'hbbb93a3d),
	.w4(32'h39319dba),
	.w5(32'h3be2a65c),
	.w6(32'hbbc97ce1),
	.w7(32'h3b0e80a5),
	.w8(32'h3b8c3c2f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b186add),
	.w1(32'hba39d075),
	.w2(32'hbb97f0ee),
	.w3(32'hbb2f5e0b),
	.w4(32'hba87713f),
	.w5(32'hbb68dcc2),
	.w6(32'hbb1774ff),
	.w7(32'h3c069726),
	.w8(32'hbba80289),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab11c),
	.w1(32'hbb32189f),
	.w2(32'h3b6aad69),
	.w3(32'h3c116856),
	.w4(32'h3b87076e),
	.w5(32'h3bad78c5),
	.w6(32'h3bc7bd6e),
	.w7(32'h3a1d1b28),
	.w8(32'hbaaa27cd),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3cbbd),
	.w1(32'hbc6ab7d2),
	.w2(32'hb95a13e8),
	.w3(32'hbd022b2a),
	.w4(32'hbc96d066),
	.w5(32'h3c23ee18),
	.w6(32'hbcf5065d),
	.w7(32'hbc6b930c),
	.w8(32'h3c9cc9a8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e0d8a),
	.w1(32'hb920ad2b),
	.w2(32'h3b133be9),
	.w3(32'hbc4fb389),
	.w4(32'hbc27d76a),
	.w5(32'h3c222f54),
	.w6(32'hbaaea26e),
	.w7(32'hbb98b296),
	.w8(32'h3c50ff55),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1636c4),
	.w1(32'h3c70c3b2),
	.w2(32'hbc0e9696),
	.w3(32'h3b85f504),
	.w4(32'h3b7b00c6),
	.w5(32'hbcc86f5f),
	.w6(32'h3c4a7121),
	.w7(32'h3a414727),
	.w8(32'hbcb80c21),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a419b),
	.w1(32'h3b999082),
	.w2(32'hbac119cd),
	.w3(32'hbc8d865a),
	.w4(32'h3be8b729),
	.w5(32'h3aa8eef9),
	.w6(32'hbbe8312a),
	.w7(32'h3c9807af),
	.w8(32'h3b4523b7),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc28753),
	.w1(32'hbb9c6af1),
	.w2(32'hbb92f213),
	.w3(32'h3ba74937),
	.w4(32'hbb9eef5d),
	.w5(32'hbbb7bed3),
	.w6(32'h3b8c6676),
	.w7(32'hbbf8bb68),
	.w8(32'hbb74c34d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f16e2),
	.w1(32'hbae4af7b),
	.w2(32'h3bea7256),
	.w3(32'hbbce8600),
	.w4(32'hbb40adc0),
	.w5(32'h3ad4409b),
	.w6(32'hbb36daf7),
	.w7(32'hb884920a),
	.w8(32'hbb961957),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc349be),
	.w1(32'hb9b54452),
	.w2(32'hba883f10),
	.w3(32'hbaadf00b),
	.w4(32'hba4c6433),
	.w5(32'hbbf2c3bd),
	.w6(32'h39f4e4fc),
	.w7(32'h3c0e60c7),
	.w8(32'hbb95b8ab),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91666),
	.w1(32'hbbbf735e),
	.w2(32'hbb5c1add),
	.w3(32'hbbe583fd),
	.w4(32'hbbbe9df0),
	.w5(32'h3b2e778a),
	.w6(32'hba05923a),
	.w7(32'h3c1565fd),
	.w8(32'hb936f16d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7715),
	.w1(32'hbbbe9085),
	.w2(32'h3c3df3f5),
	.w3(32'h3b29d9fc),
	.w4(32'hbb8ea073),
	.w5(32'h3c8ec8f2),
	.w6(32'h3af55a21),
	.w7(32'hbc082324),
	.w8(32'h3bf13e0d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dfde9),
	.w1(32'h3aa816e6),
	.w2(32'hbad9d9d4),
	.w3(32'h3cdc6a42),
	.w4(32'h3b79e268),
	.w5(32'hb8ae7c5f),
	.w6(32'h3c7e4fc7),
	.w7(32'hbc18d711),
	.w8(32'hb9da2d7c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac04f6),
	.w1(32'h3af9c5df),
	.w2(32'hbb39e457),
	.w3(32'hbb8e60b3),
	.w4(32'h3b5a6da7),
	.w5(32'hbb78c231),
	.w6(32'hbb835eb7),
	.w7(32'h3b4ed3dc),
	.w8(32'hba1b6a44),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7e892),
	.w1(32'h3baaa5e7),
	.w2(32'h3c2a1527),
	.w3(32'hbb075dc2),
	.w4(32'h3ba87d7b),
	.w5(32'h3b976692),
	.w6(32'hba3bd010),
	.w7(32'h3b8b74ee),
	.w8(32'h3b8bf1fe),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35c585),
	.w1(32'h3bde1bca),
	.w2(32'hbb9211db),
	.w3(32'h3be03ba0),
	.w4(32'h3acc18e8),
	.w5(32'hbd199ee2),
	.w6(32'h3bcf8f30),
	.w7(32'hbb6771d4),
	.w8(32'hbce1da0f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97986c),
	.w1(32'hbc5ccb5a),
	.w2(32'hbc8cc867),
	.w3(32'hbd32796d),
	.w4(32'hbd361b0b),
	.w5(32'hbccebf43),
	.w6(32'hbd0dbac7),
	.w7(32'hbcdd7ba0),
	.w8(32'hbbffbd86),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb41e20),
	.w1(32'hbabb355c),
	.w2(32'hbbc396c2),
	.w3(32'hbcd048cc),
	.w4(32'hbc498810),
	.w5(32'h3b42ef50),
	.w6(32'hbc54c1d5),
	.w7(32'h3b2dd434),
	.w8(32'h3c24675c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd75be6),
	.w1(32'h3c1a7aea),
	.w2(32'h3bc47032),
	.w3(32'h3b271249),
	.w4(32'h3be15403),
	.w5(32'h3c59c6b5),
	.w6(32'h3bfe63cf),
	.w7(32'h3aa1d848),
	.w8(32'hbb3bab8a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c286185),
	.w1(32'h3c7ae517),
	.w2(32'hbbcc6ad2),
	.w3(32'h3bb529bb),
	.w4(32'h3c44f544),
	.w5(32'hbb827f6f),
	.w6(32'h3bb98934),
	.w7(32'h3b44f1e9),
	.w8(32'hbadb0aed),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05d7f),
	.w1(32'hbc24d941),
	.w2(32'hbb93efd2),
	.w3(32'hbaa383a8),
	.w4(32'hbc4fa2f3),
	.w5(32'hbbbce618),
	.w6(32'h3aaaeda7),
	.w7(32'hbc0b977c),
	.w8(32'h3a92624e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae67e93),
	.w1(32'h3c776173),
	.w2(32'hbacecf45),
	.w3(32'h39ab36d1),
	.w4(32'h3c3cfae8),
	.w5(32'h3b1a4300),
	.w6(32'hbad4f1fe),
	.w7(32'h3c878db2),
	.w8(32'hba604e41),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6a0a3),
	.w1(32'h3c7b6c3d),
	.w2(32'hb953383b),
	.w3(32'h3b8e8c41),
	.w4(32'h3c941e0f),
	.w5(32'hbbcb1793),
	.w6(32'h3ba03dcb),
	.w7(32'h3c8860f5),
	.w8(32'hbbc8e09a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa78a),
	.w1(32'h390ebe71),
	.w2(32'h3c4c03b4),
	.w3(32'hbb8699c5),
	.w4(32'hbb852f99),
	.w5(32'hbba0555b),
	.w6(32'hbaf2db34),
	.w7(32'h3a88ebb5),
	.w8(32'hbc0a047c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add306e),
	.w1(32'h3aa2c1b4),
	.w2(32'h3c66d00e),
	.w3(32'hbc8fa580),
	.w4(32'hbb630530),
	.w5(32'h3becd0d0),
	.w6(32'hbbe2ea9b),
	.w7(32'h3bc73255),
	.w8(32'h3c5365b7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5b086),
	.w1(32'h3c219b7f),
	.w2(32'h3c3cbab1),
	.w3(32'h3b02f7f6),
	.w4(32'h3c360b45),
	.w5(32'h3b80168c),
	.w6(32'h3c54329c),
	.w7(32'h3c7bd4be),
	.w8(32'h38439c95),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb42d26),
	.w1(32'h3bf86286),
	.w2(32'hba50a29b),
	.w3(32'hbb83469d),
	.w4(32'h3c1d2207),
	.w5(32'hbbd969d4),
	.w6(32'h3b80face),
	.w7(32'h3c466b1c),
	.w8(32'hbb49e214),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d0d15),
	.w1(32'h3c6d16e2),
	.w2(32'hbb21ef50),
	.w3(32'hbbce4e0c),
	.w4(32'h3c46b6bb),
	.w5(32'h3b5dc176),
	.w6(32'hbb809e2c),
	.w7(32'h3c517acb),
	.w8(32'h3b8cd42d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25d6dc),
	.w1(32'h3c084111),
	.w2(32'hbbfa5dd8),
	.w3(32'hbc1db774),
	.w4(32'hbb0ead55),
	.w5(32'h3a18f142),
	.w6(32'hbb794a6f),
	.w7(32'hbbacc1d9),
	.w8(32'h3bf1da2f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854039),
	.w1(32'h3c60f2ce),
	.w2(32'h3c4b8d2c),
	.w3(32'h3923b9ad),
	.w4(32'h3c030cba),
	.w5(32'h3c274a4f),
	.w6(32'hba15fb4b),
	.w7(32'h3b5acd38),
	.w8(32'h3c0d49b5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3238c3),
	.w1(32'h3c896f2e),
	.w2(32'h3ab6ea89),
	.w3(32'h3c3de25d),
	.w4(32'h3caa12d1),
	.w5(32'hbb14808c),
	.w6(32'h3c46b4eb),
	.w7(32'h3cae8936),
	.w8(32'h3b8f1d76),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f3ab6),
	.w1(32'h3c286ae5),
	.w2(32'h3c017cd4),
	.w3(32'h3bd72ad2),
	.w4(32'h3c1fe4e2),
	.w5(32'h3bdb5b30),
	.w6(32'h3be8cf23),
	.w7(32'h3c5b5487),
	.w8(32'h3bf6eca1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ad4fc),
	.w1(32'h3b5a9250),
	.w2(32'h3c465136),
	.w3(32'hbb8cdfb9),
	.w4(32'h3c1fbbd2),
	.w5(32'h3c4caa6c),
	.w6(32'hbbf9b6d8),
	.w7(32'h3c5c176d),
	.w8(32'hbbfed6cd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c6ff9),
	.w1(32'hbc504509),
	.w2(32'hbb917876),
	.w3(32'hbbfc9544),
	.w4(32'hbce49290),
	.w5(32'h3b895c4c),
	.w6(32'hbc7d3a8e),
	.w7(32'hbc72bd3c),
	.w8(32'h3b1ac940),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27d542),
	.w1(32'h3c7b3a2c),
	.w2(32'hb8fc0b80),
	.w3(32'h3c1f5bc9),
	.w4(32'h3c67f161),
	.w5(32'hbc0f002f),
	.w6(32'h3c5a5681),
	.w7(32'h3ca25eab),
	.w8(32'hbc1bcad1),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae398),
	.w1(32'h3a366e40),
	.w2(32'h3b29c297),
	.w3(32'hbc27897b),
	.w4(32'hbc7132be),
	.w5(32'h3c15ab56),
	.w6(32'hbca19627),
	.w7(32'hbc2c2c19),
	.w8(32'h3c294aae),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f5d36),
	.w1(32'hbb227a38),
	.w2(32'h3b09eab6),
	.w3(32'hb9ed6a05),
	.w4(32'h3a5740ec),
	.w5(32'h3a9bf978),
	.w6(32'h3b774821),
	.w7(32'hbaa52f84),
	.w8(32'h3beea7a2),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39318f5b),
	.w1(32'hbad7abf6),
	.w2(32'h3b52bffa),
	.w3(32'hba4f2a15),
	.w4(32'h3ab9bfa0),
	.w5(32'h3aca55ef),
	.w6(32'h3bce3868),
	.w7(32'h3b75ef22),
	.w8(32'h3a8a82ce),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05fa94),
	.w1(32'h3b47aefc),
	.w2(32'hbac44947),
	.w3(32'hba89c983),
	.w4(32'h3bd87e27),
	.w5(32'hbb383721),
	.w6(32'hb93fd540),
	.w7(32'h3bd083c8),
	.w8(32'h39bd63dc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b7328),
	.w1(32'h3c379a70),
	.w2(32'hbb11309c),
	.w3(32'h3b9299f3),
	.w4(32'h3c5170c6),
	.w5(32'hb8001912),
	.w6(32'h3ab3843d),
	.w7(32'h3c64fd62),
	.w8(32'h3b7fa968),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25a17a),
	.w1(32'h3b85d348),
	.w2(32'hbc101c61),
	.w3(32'h3bed4cb6),
	.w4(32'h3c754190),
	.w5(32'hbc24be8d),
	.w6(32'h3b621bea),
	.w7(32'h3c2e7ed3),
	.w8(32'h3ba9e892),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6d947),
	.w1(32'hbab68634),
	.w2(32'h3b3c095d),
	.w3(32'hbc17a24e),
	.w4(32'hbbe10cda),
	.w5(32'h3b816fbe),
	.w6(32'h3b474b87),
	.w7(32'h3bdc3ea6),
	.w8(32'h3b9670ec),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1c956),
	.w1(32'hbab18947),
	.w2(32'hbbe09219),
	.w3(32'h3b4daf64),
	.w4(32'hbaddf6c8),
	.w5(32'hbc08b79d),
	.w6(32'h3aba929b),
	.w7(32'h39a1dd55),
	.w8(32'hbbc3e758),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb39d6),
	.w1(32'hbbb7cfef),
	.w2(32'h3bf6acc2),
	.w3(32'hbbc92719),
	.w4(32'hbbcb3f29),
	.w5(32'h3c805a64),
	.w6(32'hbb737a0a),
	.w7(32'hbb1387fc),
	.w8(32'h3c4c70bc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc474b1c),
	.w1(32'hbce98212),
	.w2(32'hbb3f4c4e),
	.w3(32'hbca8ca52),
	.w4(32'hbcf42216),
	.w5(32'hbb34ad7a),
	.w6(32'hbc32830f),
	.w7(32'hbc77f5ee),
	.w8(32'h39c5f30e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5794f8),
	.w1(32'h3b623353),
	.w2(32'h3b7cb0f4),
	.w3(32'h3bb64b2c),
	.w4(32'h3bc43b89),
	.w5(32'hbc117d3d),
	.w6(32'h3bfafd5a),
	.w7(32'h3bf0e0c0),
	.w8(32'hbbd19ab5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d929),
	.w1(32'h3b9580a4),
	.w2(32'h3be4b3e6),
	.w3(32'h3a9839db),
	.w4(32'h3b1211d5),
	.w5(32'hba1bb830),
	.w6(32'hbaae3b5e),
	.w7(32'h3bd8868b),
	.w8(32'h3b55a90e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03577b),
	.w1(32'h3bccf2ae),
	.w2(32'h3c193d1f),
	.w3(32'hbb479652),
	.w4(32'h3bb768b6),
	.w5(32'hbb5c92eb),
	.w6(32'h3c02d63f),
	.w7(32'h3c09a69f),
	.w8(32'h3b5a4e29),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae05611),
	.w1(32'hbb3bcb80),
	.w2(32'hbbf2c090),
	.w3(32'hbb8d45ef),
	.w4(32'h3a0ff52f),
	.w5(32'hbca2ed22),
	.w6(32'hba90bfcd),
	.w7(32'h3c702ead),
	.w8(32'hbc3abbcb),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule