module layer_10_featuremap_289(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b34f),
	.w1(32'hbbab660b),
	.w2(32'hbaae3206),
	.w3(32'hbb7596d5),
	.w4(32'h3aa4100a),
	.w5(32'hbbfacab4),
	.w6(32'hbc1b060e),
	.w7(32'hb9d33093),
	.w8(32'hbc1b9ab9),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a3461),
	.w1(32'hbbe54b23),
	.w2(32'hbb35e06b),
	.w3(32'hbc29dda3),
	.w4(32'hbbbcfbe6),
	.w5(32'h3b73bb67),
	.w6(32'hbc7552d4),
	.w7(32'hbc2aaa17),
	.w8(32'h3a501a6a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fd09a),
	.w1(32'hbaeca7c1),
	.w2(32'hb798990a),
	.w3(32'h398366f3),
	.w4(32'h3a80338b),
	.w5(32'h39e127e4),
	.w6(32'hbb1ac945),
	.w7(32'h3b133955),
	.w8(32'h3a3ab84a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba708cc0),
	.w1(32'h3b6c96ac),
	.w2(32'h3a6b8017),
	.w3(32'h39b6d8ca),
	.w4(32'hba604996),
	.w5(32'h3b4b336f),
	.w6(32'h3bb40f4a),
	.w7(32'h3ad1f87a),
	.w8(32'h38b430b1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23197c),
	.w1(32'h3bea5f81),
	.w2(32'h3b167681),
	.w3(32'hb9fa48e3),
	.w4(32'hb9522ae5),
	.w5(32'h3ac56811),
	.w6(32'h3a4c5ab3),
	.w7(32'hbb10e787),
	.w8(32'hbaab9e05),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba837253),
	.w1(32'hbaae8af0),
	.w2(32'hba5fa97b),
	.w3(32'h3ae3f649),
	.w4(32'h3af2c5ef),
	.w5(32'hbb61bb40),
	.w6(32'hb90f30dc),
	.w7(32'hba6d5b38),
	.w8(32'hbb97a40c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81265c),
	.w1(32'hba83b93b),
	.w2(32'hbbc7aa72),
	.w3(32'hba874c80),
	.w4(32'h3a9cf93c),
	.w5(32'hbbc83f19),
	.w6(32'hbb04ab62),
	.w7(32'hbbcaec7b),
	.w8(32'hbbac71a9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5ae5e),
	.w1(32'hbc29b465),
	.w2(32'hbc43255c),
	.w3(32'hbc679d17),
	.w4(32'hbb89a36f),
	.w5(32'h398cd58e),
	.w6(32'hbb0579be),
	.w7(32'hbba36722),
	.w8(32'hbaf22bbc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a102),
	.w1(32'hbae87b05),
	.w2(32'h3b07e92f),
	.w3(32'h3b195d98),
	.w4(32'h3b68526d),
	.w5(32'h3b3dc895),
	.w6(32'h3b280f66),
	.w7(32'h3b642cfc),
	.w8(32'hbb661023),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ab155),
	.w1(32'hba255d5b),
	.w2(32'hbae1b118),
	.w3(32'h3b8eca98),
	.w4(32'hbafcc368),
	.w5(32'hbb3890e4),
	.w6(32'h3aee97f9),
	.w7(32'hbb33e826),
	.w8(32'hbb9a7b4c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93aaaa),
	.w1(32'h3a7e235a),
	.w2(32'hba41ba33),
	.w3(32'h3b1ecb70),
	.w4(32'hbae1adb8),
	.w5(32'hbb929a3c),
	.w6(32'h3b15b478),
	.w7(32'hbaf23261),
	.w8(32'hb97676af),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6827),
	.w1(32'h3b74c74c),
	.w2(32'hbb3c2968),
	.w3(32'h3b0424ac),
	.w4(32'h3b6b6482),
	.w5(32'h3912a1e7),
	.w6(32'hbb395d80),
	.w7(32'h3b24b904),
	.w8(32'hbab41d5a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b468ee4),
	.w1(32'hbb2af1e0),
	.w2(32'hba88aa62),
	.w3(32'hbb0640be),
	.w4(32'h3a49765d),
	.w5(32'h3b9a6ee7),
	.w6(32'h39b54911),
	.w7(32'h3b35c4a9),
	.w8(32'hbb1bf0d9),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ed673),
	.w1(32'h3b7336de),
	.w2(32'h3b316e9d),
	.w3(32'h37b56264),
	.w4(32'hbbd0d341),
	.w5(32'hb9e73d74),
	.w6(32'h3b3ef73c),
	.w7(32'hbb7c07e2),
	.w8(32'h37bb02af),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb641701),
	.w1(32'h3ac54bc4),
	.w2(32'h3a5d3a7c),
	.w3(32'hbb1366c6),
	.w4(32'h3883a632),
	.w5(32'h3be2913c),
	.w6(32'h3b48fde9),
	.w7(32'h3b3cc4e3),
	.w8(32'h3c19a1f5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b2084),
	.w1(32'h3bbd8f2a),
	.w2(32'h3b68ed82),
	.w3(32'h3b3f50a9),
	.w4(32'hba24c871),
	.w5(32'hbaf70b3a),
	.w6(32'h3c0b0dfb),
	.w7(32'hbb0e49ee),
	.w8(32'hbb4a73c0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d0c51),
	.w1(32'hbbe3c8d3),
	.w2(32'hba387d79),
	.w3(32'hbbeb97ef),
	.w4(32'h3ba90450),
	.w5(32'hbb075507),
	.w6(32'hbc1f0a1d),
	.w7(32'h3a7dace1),
	.w8(32'hbaf39fc8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeef1ad),
	.w1(32'hbb904ecb),
	.w2(32'hbc1d6773),
	.w3(32'h3aa25554),
	.w4(32'hbbf51652),
	.w5(32'hbc5d049a),
	.w6(32'hb8ed7d07),
	.w7(32'hbbfdb164),
	.w8(32'hbc57f9cb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39123b54),
	.w1(32'hbb7a3574),
	.w2(32'hbb992ff7),
	.w3(32'hbb1a1fe4),
	.w4(32'hbbc49718),
	.w5(32'h3a95d364),
	.w6(32'hbb26b39d),
	.w7(32'hbc0849cd),
	.w8(32'hba9672f5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0069cc),
	.w1(32'h3ac46ab1),
	.w2(32'h3b110f6f),
	.w3(32'h3a8d3250),
	.w4(32'hba844363),
	.w5(32'h3c363127),
	.w6(32'h3ac580aa),
	.w7(32'h39f019c9),
	.w8(32'h3c2b343a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd42266),
	.w1(32'h3c15a070),
	.w2(32'h3c327002),
	.w3(32'h3c034fe9),
	.w4(32'h3b054b5f),
	.w5(32'h3bfaef8b),
	.w6(32'h3c8581f0),
	.w7(32'h3b920f86),
	.w8(32'h3be57019),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee76f),
	.w1(32'h3bc91c5a),
	.w2(32'h3b8c2260),
	.w3(32'h3bd02cae),
	.w4(32'h3b8aae82),
	.w5(32'h3a533d07),
	.w6(32'h3bd3b1b4),
	.w7(32'h3ba99847),
	.w8(32'h3ba92155),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b968a48),
	.w1(32'h3a4d7aa5),
	.w2(32'hbbec87aa),
	.w3(32'h3c1ed43d),
	.w4(32'h3bd38825),
	.w5(32'hbbc4c42d),
	.w6(32'h3b90166e),
	.w7(32'h3b304b62),
	.w8(32'hbc090952),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb031d6b),
	.w1(32'h3bfb01d3),
	.w2(32'h3b331611),
	.w3(32'h3c47642b),
	.w4(32'hbaa0a62e),
	.w5(32'h3bbd22f3),
	.w6(32'h3c72d560),
	.w7(32'h3adbeb95),
	.w8(32'h35242487),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955a7f6),
	.w1(32'h3a1948f8),
	.w2(32'hbb829ab3),
	.w3(32'hbb9290e7),
	.w4(32'h39ee3876),
	.w5(32'h3bff08ce),
	.w6(32'hbc029b25),
	.w7(32'hb9e4a40f),
	.w8(32'h3bc38a99),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac33fb1),
	.w1(32'hbaa08437),
	.w2(32'hb8811a90),
	.w3(32'hbb151a8d),
	.w4(32'h3aa65ca3),
	.w5(32'hba3fb37e),
	.w6(32'h39c008d7),
	.w7(32'h39716b4a),
	.w8(32'h3a13b350),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ad17a),
	.w1(32'hbb2fcec3),
	.w2(32'hbaebc20c),
	.w3(32'hbaaa2d70),
	.w4(32'h3b114446),
	.w5(32'h3ba26971),
	.w6(32'hba65556b),
	.w7(32'h39760de7),
	.w8(32'hbb0a0e68),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391d9543),
	.w1(32'hb8f5e7b7),
	.w2(32'h3b8b609d),
	.w3(32'h3be27867),
	.w4(32'h3bc6b8e8),
	.w5(32'h3c25930d),
	.w6(32'hba96050f),
	.w7(32'h3af9cdc9),
	.w8(32'hbabd44a2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f76b4),
	.w1(32'h3c010bc7),
	.w2(32'hba6c059a),
	.w3(32'h3b96bbe4),
	.w4(32'hbb80e753),
	.w5(32'h3ba68c6b),
	.w6(32'h3c02a7be),
	.w7(32'hbbd33340),
	.w8(32'hbb17b394),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c177),
	.w1(32'h3c0e2751),
	.w2(32'h3bc46e56),
	.w3(32'h3b8df9e1),
	.w4(32'hb9e5932d),
	.w5(32'hb9bc983d),
	.w6(32'h3bcdc145),
	.w7(32'h3aecfece),
	.w8(32'h3adef07e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadc534),
	.w1(32'hbb4dc57d),
	.w2(32'hbb138988),
	.w3(32'h3a0ceef8),
	.w4(32'h3b8d8da2),
	.w5(32'hbb0ca450),
	.w6(32'hbb89c82f),
	.w7(32'h3a687c31),
	.w8(32'hbbeeda58),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae45de),
	.w1(32'h3baa8de6),
	.w2(32'h3b0084c0),
	.w3(32'h3a301aa2),
	.w4(32'h3a1fca75),
	.w5(32'hba147f12),
	.w6(32'h39dd4358),
	.w7(32'h3b947fb0),
	.w8(32'h38411222),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac642a6),
	.w1(32'h3ac09a96),
	.w2(32'h3b0951b3),
	.w3(32'hba81071f),
	.w4(32'hbb56576c),
	.w5(32'hbb76e051),
	.w6(32'h389bac95),
	.w7(32'hba6ec288),
	.w8(32'h3a4524b9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91e279),
	.w1(32'hba3b2fd2),
	.w2(32'hba380f91),
	.w3(32'hbb134b9d),
	.w4(32'hbaa4f7df),
	.w5(32'h3b83da78),
	.w6(32'h3ae0e23b),
	.w7(32'h3a12f31f),
	.w8(32'h3b2ad05c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b949e7b),
	.w1(32'h3bd41a44),
	.w2(32'h3b745fa9),
	.w3(32'h3bb532c0),
	.w4(32'hbaf082fe),
	.w5(32'hb9ee4f7b),
	.w6(32'h3c25ed25),
	.w7(32'hb981f103),
	.w8(32'h3a188160),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e45c3),
	.w1(32'hbb117a10),
	.w2(32'h39a85981),
	.w3(32'h3a7eb29b),
	.w4(32'h3be32a9e),
	.w5(32'h39acb460),
	.w6(32'h3a276ac4),
	.w7(32'h3bb03f2e),
	.w8(32'h3a7f0c0f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc11b8b),
	.w1(32'h3c4d3f2f),
	.w2(32'hbb01bcc0),
	.w3(32'h3b2a4ec2),
	.w4(32'h3c374daf),
	.w5(32'hba45bdae),
	.w6(32'h3b0be6aa),
	.w7(32'h3c134617),
	.w8(32'hbb06b38b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bdbbb),
	.w1(32'hbae3478d),
	.w2(32'h3b86e06b),
	.w3(32'h3aa8efea),
	.w4(32'h3c343552),
	.w5(32'h3ba2e5c4),
	.w6(32'h3bb6d155),
	.w7(32'h3bdf1b9b),
	.w8(32'h3be8cfda),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64670a),
	.w1(32'hbb567ee2),
	.w2(32'hb94ea145),
	.w3(32'hbb849a07),
	.w4(32'h3b3974f3),
	.w5(32'h3c4a07fd),
	.w6(32'hbb26ec10),
	.w7(32'h3abcf07e),
	.w8(32'h3c61d8a2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bbc6f),
	.w1(32'h3c3f034f),
	.w2(32'h3baf18a7),
	.w3(32'h3b7cf140),
	.w4(32'hbb27b7ed),
	.w5(32'h3c03b22d),
	.w6(32'h3c265100),
	.w7(32'h3b382863),
	.w8(32'h3b8cef76),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f1adf5),
	.w1(32'h3c03be6e),
	.w2(32'h3b578421),
	.w3(32'h3ba18a00),
	.w4(32'hbabe9010),
	.w5(32'hbaa4694a),
	.w6(32'h3b5b48cd),
	.w7(32'hba8aa0d7),
	.w8(32'hbb4dd4cd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7dcd73),
	.w1(32'hbb8c4a62),
	.w2(32'hbbdade84),
	.w3(32'hbb70d2e1),
	.w4(32'hb99442ce),
	.w5(32'hbb6b26f3),
	.w6(32'hbb2503ab),
	.w7(32'hbb8ef684),
	.w8(32'hba9d2d61),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f97df8),
	.w1(32'h3b3cb83e),
	.w2(32'h3ad5e8f9),
	.w3(32'h3b75f635),
	.w4(32'h3adb2117),
	.w5(32'hbbb830d5),
	.w6(32'h3c1f03ea),
	.w7(32'hbab54c7e),
	.w8(32'hbb81ef45),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba818a5a),
	.w1(32'hbbc92552),
	.w2(32'hbb837d62),
	.w3(32'hbb9995ad),
	.w4(32'hbafcba6f),
	.w5(32'hbb9b88ef),
	.w6(32'hbbd0a5bb),
	.w7(32'hbc2c9591),
	.w8(32'hbba3a04c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb423bad),
	.w1(32'h3aca4cae),
	.w2(32'h3a41d6f5),
	.w3(32'hbaf4c3f1),
	.w4(32'h37aea5fd),
	.w5(32'h3b226563),
	.w6(32'h3b411e8b),
	.w7(32'h3ae6d9cb),
	.w8(32'hbb414cc4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa32edc),
	.w1(32'hbba5cc5a),
	.w2(32'hba7ffe62),
	.w3(32'hbb19cd07),
	.w4(32'h3b57a183),
	.w5(32'h3ba60500),
	.w6(32'hbc28c7a0),
	.w7(32'h399bbe3f),
	.w8(32'h3b9dade6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da605),
	.w1(32'hba0c3738),
	.w2(32'hba833194),
	.w3(32'hba9bd9ce),
	.w4(32'h3b6967e4),
	.w5(32'h3c4369e2),
	.w6(32'hb86cc7ed),
	.w7(32'h3b0916d7),
	.w8(32'h3c157899),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ace8d),
	.w1(32'h3bacaa4e),
	.w2(32'hbb0257e8),
	.w3(32'h3c72cbae),
	.w4(32'h3b95e9cd),
	.w5(32'hbc4e81cb),
	.w6(32'h3c23dbea),
	.w7(32'h3b74cb10),
	.w8(32'hbc79df3d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ed60b),
	.w1(32'hbb212583),
	.w2(32'h393e71d1),
	.w3(32'h3a139cbb),
	.w4(32'h3ba4d873),
	.w5(32'h3bd03bc8),
	.w6(32'h3ab21daf),
	.w7(32'h3bc3d8b1),
	.w8(32'h3ba3a16a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd061),
	.w1(32'h3bd62a2d),
	.w2(32'h3b47f600),
	.w3(32'h3bd8099a),
	.w4(32'h3b8b8128),
	.w5(32'hba6fb94d),
	.w6(32'h3be8cd03),
	.w7(32'h3ba6d34f),
	.w8(32'hbb78dadd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0172d5),
	.w1(32'h3914fcec),
	.w2(32'hbaf1cd27),
	.w3(32'h3b9e2236),
	.w4(32'h37a9422c),
	.w5(32'hb9e136ac),
	.w6(32'h3b7f27dd),
	.w7(32'hbb792531),
	.w8(32'h3ae3a84f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c0ea3),
	.w1(32'hbb814026),
	.w2(32'h38b1e172),
	.w3(32'hba401d03),
	.w4(32'h3a08f2cb),
	.w5(32'hbb14a98c),
	.w6(32'hbad7bb7b),
	.w7(32'h3a18ce24),
	.w8(32'hbb6ee350),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb443a41),
	.w1(32'h3accef0e),
	.w2(32'hb9188660),
	.w3(32'h3b0bc34e),
	.w4(32'hbb98c13d),
	.w5(32'h3adc67d6),
	.w6(32'hbae54282),
	.w7(32'hbb321aef),
	.w8(32'h3bceb566),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11da2f),
	.w1(32'h3b24c811),
	.w2(32'hbc1f4de3),
	.w3(32'h3bd2b774),
	.w4(32'hbb42503f),
	.w5(32'hbb21bf97),
	.w6(32'h3bc0460a),
	.w7(32'hbb293419),
	.w8(32'hbba2374c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01beae),
	.w1(32'hbb27e558),
	.w2(32'h3b0042cd),
	.w3(32'hba5348cf),
	.w4(32'h3a0f290e),
	.w5(32'h3b6577d5),
	.w6(32'hba60b2c4),
	.w7(32'hb96fc037),
	.w8(32'hbb8bcc47),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fb10),
	.w1(32'h3bb1b599),
	.w2(32'hbb00990c),
	.w3(32'h3abfe6da),
	.w4(32'hbb3b0839),
	.w5(32'h3ba73299),
	.w6(32'h3bd1962f),
	.w7(32'hbbdead9e),
	.w8(32'h3a0f7d16),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dee51),
	.w1(32'h3b8b77b8),
	.w2(32'hbb09ef8d),
	.w3(32'h3b007286),
	.w4(32'hbad35c38),
	.w5(32'h3c13f74a),
	.w6(32'h3baed8df),
	.w7(32'hbb153138),
	.w8(32'h3c110e62),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb78e3),
	.w1(32'h3baed290),
	.w2(32'h3b24f730),
	.w3(32'h3b28957a),
	.w4(32'hbb15d5d7),
	.w5(32'h3b87b598),
	.w6(32'h3bf40e47),
	.w7(32'h3aa93c28),
	.w8(32'h3b76c488),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a975446),
	.w1(32'h3bdf776f),
	.w2(32'h3bb538f0),
	.w3(32'h3ba672e3),
	.w4(32'h3b502e9b),
	.w5(32'hbbd79f6c),
	.w6(32'h3bf0a687),
	.w7(32'h3b854e19),
	.w8(32'hbc14719a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cc6c8),
	.w1(32'hbc59bc69),
	.w2(32'hbc98380e),
	.w3(32'hbc3fd61d),
	.w4(32'hbbb076a1),
	.w5(32'hba780a01),
	.w6(32'hbc743e03),
	.w7(32'hbc6deb33),
	.w8(32'hba300ebb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c54a25),
	.w1(32'h3b289bf6),
	.w2(32'hbb5dc150),
	.w3(32'h3bacb4f6),
	.w4(32'hbb387260),
	.w5(32'hbb9b52b8),
	.w6(32'h3bad649e),
	.w7(32'hba3d2dd1),
	.w8(32'hbc196e86),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8193e),
	.w1(32'hbb9c2bb7),
	.w2(32'hbb5f215f),
	.w3(32'hbba4fd59),
	.w4(32'hbb47a555),
	.w5(32'hbbd4f620),
	.w6(32'hbc1cb6e3),
	.w7(32'hbbd447af),
	.w8(32'hbba5a18c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba90667),
	.w1(32'h3b7eaf92),
	.w2(32'h3b4fd2be),
	.w3(32'hbb4db0be),
	.w4(32'hbab1fc3f),
	.w5(32'h3bea246a),
	.w6(32'hbb5972bc),
	.w7(32'hba9ee979),
	.w8(32'h3b098239),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c20130),
	.w1(32'h3b8786aa),
	.w2(32'h3ad07b07),
	.w3(32'h3b9dfd63),
	.w4(32'hbb6fd4f1),
	.w5(32'h3b8ed683),
	.w6(32'h3bcce575),
	.w7(32'hbb0bef49),
	.w8(32'h3a426bfc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fe840),
	.w1(32'h3b23b8f4),
	.w2(32'h3b309c3c),
	.w3(32'h3b346a40),
	.w4(32'hbaded761),
	.w5(32'hbaf94db7),
	.w6(32'h3bf8b860),
	.w7(32'hbab5bd6f),
	.w8(32'hbaa97449),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14de28),
	.w1(32'hbabb8872),
	.w2(32'h3b3a6110),
	.w3(32'hba8371ab),
	.w4(32'h3b0cb6a0),
	.w5(32'hbaba0d75),
	.w6(32'hbbdca1bb),
	.w7(32'h3a80d125),
	.w8(32'h3b160d15),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f6e4),
	.w1(32'hb8399f60),
	.w2(32'hbbbfd2f3),
	.w3(32'h3abb96d2),
	.w4(32'h3ae020cf),
	.w5(32'hba6e3f86),
	.w6(32'h3aec1634),
	.w7(32'hb929e2fa),
	.w8(32'hbb4e00c2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72faf99),
	.w1(32'hbbe3a891),
	.w2(32'hbb93bdef),
	.w3(32'hbb33db3f),
	.w4(32'h3b5bc16d),
	.w5(32'h3bafe41a),
	.w6(32'hbb4fa1f9),
	.w7(32'h3a65b390),
	.w8(32'hbaa1307e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba981334),
	.w1(32'h38d942ee),
	.w2(32'hbb0f822c),
	.w3(32'h3bac6819),
	.w4(32'hba504e89),
	.w5(32'hbbe40e2b),
	.w6(32'h3bf2de81),
	.w7(32'hbb2c9e97),
	.w8(32'hbbd1e5d5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3e798),
	.w1(32'hbb3fd720),
	.w2(32'h3b1b67c7),
	.w3(32'hbbd002e5),
	.w4(32'h3be146f5),
	.w5(32'h3be547cb),
	.w6(32'h39e58076),
	.w7(32'h3ba1c427),
	.w8(32'h3bed44ac),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa74059),
	.w1(32'hb9d2b817),
	.w2(32'h3b04ee54),
	.w3(32'h3aa7edc4),
	.w4(32'h3ac093ae),
	.w5(32'hbb67153d),
	.w6(32'h3b21d86a),
	.w7(32'hb8c3f461),
	.w8(32'h3b709382),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0052ed),
	.w1(32'hba207d87),
	.w2(32'hbbca0bea),
	.w3(32'hbc03d0c1),
	.w4(32'hba6194a4),
	.w5(32'hbc2ef07d),
	.w6(32'hbb56c47a),
	.w7(32'hbacaa0c2),
	.w8(32'hbc09655a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca8a35),
	.w1(32'hbc18146c),
	.w2(32'hbb5852a3),
	.w3(32'hbbaf5982),
	.w4(32'hb9a9a793),
	.w5(32'hbaab22aa),
	.w6(32'hbc3f4030),
	.w7(32'h3ae4cb9f),
	.w8(32'h3a796403),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58f56e),
	.w1(32'hbb5d6296),
	.w2(32'hbbf741c8),
	.w3(32'hbb8978a1),
	.w4(32'hbbe2c007),
	.w5(32'hbbce11fa),
	.w6(32'hba893595),
	.w7(32'hbc001782),
	.w8(32'hba5ace12),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ef81a),
	.w1(32'hba2162fb),
	.w2(32'hbabef0b2),
	.w3(32'hbb1a14f5),
	.w4(32'hbb104bcb),
	.w5(32'hbba1b4cf),
	.w6(32'h39f2f1d1),
	.w7(32'hbb00f59b),
	.w8(32'hbbc4978a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad81f3d),
	.w1(32'hbba213e2),
	.w2(32'hbbfa1b0f),
	.w3(32'hbab6b6c4),
	.w4(32'hbad61e1c),
	.w5(32'hbb9cd084),
	.w6(32'hbb29c314),
	.w7(32'hbb5e1ea1),
	.w8(32'hbb881818),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5de64),
	.w1(32'hba837a9e),
	.w2(32'hbbd7b60b),
	.w3(32'hba320672),
	.w4(32'hbae74ed5),
	.w5(32'hbc1ae909),
	.w6(32'hbbbafe9e),
	.w7(32'hbc0bdab5),
	.w8(32'hbc0d5ad4),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56a6b6),
	.w1(32'hbb74489c),
	.w2(32'h398d18f0),
	.w3(32'hbb34325d),
	.w4(32'h3925a910),
	.w5(32'hbb85fef9),
	.w6(32'hbb292879),
	.w7(32'h3a0e9ecc),
	.w8(32'hbb024458),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe84f8b),
	.w1(32'hbb91dbb6),
	.w2(32'hbbac2a1d),
	.w3(32'hbba546a9),
	.w4(32'hbba1a752),
	.w5(32'hbb93cd8b),
	.w6(32'hbba10fe2),
	.w7(32'h3884dcb1),
	.w8(32'hbbcb623b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f2c28),
	.w1(32'hbc005d6b),
	.w2(32'hbbb6163e),
	.w3(32'hbb95cddf),
	.w4(32'h3b9e0d00),
	.w5(32'h3bbd2783),
	.w6(32'hbc0f4b0b),
	.w7(32'hb91524f6),
	.w8(32'h3b3a6299),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95be5a),
	.w1(32'h3c119af5),
	.w2(32'h393b959d),
	.w3(32'h3bc24c14),
	.w4(32'hbaf22588),
	.w5(32'hbb185c78),
	.w6(32'h3c6f4a3c),
	.w7(32'h3ba50cf1),
	.w8(32'hbb08fd77),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4614a),
	.w1(32'hba2f06b4),
	.w2(32'hbb86be3d),
	.w3(32'h3a2c4945),
	.w4(32'h3aa232e0),
	.w5(32'hbba8aa14),
	.w6(32'h3abad953),
	.w7(32'hb9ff89d5),
	.w8(32'hbba30381),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb727ed5),
	.w1(32'hbb1a16d8),
	.w2(32'hbb89dc2d),
	.w3(32'h3aca2115),
	.w4(32'h3b39771a),
	.w5(32'hbaa08476),
	.w6(32'hba55c086),
	.w7(32'hbab0b80f),
	.w8(32'hbb2f5ac8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23173a),
	.w1(32'hb9edf206),
	.w2(32'h3af4e26b),
	.w3(32'hbb4bf656),
	.w4(32'hbb3a913f),
	.w5(32'hbafdb4be),
	.w6(32'hba7907ef),
	.w7(32'hbac47c69),
	.w8(32'h3a2f2af7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07718d),
	.w1(32'hbafaecf1),
	.w2(32'hbb19b0c2),
	.w3(32'h3b1d43e9),
	.w4(32'h3b9ce27b),
	.w5(32'hbafcdadc),
	.w6(32'hbb70bedd),
	.w7(32'h394030ac),
	.w8(32'hbc050945),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7faa),
	.w1(32'hbbf24b96),
	.w2(32'hbb3607bf),
	.w3(32'hbb9e8a29),
	.w4(32'h3914c97c),
	.w5(32'hba315b4e),
	.w6(32'hbc3140fa),
	.w7(32'hbb5e8838),
	.w8(32'h39c9f50c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9f7ad),
	.w1(32'hbb6fb42c),
	.w2(32'h38aae036),
	.w3(32'hbba0dadb),
	.w4(32'h3bd38418),
	.w5(32'h3b6fd955),
	.w6(32'hba9855e6),
	.w7(32'h3bbb5ad5),
	.w8(32'h3b413944),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1838f8),
	.w1(32'hba19a2fc),
	.w2(32'h398a50ba),
	.w3(32'h3aa1d369),
	.w4(32'h3b21c0a3),
	.w5(32'hb8a85b0c),
	.w6(32'hbaf434e6),
	.w7(32'h3a4c99d0),
	.w8(32'h3a45742d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada1d1e),
	.w1(32'hbb43ee6d),
	.w2(32'h39cbd2d1),
	.w3(32'hbb2eecd6),
	.w4(32'h3b38bea8),
	.w5(32'h3c357f4d),
	.w6(32'hbac5ed82),
	.w7(32'h3abff0c6),
	.w8(32'hba8c6a0f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf71937),
	.w1(32'h3bd6d675),
	.w2(32'hb9214b0f),
	.w3(32'h3af5271c),
	.w4(32'h3ab364de),
	.w5(32'hbba05b21),
	.w6(32'h3b1ed884),
	.w7(32'hbb0c9151),
	.w8(32'hbbe4efea),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb078723),
	.w1(32'h3c378f3c),
	.w2(32'h3c885550),
	.w3(32'h3c91f85d),
	.w4(32'h3b2bd1a8),
	.w5(32'h3bed2a5c),
	.w6(32'h3c4ffe7b),
	.w7(32'h3c23ef38),
	.w8(32'h3a22a443),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb819324),
	.w1(32'h3be3ade2),
	.w2(32'h3b2c5022),
	.w3(32'h3bdced38),
	.w4(32'h3bf090da),
	.w5(32'hba2ec1d3),
	.w6(32'h3be5047a),
	.w7(32'h3ba79623),
	.w8(32'hbc0d0f49),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10af41),
	.w1(32'h387baad7),
	.w2(32'h3afa8a2a),
	.w3(32'hbaef3d96),
	.w4(32'h3b492808),
	.w5(32'h3c0b62b2),
	.w6(32'hbaa425c0),
	.w7(32'hb88db3af),
	.w8(32'h3b6fc214),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af31066),
	.w1(32'h394060a2),
	.w2(32'h3a5d36f6),
	.w3(32'h3b9ad103),
	.w4(32'h3a8d3c21),
	.w5(32'hbb9c92bd),
	.w6(32'h3ba2c7e5),
	.w7(32'h39cac1f8),
	.w8(32'hbbbc5a5a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1cb08),
	.w1(32'hbb809c6d),
	.w2(32'hbb35caf7),
	.w3(32'h39bd4f62),
	.w4(32'h3b260ad3),
	.w5(32'hbb778640),
	.w6(32'h3baa6452),
	.w7(32'h3a5577c5),
	.w8(32'hba91f95e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4fe2f),
	.w1(32'hbb96d193),
	.w2(32'hbb310ed6),
	.w3(32'hb9894df3),
	.w4(32'h3a9bf573),
	.w5(32'hbac7b259),
	.w6(32'hb9b230e4),
	.w7(32'hbb2a4546),
	.w8(32'hbbad68d7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e347e),
	.w1(32'hbb62f676),
	.w2(32'hbbd340f9),
	.w3(32'hbb6782ec),
	.w4(32'hbc0c3fc8),
	.w5(32'h3bbd9dcd),
	.w6(32'hbb9c47dc),
	.w7(32'hbbd06bed),
	.w8(32'h3b01973a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69fee),
	.w1(32'h3bea0cc2),
	.w2(32'h39d105c5),
	.w3(32'h3bc536fa),
	.w4(32'h3b8029ce),
	.w5(32'hbbbf8b8a),
	.w6(32'h3c064e1c),
	.w7(32'hbaca2e20),
	.w8(32'hbbc9196a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c62fd),
	.w1(32'hba2ad7e9),
	.w2(32'hbb465a1b),
	.w3(32'h39c5447c),
	.w4(32'h3b12180a),
	.w5(32'h3b2b0106),
	.w6(32'h3a87616e),
	.w7(32'h39e66d5f),
	.w8(32'hbb692ef5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f1b78),
	.w1(32'h3ae81e7b),
	.w2(32'hbc469a16),
	.w3(32'hbac43f08),
	.w4(32'h3ac819e2),
	.w5(32'hba8893ad),
	.w6(32'hba8758ba),
	.w7(32'h3a760865),
	.w8(32'h3a87d9d7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7934),
	.w1(32'h3b67d180),
	.w2(32'h3c74b235),
	.w3(32'h38438632),
	.w4(32'h3c3035ff),
	.w5(32'h3c5229d2),
	.w6(32'h3bbce268),
	.w7(32'h3c6fb6a5),
	.w8(32'h3c02a70a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb223d0),
	.w1(32'h3be9197e),
	.w2(32'h3bdba321),
	.w3(32'hbaa98e73),
	.w4(32'h3ae883f2),
	.w5(32'h3b715496),
	.w6(32'hbb3b23d6),
	.w7(32'hba47b535),
	.w8(32'h3b9261ca),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e75d2),
	.w1(32'h3b8d31a1),
	.w2(32'hb9ba09b1),
	.w3(32'h3bb470f8),
	.w4(32'h3bed2928),
	.w5(32'h3b834aac),
	.w6(32'h3b87201c),
	.w7(32'h3ba6170a),
	.w8(32'h3bbb6667),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e189),
	.w1(32'hbb8123c2),
	.w2(32'hba1e3ad5),
	.w3(32'hb98fa8ab),
	.w4(32'h3ab9f72c),
	.w5(32'hbab9cc75),
	.w6(32'h3bb02b4a),
	.w7(32'h3bcced86),
	.w8(32'hbb2579a2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe00f6f),
	.w1(32'hbaa45265),
	.w2(32'hbbd1a0b8),
	.w3(32'hbbd87181),
	.w4(32'h3b072460),
	.w5(32'hbbb94586),
	.w6(32'hbba6f0f8),
	.w7(32'hbb06bf1e),
	.w8(32'hbc1be55e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82c1c4),
	.w1(32'hbb8d3b3c),
	.w2(32'hbb8fa265),
	.w3(32'hb975fea4),
	.w4(32'hb9be3932),
	.w5(32'hb988f7cc),
	.w6(32'hbb84adf7),
	.w7(32'hba794224),
	.w8(32'hbb1ea8d4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a801bbe),
	.w1(32'h398f53e6),
	.w2(32'hbab4e651),
	.w3(32'h3b050ca5),
	.w4(32'hba430809),
	.w5(32'h3b1e29a7),
	.w6(32'hb94ca39f),
	.w7(32'hbb5b35a6),
	.w8(32'h3b26e803),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14630e),
	.w1(32'h3ac6358e),
	.w2(32'hba88814c),
	.w3(32'h3adafab6),
	.w4(32'h39cd80f6),
	.w5(32'hbb6351a6),
	.w6(32'h3b0b06ac),
	.w7(32'h3984f11e),
	.w8(32'hbb1f17db),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acebae2),
	.w1(32'hbb247ea5),
	.w2(32'hbbad6e3c),
	.w3(32'hbb5f9b2a),
	.w4(32'hbbc36ee5),
	.w5(32'hbbac8840),
	.w6(32'hbae1ac0a),
	.w7(32'hbb7fa660),
	.w8(32'hbbe723a6),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86e43b),
	.w1(32'hbbd5a626),
	.w2(32'hba8892c9),
	.w3(32'hbbd69d4f),
	.w4(32'hbafe5bf9),
	.w5(32'h3b142938),
	.w6(32'hbbcb40cb),
	.w7(32'hba96bd47),
	.w8(32'h389cd2d9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3270),
	.w1(32'hbb17aeed),
	.w2(32'hbae558b0),
	.w3(32'hba9f3f94),
	.w4(32'hbb2d2dfe),
	.w5(32'h398136f4),
	.w6(32'h38bf45b7),
	.w7(32'hbb50529d),
	.w8(32'h3aace7ed),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf395e),
	.w1(32'hba7e1263),
	.w2(32'hb986a802),
	.w3(32'hba960c76),
	.w4(32'hbab0034c),
	.w5(32'hba99d492),
	.w6(32'hb9031ece),
	.w7(32'h38cfa026),
	.w8(32'hbb30e24a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14362c),
	.w1(32'hb96b875d),
	.w2(32'h3aa63381),
	.w3(32'hbb87fad3),
	.w4(32'h3b29eeab),
	.w5(32'hbb804f9e),
	.w6(32'hbb95a4c4),
	.w7(32'h3b5fa654),
	.w8(32'hb9ead13e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18bc45),
	.w1(32'hbb595586),
	.w2(32'hbb417daf),
	.w3(32'hbb266191),
	.w4(32'hbac63877),
	.w5(32'h39ffacae),
	.w6(32'hbadeb44e),
	.w7(32'hbb7a3621),
	.w8(32'hbb9e8a30),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb802419),
	.w1(32'hbb27dc35),
	.w2(32'hbb2f2b3a),
	.w3(32'h38c7e6b9),
	.w4(32'hbaa56ba4),
	.w5(32'hba8346be),
	.w6(32'hbb1f15a9),
	.w7(32'hbb4a5742),
	.w8(32'h3a3a0341),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acac520),
	.w1(32'h39ddcbce),
	.w2(32'h38abc0e5),
	.w3(32'hbb3a846c),
	.w4(32'hbb7c5877),
	.w5(32'hb97c904e),
	.w6(32'hbb6202b1),
	.w7(32'hbb5a4601),
	.w8(32'hbabfd65d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189027),
	.w1(32'hbb673434),
	.w2(32'hbb4ede49),
	.w3(32'hbaf124f4),
	.w4(32'hbb07aa1a),
	.w5(32'h3b04e4e4),
	.w6(32'hbaf869f1),
	.w7(32'hbaba1ce5),
	.w8(32'h3b159aff),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfda520),
	.w1(32'h3c43ad10),
	.w2(32'h3c221f8f),
	.w3(32'h3b60177d),
	.w4(32'h3b2b5b34),
	.w5(32'hb942c8f6),
	.w6(32'h36dd2e06),
	.w7(32'hb981bc62),
	.w8(32'hbb039012),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736d0e),
	.w1(32'hbb8dfea1),
	.w2(32'hbaaa253a),
	.w3(32'hbacc59e9),
	.w4(32'h3a4c5180),
	.w5(32'hbb1cb72e),
	.w6(32'hbb745975),
	.w7(32'hbaa06243),
	.w8(32'hbad38d4e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd604b3),
	.w1(32'hbc420218),
	.w2(32'hbbf258c7),
	.w3(32'hbbddb406),
	.w4(32'hbb067878),
	.w5(32'h3affd004),
	.w6(32'hbba0a95e),
	.w7(32'hbad0a41e),
	.w8(32'h3ba8a2c3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43a33f),
	.w1(32'h3af4fdc9),
	.w2(32'h3ab71a12),
	.w3(32'hba7062e7),
	.w4(32'h3a1a250f),
	.w5(32'hb8fe44c1),
	.w6(32'h3b0a7726),
	.w7(32'h3a04822c),
	.w8(32'hba31755c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6d979),
	.w1(32'hba82eba9),
	.w2(32'hbb56b5d2),
	.w3(32'h3ab08d26),
	.w4(32'h3a22cedf),
	.w5(32'h38f2af8c),
	.w6(32'hbb26facb),
	.w7(32'hb8d6fd5e),
	.w8(32'hbb274c86),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3208),
	.w1(32'h3b83eb20),
	.w2(32'h3bad053d),
	.w3(32'h3b0b6ae6),
	.w4(32'h3b8d89ff),
	.w5(32'h3bc60ff5),
	.w6(32'h3a9060ab),
	.w7(32'hba4307c7),
	.w8(32'h3ba37931),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f4106),
	.w1(32'h3a9ad966),
	.w2(32'h3a7d4053),
	.w3(32'h3a885870),
	.w4(32'hba9c51cc),
	.w5(32'h3a8b6add),
	.w6(32'h3a83c8be),
	.w7(32'h3acaa90b),
	.w8(32'h3a8788e8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd0ae),
	.w1(32'h3b12e062),
	.w2(32'hbadca3c5),
	.w3(32'h3aee1fae),
	.w4(32'h3b2b8746),
	.w5(32'hba341457),
	.w6(32'h3a4ad610),
	.w7(32'hbaa84b42),
	.w8(32'h3a12c6fb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9d5a),
	.w1(32'h3b297bfe),
	.w2(32'h3a8eb06d),
	.w3(32'hb9b029fe),
	.w4(32'h3a2ae262),
	.w5(32'hbaa64a30),
	.w6(32'h3a09a6ff),
	.w7(32'hb7af828a),
	.w8(32'hbae1cf52),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56b4e1),
	.w1(32'hbad1a735),
	.w2(32'hb9ec6d07),
	.w3(32'hba8c9b52),
	.w4(32'hb99b5165),
	.w5(32'h39410537),
	.w6(32'hba3bb69b),
	.w7(32'hba9e8341),
	.w8(32'hb95024d2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0991a8),
	.w1(32'hbb20eeed),
	.w2(32'hbb4d8de1),
	.w3(32'h3b1a39f2),
	.w4(32'h3ae4cf61),
	.w5(32'hbc0f8f08),
	.w6(32'h3b15d278),
	.w7(32'h399a2ff7),
	.w8(32'hbc14b4f2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8c9ec),
	.w1(32'hbbc882fa),
	.w2(32'hbb3576ef),
	.w3(32'hbbaa94c5),
	.w4(32'hbb2c5984),
	.w5(32'hbb46ec6a),
	.w6(32'hbc01d3d9),
	.w7(32'hbb9d48c8),
	.w8(32'hbb5cb5dd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b2a7a),
	.w1(32'h3b672b08),
	.w2(32'h3aecd51b),
	.w3(32'h3b4d82e3),
	.w4(32'h3b7d7dd3),
	.w5(32'h3a1ee291),
	.w6(32'h3a8aa6dc),
	.w7(32'h3a7eae92),
	.w8(32'h3ac8cbe3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed9e0),
	.w1(32'h3be026a8),
	.w2(32'h3c116d99),
	.w3(32'h3b38acf9),
	.w4(32'h3b39c87a),
	.w5(32'hb98a7c26),
	.w6(32'h37a10025),
	.w7(32'h399763c3),
	.w8(32'h3987b8b2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54ecea),
	.w1(32'h3a1ece4b),
	.w2(32'hba295346),
	.w3(32'h39d6cfbb),
	.w4(32'h39ea89a1),
	.w5(32'hbaa9c415),
	.w6(32'h3b680658),
	.w7(32'h3b2ef92b),
	.w8(32'hbbe32c2c),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c113806),
	.w1(32'h3bdffd04),
	.w2(32'h3c8477ba),
	.w3(32'hbaa03be3),
	.w4(32'h3bd92cfa),
	.w5(32'hbb84856e),
	.w6(32'hbbf4f45b),
	.w7(32'h393ad130),
	.w8(32'hbb43ab85),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f6daa),
	.w1(32'hbb93065c),
	.w2(32'hbafaa3e6),
	.w3(32'hbb95af3d),
	.w4(32'hbb05d74a),
	.w5(32'hbafbdb4a),
	.w6(32'hbb3cb7be),
	.w7(32'hba80b891),
	.w8(32'hbad72cee),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a095b8a),
	.w1(32'hbb46d557),
	.w2(32'hbbc7e514),
	.w3(32'hb9191668),
	.w4(32'hbb0504d5),
	.w5(32'hbbf76aab),
	.w6(32'hbaec2098),
	.w7(32'hbb9fd7e7),
	.w8(32'hbc274a4d),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b354b),
	.w1(32'hbb8b2427),
	.w2(32'hba156125),
	.w3(32'hbb7e4226),
	.w4(32'h37d6076f),
	.w5(32'hbabb23ee),
	.w6(32'hbb8ba1af),
	.w7(32'hbac22349),
	.w8(32'hbb0542e4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24e114),
	.w1(32'hbbb430c6),
	.w2(32'hbb8b2646),
	.w3(32'hbb3637cb),
	.w4(32'hbaa910d4),
	.w5(32'hbb29dfd4),
	.w6(32'hbb944339),
	.w7(32'hbb053120),
	.w8(32'hbb1c8bec),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06ba0f),
	.w1(32'hbae3a4e2),
	.w2(32'hbb6bfb33),
	.w3(32'hba805fd2),
	.w4(32'hbabd9d9e),
	.w5(32'hbb6484ac),
	.w6(32'hba84c76f),
	.w7(32'hbad67e41),
	.w8(32'hbb455229),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad88d37),
	.w1(32'h3a13f6ae),
	.w2(32'h3ab557c5),
	.w3(32'hbb1d70d1),
	.w4(32'h3a1c9dfc),
	.w5(32'hbabf11bf),
	.w6(32'h39c1c25a),
	.w7(32'h3b8802db),
	.w8(32'h38d60279),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07e49e),
	.w1(32'h39c1e554),
	.w2(32'hba6272e8),
	.w3(32'h3af1fc99),
	.w4(32'h3b73b144),
	.w5(32'hbaca8441),
	.w6(32'h39dba66a),
	.w7(32'hbb259341),
	.w8(32'hbbab5e9d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26cc4),
	.w1(32'hbb3e9b3e),
	.w2(32'hba8674e9),
	.w3(32'h38ff6621),
	.w4(32'h3ac82d53),
	.w5(32'hbb368cc8),
	.w6(32'hbafb3197),
	.w7(32'hbb037619),
	.w8(32'hbb7e56cf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a388d),
	.w1(32'hbab468db),
	.w2(32'h3b8f88cd),
	.w3(32'hb53e3fe0),
	.w4(32'h3b6415aa),
	.w5(32'h3bbc9259),
	.w6(32'hbb2f0f06),
	.w7(32'h3ac0240d),
	.w8(32'h3bba7f1f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0024d),
	.w1(32'hb9716ed3),
	.w2(32'hbb06d917),
	.w3(32'h3ae53aa5),
	.w4(32'h3ab379b1),
	.w5(32'h3902c331),
	.w6(32'h3b36419f),
	.w7(32'h3a9afa71),
	.w8(32'h39faa42a),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47247e),
	.w1(32'h3b2cc983),
	.w2(32'h3bc4b8ab),
	.w3(32'hb8151751),
	.w4(32'h3b1c89ae),
	.w5(32'hbb71760a),
	.w6(32'h388785e5),
	.w7(32'h3ad6bf08),
	.w8(32'hbb299f2a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba816c0e),
	.w1(32'hbae1ed2f),
	.w2(32'hba94d35b),
	.w3(32'hbb06bfa3),
	.w4(32'hbae29b3a),
	.w5(32'hbb1e8399),
	.w6(32'hbabcbe86),
	.w7(32'hbb0831e3),
	.w8(32'hbb25da5a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d0edc),
	.w1(32'hbaebd057),
	.w2(32'hbb63604f),
	.w3(32'hbacf1b3c),
	.w4(32'hbb59bf01),
	.w5(32'hbb0d035f),
	.w6(32'hba3d14ce),
	.w7(32'hba04d65d),
	.w8(32'h3a44b5f8),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd10fe3),
	.w1(32'h3c001a86),
	.w2(32'h3bc36eea),
	.w3(32'hbaa057ec),
	.w4(32'h3b0737d7),
	.w5(32'h3b0d800c),
	.w6(32'h3b60ee9f),
	.w7(32'h3bd3c19e),
	.w8(32'h38a9bb11),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7967e),
	.w1(32'hbb100f75),
	.w2(32'hbae7c501),
	.w3(32'hb9cf7375),
	.w4(32'hbb1212d2),
	.w5(32'h38175d29),
	.w6(32'hbaa2a3d0),
	.w7(32'hbb32a56e),
	.w8(32'hb9458d7d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b741425),
	.w1(32'h3b0c803e),
	.w2(32'h3b91a959),
	.w3(32'h3a0c761e),
	.w4(32'h39aca254),
	.w5(32'h3b48be36),
	.w6(32'hb895183b),
	.w7(32'h3aa85a29),
	.w8(32'h3b050792),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f2ad4),
	.w1(32'hbb3eb40c),
	.w2(32'hbb7a766f),
	.w3(32'h3b7bd588),
	.w4(32'h3ade0bc6),
	.w5(32'hbb371cf1),
	.w6(32'h3b4b14fc),
	.w7(32'h39ab37d7),
	.w8(32'hba9b80e0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b6794),
	.w1(32'h3a0bd597),
	.w2(32'h3a944b99),
	.w3(32'h3a3b2dc5),
	.w4(32'h399fc3b6),
	.w5(32'h3a96587c),
	.w6(32'h3a17a7d1),
	.w7(32'hba1d21bd),
	.w8(32'h3ad69f79),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e280a),
	.w1(32'h3b74d51d),
	.w2(32'h3a174b3d),
	.w3(32'h3b2ef355),
	.w4(32'h3a87a893),
	.w5(32'hbc1c8565),
	.w6(32'hb905811f),
	.w7(32'h390a7c6b),
	.w8(32'hbbf2048c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2f4dc),
	.w1(32'hba8b38a0),
	.w2(32'h3b07d521),
	.w3(32'hbbae8fcc),
	.w4(32'hbbd0314a),
	.w5(32'hb9be97ce),
	.w6(32'hbb9ea06b),
	.w7(32'hbbce9da2),
	.w8(32'hba327078),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a923dc5),
	.w1(32'h3a5791fe),
	.w2(32'h3ae531cd),
	.w3(32'hb9d6041d),
	.w4(32'h39b5480f),
	.w5(32'hb99f20f9),
	.w6(32'h3b24dcad),
	.w7(32'h3ad3d391),
	.w8(32'h38f91926),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e790b),
	.w1(32'hba0465ec),
	.w2(32'h3a2ebdab),
	.w3(32'hbaaf73c1),
	.w4(32'h39ee552c),
	.w5(32'hbb5aa8b5),
	.w6(32'h39c475dc),
	.w7(32'h3ad199ea),
	.w8(32'hbbb86057),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7a6d9),
	.w1(32'hbc179deb),
	.w2(32'hbb5f97a0),
	.w3(32'hbc0eecda),
	.w4(32'hbb84fefe),
	.w5(32'hbacc7e7c),
	.w6(32'hbc267a6c),
	.w7(32'hbb941f63),
	.w8(32'h3a24bc2a),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf9e62),
	.w1(32'h3b7ea7f2),
	.w2(32'h3addb5cc),
	.w3(32'h39cdf3f1),
	.w4(32'h3afa61ec),
	.w5(32'h3b5b86fd),
	.w6(32'h3b1bf49e),
	.w7(32'h3b4d8012),
	.w8(32'h3b100d1b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8e27),
	.w1(32'hb8448af2),
	.w2(32'h3aa4ac88),
	.w3(32'hba7f9966),
	.w4(32'h39af2eb5),
	.w5(32'h3c015c43),
	.w6(32'hbb4d2a8f),
	.w7(32'hb9be5365),
	.w8(32'h3a16e26b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884838),
	.w1(32'h38bd21d8),
	.w2(32'hbad9708f),
	.w3(32'h3bb55b00),
	.w4(32'h3b4990bc),
	.w5(32'h3b14267a),
	.w6(32'hbaa8214a),
	.w7(32'hbafb18b3),
	.w8(32'hba34f40d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66e021),
	.w1(32'h3ab2d852),
	.w2(32'h3aa271a1),
	.w3(32'h3bbc4201),
	.w4(32'h3b1d9b39),
	.w5(32'hba878804),
	.w6(32'h3ad5e60f),
	.w7(32'hbadc9174),
	.w8(32'h3a5c4050),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e63f),
	.w1(32'h394c9d34),
	.w2(32'hbb89c242),
	.w3(32'hb9ad9e2c),
	.w4(32'hbad8c6a5),
	.w5(32'hbb59f3c3),
	.w6(32'h3b4159af),
	.w7(32'h3b6b75d5),
	.w8(32'hbbbdd8c8),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700390),
	.w1(32'hbbaa5c57),
	.w2(32'hbbe636d6),
	.w3(32'hba9b9c74),
	.w4(32'hbb84808c),
	.w5(32'hb9ca4bba),
	.w6(32'hbb245643),
	.w7(32'hbb5a8afa),
	.w8(32'h3b21e2f7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45ae17),
	.w1(32'h39ae1e56),
	.w2(32'h3a7f5b2d),
	.w3(32'hb8f1b27c),
	.w4(32'h39ac81f3),
	.w5(32'hba8fdccb),
	.w6(32'h3b0d1d64),
	.w7(32'h3b4a4259),
	.w8(32'hb98972d4),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef8e37),
	.w1(32'h3aaf2b7a),
	.w2(32'h3b042c5d),
	.w3(32'hbab5f201),
	.w4(32'hbb2da64e),
	.w5(32'h3a820909),
	.w6(32'hbb40d69e),
	.w7(32'hba99fa62),
	.w8(32'h3b8da475),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e9413),
	.w1(32'h3bcb5b1e),
	.w2(32'h3b786a42),
	.w3(32'h3b4a964b),
	.w4(32'h3b3cf7ed),
	.w5(32'hbbd8a0b0),
	.w6(32'h3b85575b),
	.w7(32'h3aac782f),
	.w8(32'hbb9e7a87),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d46d3),
	.w1(32'hbacb47c6),
	.w2(32'h3b8ba1ce),
	.w3(32'hbc0b020c),
	.w4(32'hbb456d54),
	.w5(32'hba277907),
	.w6(32'hbba98691),
	.w7(32'hba2368c8),
	.w8(32'h3b189309),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0adfe9),
	.w1(32'h3b268292),
	.w2(32'h3b490a33),
	.w3(32'h3a470e33),
	.w4(32'hba8d321a),
	.w5(32'hba1f0bba),
	.w6(32'h3b626fed),
	.w7(32'h3b292fef),
	.w8(32'h3aa03c76),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0035e6),
	.w1(32'hbc1d94a4),
	.w2(32'hbb2ab807),
	.w3(32'hbb404f12),
	.w4(32'h3a8333f4),
	.w5(32'hbadb24ad),
	.w6(32'h3accbca3),
	.w7(32'h3bb3a526),
	.w8(32'hb9519f4e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71d6e8),
	.w1(32'h38fc1667),
	.w2(32'hbbe33be5),
	.w3(32'h3a125ed7),
	.w4(32'h397007bc),
	.w5(32'hbba01050),
	.w6(32'hbb1fb8a9),
	.w7(32'hbb7db4ba),
	.w8(32'hbbc136d6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1e511),
	.w1(32'hbae3979e),
	.w2(32'h38b5f846),
	.w3(32'hbb4e63cc),
	.w4(32'hba8c8800),
	.w5(32'hbaf3b329),
	.w6(32'hbae3c963),
	.w7(32'hbab2d5c0),
	.w8(32'hba812745),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd855b5),
	.w1(32'h3c200ed1),
	.w2(32'h3c60b953),
	.w3(32'hbb3a1df4),
	.w4(32'hba8d2bee),
	.w5(32'h3b31086c),
	.w6(32'hbb9c0655),
	.w7(32'h3b17d411),
	.w8(32'h3a99a5d3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78c50f),
	.w1(32'h3b91d5c6),
	.w2(32'h3b1075d1),
	.w3(32'h3b7d4053),
	.w4(32'h3b822297),
	.w5(32'h3aa1de9e),
	.w6(32'h3ab86ca9),
	.w7(32'h398dd790),
	.w8(32'h3b9c2a6a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e6e627),
	.w1(32'hbb806ff4),
	.w2(32'hbb09052a),
	.w3(32'hb98b47ea),
	.w4(32'hbb41e1d0),
	.w5(32'h3a16360e),
	.w6(32'h3ac7664c),
	.w7(32'hbb126dea),
	.w8(32'h3a141e62),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a0ad2),
	.w1(32'hbb30d21b),
	.w2(32'hbb697179),
	.w3(32'h3b7aabcd),
	.w4(32'h3af95e8f),
	.w5(32'hbb3b1950),
	.w6(32'h3b804eab),
	.w7(32'h38f3bfbf),
	.w8(32'hbb5739ac),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2687ae),
	.w1(32'hbbbea9e1),
	.w2(32'hbc0c7aeb),
	.w3(32'hbb345998),
	.w4(32'hbb94e5e9),
	.w5(32'h3a237285),
	.w6(32'hbb32644a),
	.w7(32'hbbba0f53),
	.w8(32'hba8575d7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f1b4),
	.w1(32'h3b5af987),
	.w2(32'h3b83b3cf),
	.w3(32'h3b2b6d02),
	.w4(32'h3b6d8964),
	.w5(32'h3a1ec796),
	.w6(32'h3b098c71),
	.w7(32'h3b716e04),
	.w8(32'hbaaf2e8a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7008d8),
	.w1(32'hbb48ce51),
	.w2(32'hbb84641b),
	.w3(32'h3ae45ebb),
	.w4(32'hba33abcc),
	.w5(32'h3972b783),
	.w6(32'hba17b02a),
	.w7(32'hba79d18f),
	.w8(32'h3aa5464b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae83aac),
	.w1(32'hbb5c0e10),
	.w2(32'h3a842a7e),
	.w3(32'hbadb7f5e),
	.w4(32'h3aee9fcd),
	.w5(32'hbabd6b06),
	.w6(32'hb9588597),
	.w7(32'h3b2b4821),
	.w8(32'hbb876236),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2fa5f),
	.w1(32'hba3442de),
	.w2(32'hba817a46),
	.w3(32'hb86e88e9),
	.w4(32'h3a5c34dc),
	.w5(32'hb9f70c76),
	.w6(32'hbb81a41e),
	.w7(32'hbb178f79),
	.w8(32'hbb28c688),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830ffb),
	.w1(32'h3bf1deb8),
	.w2(32'h3bcf2fae),
	.w3(32'h3af12a8a),
	.w4(32'h3a27bca2),
	.w5(32'hba717ff3),
	.w6(32'h386d1bfa),
	.w7(32'hb9aed1e7),
	.w8(32'hb90df866),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a619),
	.w1(32'hbb8bd40f),
	.w2(32'hbbb9e63f),
	.w3(32'hbabe894b),
	.w4(32'h392b2de6),
	.w5(32'hbb7c45f9),
	.w6(32'hbab1cfa2),
	.w7(32'hbb0db85c),
	.w8(32'hbb672513),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77c1d6),
	.w1(32'hbb7979e8),
	.w2(32'hbaf5a527),
	.w3(32'hbad0f37c),
	.w4(32'h3b2b8844),
	.w5(32'hbb197d9d),
	.w6(32'hbbb16d38),
	.w7(32'hba33959a),
	.w8(32'hbb661e10),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb359cd3),
	.w1(32'hbabc5e2d),
	.w2(32'hba284bb0),
	.w3(32'h39af0e5d),
	.w4(32'hbaabe727),
	.w5(32'hbaa0cb78),
	.w6(32'hba225015),
	.w7(32'hba7b99c4),
	.w8(32'h3a0b89a4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3612a6),
	.w1(32'h3b3189a0),
	.w2(32'h3b0c4acb),
	.w3(32'hba97ef5c),
	.w4(32'hb987c1e3),
	.w5(32'hbad6b685),
	.w6(32'hbafa443a),
	.w7(32'hbadf3201),
	.w8(32'hbb26f3b6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bc27e),
	.w1(32'hbac569c3),
	.w2(32'hbb7a3d09),
	.w3(32'h38ab832c),
	.w4(32'h3aea4a40),
	.w5(32'hba2cd92d),
	.w6(32'hbab69465),
	.w7(32'hba9c41a7),
	.w8(32'hbaff49b8),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba689757),
	.w1(32'h3b7ba474),
	.w2(32'h39aede28),
	.w3(32'h3aaabc55),
	.w4(32'h3b91b68a),
	.w5(32'hbaa1cd4e),
	.w6(32'hba33c6de),
	.w7(32'h3b475e31),
	.w8(32'hbb1eb98a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c31be),
	.w1(32'hbb9e0001),
	.w2(32'h355d6835),
	.w3(32'hbbc12945),
	.w4(32'hbb2a22d2),
	.w5(32'h3b99796d),
	.w6(32'hbb8edbec),
	.w7(32'hba92292e),
	.w8(32'h3bd4503c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab775b),
	.w1(32'hbb77b617),
	.w2(32'hbbf9ea5b),
	.w3(32'h3b4b5dab),
	.w4(32'hb9f30816),
	.w5(32'hbc231889),
	.w6(32'h3c2da3fe),
	.w7(32'hbaac0ac8),
	.w8(32'hbc2584e7),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a7a82),
	.w1(32'hbb0296af),
	.w2(32'h3b19e447),
	.w3(32'h3b5bfdfc),
	.w4(32'h3b463d93),
	.w5(32'h3b380256),
	.w6(32'h3b501492),
	.w7(32'h3ae73795),
	.w8(32'h3aee2ad0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d94d2),
	.w1(32'h399d2997),
	.w2(32'hbb028688),
	.w3(32'hb6f87754),
	.w4(32'hba5cec8a),
	.w5(32'h3a3ee3a1),
	.w6(32'h3b0f7aa9),
	.w7(32'hba4ab274),
	.w8(32'h38fdb837),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24890),
	.w1(32'h3b4bab12),
	.w2(32'h3ba3eec6),
	.w3(32'h3b2de129),
	.w4(32'h3b9997d2),
	.w5(32'hbb4e6821),
	.w6(32'h3b187501),
	.w7(32'h3b3e6a02),
	.w8(32'hbb226e9e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fecbb),
	.w1(32'hbb06409c),
	.w2(32'hbb3692ff),
	.w3(32'hbaf8ea3a),
	.w4(32'hbb11cd70),
	.w5(32'h3acb8209),
	.w6(32'hbb442ce0),
	.w7(32'hbb214630),
	.w8(32'hba116eca),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36f86c),
	.w1(32'hb9903938),
	.w2(32'hba57b287),
	.w3(32'h3b248dba),
	.w4(32'h3b07e7b8),
	.w5(32'hbb0a060a),
	.w6(32'hb91f69b7),
	.w7(32'h3aba8136),
	.w8(32'hb9fe203f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd28a57),
	.w1(32'h3ba8874a),
	.w2(32'h3b377f47),
	.w3(32'h3b162c22),
	.w4(32'h3b5f93c4),
	.w5(32'hba7268d5),
	.w6(32'h3b89774e),
	.w7(32'h3acb5693),
	.w8(32'hbb129df8),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa933b),
	.w1(32'h397e76cd),
	.w2(32'h3a17bfe5),
	.w3(32'h3b130ed9),
	.w4(32'h3b455dd6),
	.w5(32'h37a2a53b),
	.w6(32'h3b01aea4),
	.w7(32'h3ac698db),
	.w8(32'h392ab284),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16c83e),
	.w1(32'hb9e7298e),
	.w2(32'h39643940),
	.w3(32'hbb12e7ff),
	.w4(32'h3ab41047),
	.w5(32'h3af208b9),
	.w6(32'hbb31bfd5),
	.w7(32'hb9b09ba6),
	.w8(32'h3a9d36b6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa31e27),
	.w1(32'hba3e0ccc),
	.w2(32'hb9917469),
	.w3(32'hb9884752),
	.w4(32'hba0cc4bc),
	.w5(32'hb9c05d34),
	.w6(32'hbb1b8ee0),
	.w7(32'h3aea4777),
	.w8(32'hb9f6a27c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0b11),
	.w1(32'hba8be0c2),
	.w2(32'hbb5a9a7d),
	.w3(32'hb91d6337),
	.w4(32'hbb61d77f),
	.w5(32'hbb42be79),
	.w6(32'h3b0d068e),
	.w7(32'hbb2fa209),
	.w8(32'h3a0e865a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70aca4),
	.w1(32'h3bbe51f4),
	.w2(32'h3bd39083),
	.w3(32'hbaabf69a),
	.w4(32'h3b04bd39),
	.w5(32'hba53ae95),
	.w6(32'h3b3b8acc),
	.w7(32'h3bf71181),
	.w8(32'hba4bbc71),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7d29c),
	.w1(32'hba140727),
	.w2(32'hba8fccd0),
	.w3(32'h3999a0c4),
	.w4(32'hbaca7037),
	.w5(32'hbb282cd7),
	.w6(32'hb9a0b440),
	.w7(32'hbb48becf),
	.w8(32'hba01710d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd03656),
	.w1(32'h3c08740a),
	.w2(32'h3be229f9),
	.w3(32'hbac4be44),
	.w4(32'hbaccfae3),
	.w5(32'hbb7b833d),
	.w6(32'h3a11da8e),
	.w7(32'h3a8f7e03),
	.w8(32'hbb938860),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba88a2d),
	.w1(32'hbb989e9b),
	.w2(32'hbb4bc67a),
	.w3(32'hba1d1860),
	.w4(32'hbacffcca),
	.w5(32'hbaec875e),
	.w6(32'hbb7fda01),
	.w7(32'hbb4000a3),
	.w8(32'hb9b80887),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92113e9),
	.w1(32'hbad17daf),
	.w2(32'h3aa9c2ea),
	.w3(32'hbafc9d5c),
	.w4(32'h3ab7ec52),
	.w5(32'hba35d3a8),
	.w6(32'hbada1add),
	.w7(32'h3a8947d9),
	.w8(32'hbb52fe63),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7026219),
	.w1(32'h3a9a10a8),
	.w2(32'h3ac81576),
	.w3(32'h3b24214e),
	.w4(32'h3b334650),
	.w5(32'h3b1222f6),
	.w6(32'hb834ef10),
	.w7(32'h3af461b2),
	.w8(32'h3b1a5635),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952939f),
	.w1(32'hb9b337e3),
	.w2(32'hb9f2e3f5),
	.w3(32'hbab348ac),
	.w4(32'h3aaa1613),
	.w5(32'h39a3a6db),
	.w6(32'hba2d7396),
	.w7(32'hb9ce402b),
	.w8(32'h39b6921a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6368ee),
	.w1(32'h3a8c6a8d),
	.w2(32'h3aeaffeb),
	.w3(32'hb983461e),
	.w4(32'hb9829f5d),
	.w5(32'hb97688f3),
	.w6(32'h3950ff27),
	.w7(32'h38386d4a),
	.w8(32'hbb339182),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb708e7),
	.w1(32'hbbcd8ef1),
	.w2(32'hbb6f1a82),
	.w3(32'hbac5c9f8),
	.w4(32'hba4cde5c),
	.w5(32'h3a7738ee),
	.w6(32'hb965aed9),
	.w7(32'hb99bf126),
	.w8(32'h39770023),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04cc9),
	.w1(32'hbb85aa6c),
	.w2(32'hbb848e86),
	.w3(32'hbaebf941),
	.w4(32'hbb055b9d),
	.w5(32'h3ae1013f),
	.w6(32'hbb0b1c1c),
	.w7(32'hbb6ca4a0),
	.w8(32'hbb9222cc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2920),
	.w1(32'hbc0111ef),
	.w2(32'hbbc4227f),
	.w3(32'hb94bb987),
	.w4(32'h3a29bf1d),
	.w5(32'hbb2da6c5),
	.w6(32'hbbd579e5),
	.w7(32'hbb984b1c),
	.w8(32'hbbbef232),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba52a93),
	.w1(32'hbb2dccec),
	.w2(32'hbb0ec51f),
	.w3(32'hbaf6598e),
	.w4(32'hbb3a9b97),
	.w5(32'h3aad34f1),
	.w6(32'hbb7877ed),
	.w7(32'hbad3fbba),
	.w8(32'h3a035763),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d5f61),
	.w1(32'h3a2a60eb),
	.w2(32'hb9b4a312),
	.w3(32'h3a50a14b),
	.w4(32'hba40fba9),
	.w5(32'hbb6b1f08),
	.w6(32'hba900d71),
	.w7(32'hba8a463a),
	.w8(32'h3b43b1ad),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c126a1c),
	.w1(32'h3b99b449),
	.w2(32'h3a9d0739),
	.w3(32'hba880ed7),
	.w4(32'hbb6d9972),
	.w5(32'hbadd9ec4),
	.w6(32'h3bba72d9),
	.w7(32'h3b6ff303),
	.w8(32'hbab4e813),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13bc04),
	.w1(32'hb79ac058),
	.w2(32'hbb682ffa),
	.w3(32'h3ac62f59),
	.w4(32'hba4bbb22),
	.w5(32'h38919d18),
	.w6(32'hb9b43728),
	.w7(32'hbb214516),
	.w8(32'hbb28a526),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd3414),
	.w1(32'h3b76688b),
	.w2(32'h3ab91476),
	.w3(32'h3a861ef6),
	.w4(32'h3a674882),
	.w5(32'hbae5a4a6),
	.w6(32'h3b5c4a15),
	.w7(32'h39e0e22f),
	.w8(32'hb8816410),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9091aa),
	.w1(32'h3ba8a377),
	.w2(32'h3b112203),
	.w3(32'h3b206c69),
	.w4(32'h3baf80bd),
	.w5(32'hb9baf1c0),
	.w6(32'h3aeae3e5),
	.w7(32'hb82d16ce),
	.w8(32'hbaffb153),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51e40e),
	.w1(32'h3b3e529a),
	.w2(32'h3b7c9e9a),
	.w3(32'h3a4ba5e3),
	.w4(32'h3a8dbe25),
	.w5(32'hbb8f36e9),
	.w6(32'h3a033cec),
	.w7(32'hb8fcb686),
	.w8(32'hbb9a376e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7cff7),
	.w1(32'hbbe93c5f),
	.w2(32'hbba20cea),
	.w3(32'hbbb3f549),
	.w4(32'hbb62202f),
	.w5(32'h3b46f88b),
	.w6(32'hbb8f773a),
	.w7(32'hbb4471c0),
	.w8(32'h3a450ff9),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b798794),
	.w1(32'h3bf7ac74),
	.w2(32'hbb2077cc),
	.w3(32'h3af7a53a),
	.w4(32'h3bb9081d),
	.w5(32'hbb747e2d),
	.w6(32'hb8b295be),
	.w7(32'h3bcebbfa),
	.w8(32'hbb870bc4),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91220e),
	.w1(32'hb9e8ea10),
	.w2(32'hbba819e0),
	.w3(32'hba641b78),
	.w4(32'hbb9c4e1d),
	.w5(32'hbba6ea3a),
	.w6(32'hba9779f6),
	.w7(32'hbbab6285),
	.w8(32'hbc018c46),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae56a9a),
	.w1(32'h3ab868b2),
	.w2(32'hbb81da25),
	.w3(32'h3b2c5128),
	.w4(32'h3a461ee6),
	.w5(32'hbb8737dc),
	.w6(32'hbaff114f),
	.w7(32'hbad89935),
	.w8(32'hbbfd073a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24047a),
	.w1(32'h3b435487),
	.w2(32'h3c170946),
	.w3(32'hba4c2ce7),
	.w4(32'h3ba2bca1),
	.w5(32'h3bca510a),
	.w6(32'hbb881513),
	.w7(32'h3b5253be),
	.w8(32'h3baf7de3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb437dea),
	.w1(32'hba518893),
	.w2(32'h3b512870),
	.w3(32'h3a4c9eda),
	.w4(32'h3b8ff3d1),
	.w5(32'h3af46569),
	.w6(32'hba742d39),
	.w7(32'h3ad2f482),
	.w8(32'h3b06ff2a),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a815e43),
	.w1(32'h3a9e7ad5),
	.w2(32'h3b8ad2fe),
	.w3(32'hbb3f2e0c),
	.w4(32'hb9b2dc8c),
	.w5(32'hba75d320),
	.w6(32'hbb05c988),
	.w7(32'h3ac371c4),
	.w8(32'h3a46ccb4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c013cb0),
	.w1(32'h3bb3a8fc),
	.w2(32'h3c2b0077),
	.w3(32'h3b836214),
	.w4(32'h3b877236),
	.w5(32'h3ba0e299),
	.w6(32'h3a86795d),
	.w7(32'h3b6cea19),
	.w8(32'h3bfcf7e3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934bb98),
	.w1(32'hba83211f),
	.w2(32'h3a1ee609),
	.w3(32'h3b7d9d9f),
	.w4(32'h3b3e12ec),
	.w5(32'h3ad3e5c5),
	.w6(32'h3c224bba),
	.w7(32'h3bf25ac2),
	.w8(32'h3b77588d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78a8da),
	.w1(32'h3ae08d28),
	.w2(32'h3abe038d),
	.w3(32'h3ae10034),
	.w4(32'h3b537222),
	.w5(32'hb917aba9),
	.w6(32'h3b4adb67),
	.w7(32'h3bce3591),
	.w8(32'h3b268411),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9328fb),
	.w1(32'h3b9e530e),
	.w2(32'h3bfa5776),
	.w3(32'h3b2cc243),
	.w4(32'h3baf9497),
	.w5(32'hba161cf0),
	.w6(32'h3c37c8ff),
	.w7(32'h3bf997d0),
	.w8(32'hbb4851a1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7bb19),
	.w1(32'hbc1e538d),
	.w2(32'hbaba22b5),
	.w3(32'hbc5f4d12),
	.w4(32'hbb0f4b08),
	.w5(32'h3b1b8fb8),
	.w6(32'hbbe7e1de),
	.w7(32'hba3741a1),
	.w8(32'hbb68a9a6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d46c8),
	.w1(32'hbad5646a),
	.w2(32'h3b8eee2e),
	.w3(32'h3bcb21a5),
	.w4(32'h3c034063),
	.w5(32'h3b98be0d),
	.w6(32'hbcaf5ba8),
	.w7(32'h3c212e25),
	.w8(32'h3b98e42d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28d848),
	.w1(32'hbc37c887),
	.w2(32'hbb609ebc),
	.w3(32'hbb6a8291),
	.w4(32'h3a2019c0),
	.w5(32'h3bbed126),
	.w6(32'hbc546759),
	.w7(32'h3ae7278d),
	.w8(32'h3a6100a2),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc347e),
	.w1(32'h3b8feec0),
	.w2(32'hb9b05c73),
	.w3(32'h3c0749dd),
	.w4(32'h3c0e5bb3),
	.w5(32'hbc8bf796),
	.w6(32'h3a494f6e),
	.w7(32'h3aa2ca97),
	.w8(32'hbcbb3d35),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8616ec),
	.w1(32'hbc07c909),
	.w2(32'hbc93c3dd),
	.w3(32'hbc872fce),
	.w4(32'hbc5af5ef),
	.w5(32'h3b046d9a),
	.w6(32'h3cfb7010),
	.w7(32'hbca1a47f),
	.w8(32'h3bfaa73e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5321fd),
	.w1(32'h3a37fa4a),
	.w2(32'h3c28da03),
	.w3(32'hbb8224f9),
	.w4(32'h3c4ec056),
	.w5(32'h3b464562),
	.w6(32'hbc94528e),
	.w7(32'h3c478770),
	.w8(32'h3b227f10),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2444),
	.w1(32'h39798dd1),
	.w2(32'h3b242e74),
	.w3(32'h3ae11b2c),
	.w4(32'h3b1bacfd),
	.w5(32'h3baf497e),
	.w6(32'hbb867a18),
	.w7(32'h3b99ada1),
	.w8(32'h3bbab658),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61d73),
	.w1(32'hbc5d3828),
	.w2(32'hbaf6b6d3),
	.w3(32'hbb4e9493),
	.w4(32'hbc29c8f4),
	.w5(32'h3b19aeee),
	.w6(32'hbc17b324),
	.w7(32'hbc10ec56),
	.w8(32'h3a56dfba),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb454e6),
	.w1(32'h3b16cb76),
	.w2(32'h3b65a5b3),
	.w3(32'h3a6c10a2),
	.w4(32'h3c347f42),
	.w5(32'hbbed327c),
	.w6(32'hbc90cdd0),
	.w7(32'hbc2f5b7c),
	.w8(32'h3a150948),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad596ff),
	.w1(32'h3becc110),
	.w2(32'h3c1d4208),
	.w3(32'h3b3481dc),
	.w4(32'h3b614f53),
	.w5(32'h3c85e6b3),
	.w6(32'h3ca7b103),
	.w7(32'h3c27d935),
	.w8(32'hbb53dcff),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c082f0e),
	.w1(32'hba375bd7),
	.w2(32'h3c4cc7a4),
	.w3(32'h3bf12e5f),
	.w4(32'h3c8c5704),
	.w5(32'h3c10a8f5),
	.w6(32'hbc6655e1),
	.w7(32'hb8e93a51),
	.w8(32'hbb922d0b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc680be8),
	.w1(32'hbb974694),
	.w2(32'h3c4368e4),
	.w3(32'hbc12570f),
	.w4(32'hbc52be7e),
	.w5(32'h3be0bce5),
	.w6(32'hbc8bc2ca),
	.w7(32'h39e89a8d),
	.w8(32'hbb4f535c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9c905),
	.w1(32'h3b9194b0),
	.w2(32'hbb260368),
	.w3(32'h3b731940),
	.w4(32'h3c10f920),
	.w5(32'h3a6aeea5),
	.w6(32'hb993cbf3),
	.w7(32'hbafedc10),
	.w8(32'hbb740080),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac6ffc),
	.w1(32'h3b771e2a),
	.w2(32'h3bbd48ab),
	.w3(32'h3b1b64f5),
	.w4(32'h3ba8b88a),
	.w5(32'hbb80bd39),
	.w6(32'hbbb2e6e1),
	.w7(32'h3c4e2b54),
	.w8(32'h3b4e9625),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe65e5c),
	.w1(32'hbc1bf43e),
	.w2(32'hbc07b7ce),
	.w3(32'hbc0a6825),
	.w4(32'hbbb458b2),
	.w5(32'hbc9193a1),
	.w6(32'hbbd68d04),
	.w7(32'hbb5b3709),
	.w8(32'hbc46c698),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e17fa),
	.w1(32'hbc49bea7),
	.w2(32'hbc0de8c5),
	.w3(32'h3addc10d),
	.w4(32'h3b4a9c16),
	.w5(32'hbace9205),
	.w6(32'hbc1008b5),
	.w7(32'hb74b9569),
	.w8(32'hbc3315d4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8574cf),
	.w1(32'hbbfdeb10),
	.w2(32'hbbc331be),
	.w3(32'hbad83a16),
	.w4(32'h3b7f7187),
	.w5(32'h3ca1ba29),
	.w6(32'hbc2c6abc),
	.w7(32'hbaf3d93b),
	.w8(32'h3c9fa880),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4294da),
	.w1(32'h3b300367),
	.w2(32'hba99b566),
	.w3(32'h3c863617),
	.w4(32'h3bda8e39),
	.w5(32'hbb17fcc5),
	.w6(32'h3bb6d081),
	.w7(32'hbbbf69e8),
	.w8(32'hbb7e1ba4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30e443),
	.w1(32'hbaf76b59),
	.w2(32'h3a0f19e8),
	.w3(32'hbba7980e),
	.w4(32'h3a9d528e),
	.w5(32'hbbf1e8d0),
	.w6(32'hbc0ee635),
	.w7(32'hbb038798),
	.w8(32'h392f52db),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08b94c),
	.w1(32'hbc01dc99),
	.w2(32'hbc2dbfcf),
	.w3(32'hbc0255f6),
	.w4(32'hbbf709df),
	.w5(32'hbc8024fb),
	.w6(32'h39a84b7a),
	.w7(32'hbb4f259f),
	.w8(32'hbbe49aee),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed925a),
	.w1(32'h3c1dae12),
	.w2(32'hb8b0d4d2),
	.w3(32'hbb8affe2),
	.w4(32'hbc30d2ee),
	.w5(32'h3c1fe07d),
	.w6(32'h3ce9e22c),
	.w7(32'h3b15e177),
	.w8(32'hbb6bce1a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab1c7),
	.w1(32'hbbd2d953),
	.w2(32'hbb061205),
	.w3(32'h3aadef48),
	.w4(32'h3b8d8dd5),
	.w5(32'hbb0c5e6f),
	.w6(32'h39cda784),
	.w7(32'hbb8dec15),
	.w8(32'hbbc2b581),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133650),
	.w1(32'hbb0ba4a3),
	.w2(32'hbbb03fc6),
	.w3(32'hbc145976),
	.w4(32'h3b417ccc),
	.w5(32'hbac22380),
	.w6(32'hbbead2c1),
	.w7(32'h399fca8c),
	.w8(32'hbb80f439),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c167797),
	.w1(32'hbbcc5df5),
	.w2(32'hbbb32c13),
	.w3(32'hbc844dcd),
	.w4(32'hbaed3d63),
	.w5(32'hbb64c446),
	.w6(32'hbc7ed9ff),
	.w7(32'hba5de23b),
	.w8(32'h3b1f0e50),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51f252),
	.w1(32'hba99393e),
	.w2(32'h3b72966b),
	.w3(32'hbabfe138),
	.w4(32'hbb2f36d6),
	.w5(32'hbb1fe996),
	.w6(32'hbc43e8e4),
	.w7(32'h3b28d429),
	.w8(32'hbc170960),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04ce69),
	.w1(32'hbc7cc570),
	.w2(32'hbb939fd8),
	.w3(32'hbaafa864),
	.w4(32'hbb3d33f9),
	.w5(32'hbb0693a0),
	.w6(32'hbd006be8),
	.w7(32'hbc01e564),
	.w8(32'hbbd2fbf6),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43ac43),
	.w1(32'hbbc45b3f),
	.w2(32'hbb07f057),
	.w3(32'hb87009e6),
	.w4(32'hb818756f),
	.w5(32'h3a4f4d7e),
	.w6(32'hbb4efe5f),
	.w7(32'hbb814f05),
	.w8(32'hbbdd4328),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c499f17),
	.w1(32'hbb52d5d3),
	.w2(32'h3c08f0b7),
	.w3(32'h3bfdb028),
	.w4(32'h3c8fe2cf),
	.w5(32'hbbbc0d6f),
	.w6(32'hbd092e8d),
	.w7(32'h3b3154cd),
	.w8(32'hbc1f1fe4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf324b7),
	.w1(32'hbb1bbc4d),
	.w2(32'hbb84b8d0),
	.w3(32'h3b12e67d),
	.w4(32'h3c07d2bf),
	.w5(32'h3c02088d),
	.w6(32'hbb2bffd0),
	.w7(32'h3ae025ed),
	.w8(32'hbc11b009),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule