module layer_8_featuremap_2(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2b16cf),
	.w1(32'h3b92f639),
	.w2(32'h3a4d2132),
	.w3(32'h3d71a4af),
	.w4(32'h3accf6dd),
	.w5(32'h3ac27b15),
	.w6(32'hbd12ee90),
	.w7(32'h3bd6f9c7),
	.w8(32'h3b0a5cd1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceeee4),
	.w1(32'h3b276eba),
	.w2(32'h3aa512ec),
	.w3(32'h37292ec8),
	.w4(32'h3a14ff20),
	.w5(32'h3bde795f),
	.w6(32'h398ad64f),
	.w7(32'h3b0b07d7),
	.w8(32'h3bf0419b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18fc1),
	.w1(32'hbb2ee372),
	.w2(32'hbb37c165),
	.w3(32'h3b80914e),
	.w4(32'h3a33430f),
	.w5(32'hbb1582dd),
	.w6(32'h3bd19819),
	.w7(32'h3b0db4ea),
	.w8(32'hbb02b6c9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd91ee),
	.w1(32'h3991b864),
	.w2(32'hbbbd9a14),
	.w3(32'hbb94a037),
	.w4(32'h3b4d2f4d),
	.w5(32'h3a7e6f0e),
	.w6(32'h3820e086),
	.w7(32'h3c04c6cd),
	.w8(32'h3bee2653),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb620ba2),
	.w1(32'h3b3785c8),
	.w2(32'hba174640),
	.w3(32'hbb28e797),
	.w4(32'h3b849fcc),
	.w5(32'h3b9b93f4),
	.w6(32'h3a2383ec),
	.w7(32'h3bc7b392),
	.w8(32'h39b8a4ed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ae4de),
	.w1(32'hbcde2e29),
	.w2(32'hbd0878c5),
	.w3(32'h3ab0fece),
	.w4(32'hbcbcfd44),
	.w5(32'h3c1cdf28),
	.w6(32'h3a96e20c),
	.w7(32'h3c83c47b),
	.w8(32'h3d2ebcee),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd09b8a9),
	.w1(32'h3bc25c05),
	.w2(32'h3b686560),
	.w3(32'h3d05409d),
	.w4(32'h3b0f9dc8),
	.w5(32'hbb7dd436),
	.w6(32'h3d315fe8),
	.w7(32'h3b023dc2),
	.w8(32'h3aba734d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a789d),
	.w1(32'hbaa09435),
	.w2(32'hba1220ab),
	.w3(32'hbbd47773),
	.w4(32'h3c88d140),
	.w5(32'h3c31aead),
	.w6(32'h3abecd31),
	.w7(32'h3bba2b89),
	.w8(32'h3c35df62),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefab3b),
	.w1(32'h3b5a6579),
	.w2(32'h3b67ce03),
	.w3(32'hbb54012b),
	.w4(32'h3aa3aabd),
	.w5(32'h3a8c351c),
	.w6(32'h3caf8aa4),
	.w7(32'hbb7f7fd6),
	.w8(32'hbc01b715),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17ba64),
	.w1(32'hbc5500af),
	.w2(32'hbcf36375),
	.w3(32'hbb13a91a),
	.w4(32'hbbaf8d25),
	.w5(32'h3d1ad72a),
	.w6(32'hbc272011),
	.w7(32'h3ca667d9),
	.w8(32'hbac863f6),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eff0f),
	.w1(32'hbb0cdd6c),
	.w2(32'hbaa70ec4),
	.w3(32'h3cf92660),
	.w4(32'h3a83e50c),
	.w5(32'h3ae54bf7),
	.w6(32'hbd001176),
	.w7(32'hbbd55c23),
	.w8(32'hbc3ae487),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89a36f1),
	.w1(32'h3bd717b0),
	.w2(32'h3c23d460),
	.w3(32'hbb05fc35),
	.w4(32'h3b232ad0),
	.w5(32'hbc07480f),
	.w6(32'hbbe8013d),
	.w7(32'h3bb7eecb),
	.w8(32'h3c71ac3d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8634f2),
	.w1(32'h3c25a80a),
	.w2(32'h3c008b7c),
	.w3(32'hbc8ba47f),
	.w4(32'hbbe4258a),
	.w5(32'hbd4d2703),
	.w6(32'h3c885256),
	.w7(32'h3b850972),
	.w8(32'h3cf035c5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31b170),
	.w1(32'hbaa5a27a),
	.w2(32'h3acdc4f4),
	.w3(32'hbd6c4b50),
	.w4(32'hbb717c54),
	.w5(32'h3be79887),
	.w6(32'h3d392e91),
	.w7(32'hbbbed96d),
	.w8(32'hbc6add2d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933845),
	.w1(32'hbb7d3fdc),
	.w2(32'hbbdd8e9b),
	.w3(32'h3c141956),
	.w4(32'hbb473499),
	.w5(32'hbbb360d2),
	.w6(32'hbc9d3019),
	.w7(32'h3bc86feb),
	.w8(32'h3c42b111),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac1c7),
	.w1(32'hbb223cb2),
	.w2(32'hbbab7136),
	.w3(32'hbb1dcf5c),
	.w4(32'hbc5bb34c),
	.w5(32'hbb08d080),
	.w6(32'h3c97f23b),
	.w7(32'h3b5c89c7),
	.w8(32'h3acc13e7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc6d2),
	.w1(32'h3b4e5de0),
	.w2(32'h3cbf25bf),
	.w3(32'h3ace90ef),
	.w4(32'hbca2037d),
	.w5(32'hbd2ef273),
	.w6(32'hbb2bc4c8),
	.w7(32'hbc8289cc),
	.w8(32'hba42338d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135a21),
	.w1(32'hbb71242b),
	.w2(32'hbb196241),
	.w3(32'hbd1b9029),
	.w4(32'hbb2ef9cd),
	.w5(32'h3a57b7f9),
	.w6(32'h3cc239e9),
	.w7(32'hbb13a6f4),
	.w8(32'h3a80a071),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14999d),
	.w1(32'hbac96549),
	.w2(32'h3c355c0f),
	.w3(32'h3b29d34b),
	.w4(32'h3b410116),
	.w5(32'hbc870010),
	.w6(32'hb903ef88),
	.w7(32'hbc241420),
	.w8(32'hbc501de7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660c96),
	.w1(32'h3bf3d620),
	.w2(32'h3bc77acf),
	.w3(32'hbd05bc7c),
	.w4(32'h3b9c6809),
	.w5(32'hbb5befa6),
	.w6(32'h3bb0d9dd),
	.w7(32'hbac049b0),
	.w8(32'hbb587d0b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94e260),
	.w1(32'hba425137),
	.w2(32'h3a81e2a9),
	.w3(32'hbc11c9ac),
	.w4(32'hbb9b3a86),
	.w5(32'h3bd738f3),
	.w6(32'h39885adb),
	.w7(32'hba95e50b),
	.w8(32'hbb7a9efc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf6ffb),
	.w1(32'hbc451acf),
	.w2(32'hbc2b1172),
	.w3(32'h3c34f116),
	.w4(32'h3bd45190),
	.w5(32'h3cd075f8),
	.w6(32'hbbda9daa),
	.w7(32'h3bde8bce),
	.w8(32'hbc1200e0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c2d0b),
	.w1(32'h3a8afd81),
	.w2(32'hbc29a64c),
	.w3(32'h3c932010),
	.w4(32'hbc6234a5),
	.w5(32'hbccbca98),
	.w6(32'hbcedb802),
	.w7(32'hbafee5c6),
	.w8(32'h3ca14f44),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c075f),
	.w1(32'h3c0ae60a),
	.w2(32'h3b85e8af),
	.w3(32'hbb597134),
	.w4(32'h3b62d922),
	.w5(32'hba8c0983),
	.w6(32'h3d3ee4ea),
	.w7(32'hba686c5a),
	.w8(32'h3bb5cdff),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26da57),
	.w1(32'h3a8feb3a),
	.w2(32'hbc6207fc),
	.w3(32'hbb6568b7),
	.w4(32'hbc6c6f10),
	.w5(32'hbc9536f9),
	.w6(32'h3c066dd2),
	.w7(32'hbc5a2493),
	.w8(32'h3b5878b2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49e51b),
	.w1(32'h3a846a3a),
	.w2(32'hbba0d868),
	.w3(32'hbbba669d),
	.w4(32'hbc260ba9),
	.w5(32'hbc080a9a),
	.w6(32'h3ca5a0f0),
	.w7(32'hba89bae8),
	.w8(32'h3c801662),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d1601),
	.w1(32'h3b9e7fb3),
	.w2(32'h3bd771cb),
	.w3(32'h3bcbd844),
	.w4(32'hbaa8a8e5),
	.w5(32'h3b5816e4),
	.w6(32'h3cbca99b),
	.w7(32'hbb754026),
	.w8(32'hbab09e09),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46e8d7),
	.w1(32'hbb86b63e),
	.w2(32'h39dabe28),
	.w3(32'hbb2992ba),
	.w4(32'hbb9d2b28),
	.w5(32'hbc91fe3f),
	.w6(32'hbbad4992),
	.w7(32'hb9e805d8),
	.w8(32'hb85e4c28),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a0961),
	.w1(32'hbadf6e31),
	.w2(32'h3b1e05ac),
	.w3(32'hbc9d1530),
	.w4(32'h3b8c2dbf),
	.w5(32'hb96b69bf),
	.w6(32'h3bb49f86),
	.w7(32'h3c35eec1),
	.w8(32'h3c06d5a4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b023),
	.w1(32'h3a031ec4),
	.w2(32'hbb6972bd),
	.w3(32'h3af0ecf4),
	.w4(32'hbb4f206d),
	.w5(32'hbbbb539d),
	.w6(32'h3c0da30a),
	.w7(32'hbb42cdcd),
	.w8(32'hbbac0c13),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8e275),
	.w1(32'h3b109e01),
	.w2(32'h387b6951),
	.w3(32'hbba6a399),
	.w4(32'h39468e87),
	.w5(32'hbbfa1346),
	.w6(32'hbb6a3b3b),
	.w7(32'h3ad9228f),
	.w8(32'h3c544168),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc7b9),
	.w1(32'h3be0e9c0),
	.w2(32'h3ba128b9),
	.w3(32'hbc112f49),
	.w4(32'h3b85cce5),
	.w5(32'h3a9e6739),
	.w6(32'hbc497dee),
	.w7(32'h3b9f07ca),
	.w8(32'h3b942913),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ee67),
	.w1(32'h3c27f23e),
	.w2(32'h3c22d614),
	.w3(32'h3b00a799),
	.w4(32'h3c15bc01),
	.w5(32'h3bd29cd9),
	.w6(32'h3bce1708),
	.w7(32'h3a0573bc),
	.w8(32'hbbd0f62d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc8295),
	.w1(32'h3c02105c),
	.w2(32'h3bda9ae3),
	.w3(32'h3a85eca2),
	.w4(32'h3c5461b5),
	.w5(32'hbbf30b26),
	.w6(32'hbbf077b9),
	.w7(32'hbba48880),
	.w8(32'hbc3234c8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace95b4),
	.w1(32'h385dbe5e),
	.w2(32'h38e48d78),
	.w3(32'hbca67fd4),
	.w4(32'h3af8a6e9),
	.w5(32'h3b1ba37c),
	.w6(32'hbb8790c1),
	.w7(32'h3b508ca5),
	.w8(32'h3b446224),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60a79e),
	.w1(32'hbc4745a8),
	.w2(32'hbc4a8ae2),
	.w3(32'h3b93b6bf),
	.w4(32'hbc1d8fd0),
	.w5(32'hbb81188b),
	.w6(32'h3b47580e),
	.w7(32'hb9358cfb),
	.w8(32'h3c45686d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5a2f),
	.w1(32'h3bac028b),
	.w2(32'hbb43695d),
	.w3(32'hba20f1e1),
	.w4(32'hbc6f8b89),
	.w5(32'hbca27cee),
	.w6(32'h3bbed868),
	.w7(32'h3cadd28b),
	.w8(32'h3cc84686),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c7418),
	.w1(32'hbcaab5b7),
	.w2(32'hbc686256),
	.w3(32'hbc70b940),
	.w4(32'hbc726232),
	.w5(32'hbc13e8c0),
	.w6(32'h3d0be982),
	.w7(32'hbad24c55),
	.w8(32'hbc1982bd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2580e),
	.w1(32'hbcb0b4a7),
	.w2(32'hbca449ec),
	.w3(32'hbb1b6df9),
	.w4(32'hbcdf254a),
	.w5(32'hbcd003d4),
	.w6(32'hbc6271de),
	.w7(32'hbb707b6d),
	.w8(32'hba8f1c8a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ac6b0),
	.w1(32'hbb8aaee5),
	.w2(32'h389cc00a),
	.w3(32'hb8f4e34a),
	.w4(32'h3ba06a86),
	.w5(32'hbb2ab3de),
	.w6(32'h3c640540),
	.w7(32'h3b91294a),
	.w8(32'hbbbda65d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae444da),
	.w1(32'hbbe87453),
	.w2(32'hbbe828a2),
	.w3(32'hbbc233b1),
	.w4(32'hbc1c3d9f),
	.w5(32'hbb4bd1b0),
	.w6(32'hbc618cf3),
	.w7(32'hbc517a8b),
	.w8(32'h3a94b4aa),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b360),
	.w1(32'hb9a83fd7),
	.w2(32'h3b530eff),
	.w3(32'hbb93d511),
	.w4(32'hb9450f07),
	.w5(32'h3b4ef2b6),
	.w6(32'h3c0bdce0),
	.w7(32'hbba1ad0e),
	.w8(32'hbc41b7a6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8882df),
	.w1(32'hba2f5527),
	.w2(32'hba8df1e6),
	.w3(32'h3b04aabb),
	.w4(32'h3a8287e5),
	.w5(32'h3b05b4c5),
	.w6(32'hbc808702),
	.w7(32'h3ad7c94d),
	.w8(32'h3a8e9b45),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2430c),
	.w1(32'h3aeaabd8),
	.w2(32'hbc882e58),
	.w3(32'h3b78e146),
	.w4(32'hbb3104b3),
	.w5(32'hbae30fe7),
	.w6(32'h3a322583),
	.w7(32'hbc34cc5f),
	.w8(32'hbb622d50),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d9085),
	.w1(32'h3c24a556),
	.w2(32'h3c5ff015),
	.w3(32'hb95bffc1),
	.w4(32'hbc0ebdad),
	.w5(32'hbc7e3650),
	.w6(32'h3ca4cf1c),
	.w7(32'hbb7e44d6),
	.w8(32'hbc8a329d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ffd55),
	.w1(32'hbb38d487),
	.w2(32'h3c0bfc05),
	.w3(32'hbbbffbe1),
	.w4(32'hbb9aece7),
	.w5(32'hbc747417),
	.w6(32'hbd365bda),
	.w7(32'hbc9e2e43),
	.w8(32'hbd1b2349),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4742b4),
	.w1(32'h3c1bb80c),
	.w2(32'h3c108adb),
	.w3(32'hbca4b653),
	.w4(32'hbb7e7866),
	.w5(32'hbc54c8b6),
	.w6(32'hbcadb3f0),
	.w7(32'hbc16e051),
	.w8(32'hbbed6c7b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9a8ba),
	.w1(32'h3be9b5d3),
	.w2(32'h3c38a006),
	.w3(32'hbcd7426e),
	.w4(32'h3bbcec99),
	.w5(32'hbba6b747),
	.w6(32'hbcac6a95),
	.w7(32'h3b1f89bd),
	.w8(32'h3b7e8c4a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ea15d),
	.w1(32'h3a68521f),
	.w2(32'hbac1b761),
	.w3(32'hbbec5bd2),
	.w4(32'h3b32ff8d),
	.w5(32'h3a9c4c4f),
	.w6(32'h3c54c3b3),
	.w7(32'h3c2f8944),
	.w8(32'h3c9d1b65),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb057766),
	.w1(32'hba235945),
	.w2(32'h3b8ecf53),
	.w3(32'h3ad398f8),
	.w4(32'hbb34b044),
	.w5(32'h3a438cd9),
	.w6(32'h3c42ae69),
	.w7(32'hbc0ad29b),
	.w8(32'hbbc7a64f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e37a),
	.w1(32'h3b94b512),
	.w2(32'h3b4c45c6),
	.w3(32'hbb96b9a1),
	.w4(32'hbaeabf0f),
	.w5(32'hbbd4f165),
	.w6(32'h3b994c31),
	.w7(32'h3bb940ac),
	.w8(32'h3a6de6a0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58af4c),
	.w1(32'hbb417f3e),
	.w2(32'hba80be4a),
	.w3(32'hbbe5ff73),
	.w4(32'h39eb8ac5),
	.w5(32'h3af3ebc6),
	.w6(32'h3bac9630),
	.w7(32'h3aac4f51),
	.w8(32'hb8d3c040),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf209b),
	.w1(32'h3ade2089),
	.w2(32'hbc055a67),
	.w3(32'h3b63599b),
	.w4(32'hbcb9fb72),
	.w5(32'hbc0d4bb8),
	.w6(32'hbb2dac05),
	.w7(32'h3bb711c0),
	.w8(32'h3d0685c9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8df98a),
	.w1(32'hbaaca32d),
	.w2(32'h3b0d08b5),
	.w3(32'h3d00d6a3),
	.w4(32'hbb71324d),
	.w5(32'h3a4e993f),
	.w6(32'h3cd6c53e),
	.w7(32'hbb3fece0),
	.w8(32'hbbccd931),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba47a2c),
	.w1(32'h3c47a622),
	.w2(32'hbc8d53d7),
	.w3(32'hbc8b5202),
	.w4(32'h3c59f469),
	.w5(32'h3cc94a8c),
	.w6(32'hbabd7227),
	.w7(32'h3b349564),
	.w8(32'h3c0b3ab1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5e859),
	.w1(32'hbb3de299),
	.w2(32'hba70dfc9),
	.w3(32'h3d4b7af2),
	.w4(32'h395b0271),
	.w5(32'h3b450f09),
	.w6(32'hbadba32c),
	.w7(32'h3894e9da),
	.w8(32'h3b44f9f6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9185b42),
	.w1(32'hbb5cb66c),
	.w2(32'hbbdf7585),
	.w3(32'h3b856972),
	.w4(32'hbb9d1546),
	.w5(32'hbc6029d5),
	.w6(32'hb92d9bdd),
	.w7(32'h3b7da99d),
	.w8(32'h3baec139),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2eb51),
	.w1(32'hbcba819c),
	.w2(32'hbc96d959),
	.w3(32'hbbce219c),
	.w4(32'hbc5c1cbd),
	.w5(32'hbb46f4a0),
	.w6(32'h3c950b9b),
	.w7(32'hbae567fb),
	.w8(32'hbbef5394),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b4bb2),
	.w1(32'h3a58831b),
	.w2(32'hbb0a3aea),
	.w3(32'hbbda8cb4),
	.w4(32'hbb340ac6),
	.w5(32'hba9ceeda),
	.w6(32'hbc43d478),
	.w7(32'hbac7b84f),
	.w8(32'h3bbb6834),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e0c59),
	.w1(32'hbceb9cea),
	.w2(32'hbd29d4f1),
	.w3(32'hba4be9cf),
	.w4(32'hbd299ab9),
	.w5(32'hbcf142cf),
	.w6(32'h3c084544),
	.w7(32'h3c97aaa6),
	.w8(32'h3d6dfcc5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce04cd),
	.w1(32'h3b66edfb),
	.w2(32'h3bee2859),
	.w3(32'h3c37e5ce),
	.w4(32'h39f355f1),
	.w5(32'h3c5f7712),
	.w6(32'h3d2da98b),
	.w7(32'hbb31c881),
	.w8(32'hbc419f48),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d194c),
	.w1(32'h3bcd8465),
	.w2(32'h3c8aa7ac),
	.w3(32'h3cb6df28),
	.w4(32'hba4e3668),
	.w5(32'hbcbebf57),
	.w6(32'hbcf85672),
	.w7(32'hbb8df1fc),
	.w8(32'h3ba94793),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd3e0f),
	.w1(32'h3bac1d24),
	.w2(32'h3b81f79e),
	.w3(32'hbc8b681c),
	.w4(32'h3b2df90f),
	.w5(32'h3b6e6f5a),
	.w6(32'h3a8ee826),
	.w7(32'h3a3efba0),
	.w8(32'h3a8fb556),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2f7df),
	.w1(32'h3c1220d9),
	.w2(32'h3c19a5e0),
	.w3(32'h3b16e73e),
	.w4(32'hb9f2498c),
	.w5(32'h3c6831cf),
	.w6(32'h39c0c22e),
	.w7(32'hbb72b3dc),
	.w8(32'hbcff7c58),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb587c47),
	.w1(32'hbb83b723),
	.w2(32'h3b551d5e),
	.w3(32'h3c9f1ed0),
	.w4(32'hbb77b040),
	.w5(32'h3b8ef11e),
	.w6(32'h3b50c003),
	.w7(32'h37ef668a),
	.w8(32'h3c1578d1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d13f),
	.w1(32'h3b0829e6),
	.w2(32'h3ac18804),
	.w3(32'hba83a89a),
	.w4(32'hb8325a44),
	.w5(32'h3ade1fdd),
	.w6(32'h3b25d3d5),
	.w7(32'h3adc0ad3),
	.w8(32'h3b938c5b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8afb84),
	.w1(32'h3a753f62),
	.w2(32'hbac2e220),
	.w3(32'h3c37c0f3),
	.w4(32'h39c75dd5),
	.w5(32'h3b5dcc5a),
	.w6(32'h3c122f57),
	.w7(32'h3b5470be),
	.w8(32'hba94fd50),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116bed),
	.w1(32'hbc1cca05),
	.w2(32'hbbf49649),
	.w3(32'h3c140621),
	.w4(32'hbc2700ec),
	.w5(32'hba81a371),
	.w6(32'hbaff8ae1),
	.w7(32'h3b907c89),
	.w8(32'h3c0f60b0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebb1fc),
	.w1(32'hbb96e05f),
	.w2(32'hbac7e810),
	.w3(32'h3c19f215),
	.w4(32'hbc17f63b),
	.w5(32'hbb6a6328),
	.w6(32'h3be89d04),
	.w7(32'hbb9ada2d),
	.w8(32'h3a1d08ce),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ea7a),
	.w1(32'h3c00fd88),
	.w2(32'hbc83c0a5),
	.w3(32'hbb6e7001),
	.w4(32'h3c5bf902),
	.w5(32'hbb691a42),
	.w6(32'hbaef8066),
	.w7(32'h3c8b615c),
	.w8(32'h3b5d769d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0b2ae),
	.w1(32'hbc0e220d),
	.w2(32'hbb61474a),
	.w3(32'hbc95de2d),
	.w4(32'hbbf4c2c9),
	.w5(32'hbb920765),
	.w6(32'hbc9d4f8e),
	.w7(32'hbb9c4e77),
	.w8(32'hba31b779),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05b38b),
	.w1(32'h3bb07243),
	.w2(32'h3abc979b),
	.w3(32'h3bec733b),
	.w4(32'h3bd153ca),
	.w5(32'hbadcf95d),
	.w6(32'h3bd6ff68),
	.w7(32'h3c761e66),
	.w8(32'h3c73c534),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc679dab),
	.w1(32'h3b173e03),
	.w2(32'h3ae43e8a),
	.w3(32'hbc9257e3),
	.w4(32'h3b822763),
	.w5(32'h3b201949),
	.w6(32'hbc2ed01b),
	.w7(32'h3b073e79),
	.w8(32'h392c368b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ff4ee),
	.w1(32'hbc81fc4b),
	.w2(32'hbc874219),
	.w3(32'h3a6fed1d),
	.w4(32'hbca21ecb),
	.w5(32'hba942c08),
	.w6(32'h3a12fc64),
	.w7(32'hbc7711e7),
	.w8(32'h3b8c8d42),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c937c99),
	.w1(32'h3ad1f02b),
	.w2(32'hbc063e19),
	.w3(32'h3c5b1289),
	.w4(32'h39307b75),
	.w5(32'hbc1a04c9),
	.w6(32'h3c0b4248),
	.w7(32'hbb8d9f18),
	.w8(32'hbc294d7c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c629bb6),
	.w1(32'hbd084df0),
	.w2(32'hbd0a1652),
	.w3(32'h3c025a61),
	.w4(32'hbcce7cce),
	.w5(32'hbd0b06a7),
	.w6(32'h3c253aeb),
	.w7(32'hbd171df1),
	.w8(32'hbd272d45),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d40b1b1),
	.w1(32'hbc9cb855),
	.w2(32'h3d1c63e6),
	.w3(32'h3d6fb15a),
	.w4(32'hbca6ab1d),
	.w5(32'h3d01ce7f),
	.w6(32'h3d368aa3),
	.w7(32'hbccde53b),
	.w8(32'h3be4f9de),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9db62b),
	.w1(32'hbbed0543),
	.w2(32'hbb3f86a1),
	.w3(32'hba89f281),
	.w4(32'hbc4b557e),
	.w5(32'hbbf7f091),
	.w6(32'hbc31a80a),
	.w7(32'hbc3fa0e6),
	.w8(32'hbbfe3332),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3905d5),
	.w1(32'hbacaff8e),
	.w2(32'hbb6dbe03),
	.w3(32'h3c5297d7),
	.w4(32'h3a091b19),
	.w5(32'hb9067997),
	.w6(32'h3c1eb324),
	.w7(32'hb9d6654f),
	.w8(32'hba879a1d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c61288),
	.w1(32'h3c37e7e2),
	.w2(32'h3c070ee4),
	.w3(32'h3aa76a86),
	.w4(32'h3c236a23),
	.w5(32'h3c155033),
	.w6(32'h3b8b81ee),
	.w7(32'h3c99749f),
	.w8(32'h3c1dc084),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951e80),
	.w1(32'hbc10d26f),
	.w2(32'hbd05d787),
	.w3(32'h3b6be680),
	.w4(32'hbc1c5871),
	.w5(32'hbd07330c),
	.w6(32'h3bf0bbb9),
	.w7(32'hbca683e4),
	.w8(32'hbc7f1a40),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d272b04),
	.w1(32'h3a819a81),
	.w2(32'h3a016fec),
	.w3(32'h3d9d1b1f),
	.w4(32'hbb0264c8),
	.w5(32'hbb218452),
	.w6(32'h3d7ffa47),
	.w7(32'hbb53cea5),
	.w8(32'hbaf4e599),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85aaaa),
	.w1(32'h3b8be806),
	.w2(32'h3b8af73a),
	.w3(32'h3ad69694),
	.w4(32'h3c46c8b7),
	.w5(32'h3bbb61c1),
	.w6(32'hb7bbfcfc),
	.w7(32'h3bff6329),
	.w8(32'h3c43da42),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44f572),
	.w1(32'hbba78dd6),
	.w2(32'h3a9c9012),
	.w3(32'hbc1a823a),
	.w4(32'hbb12cb36),
	.w5(32'h3aeff48e),
	.w6(32'hbba53296),
	.w7(32'hba40c7ac),
	.w8(32'h3b400515),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50681),
	.w1(32'h3b612308),
	.w2(32'h3b64285b),
	.w3(32'hba57f972),
	.w4(32'hba3bcaa7),
	.w5(32'h3b9de256),
	.w6(32'h391d667c),
	.w7(32'hbb3f4906),
	.w8(32'hba816d7b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2a29),
	.w1(32'hbba66d8c),
	.w2(32'h3c9279b6),
	.w3(32'hbb594151),
	.w4(32'hbc771929),
	.w5(32'h3c5e4efb),
	.w6(32'hbb854765),
	.w7(32'hbc05ee30),
	.w8(32'h3ab6bf61),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f755),
	.w1(32'h3b9f265e),
	.w2(32'h3ab89832),
	.w3(32'hbc8b6eea),
	.w4(32'h3c66f20d),
	.w5(32'hbaf2dc7b),
	.w6(32'hbbacceea),
	.w7(32'h3c06d5ad),
	.w8(32'hbacbd6b1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc852b65),
	.w1(32'hbb189af7),
	.w2(32'h3b4266d9),
	.w3(32'hbbca6379),
	.w4(32'hba64e70d),
	.w5(32'h3aabf21e),
	.w6(32'h3a5120d9),
	.w7(32'hb983798b),
	.w8(32'h3a0f88aa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abda883),
	.w1(32'hbc3aef52),
	.w2(32'hbd123f11),
	.w3(32'h3a4ffdb9),
	.w4(32'hbcc6bce2),
	.w5(32'hbc7661c5),
	.w6(32'hb98c9a30),
	.w7(32'hbc976831),
	.w8(32'h3c1a3031),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca7e42d),
	.w1(32'h3acac040),
	.w2(32'h3c11a756),
	.w3(32'h3d2a55f9),
	.w4(32'hbb0eb685),
	.w5(32'h3aebb8c0),
	.w6(32'h3cbfaed5),
	.w7(32'h3bed13b3),
	.w8(32'h3c01147c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8dcc),
	.w1(32'h3a17e781),
	.w2(32'h3ba5b294),
	.w3(32'h3b5c732d),
	.w4(32'hbb0d2b2b),
	.w5(32'h3b94f4a6),
	.w6(32'h3c2aed8c),
	.w7(32'hba878074),
	.w8(32'h3bb6c762),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e1d85),
	.w1(32'h39fc4a0d),
	.w2(32'h3bb2d27a),
	.w3(32'hbc0b6ba8),
	.w4(32'h3bdc5887),
	.w5(32'h3c5d99fe),
	.w6(32'hbbc6c759),
	.w7(32'h3bc299af),
	.w8(32'h3c0d7df2),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999bc3c),
	.w1(32'h3bb073d0),
	.w2(32'h3b141865),
	.w3(32'hba91c4a4),
	.w4(32'hbb3b6870),
	.w5(32'hbbb9f791),
	.w6(32'hbbcedaee),
	.w7(32'h3c003963),
	.w8(32'hbb0bfa8d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38941c),
	.w1(32'h3a6dbf09),
	.w2(32'h3a457829),
	.w3(32'hbb618642),
	.w4(32'hbb0e1a1d),
	.w5(32'hba9dcf37),
	.w6(32'hbb9b4c8b),
	.w7(32'h39f2056a),
	.w8(32'h397793f1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a2b611),
	.w1(32'hbbfe757e),
	.w2(32'hbd03e109),
	.w3(32'h3bb6dce3),
	.w4(32'hbc111568),
	.w5(32'hbd00a9b0),
	.w6(32'h3b9a8ccc),
	.w7(32'hbc351978),
	.w8(32'hbc6fbcaa),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc111ea),
	.w1(32'h3a7c3804),
	.w2(32'h3ba61f1a),
	.w3(32'h3d31b84f),
	.w4(32'h3bc76016),
	.w5(32'h3bb46390),
	.w6(32'h3d040bde),
	.w7(32'h3bda06f0),
	.w8(32'h3b86ea9e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93befa),
	.w1(32'hbbfd06c6),
	.w2(32'hbb2990f9),
	.w3(32'hbad917cf),
	.w4(32'hbc09b03b),
	.w5(32'hbbb085e0),
	.w6(32'hbb9846ad),
	.w7(32'hbbf713ba),
	.w8(32'hbb64e0fe),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c194634),
	.w1(32'hbd014bf2),
	.w2(32'h3b375ba4),
	.w3(32'h3c1cc845),
	.w4(32'hbd12a40b),
	.w5(32'h3b883724),
	.w6(32'h3c0ca434),
	.w7(32'hbd263e5c),
	.w8(32'hb955c114),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90c798),
	.w1(32'h39a3dfde),
	.w2(32'h3b60b504),
	.w3(32'h3ce9145e),
	.w4(32'h398c4d4a),
	.w5(32'h3b4cc474),
	.w6(32'h3cbd5b0b),
	.w7(32'h3afdbea3),
	.w8(32'h3b5fb355),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89316d),
	.w1(32'hbaab3250),
	.w2(32'hbb88e710),
	.w3(32'hbae4c110),
	.w4(32'hbc461aee),
	.w5(32'hbbebdc10),
	.w6(32'hbb4f8126),
	.w7(32'hbc287f4d),
	.w8(32'hbbb59cc1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97857a),
	.w1(32'h3b76c216),
	.w2(32'hbc10794e),
	.w3(32'h3c7a500d),
	.w4(32'h3bc89e18),
	.w5(32'hbcc6d017),
	.w6(32'h3b9f3476),
	.w7(32'hbbd35a85),
	.w8(32'hbc94ae8c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87068a),
	.w1(32'h3b9cf23c),
	.w2(32'h3c5d0980),
	.w3(32'h3bfb7361),
	.w4(32'h3aabb85b),
	.w5(32'h3c56898a),
	.w6(32'h3b63bc8c),
	.w7(32'hbc114e18),
	.w8(32'h3b60d9da),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ae79e),
	.w1(32'hbb5e4d8d),
	.w2(32'h3c96f900),
	.w3(32'hbd20e89c),
	.w4(32'h3b83246e),
	.w5(32'h3cc9e8f4),
	.w6(32'hbd186cfe),
	.w7(32'h3c19d048),
	.w8(32'h3ca2fd3f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf03e32),
	.w1(32'hbcfc13d2),
	.w2(32'hbcc70d27),
	.w3(32'hbccdbc97),
	.w4(32'hbccdef93),
	.w5(32'hbc8bb76f),
	.w6(32'hbce9b8fb),
	.w7(32'hbc8a6969),
	.w8(32'hbc74765f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc203454),
	.w1(32'h3c048278),
	.w2(32'h3bf1fb71),
	.w3(32'h3b9d16b3),
	.w4(32'h3bed614f),
	.w5(32'h3ba4ae9e),
	.w6(32'hbbf08748),
	.w7(32'h3a040a6c),
	.w8(32'h3ba6d495),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba997fc2),
	.w1(32'hbbe466e1),
	.w2(32'hbadfec24),
	.w3(32'h3bdf8a9e),
	.w4(32'hbbefe49c),
	.w5(32'hbae5e3ce),
	.w6(32'hbaf86922),
	.w7(32'hbbcc9516),
	.w8(32'hbb09ee94),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add449f),
	.w1(32'hbac939c9),
	.w2(32'hbaf19ab3),
	.w3(32'h3b0feade),
	.w4(32'hbb39da20),
	.w5(32'hbaf32e3d),
	.w6(32'h3ae94b6d),
	.w7(32'hba872d5e),
	.w8(32'hba07036f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af109ab),
	.w1(32'hbbe1c409),
	.w2(32'hbbce08e5),
	.w3(32'h3b05c8bc),
	.w4(32'hbbce4bea),
	.w5(32'hbc6ddb20),
	.w6(32'h3b8f95b9),
	.w7(32'hbbb1a604),
	.w8(32'hbbdbbadc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8337),
	.w1(32'h3c3d9542),
	.w2(32'h3c2c2e1c),
	.w3(32'hbc1bbd21),
	.w4(32'hbaf314cf),
	.w5(32'h3ccba8f4),
	.w6(32'h3b89ed40),
	.w7(32'hbbea2c54),
	.w8(32'h3cb27d5f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3656f4),
	.w1(32'hbcd53aaa),
	.w2(32'h3cc6fb07),
	.w3(32'hbc071ea0),
	.w4(32'hbccca09a),
	.w5(32'h3d09d18f),
	.w6(32'hbcad5094),
	.w7(32'hbc818f5a),
	.w8(32'h3d2739f5),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2d1845),
	.w1(32'hbca3df18),
	.w2(32'hbd5aa981),
	.w3(32'hbd63f740),
	.w4(32'hbc4f480b),
	.w5(32'hbd1c3ea6),
	.w6(32'hbd3e8a5c),
	.w7(32'hbc96e1e4),
	.w8(32'hbd0bad6d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd23f7),
	.w1(32'hbc8ed2f9),
	.w2(32'hbc103fbc),
	.w3(32'h3d61086c),
	.w4(32'hbc6df4d4),
	.w5(32'hbce40ddd),
	.w6(32'h3cae0ec9),
	.w7(32'hbc036abf),
	.w8(32'hbd06fae4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c893a68),
	.w1(32'hbac08a7b),
	.w2(32'h3984daa4),
	.w3(32'h3c956aae),
	.w4(32'h3a31b41d),
	.w5(32'h3b1228b1),
	.w6(32'h3c3e5469),
	.w7(32'h3b53bf32),
	.w8(32'h3ae96eb6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241ebc),
	.w1(32'h3bf675b5),
	.w2(32'hbc2c83d5),
	.w3(32'h3b9d2d84),
	.w4(32'h3c0d6315),
	.w5(32'hbbcae658),
	.w6(32'h3b9a84b9),
	.w7(32'h3c0185fe),
	.w8(32'h3a83425a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb933e18),
	.w1(32'hbb47f6ef),
	.w2(32'hbae22685),
	.w3(32'hbb9ee799),
	.w4(32'h3b6896a5),
	.w5(32'h3bc65f5d),
	.w6(32'hbac6e87a),
	.w7(32'h3a82fde0),
	.w8(32'h3c2d3f44),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2493ab),
	.w1(32'hbb597ddb),
	.w2(32'hbb1181fd),
	.w3(32'hbc01ab50),
	.w4(32'hbba8cf37),
	.w5(32'hbab17a42),
	.w6(32'hbc2de7b8),
	.w7(32'hbb551e6d),
	.w8(32'hba63df77),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cc971),
	.w1(32'h3bca718a),
	.w2(32'h3c22e57e),
	.w3(32'h3b5475da),
	.w4(32'h3c1b0d6b),
	.w5(32'h3c934a6a),
	.w6(32'h3b976e24),
	.w7(32'h3bde9188),
	.w8(32'h3ca30c14),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefca8),
	.w1(32'h3c2c4ac0),
	.w2(32'hbba101fb),
	.w3(32'h3bed1276),
	.w4(32'h3c130620),
	.w5(32'hbaccd84c),
	.w6(32'hba8c3f1e),
	.w7(32'h3bf8f728),
	.w8(32'hbc22d11f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7f3a6),
	.w1(32'hbcda81e8),
	.w2(32'h3c9fbfd6),
	.w3(32'h3c073aed),
	.w4(32'hbd30befe),
	.w5(32'h3d02e16a),
	.w6(32'h3c315690),
	.w7(32'hbd20e4c2),
	.w8(32'h3cc9e340),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ba1e),
	.w1(32'hbb0183e5),
	.w2(32'h395cbd4c),
	.w3(32'h3b6c115d),
	.w4(32'hbb731eb3),
	.w5(32'hba76e35b),
	.w6(32'hbc30acb6),
	.w7(32'hbb560e11),
	.w8(32'hb8bd649f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e7a4),
	.w1(32'hbc01417b),
	.w2(32'hbaf074ff),
	.w3(32'h3b36e6d9),
	.w4(32'hbb4af09a),
	.w5(32'hba7a8b15),
	.w6(32'h3b56e322),
	.w7(32'hbbe5dd4d),
	.w8(32'h3b0e531a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812f35),
	.w1(32'hb9acd1a7),
	.w2(32'hbb2253c7),
	.w3(32'h3c0667fd),
	.w4(32'h3b5134f6),
	.w5(32'h39b2c47c),
	.w6(32'h3c24c80b),
	.w7(32'h3b2c541b),
	.w8(32'h3b023510),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb248da9),
	.w1(32'h3b361786),
	.w2(32'hbace0013),
	.w3(32'hbc13c9d3),
	.w4(32'h3b462596),
	.w5(32'hba3f435d),
	.w6(32'hbc5995ff),
	.w7(32'h3afac567),
	.w8(32'hba0a7f1b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77c8c),
	.w1(32'hbcd08b93),
	.w2(32'hbcce726a),
	.w3(32'hbb95531e),
	.w4(32'hbd02b341),
	.w5(32'hbc75937b),
	.w6(32'hbadb7ce9),
	.w7(32'hbcd9fa09),
	.w8(32'hbb3fe519),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a64c8),
	.w1(32'h3c0f8a3e),
	.w2(32'h3b83e9d8),
	.w3(32'h3be57e0d),
	.w4(32'h3a019365),
	.w5(32'hb9452a4e),
	.w6(32'hbc5309d6),
	.w7(32'h3ba38045),
	.w8(32'h3894ea7d),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc165),
	.w1(32'hbd2a5c20),
	.w2(32'hbb9de89f),
	.w3(32'h3bec9961),
	.w4(32'hbd1ab0f4),
	.w5(32'hbb5cdad4),
	.w6(32'h3bba3853),
	.w7(32'hbd1a0cdf),
	.w8(32'hbb81367e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d203adf),
	.w1(32'h3ac3b6e5),
	.w2(32'hbb4b8035),
	.w3(32'h3d659460),
	.w4(32'h3b47f966),
	.w5(32'hbacf18d2),
	.w6(32'h3d200327),
	.w7(32'h39a5ea83),
	.w8(32'hbb81eeb1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c920a),
	.w1(32'hbc29b4e7),
	.w2(32'h3a6d06ba),
	.w3(32'h39cfac78),
	.w4(32'hbc5441b0),
	.w5(32'h3b9bc530),
	.w6(32'h3af1aec7),
	.w7(32'hbc5062ff),
	.w8(32'h3b9a16d7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule