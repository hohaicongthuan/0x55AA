module layer_8_featuremap_80(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba49321),
	.w1(32'h3aa51d80),
	.w2(32'hbaab11ef),
	.w3(32'h3bc198a5),
	.w4(32'h3af2fa4b),
	.w5(32'hbb0729b6),
	.w6(32'h3bbc7a15),
	.w7(32'h3b2e0c82),
	.w8(32'hba4a6c66),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019152),
	.w1(32'h3aabae43),
	.w2(32'h3abff913),
	.w3(32'h3b09c51b),
	.w4(32'h3ac31a16),
	.w5(32'h3ae39d36),
	.w6(32'h3a96fcb0),
	.w7(32'h3a949961),
	.w8(32'h3aaf4b9f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ed28c),
	.w1(32'h3ae89eac),
	.w2(32'h3a94563d),
	.w3(32'h3b446288),
	.w4(32'h3b31808c),
	.w5(32'h3b01a627),
	.w6(32'h3b487808),
	.w7(32'h3b311b6d),
	.w8(32'h3b140447),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c1411),
	.w1(32'hbb2ef8b7),
	.w2(32'hbb2544b4),
	.w3(32'h3a9ddcd4),
	.w4(32'h39d7b8a0),
	.w5(32'h3a877c29),
	.w6(32'h3af5dde7),
	.w7(32'h3b1c18b3),
	.w8(32'h3af326af),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a207a2c),
	.w1(32'h3b1fbcd5),
	.w2(32'h3aee2cc9),
	.w3(32'h3a710c7c),
	.w4(32'h3b308abe),
	.w5(32'h3b1ca1e8),
	.w6(32'hba7482cf),
	.w7(32'h3a6b9936),
	.w8(32'hbbaffa8b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c78d6),
	.w1(32'hbbe105d6),
	.w2(32'hbb70dd0c),
	.w3(32'hbc1db126),
	.w4(32'hbbb394c0),
	.w5(32'hbaa123cd),
	.w6(32'hbbf071e8),
	.w7(32'hbbb703dc),
	.w8(32'h3b8e1d74),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7cd14),
	.w1(32'h39f869af),
	.w2(32'h3a220e0b),
	.w3(32'h3a6c09fb),
	.w4(32'h3a177b2e),
	.w5(32'h39cb1a5b),
	.w6(32'h39b934a9),
	.w7(32'h3a58a86c),
	.w8(32'h3a8d43bd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1b52),
	.w1(32'h39cf28e0),
	.w2(32'hbac785b7),
	.w3(32'h3bb27692),
	.w4(32'h3b061cd6),
	.w5(32'hba23425c),
	.w6(32'h3b9e848c),
	.w7(32'h3b1be28a),
	.w8(32'hb9b5c2a8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b751f76),
	.w1(32'h3b659507),
	.w2(32'h3af89e91),
	.w3(32'h3b56378f),
	.w4(32'h3b7d0980),
	.w5(32'h3b00a704),
	.w6(32'h3a902b7a),
	.w7(32'h3acc0a01),
	.w8(32'h386e2d5b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d535),
	.w1(32'hbb18e466),
	.w2(32'hbbc78b2e),
	.w3(32'h3ad1c944),
	.w4(32'hbaa73b03),
	.w5(32'hbba27cd0),
	.w6(32'h3bae2d53),
	.w7(32'hb94ff963),
	.w8(32'hbb35f17c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fc13a),
	.w1(32'h3b3150e4),
	.w2(32'h392bcc12),
	.w3(32'h3bda3f4d),
	.w4(32'h3b8bd6fa),
	.w5(32'hba5e6220),
	.w6(32'h3b8bc61b),
	.w7(32'h3a5eb967),
	.w8(32'hba82a992),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5384f5),
	.w1(32'hbb3e8c88),
	.w2(32'hbb842827),
	.w3(32'h3b36f7af),
	.w4(32'hb907bf8d),
	.w5(32'hbb034fb1),
	.w6(32'h3b35c870),
	.w7(32'h3a1d0446),
	.w8(32'h399bbd4f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3242c),
	.w1(32'h3aa6b451),
	.w2(32'h39bc256b),
	.w3(32'h3b0480c9),
	.w4(32'h3b11ae23),
	.w5(32'h3b035693),
	.w6(32'h3a3307ad),
	.w7(32'h3a8b8cc9),
	.w8(32'hbbc1dc52),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35ee6),
	.w1(32'hbb5bd558),
	.w2(32'hbb4cfa54),
	.w3(32'hbb85c0fb),
	.w4(32'hbb4553b1),
	.w5(32'hbb4f0d10),
	.w6(32'hbb920bea),
	.w7(32'hbb8a877b),
	.w8(32'hbb75ceed),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405399),
	.w1(32'hbb1c7ce0),
	.w2(32'hbb0a76dc),
	.w3(32'hbb2e4f1c),
	.w4(32'hbb1c6c25),
	.w5(32'hbb169ac3),
	.w6(32'hbb3d79f1),
	.w7(32'hbb2581d3),
	.w8(32'h3547d63c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399764f6),
	.w1(32'h37be1d51),
	.w2(32'hb7918d14),
	.w3(32'hb933db70),
	.w4(32'hb95408a4),
	.w5(32'hb940d304),
	.w6(32'hb621adfc),
	.w7(32'h3933920f),
	.w8(32'hba07bb64),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68b939),
	.w1(32'hb9ab3c66),
	.w2(32'hbac98244),
	.w3(32'h3a99efb6),
	.w4(32'h3a76d326),
	.w5(32'hbadb2f32),
	.w6(32'hb991abe4),
	.w7(32'h379fc247),
	.w8(32'hb8da1f56),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb389),
	.w1(32'h3a938e8d),
	.w2(32'hbae0f9bf),
	.w3(32'h3bb4804d),
	.w4(32'h3b87250b),
	.w5(32'h3b117cf0),
	.w6(32'h3b8b05ba),
	.w7(32'h3ac82184),
	.w8(32'h3b7ac79a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53b43c),
	.w1(32'hbaf00d51),
	.w2(32'hbc7292f3),
	.w3(32'h3c48b6ec),
	.w4(32'hbb36c446),
	.w5(32'hbc7a8e14),
	.w6(32'h3c7cfda3),
	.w7(32'h3b35cbca),
	.w8(32'hbc3e98b8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d30a),
	.w1(32'h3b657c1f),
	.w2(32'hbaa7bd62),
	.w3(32'h3b8cece2),
	.w4(32'h3b5cb202),
	.w5(32'h3b393b14),
	.w6(32'h3a3079b5),
	.w7(32'hba9c977d),
	.w8(32'h3a66ec79),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e4763),
	.w1(32'hb9271c2a),
	.w2(32'h3a0aeb9b),
	.w3(32'hbaef35b0),
	.w4(32'hbad14318),
	.w5(32'h3b4b99c0),
	.w6(32'hbaedf964),
	.w7(32'hbac197b4),
	.w8(32'h39025240),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef7f1b),
	.w1(32'hbaee8b56),
	.w2(32'hba90ed2c),
	.w3(32'hbad15d8c),
	.w4(32'hbad2c57c),
	.w5(32'hba995370),
	.w6(32'hbac81e70),
	.w7(32'hbb420a6a),
	.w8(32'h3a5e85c3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6eda4e),
	.w1(32'h3c0189f4),
	.w2(32'hbb92058b),
	.w3(32'h3ca709ee),
	.w4(32'h3c6999a7),
	.w5(32'hbb10c254),
	.w6(32'h3c8d2b18),
	.w7(32'h3bfe5180),
	.w8(32'hbba8134b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e9100),
	.w1(32'h39011b35),
	.w2(32'h3ac1192a),
	.w3(32'hb9d71d86),
	.w4(32'h39d8b5a4),
	.w5(32'h3af43c8e),
	.w6(32'hba6ee1ba),
	.w7(32'hb9d61e08),
	.w8(32'h3af80cb9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1cf09),
	.w1(32'h3b89d059),
	.w2(32'h3a3d7715),
	.w3(32'h3a72c29a),
	.w4(32'h3b56cbe0),
	.w5(32'h3ab29f74),
	.w6(32'h3b91d158),
	.w7(32'h3b4dc97a),
	.w8(32'h3b7231fe),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bf0b),
	.w1(32'h3b61d803),
	.w2(32'h3a2c7dc6),
	.w3(32'h3bcbdefa),
	.w4(32'h3bc0e16c),
	.w5(32'h3ac1c1a9),
	.w6(32'h3b9b2364),
	.w7(32'h3a8e6d98),
	.w8(32'hb9cdeb42),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2c5bb),
	.w1(32'h3ad914f5),
	.w2(32'h3b0a0982),
	.w3(32'h3ae0a2a4),
	.w4(32'h3b2339ec),
	.w5(32'h3b3317f1),
	.w6(32'h3ae4e52b),
	.w7(32'h3ae1c413),
	.w8(32'h3ad8aaca),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cda7472),
	.w1(32'h3a1cb577),
	.w2(32'hbcbb432b),
	.w3(32'h3cce7ad5),
	.w4(32'h3b9d559d),
	.w5(32'hbca9dc59),
	.w6(32'h3c7b80d2),
	.w7(32'hbb84ced2),
	.w8(32'hbc52e736),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199894),
	.w1(32'hba8bbc80),
	.w2(32'hbb1f996a),
	.w3(32'h3b6ffac3),
	.w4(32'h397079d0),
	.w5(32'hbb08a588),
	.w6(32'h3af3626c),
	.w7(32'hba2f78c0),
	.w8(32'hbab42474),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a659945),
	.w1(32'h3a4f5794),
	.w2(32'h3a4da4e5),
	.w3(32'h3a80083b),
	.w4(32'h3a357b22),
	.w5(32'h3a0e83a6),
	.w6(32'h3a3c7f4f),
	.w7(32'h3a161730),
	.w8(32'h3aef18fe),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aa894),
	.w1(32'hbb483c1f),
	.w2(32'hbb5fc623),
	.w3(32'hbb0699dd),
	.w4(32'hbb415159),
	.w5(32'hbb039822),
	.w6(32'hb8da6817),
	.w7(32'hba5a335a),
	.w8(32'h3b316303),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841354),
	.w1(32'h3b9aa7e7),
	.w2(32'h3b99e509),
	.w3(32'h3aedca7d),
	.w4(32'h3b180189),
	.w5(32'h3b8cb495),
	.w6(32'h3b1354bf),
	.w7(32'h3a79acd6),
	.w8(32'h3b1ec2a6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba316ea7),
	.w1(32'hbb1840bf),
	.w2(32'hba6fd9f7),
	.w3(32'h39a50d85),
	.w4(32'hb963b3b8),
	.w5(32'hb98c8dd9),
	.w6(32'h3a0af6c6),
	.w7(32'h3aba7d29),
	.w8(32'h3923a306),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a752f49),
	.w1(32'h3ab90a2e),
	.w2(32'hb8126dd0),
	.w3(32'hb97d35e8),
	.w4(32'hba68a1a2),
	.w5(32'h3a0ea306),
	.w6(32'h3aa120ae),
	.w7(32'hb9b8b1e1),
	.w8(32'hbbcb2e2a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d5df2),
	.w1(32'hbb938b02),
	.w2(32'hbb84e992),
	.w3(32'hbbd9b719),
	.w4(32'hbb42d482),
	.w5(32'hbb05b7f5),
	.w6(32'hbbee73eb),
	.w7(32'hbb89158b),
	.w8(32'h3ad312da),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b700427),
	.w1(32'h3a915b9d),
	.w2(32'hbb6c3e5c),
	.w3(32'h3b807c01),
	.w4(32'h39212f7d),
	.w5(32'hbb7e8f55),
	.w6(32'h3b34515d),
	.w7(32'hb924fab4),
	.w8(32'hbad117c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e511),
	.w1(32'h3b06febc),
	.w2(32'h3942f569),
	.w3(32'h3b059dc7),
	.w4(32'h3afc9cee),
	.w5(32'h3a85fb4c),
	.w6(32'h3b254ba7),
	.w7(32'h3a1d62f9),
	.w8(32'h39695873),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16819d),
	.w1(32'h3b0f546b),
	.w2(32'h3af09845),
	.w3(32'h3abfa7e3),
	.w4(32'h3aa2ed7a),
	.w5(32'h3a831913),
	.w6(32'hb994ea7d),
	.w7(32'hba558659),
	.w8(32'hbbd19304),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5a60a),
	.w1(32'hbb8d39d2),
	.w2(32'hbb780a5a),
	.w3(32'hbb8779c8),
	.w4(32'hbb79d337),
	.w5(32'hbb6d9428),
	.w6(32'hbb9c91c6),
	.w7(32'hbb73b263),
	.w8(32'h3b1bffff),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e106d),
	.w1(32'h3a14b780),
	.w2(32'h39eec796),
	.w3(32'h3aa3dbb2),
	.w4(32'h3a5d79ed),
	.w5(32'h3a801561),
	.w6(32'h3acba8f2),
	.w7(32'h3a58ac5e),
	.w8(32'h3a854c4a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a57bd),
	.w1(32'hbbcdb844),
	.w2(32'hbbc1c372),
	.w3(32'h3c079c31),
	.w4(32'h3b7f434e),
	.w5(32'h3aec135a),
	.w6(32'h3bc05a1d),
	.w7(32'h39ecc15a),
	.w8(32'hb954f320),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9a8fc),
	.w1(32'hb940382e),
	.w2(32'hbb4247f3),
	.w3(32'h3ade90d7),
	.w4(32'hba002260),
	.w5(32'hbb3796ce),
	.w6(32'h3a859592),
	.w7(32'h38d9e83a),
	.w8(32'hbb10404e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0659b0),
	.w1(32'hba06d830),
	.w2(32'hb9a6a3b8),
	.w3(32'hba5968f0),
	.w4(32'hba28e0ab),
	.w5(32'hb9806a94),
	.w6(32'hba494667),
	.w7(32'hb9fce11d),
	.w8(32'hb956adab),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00e854),
	.w1(32'h3a4289c0),
	.w2(32'hba08bfde),
	.w3(32'h3b619730),
	.w4(32'h3a8e083d),
	.w5(32'hba7e8969),
	.w6(32'h3b2c064a),
	.w7(32'h398dad2a),
	.w8(32'hba18fb3e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda84ca),
	.w1(32'h3a50b26e),
	.w2(32'hbba4483c),
	.w3(32'h3c04184b),
	.w4(32'h3a323db1),
	.w5(32'hbbef6933),
	.w6(32'h3bb35733),
	.w7(32'hba1bc4a2),
	.w8(32'hbbd9037b),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadac3e),
	.w1(32'hbb1760c2),
	.w2(32'hbba540da),
	.w3(32'h3a2bfed9),
	.w4(32'hbb4d880d),
	.w5(32'hbba4bab8),
	.w6(32'h3aad7572),
	.w7(32'hb99461f9),
	.w8(32'hbb446e13),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367d27f4),
	.w1(32'h374945ce),
	.w2(32'hb63242a5),
	.w3(32'h376c618c),
	.w4(32'h37b9a691),
	.w5(32'h368930a4),
	.w6(32'h375326e9),
	.w7(32'h37c2a6c1),
	.w8(32'h36947746),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05fd9e),
	.w1(32'h3b89bc66),
	.w2(32'hbaced4c8),
	.w3(32'h3bdde7e5),
	.w4(32'h3afb3ce2),
	.w5(32'hbbaa2985),
	.w6(32'h3bd4855a),
	.w7(32'h3afd6ab2),
	.w8(32'hbb6b602b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab99353),
	.w1(32'h399d5768),
	.w2(32'hb992604e),
	.w3(32'h3ad8744c),
	.w4(32'h3a59800e),
	.w5(32'h3a34edf2),
	.w6(32'h3ac6c038),
	.w7(32'h3a64de63),
	.w8(32'h3a079f6c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09942a),
	.w1(32'hb9cfb17d),
	.w2(32'hbb1e3dfa),
	.w3(32'h3ba47820),
	.w4(32'h3b5a7dfb),
	.w5(32'h3935bffa),
	.w6(32'h3b4c4e87),
	.w7(32'h3b4687b9),
	.w8(32'hba2cbf73),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f95e39),
	.w1(32'hbb3573b8),
	.w2(32'h3ad3bf1a),
	.w3(32'hbaf841ab),
	.w4(32'hbb4d63f3),
	.w5(32'h3b62dcbc),
	.w6(32'hbb4cecca),
	.w7(32'hbb978c27),
	.w8(32'h3b02a30c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8be5b),
	.w1(32'h3b088d82),
	.w2(32'hb9d94048),
	.w3(32'h3c7ab8ed),
	.w4(32'h3bc2c2d4),
	.w5(32'hbb3ead2e),
	.w6(32'h3c60976d),
	.w7(32'h3bd8c871),
	.w8(32'hbb5c5dde),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31e29d),
	.w1(32'h3ab0b8da),
	.w2(32'h3972d278),
	.w3(32'h3bb9bad2),
	.w4(32'h3b3ee383),
	.w5(32'h3a882359),
	.w6(32'h3b2e0e54),
	.w7(32'h3aa6ba7f),
	.w8(32'hba33c970),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77bdca),
	.w1(32'h3ad07d2d),
	.w2(32'hbb02ca1b),
	.w3(32'h3b91524c),
	.w4(32'h3b61fbdd),
	.w5(32'hb9b6338b),
	.w6(32'h3bd5322c),
	.w7(32'h3b38d974),
	.w8(32'hbab3eed1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370da7f9),
	.w1(32'h38550ad4),
	.w2(32'h373563bf),
	.w3(32'hb6de1c6e),
	.w4(32'h37e8ba37),
	.w5(32'h3682c6b1),
	.w6(32'h35aaf29d),
	.w7(32'h3797f677),
	.w8(32'h36d7f46c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4bff0),
	.w1(32'hba973928),
	.w2(32'hbc1e83fb),
	.w3(32'h3b513cf1),
	.w4(32'hba42c960),
	.w5(32'hbc299b08),
	.w6(32'h3beec39c),
	.w7(32'hb9aee54a),
	.w8(32'hbb8c7eab),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1af400),
	.w1(32'hbb1dc724),
	.w2(32'hbb72f382),
	.w3(32'h3ae82cd5),
	.w4(32'h38d7f593),
	.w5(32'hba75ed95),
	.w6(32'h3a0ed613),
	.w7(32'hba3c55e5),
	.w8(32'hb9e31ce4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a805906),
	.w1(32'hbb20d356),
	.w2(32'hbb8618e0),
	.w3(32'h3b8e00ce),
	.w4(32'hba971896),
	.w5(32'hbb7fe56c),
	.w6(32'h3b3ff8cd),
	.w7(32'h39c161b0),
	.w8(32'hbb47412b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093780),
	.w1(32'h3af48af4),
	.w2(32'h37cfe720),
	.w3(32'h3b6990b1),
	.w4(32'h3b099bb4),
	.w5(32'hba5ed991),
	.w6(32'h3b173b6f),
	.w7(32'h3a57cd0e),
	.w8(32'hbac9ac62),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965e1f9),
	.w1(32'h3a505475),
	.w2(32'h3a849dba),
	.w3(32'h3b66a309),
	.w4(32'h3b2d6bc8),
	.w5(32'h3aacce78),
	.w6(32'h3aba8581),
	.w7(32'h3b226b27),
	.w8(32'h3a636778),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5127d),
	.w1(32'hb9a28dd5),
	.w2(32'hb9ed6f8c),
	.w3(32'h39e7c4cb),
	.w4(32'hb89f98d2),
	.w5(32'hb9568cb3),
	.w6(32'h3a068cd3),
	.w7(32'h39909bfc),
	.w8(32'hb68f1ef1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db8fc2),
	.w1(32'h383069f6),
	.w2(32'h3927470d),
	.w3(32'h3916d088),
	.w4(32'h39241e5b),
	.w5(32'h398239f5),
	.w6(32'h39292ae5),
	.w7(32'h394b11e8),
	.w8(32'h39489b87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f20ac),
	.w1(32'hbbb48800),
	.w2(32'hbbdda3ce),
	.w3(32'h3ac322d6),
	.w4(32'hbb0b336e),
	.w5(32'hbb4b10d6),
	.w6(32'h3b6a2cf8),
	.w7(32'hba94ac9a),
	.w8(32'hba6e5b92),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61d36a),
	.w1(32'h3a5bebdc),
	.w2(32'h386d4812),
	.w3(32'h3af4a938),
	.w4(32'h3b028109),
	.w5(32'h3a5189cb),
	.w6(32'h3b115be7),
	.w7(32'h3b1ebd6e),
	.w8(32'h3a7dd3f6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35831df7),
	.w1(32'hb94382c0),
	.w2(32'hba5c56f2),
	.w3(32'hb70716d4),
	.w4(32'h39075450),
	.w5(32'hba3eac7a),
	.w6(32'h38a56245),
	.w7(32'h39bfe7dc),
	.w8(32'hba54f78d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32df1d),
	.w1(32'hba44d335),
	.w2(32'hbb4b26a1),
	.w3(32'h3a9234b3),
	.w4(32'hba0175b9),
	.w5(32'hbb071a9f),
	.w6(32'h3a6cc4c0),
	.w7(32'hb8599833),
	.w8(32'hba9785d9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2aef82),
	.w1(32'h3b050fbe),
	.w2(32'h3b247f2d),
	.w3(32'h3abd3f3e),
	.w4(32'h3b3fa796),
	.w5(32'h3b81c08c),
	.w6(32'h3a46f8a2),
	.w7(32'h3b0bb97a),
	.w8(32'h3b2abb6b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d19019),
	.w1(32'hbb4f91f5),
	.w2(32'hbb9d9410),
	.w3(32'hbb0386fb),
	.w4(32'hbb82139c),
	.w5(32'hbb870755),
	.w6(32'hb9681b02),
	.w7(32'hbb13f3fd),
	.w8(32'hbb0984a4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e193d8),
	.w1(32'h37db04b7),
	.w2(32'hb9c54709),
	.w3(32'hb8b8e3c8),
	.w4(32'hb839bd8d),
	.w5(32'hb9e1a3b4),
	.w6(32'hb8ec51f2),
	.w7(32'h37ae49e3),
	.w8(32'hba094731),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b513b34),
	.w1(32'h3c02d9be),
	.w2(32'h3b291151),
	.w3(32'h3c1d77df),
	.w4(32'h3bc3a511),
	.w5(32'hb9bfd819),
	.w6(32'h3bc6e147),
	.w7(32'h3ba509e4),
	.w8(32'hb91833df),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978abb3),
	.w1(32'hb991064a),
	.w2(32'hb8fff924),
	.w3(32'hb9a1d97e),
	.w4(32'hb9a17e48),
	.w5(32'hb916f2ee),
	.w6(32'hb981a39f),
	.w7(32'hb978ec56),
	.w8(32'hb8f6a26d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b375fe0),
	.w1(32'h3b423544),
	.w2(32'h3a7376ae),
	.w3(32'h3b8172b0),
	.w4(32'h3b598f49),
	.w5(32'h3a988a87),
	.w6(32'h3ad84aa6),
	.w7(32'h3a91943c),
	.w8(32'h393110c7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e6ac1f),
	.w1(32'hb960d9d8),
	.w2(32'hb98f59e7),
	.w3(32'hb8bbc652),
	.w4(32'hb9a4440d),
	.w5(32'hb9d61a95),
	.w6(32'h39686505),
	.w7(32'hb91ca0bf),
	.w8(32'hb985bf8d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17bb0e),
	.w1(32'hba82e504),
	.w2(32'hbb98e87f),
	.w3(32'h3b82a644),
	.w4(32'h3a42ef57),
	.w5(32'hbb4f2667),
	.w6(32'h3b8670f9),
	.w7(32'hb993ef5e),
	.w8(32'hba31a39e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378b81bf),
	.w1(32'h37e62cf1),
	.w2(32'h3780bb3e),
	.w3(32'h3704cf42),
	.w4(32'h37c15c0b),
	.w5(32'h3752b370),
	.w6(32'hb7157a7d),
	.w7(32'h3604817f),
	.w8(32'hb6825817),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade174f),
	.w1(32'hba9b6b82),
	.w2(32'hba9b8e6d),
	.w3(32'hba8fe141),
	.w4(32'hba590c11),
	.w5(32'hba87a3f8),
	.w6(32'hbadf1d77),
	.w7(32'hba96f90c),
	.w8(32'hba1c3102),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390abb54),
	.w1(32'h38e133c1),
	.w2(32'hb7677039),
	.w3(32'h391951f9),
	.w4(32'h39029263),
	.w5(32'hb7165aae),
	.w6(32'h3952f9cf),
	.w7(32'h3911a3f8),
	.w8(32'hb82e1f70),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8979e4),
	.w1(32'h3aaaea0b),
	.w2(32'hbb11de9e),
	.w3(32'h3b9cb804),
	.w4(32'h3a9c09e5),
	.w5(32'hbb3e425a),
	.w6(32'h3b7dc921),
	.w7(32'hba31e765),
	.w8(32'hbabb956e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35fb29),
	.w1(32'hbb074cd3),
	.w2(32'hbc0a1fd8),
	.w3(32'h3b421284),
	.w4(32'hbb3bbc53),
	.w5(32'hbc07eb24),
	.w6(32'h3b8e1805),
	.w7(32'hba51bc19),
	.w8(32'hbba5462d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14822f),
	.w1(32'h3a0874db),
	.w2(32'h3a4c6e91),
	.w3(32'h39d8f376),
	.w4(32'h3a04fdd5),
	.w5(32'h39db78cf),
	.w6(32'h39aedbab),
	.w7(32'h39c8023f),
	.w8(32'h39b01037),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f6e3a9),
	.w1(32'hb8bdbc71),
	.w2(32'hb897dab7),
	.w3(32'hb6def613),
	.w4(32'hb88a42c7),
	.w5(32'hb886ea43),
	.w6(32'h374215a1),
	.w7(32'hb7ddae26),
	.w8(32'hb7eec984),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998a39d),
	.w1(32'h3af37bf4),
	.w2(32'h3a9e76c0),
	.w3(32'h3b93a65e),
	.w4(32'h3b94b80a),
	.w5(32'h3b08b03a),
	.w6(32'h395bc3cf),
	.w7(32'h3a30a207),
	.w8(32'hba95cadf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11d429),
	.w1(32'hbabd1724),
	.w2(32'hbb5d72d2),
	.w3(32'h3b80fb2e),
	.w4(32'h39a26d1f),
	.w5(32'hbb526b86),
	.w6(32'h3b2930e0),
	.w7(32'hbab17832),
	.w8(32'hbb485ba7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2db4d8),
	.w1(32'hbc01b1a7),
	.w2(32'hbb02230a),
	.w3(32'h3b559094),
	.w4(32'hbbb2b658),
	.w5(32'h3b22ce92),
	.w6(32'h3b7f40e3),
	.w7(32'h3bb58df4),
	.w8(32'h3b86002f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0af32),
	.w1(32'hb9a50249),
	.w2(32'hbbdc3e78),
	.w3(32'h3c26d62c),
	.w4(32'h3b0fce38),
	.w5(32'hbbbcdb66),
	.w6(32'h3c00e603),
	.w7(32'h399a9dbc),
	.w8(32'hbb8988a3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa70056),
	.w1(32'h3aaf9e7b),
	.w2(32'h3921a8eb),
	.w3(32'h3be78203),
	.w4(32'h3bb893aa),
	.w5(32'h3b14617d),
	.w6(32'h3b3f572c),
	.w7(32'h3b65d17d),
	.w8(32'h39483a88),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d81013),
	.w1(32'h388efc75),
	.w2(32'h389b14f3),
	.w3(32'hb8f8661a),
	.w4(32'hb835ec08),
	.w5(32'hb7cc5d81),
	.w6(32'hb91cc74b),
	.w7(32'hb81c59ad),
	.w8(32'hb79538b0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d92f4f),
	.w1(32'hb7521709),
	.w2(32'hb84524ea),
	.w3(32'hb7937405),
	.w4(32'hb719545e),
	.w5(32'hb823ac1e),
	.w6(32'hb6d2c04d),
	.w7(32'h37014038),
	.w8(32'hb78b4501),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60c0b12),
	.w1(32'hb8346016),
	.w2(32'hb95a21c4),
	.w3(32'hb6926d68),
	.w4(32'hb84d297a),
	.w5(32'hb92aba73),
	.w6(32'h38d92ed0),
	.w7(32'h37d82be6),
	.w8(32'hb86fde4d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ccd81),
	.w1(32'h3a47f015),
	.w2(32'h3a7f611f),
	.w3(32'hb9e719be),
	.w4(32'h3a8ecf81),
	.w5(32'h3abcc7e6),
	.w6(32'hb9aed201),
	.w7(32'h3a5899c7),
	.w8(32'h3a4816f0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba501248),
	.w1(32'hba9d18e9),
	.w2(32'h3a3b10d5),
	.w3(32'h39d6c5e3),
	.w4(32'h3a7b5ed8),
	.w5(32'h3b170144),
	.w6(32'h3a8175e1),
	.w7(32'h3a790d88),
	.w8(32'h3b1ea4b2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12f0d0),
	.w1(32'hbacb8c4a),
	.w2(32'hba374682),
	.w3(32'hbb147b85),
	.w4(32'hbaa7e80d),
	.w5(32'hb83fb021),
	.w6(32'hba156291),
	.w7(32'hb7af72a9),
	.w8(32'h3a948c18),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2bc6),
	.w1(32'hba9bed43),
	.w2(32'h3a934062),
	.w3(32'h3b167712),
	.w4(32'h3b06138d),
	.w5(32'h3b2b16d3),
	.w6(32'h38cb920d),
	.w7(32'h394b931f),
	.w8(32'h39228a85),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18b749),
	.w1(32'h3a3cf404),
	.w2(32'hb9be6f43),
	.w3(32'h3b38af17),
	.w4(32'h3a8a185a),
	.w5(32'hb99b7e64),
	.w6(32'h3b06a105),
	.w7(32'hb8821e25),
	.w8(32'hba53fcb1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f3eb8),
	.w1(32'hba8665d7),
	.w2(32'hbb114781),
	.w3(32'hbaddeef5),
	.w4(32'hbb036e7b),
	.w5(32'hbb2b74de),
	.w6(32'hba960b9d),
	.w7(32'hbb13e37e),
	.w8(32'hbb2ee5ef),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcdd72),
	.w1(32'hbb80ab60),
	.w2(32'hbbb652db),
	.w3(32'hba300518),
	.w4(32'hbb8b6108),
	.w5(32'hbbba3329),
	.w6(32'hba47c2e8),
	.w7(32'hbaef4c1a),
	.w8(32'hbb6ba53a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75d3a7),
	.w1(32'h3b1d58eb),
	.w2(32'h3a80cc10),
	.w3(32'h3bc0dad3),
	.w4(32'h3b5abe81),
	.w5(32'h3a90ece9),
	.w6(32'h3abd3f0a),
	.w7(32'hb9a72fb3),
	.w8(32'hbad594ea),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373eaa85),
	.w1(32'h37802935),
	.w2(32'hb7f5aef9),
	.w3(32'h375eee1a),
	.w4(32'h37ea608f),
	.w5(32'hb797fbc6),
	.w6(32'h36a32822),
	.w7(32'h372c6298),
	.w8(32'hb7c12a76),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c24474),
	.w1(32'h37308095),
	.w2(32'hb80fab42),
	.w3(32'hb882a820),
	.w4(32'h386c1586),
	.w5(32'hb76e0399),
	.w6(32'hb7d8a8e9),
	.w7(32'h38b43631),
	.w8(32'h36ba657a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8051d4b),
	.w1(32'h36d43c70),
	.w2(32'hb75ab9b1),
	.w3(32'hb81b17cd),
	.w4(32'hb77f5dba),
	.w5(32'hb7abbd14),
	.w6(32'hb6fc8e22),
	.w7(32'h36960612),
	.w8(32'hb6855d5f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b211dc),
	.w1(32'hb96f786e),
	.w2(32'h395332dd),
	.w3(32'hb927856d),
	.w4(32'h38c38605),
	.w5(32'h39a4d351),
	.w6(32'hb88ad25f),
	.w7(32'h393a4270),
	.w8(32'h39c05ecf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f647d),
	.w1(32'h3ab37350),
	.w2(32'h3a9011f0),
	.w3(32'hb89e4e64),
	.w4(32'h3a48d614),
	.w5(32'h3a9bccd4),
	.w6(32'hb9f2de91),
	.w7(32'h38eb32da),
	.w8(32'h3a10adbf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b79e),
	.w1(32'hba6d7621),
	.w2(32'hbab8e048),
	.w3(32'hba89c2c4),
	.w4(32'hb9cd9849),
	.w5(32'hba701630),
	.w6(32'h38690f11),
	.w7(32'h3a975faf),
	.w8(32'h3a47b759),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a224b29),
	.w1(32'hba91cbd2),
	.w2(32'hb7d8a36d),
	.w3(32'h3b78be41),
	.w4(32'h3a6dd83c),
	.w5(32'h3ac24e63),
	.w6(32'h3948afc1),
	.w7(32'hba76b4df),
	.w8(32'hb94d47e5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba066872),
	.w1(32'hb95d947c),
	.w2(32'h390ef790),
	.w3(32'hba4b1983),
	.w4(32'hb978603e),
	.w5(32'h39e3f581),
	.w6(32'hb9c901a8),
	.w7(32'h399ce5b5),
	.w8(32'h39e20622),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7159aa),
	.w1(32'h3b6b1c62),
	.w2(32'hbb23726e),
	.w3(32'h3c004036),
	.w4(32'h3b860169),
	.w5(32'hbb94ae73),
	.w6(32'h3bf1a868),
	.w7(32'h3b82afde),
	.w8(32'hbb4aa15a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55e8c3),
	.w1(32'h3b3265dd),
	.w2(32'h3abb4f62),
	.w3(32'h39c775c0),
	.w4(32'h3abfaef6),
	.w5(32'h38880cc4),
	.w6(32'hba0cec87),
	.w7(32'h36b9d809),
	.w8(32'hba569d0b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33778f),
	.w1(32'h39a2702b),
	.w2(32'h39da3051),
	.w3(32'hb9e12cf1),
	.w4(32'h3a1ca3a0),
	.w5(32'h3a59faa7),
	.w6(32'hba360b22),
	.w7(32'hb97f0803),
	.w8(32'h38d2a9d8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72a912),
	.w1(32'hba5a12ec),
	.w2(32'h3a220c76),
	.w3(32'hba83d1a6),
	.w4(32'hbaa0b11f),
	.w5(32'h39edec55),
	.w6(32'hb9f456c0),
	.w7(32'hba0c5ae4),
	.w8(32'h3a0b48b0),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e1447),
	.w1(32'h3b379570),
	.w2(32'h3a9dba3d),
	.w3(32'h3ad20326),
	.w4(32'h3b0390c8),
	.w5(32'h3a038794),
	.w6(32'h3881917a),
	.w7(32'hb8c54374),
	.w8(32'hb9e590c8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89ab9a),
	.w1(32'hba7d92d8),
	.w2(32'hbb1a8cd1),
	.w3(32'hba99e06e),
	.w4(32'hbb5c0a48),
	.w5(32'hbb3b9393),
	.w6(32'hbafbac6b),
	.w7(32'hbb80b826),
	.w8(32'hbb63a455),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2c09a),
	.w1(32'hba12532b),
	.w2(32'h39fb8269),
	.w3(32'h3a091ab8),
	.w4(32'hbabb2eac),
	.w5(32'h39ad98e9),
	.w6(32'h3a8a891e),
	.w7(32'hb9cce6af),
	.w8(32'h3a4487c4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac296c0),
	.w1(32'hbab6d2ae),
	.w2(32'hb9829267),
	.w3(32'hbb17596f),
	.w4(32'hbad15c1e),
	.w5(32'h38031a20),
	.w6(32'hbad7943e),
	.w7(32'hb9e5d83c),
	.w8(32'h3a804046),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9787b50),
	.w1(32'h38402977),
	.w2(32'h3693d437),
	.w3(32'hb952d3e0),
	.w4(32'h37f9f70a),
	.w5(32'h391db64d),
	.w6(32'hb8fea904),
	.w7(32'h393d6b74),
	.w8(32'h396694c3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae9766),
	.w1(32'h3a6e40da),
	.w2(32'hba36345e),
	.w3(32'h3a9d9ba4),
	.w4(32'h3a882875),
	.w5(32'h39a9a64f),
	.w6(32'h3aa7bb85),
	.w7(32'h3ad55029),
	.w8(32'h391c9567),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d27290),
	.w1(32'hb8366e75),
	.w2(32'h3910fb61),
	.w3(32'h38ae7fce),
	.w4(32'h38005b8c),
	.w5(32'h39c2b308),
	.w6(32'h38885063),
	.w7(32'h38c8f2a6),
	.w8(32'h3a1fdb36),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7b2be),
	.w1(32'hba53801f),
	.w2(32'hba062242),
	.w3(32'h39110abc),
	.w4(32'hba344d87),
	.w5(32'hb7fb2924),
	.w6(32'hb9968783),
	.w7(32'hba0cd529),
	.w8(32'hb7eedf86),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b40e7f),
	.w1(32'hbad94072),
	.w2(32'hbb11f0b1),
	.w3(32'h3ad00ca4),
	.w4(32'hba553594),
	.w5(32'hbb0cfbb0),
	.w6(32'h3b23dedd),
	.w7(32'hb99a513c),
	.w8(32'hba2cf1de),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79b9b75),
	.w1(32'hb71546af),
	.w2(32'hb6993eb4),
	.w3(32'hb79a2e70),
	.w4(32'hb743e81b),
	.w5(32'hb72b2217),
	.w6(32'hb7cc19de),
	.w7(32'hb62b7a47),
	.w8(32'hb7471df4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a090969),
	.w1(32'hb985a1cb),
	.w2(32'hba89ddb4),
	.w3(32'h39a4036c),
	.w4(32'hb9d0030e),
	.w5(32'hba5501de),
	.w6(32'h39d1c3f2),
	.w7(32'hb98d06dc),
	.w8(32'hba4b453d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e5265),
	.w1(32'hbb85edd9),
	.w2(32'hbb8f4de5),
	.w3(32'h3af940b2),
	.w4(32'h3ad6a083),
	.w5(32'hb99f90fc),
	.w6(32'h369f1744),
	.w7(32'hba0c6cac),
	.w8(32'hbab5a417),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1128b5),
	.w1(32'h3acf486e),
	.w2(32'hb928dac2),
	.w3(32'h3b016c9c),
	.w4(32'h3a9a923e),
	.w5(32'hb9d74163),
	.w6(32'h3a9925ec),
	.w7(32'h3a0fcaab),
	.w8(32'hb9e6dbd5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39190933),
	.w1(32'hb8ceec70),
	.w2(32'h380a6d50),
	.w3(32'hb8d92693),
	.w4(32'hba328ef0),
	.w5(32'hb9d6fac8),
	.w6(32'h37947afa),
	.w7(32'hba013a8e),
	.w8(32'hb9abb11c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bbbb9),
	.w1(32'hbb42ed5d),
	.w2(32'hbac911b4),
	.w3(32'hbb0b85b8),
	.w4(32'hbb286e9e),
	.w5(32'hba84e822),
	.w6(32'hba37e35c),
	.w7(32'hba62a191),
	.w8(32'h39b86ced),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad3686),
	.w1(32'h3a4064d1),
	.w2(32'h3a810c8a),
	.w3(32'h3a00fa9b),
	.w4(32'hb7ae366d),
	.w5(32'h39852be0),
	.w6(32'hb89eb4b6),
	.w7(32'hba378eaf),
	.w8(32'hb9681131),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7fdc),
	.w1(32'h39a2a3f8),
	.w2(32'hba5c9769),
	.w3(32'h3aa1be0b),
	.w4(32'h3a468486),
	.w5(32'hba000216),
	.w6(32'h3a432e90),
	.w7(32'h3a383f56),
	.w8(32'hba7d05db),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e95c7),
	.w1(32'hba922ade),
	.w2(32'hbb4860da),
	.w3(32'hba632d54),
	.w4(32'hbb08eb3c),
	.w5(32'hbb29857a),
	.w6(32'hba87b048),
	.w7(32'hbb4b12e3),
	.w8(32'hbb0be809),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14dadb),
	.w1(32'h3ab255d8),
	.w2(32'hba1fcfd3),
	.w3(32'h3b022817),
	.w4(32'h39caa79a),
	.w5(32'hbaeb1bf5),
	.w6(32'h3a9c009b),
	.w7(32'h397e08bc),
	.w8(32'hbb180b05),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule