module layer_10_featuremap_325(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de529),
	.w1(32'hba522481),
	.w2(32'hbb5bc834),
	.w3(32'hbb0844f8),
	.w4(32'hbb97467a),
	.w5(32'hb91c2078),
	.w6(32'hbad5bd6a),
	.w7(32'hbb99a672),
	.w8(32'hba001375),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75f6f2),
	.w1(32'hb99bb8b5),
	.w2(32'h3a15b762),
	.w3(32'h3aa5d767),
	.w4(32'h3b35accd),
	.w5(32'h3ac38e58),
	.w6(32'hb9f280b7),
	.w7(32'h3b13fae6),
	.w8(32'h39cd27c2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945fd6),
	.w1(32'h3acd7174),
	.w2(32'h3abc4604),
	.w3(32'hbaa05f96),
	.w4(32'hba465d62),
	.w5(32'hba0413ab),
	.w6(32'hb61f9404),
	.w7(32'hba815cec),
	.w8(32'h3917bcc2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950efb3),
	.w1(32'h3ae8e5f5),
	.w2(32'h3afb66dc),
	.w3(32'h3adb07a2),
	.w4(32'h3adee1b3),
	.w5(32'h3a69d63d),
	.w6(32'h3b1144a3),
	.w7(32'h3b25bcec),
	.w8(32'hbbae5dd5),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f03338),
	.w1(32'hbada2116),
	.w2(32'h3890f3b3),
	.w3(32'hba5a4da9),
	.w4(32'h3a10236f),
	.w5(32'h3b038118),
	.w6(32'hbc06e115),
	.w7(32'hbbd1cfef),
	.w8(32'h3aedba67),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48c124),
	.w1(32'h3aa442e4),
	.w2(32'hb9e0eec3),
	.w3(32'h3aea65f6),
	.w4(32'hb9c786ec),
	.w5(32'h3a81d4cc),
	.w6(32'h3a93a887),
	.w7(32'hba90659f),
	.w8(32'h3a0ab4c7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ccdd),
	.w1(32'h3ac0b3c9),
	.w2(32'h3a087e06),
	.w3(32'h39e539a0),
	.w4(32'h3a82cc9c),
	.w5(32'h3a254ece),
	.w6(32'h3a88aeed),
	.w7(32'h39cf74fc),
	.w8(32'h3a2170f5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d6fc7),
	.w1(32'h39572d34),
	.w2(32'hbbe1b45e),
	.w3(32'hbb4103e9),
	.w4(32'hbbf4ad9e),
	.w5(32'hbb8b1aba),
	.w6(32'hba8caecc),
	.w7(32'hbc134153),
	.w8(32'hbb4a98b7),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea7261),
	.w1(32'hbaa11a17),
	.w2(32'hbb199ac6),
	.w3(32'hbaa8f781),
	.w4(32'hbb532cbd),
	.w5(32'h3b285b2d),
	.w6(32'hbb0d1ace),
	.w7(32'hbb7cf13d),
	.w8(32'h3b2ad088),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc37a88),
	.w1(32'h3b5907c3),
	.w2(32'h3b55f697),
	.w3(32'h3ba01b24),
	.w4(32'h3b4b6102),
	.w5(32'h3b8e38f4),
	.w6(32'h3a55b699),
	.w7(32'hba872b5d),
	.w8(32'h3b42b139),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac29c),
	.w1(32'h387439dd),
	.w2(32'hba3a605f),
	.w3(32'hb9e17a4d),
	.w4(32'hbabb3813),
	.w5(32'h3924d62a),
	.w6(32'hb9924925),
	.w7(32'hba923043),
	.w8(32'hb9bb4392),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ed69b),
	.w1(32'h3b2247c4),
	.w2(32'h3a99b8b4),
	.w3(32'hbad7c0d7),
	.w4(32'h3a6c9e61),
	.w5(32'h3aa9d1ed),
	.w6(32'hb964fdfa),
	.w7(32'h3a353dfb),
	.w8(32'hbb3bfb48),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d111ce),
	.w1(32'hbae283f7),
	.w2(32'h3acbd595),
	.w3(32'h3b047e73),
	.w4(32'h3b9c8cc8),
	.w5(32'h3b8d593d),
	.w6(32'hbb3e21f4),
	.w7(32'hba084958),
	.w8(32'h3b8986e7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edbefb),
	.w1(32'hbb814683),
	.w2(32'hbb218f3d),
	.w3(32'hba7cfc55),
	.w4(32'h38627860),
	.w5(32'hbb03d1b9),
	.w6(32'hba98d3fb),
	.w7(32'hb98aaadd),
	.w8(32'hb97a9961),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c1023),
	.w1(32'h3b75a86f),
	.w2(32'h3b5002c6),
	.w3(32'h3b2c1956),
	.w4(32'h3b5e9833),
	.w5(32'h3aae4ab4),
	.w6(32'h3b1f3c8a),
	.w7(32'h3b05e19d),
	.w8(32'h3a142a7f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae142b),
	.w1(32'hba6be960),
	.w2(32'h3b2e7595),
	.w3(32'h3ace5c1b),
	.w4(32'h3b0605b9),
	.w5(32'h3b24b4dd),
	.w6(32'hba34e5eb),
	.w7(32'h379d8459),
	.w8(32'h39ca7cdc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ce2df),
	.w1(32'hb98e73c3),
	.w2(32'hb9877c02),
	.w3(32'h3a5944a3),
	.w4(32'hbaab774e),
	.w5(32'hbaa4432c),
	.w6(32'h38cd8780),
	.w7(32'hbac519b6),
	.w8(32'hbb087061),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcaf2f),
	.w1(32'hbbaf0330),
	.w2(32'hbb9c0d6d),
	.w3(32'hbb6f3362),
	.w4(32'hbbb4bdae),
	.w5(32'hbc049a6b),
	.w6(32'hbba6dabc),
	.w7(32'hbc145bcb),
	.w8(32'hbc26cdf5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3873b8c6),
	.w1(32'h397bd445),
	.w2(32'hb9cfda93),
	.w3(32'hbb37cd23),
	.w4(32'hbb16a6e0),
	.w5(32'hba75a0b5),
	.w6(32'hbb37b92a),
	.w7(32'hbb4ffcb5),
	.w8(32'hbb189b7e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7872d2),
	.w1(32'hbaa97901),
	.w2(32'hba4563d6),
	.w3(32'hba4c662c),
	.w4(32'hb9fd75ea),
	.w5(32'hbad7c841),
	.w6(32'hbac40778),
	.w7(32'hb9939696),
	.w8(32'hbaf24dae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15b377),
	.w1(32'hbb1b813a),
	.w2(32'h3a4099fc),
	.w3(32'hba60c2c3),
	.w4(32'h3a7de0e3),
	.w5(32'hb8d0f43a),
	.w6(32'hbb0ed027),
	.w7(32'h3a8f4003),
	.w8(32'h39b14136),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa422b),
	.w1(32'h3aae6a2b),
	.w2(32'h39bb5cac),
	.w3(32'h3a8cbc5d),
	.w4(32'h395c4375),
	.w5(32'h3a32fac6),
	.w6(32'h3b076814),
	.w7(32'h3aac1eb0),
	.w8(32'h37524daf),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a0c5),
	.w1(32'hbb0041d5),
	.w2(32'hbbaaadc4),
	.w3(32'h3a6e7491),
	.w4(32'hbba1eb69),
	.w5(32'hbbec9417),
	.w6(32'hbb25fbca),
	.w7(32'hbbfa870c),
	.w8(32'hbc57ad71),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ea22),
	.w1(32'h3b28f011),
	.w2(32'h3b8af3a3),
	.w3(32'h3b27993f),
	.w4(32'h3b6f0a69),
	.w5(32'h3af54dba),
	.w6(32'hba898d28),
	.w7(32'h3b0c1bd1),
	.w8(32'h3a3b5c69),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1f831),
	.w1(32'h3ad6a65e),
	.w2(32'h3b843c7f),
	.w3(32'hbab22576),
	.w4(32'h3af19d9b),
	.w5(32'h3bd320d8),
	.w6(32'hbb12766a),
	.w7(32'h3b0fb539),
	.w8(32'h3c171dfd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0cd9),
	.w1(32'h3b32edba),
	.w2(32'h3aa5a335),
	.w3(32'h3b84f4d7),
	.w4(32'h3b2ccdd2),
	.w5(32'h3b29c86e),
	.w6(32'h3b965216),
	.w7(32'h3ac9c9ef),
	.w8(32'h3b0e3924),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b660cfb),
	.w1(32'h3b642c9a),
	.w2(32'h3b80fc05),
	.w3(32'h3b3d545a),
	.w4(32'h3b5f741e),
	.w5(32'h3b4d0efa),
	.w6(32'h3b841be9),
	.w7(32'h3b78bf22),
	.w8(32'h3b2dcb4f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0402),
	.w1(32'hbb0072f2),
	.w2(32'hba34f491),
	.w3(32'hbac8d110),
	.w4(32'hbb1ce106),
	.w5(32'h3b3d3b73),
	.w6(32'hbb17332e),
	.w7(32'hbbb493ed),
	.w8(32'h3b1b8212),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3211bd),
	.w1(32'hb991fe52),
	.w2(32'hb8b68436),
	.w3(32'h39638535),
	.w4(32'hb99f4825),
	.w5(32'hbb0a8cf8),
	.w6(32'hba7053ea),
	.w7(32'h38b31663),
	.w8(32'hba5e907b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b374574),
	.w1(32'h3a47332b),
	.w2(32'h3b06cafc),
	.w3(32'hb9e4c30f),
	.w4(32'hba3a8dde),
	.w5(32'h3a8487fc),
	.w6(32'hbab256de),
	.w7(32'hbaecf818),
	.w8(32'h3b7342c8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45ad08),
	.w1(32'hb8931ceb),
	.w2(32'hb962b9a4),
	.w3(32'hba8ce5de),
	.w4(32'h388d4773),
	.w5(32'hbb04417d),
	.w6(32'hbab4883e),
	.w7(32'h3a6c9f49),
	.w8(32'hbad3b92d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e7f5e),
	.w1(32'h3a5bcdc7),
	.w2(32'h3969d813),
	.w3(32'hba4ce502),
	.w4(32'hba9b6ec3),
	.w5(32'hbb1ca322),
	.w6(32'hb9612ac3),
	.w7(32'h39d0dfc0),
	.w8(32'hbafa583d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391fc1c4),
	.w1(32'h3b49cee1),
	.w2(32'h3bb00f66),
	.w3(32'h3a7507ff),
	.w4(32'h3aa51b34),
	.w5(32'h3a358f67),
	.w6(32'h3b0a5234),
	.w7(32'h3b35b8ad),
	.w8(32'hbaba0eb1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bc9568),
	.w1(32'hba7c10e9),
	.w2(32'h3999ab8a),
	.w3(32'hb92f4af1),
	.w4(32'h39f191e0),
	.w5(32'h39aeb406),
	.w6(32'hbaeaedcf),
	.w7(32'h39cd4f3a),
	.w8(32'h3a9a7881),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65f755),
	.w1(32'hba80a425),
	.w2(32'hb942f94b),
	.w3(32'hb9aab3f2),
	.w4(32'h3a8262a2),
	.w5(32'hbb856f89),
	.w6(32'h386edd4e),
	.w7(32'h3a71e422),
	.w8(32'hbb968799),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb297207),
	.w1(32'hba8d700f),
	.w2(32'h3a73f5c9),
	.w3(32'hbb49d835),
	.w4(32'h398b7fe6),
	.w5(32'hba181a96),
	.w6(32'hbb6846a2),
	.w7(32'h39d24b33),
	.w8(32'hbab13b49),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a494641),
	.w1(32'h3abb1489),
	.w2(32'hbb9aafc5),
	.w3(32'hba966c56),
	.w4(32'hba728199),
	.w5(32'h3be5ca24),
	.w6(32'hba9875b7),
	.w7(32'hba9ae570),
	.w8(32'h3b8f2c4a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d83c2),
	.w1(32'h3bb61eb9),
	.w2(32'h3bf46dd9),
	.w3(32'h3b813686),
	.w4(32'h3b8d5151),
	.w5(32'h3bb0b174),
	.w6(32'h3b7b024c),
	.w7(32'h3baf7c7d),
	.w8(32'h3bbfa5b4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d4af5),
	.w1(32'h3b166ce4),
	.w2(32'h3b8d16d5),
	.w3(32'hbac89a22),
	.w4(32'h3a8ec1f6),
	.w5(32'h3ba4bd27),
	.w6(32'hbb39ec84),
	.w7(32'h3811dbe9),
	.w8(32'h3b9d83f5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b3916),
	.w1(32'h3a941811),
	.w2(32'h3a3bad2b),
	.w3(32'hbad012b1),
	.w4(32'hbb692c5a),
	.w5(32'h3a8ca4c6),
	.w6(32'hbabedc5f),
	.w7(32'hbb15d746),
	.w8(32'h3a96e649),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98897be),
	.w1(32'hbaa060dc),
	.w2(32'hba848373),
	.w3(32'hba273e8b),
	.w4(32'hba6841ff),
	.w5(32'h3b9be413),
	.w6(32'hba53f167),
	.w7(32'hbaa32c2e),
	.w8(32'h3b840901),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f8e2),
	.w1(32'h3b6b08de),
	.w2(32'h3acef632),
	.w3(32'h3b9be2cf),
	.w4(32'h3b3dfdda),
	.w5(32'hbb260ea4),
	.w6(32'h3b8a5f1e),
	.w7(32'h3a25cabd),
	.w8(32'hbb1256fb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf99ca),
	.w1(32'hbb029473),
	.w2(32'hbac31ef0),
	.w3(32'hbb6b2235),
	.w4(32'hbaa5ed0c),
	.w5(32'hbb4fba43),
	.w6(32'hbb4efe40),
	.w7(32'hba497e73),
	.w8(32'hbb2cb37a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa089bb),
	.w1(32'h3a1088e9),
	.w2(32'h3b90b954),
	.w3(32'hba664296),
	.w4(32'h39e727e0),
	.w5(32'h39907517),
	.w6(32'hbb9f686c),
	.w7(32'hbb81514e),
	.w8(32'hbaf64e6b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91396d),
	.w1(32'h3be598fc),
	.w2(32'h3bd41b5a),
	.w3(32'h3b0e11d3),
	.w4(32'h3aa92054),
	.w5(32'h3bc74c1c),
	.w6(32'h3b0a56b5),
	.w7(32'h3ae36fe7),
	.w8(32'h3bbc6269),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46047b),
	.w1(32'h3b858f86),
	.w2(32'h3b7d5591),
	.w3(32'h3b824db4),
	.w4(32'h3b353e1a),
	.w5(32'h3bc1192f),
	.w6(32'h3a0bc679),
	.w7(32'h39333453),
	.w8(32'h3bc538ea),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40a27e),
	.w1(32'h3b3cb50d),
	.w2(32'h3a9d8c5e),
	.w3(32'h3b36ae7d),
	.w4(32'h3aa2e64c),
	.w5(32'h3b64b4d3),
	.w6(32'h3b346ac3),
	.w7(32'h3a1141ae),
	.w8(32'h3ad1c0d1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae82934),
	.w1(32'hbb009d4b),
	.w2(32'hbbb26cad),
	.w3(32'h3b40738c),
	.w4(32'hbb054e31),
	.w5(32'hbbe97c22),
	.w6(32'h3b1d0e53),
	.w7(32'hbb905410),
	.w8(32'hbc3b6d76),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6b97a),
	.w1(32'hba0812c1),
	.w2(32'h3a2b2af9),
	.w3(32'hb939ddbb),
	.w4(32'h3af16e8b),
	.w5(32'h3abc5c91),
	.w6(32'hbaeeb182),
	.w7(32'h391372d5),
	.w8(32'h3a97e267),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b542ba7),
	.w1(32'h3b16b8c4),
	.w2(32'h39ab547f),
	.w3(32'h3ae40578),
	.w4(32'h3a48d2df),
	.w5(32'h3bee7597),
	.w6(32'h3b1d5e51),
	.w7(32'hb99b20bc),
	.w8(32'h3bf24bd5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba01c7c),
	.w1(32'hbb7c9e61),
	.w2(32'hba8321f3),
	.w3(32'hba927eed),
	.w4(32'hb9a1b5f9),
	.w5(32'hb9b4e50a),
	.w6(32'hbb7039dc),
	.w7(32'hba902d7c),
	.w8(32'hba76157e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0c5b6),
	.w1(32'hba35d7e1),
	.w2(32'hb8fd5d74),
	.w3(32'hbaec86aa),
	.w4(32'hba7b0828),
	.w5(32'h3a98264b),
	.w6(32'hbb883da3),
	.w7(32'hbb599cbc),
	.w8(32'h3a546083),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a892787),
	.w1(32'h3a6c5fbd),
	.w2(32'hbaf00ef5),
	.w3(32'hb97e2586),
	.w4(32'hbb2667fc),
	.w5(32'h3b8b4821),
	.w6(32'h3a1b5204),
	.w7(32'hbb0de555),
	.w8(32'h3b16fe03),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d0a13),
	.w1(32'h3a18e2c5),
	.w2(32'hbb019f42),
	.w3(32'h3b024d33),
	.w4(32'hbaeefe18),
	.w5(32'hbbaab2c9),
	.w6(32'h3a2d81df),
	.w7(32'hbba283da),
	.w8(32'hbbea8a60),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf424a2),
	.w1(32'hbad75c17),
	.w2(32'hbae1aede),
	.w3(32'hba785a65),
	.w4(32'h3965d7b1),
	.w5(32'h390849b8),
	.w6(32'hbb095de6),
	.w7(32'hba5d40b2),
	.w8(32'hba0dba88),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a999dff),
	.w1(32'hbad0ba9c),
	.w2(32'hba2f5c64),
	.w3(32'hb9e36893),
	.w4(32'h3a027bcf),
	.w5(32'hb94c1843),
	.w6(32'hbafae724),
	.w7(32'h388de8e4),
	.w8(32'hba21f10a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab4e24),
	.w1(32'hba600083),
	.w2(32'hb990388e),
	.w3(32'hb98988dd),
	.w4(32'h39c03430),
	.w5(32'h3b2c4ee8),
	.w6(32'hba2b160a),
	.w7(32'h392ecda7),
	.w8(32'h3b31eab0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39333f),
	.w1(32'hba0b3815),
	.w2(32'hba20a37d),
	.w3(32'hba296dd6),
	.w4(32'hba882c95),
	.w5(32'h3b20b1d5),
	.w6(32'hba636ed5),
	.w7(32'hb9b4042d),
	.w8(32'h3b1dd977),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3669ce),
	.w1(32'h3a81efe7),
	.w2(32'hba48de5c),
	.w3(32'h3a9870ad),
	.w4(32'h393a849d),
	.w5(32'h3a1b66fd),
	.w6(32'h3af94a55),
	.w7(32'hba3d59fc),
	.w8(32'hbaae0308),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e9b28),
	.w1(32'h3a90b71a),
	.w2(32'hbad839d4),
	.w3(32'h3a003564),
	.w4(32'hbac13172),
	.w5(32'hbaebab55),
	.w6(32'h388cd79e),
	.w7(32'hbb55d0a1),
	.w8(32'hbae702b0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b0c8f),
	.w1(32'hbaf86aad),
	.w2(32'hbb287c2d),
	.w3(32'hbb086aad),
	.w4(32'hbac1ca43),
	.w5(32'h3b42ffcf),
	.w6(32'hbb61ab89),
	.w7(32'hbb6e1528),
	.w8(32'h3ace2078),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02fb2c),
	.w1(32'hb936cdd6),
	.w2(32'hbaeaefd5),
	.w3(32'h3b3a1409),
	.w4(32'hb85526ee),
	.w5(32'hbb1baf91),
	.w6(32'h3aadaa6e),
	.w7(32'hbb320649),
	.w8(32'hbbd565f5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35ecd),
	.w1(32'hba4fc294),
	.w2(32'hba511065),
	.w3(32'h3adcd821),
	.w4(32'h3b1e6db8),
	.w5(32'h3b34b048),
	.w6(32'hbb0bf682),
	.w7(32'hbb064ed0),
	.w8(32'h3b09d3cc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1abc0f),
	.w1(32'hb9015705),
	.w2(32'hba1bbf09),
	.w3(32'h3a3c16b7),
	.w4(32'h3905a36e),
	.w5(32'h3a9c9a30),
	.w6(32'h39b17e53),
	.w7(32'hb9b6762d),
	.w8(32'h3ac2045d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab67d68),
	.w1(32'hb9935c6d),
	.w2(32'hbafbb767),
	.w3(32'hba137450),
	.w4(32'hba9676d3),
	.w5(32'hb845d2c2),
	.w6(32'hba83e2f0),
	.w7(32'hbaa1637a),
	.w8(32'hbaf936ad),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47bd9d),
	.w1(32'h37bfb365),
	.w2(32'hb947f80c),
	.w3(32'h3aa26a16),
	.w4(32'h3b10d447),
	.w5(32'hba929db9),
	.w6(32'hbaf8aa3f),
	.w7(32'hba919af7),
	.w8(32'hb8ee417c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f349c),
	.w1(32'h3b2334dd),
	.w2(32'h36e30c80),
	.w3(32'h3813a3d0),
	.w4(32'h3b0a5162),
	.w5(32'h3b85fbfe),
	.w6(32'hb76023a8),
	.w7(32'hbb198f59),
	.w8(32'hba5cb426),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dd927),
	.w1(32'h3ac7eedc),
	.w2(32'h3bc39afb),
	.w3(32'h3b612dbc),
	.w4(32'h3bdbf7d7),
	.w5(32'h3b9746ad),
	.w6(32'h3a8b2385),
	.w7(32'h3bce1cde),
	.w8(32'h3b94af00),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0cf5c),
	.w1(32'hbb00d198),
	.w2(32'hb943b19f),
	.w3(32'hbb5ad9e8),
	.w4(32'hba1a03c0),
	.w5(32'hbc172a07),
	.w6(32'hbb42f1a6),
	.w7(32'hb9edb7b3),
	.w8(32'hbc304230),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac92c0b),
	.w1(32'h3b17b132),
	.w2(32'h3ba8b899),
	.w3(32'hba9e8838),
	.w4(32'h3b297b6e),
	.w5(32'h3bc3a689),
	.w6(32'hbb8b7bd1),
	.w7(32'h38a2bd22),
	.w8(32'h3c024a22),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41eb76),
	.w1(32'h3afb4278),
	.w2(32'h3adae0bc),
	.w3(32'hb9569896),
	.w4(32'h3a8367b4),
	.w5(32'hba91a454),
	.w6(32'h3a84d9db),
	.w7(32'h3aa1aebd),
	.w8(32'hba6249f9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ecced),
	.w1(32'hb799eb3e),
	.w2(32'h3a683337),
	.w3(32'hb971fbd3),
	.w4(32'h39017f1c),
	.w5(32'h3832fa9f),
	.w6(32'hba31896b),
	.w7(32'hb9e69d1f),
	.w8(32'hba2b6077),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae278a2),
	.w1(32'hbabce2f9),
	.w2(32'hba3279e0),
	.w3(32'hb8d81d8e),
	.w4(32'hb9fb8c82),
	.w5(32'h3ac1b209),
	.w6(32'hbb03e182),
	.w7(32'hba834a95),
	.w8(32'h3a4d60d9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6062a3),
	.w1(32'hba59be2b),
	.w2(32'hba9c1c43),
	.w3(32'h39053605),
	.w4(32'h37cf9144),
	.w5(32'hba1f4bba),
	.w6(32'hbae47b68),
	.w7(32'hbb09d708),
	.w8(32'h39f51134),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf9d2),
	.w1(32'h3aa92c77),
	.w2(32'h3ac2e754),
	.w3(32'hba048638),
	.w4(32'hb93831d8),
	.w5(32'hb98c989b),
	.w6(32'h39eb4ce7),
	.w7(32'h3a6e1917),
	.w8(32'hbadf164d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b37f1),
	.w1(32'hbafce487),
	.w2(32'hbad683ca),
	.w3(32'hbaaaed62),
	.w4(32'hba0179db),
	.w5(32'hbad0eab1),
	.w6(32'hbb5f2a3e),
	.w7(32'hbb319f3c),
	.w8(32'hbb726dbd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81adb7),
	.w1(32'hbab09ac7),
	.w2(32'hbb4e9535),
	.w3(32'hbb3fb66f),
	.w4(32'hbb487a27),
	.w5(32'hbbb4be85),
	.w6(32'hbb00b59b),
	.w7(32'hbbce1f1d),
	.w8(32'hbbecf050),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cd3d8),
	.w1(32'hba113c65),
	.w2(32'h3a80469a),
	.w3(32'hbb236a1d),
	.w4(32'hba9f9a9e),
	.w5(32'h3b4d7867),
	.w6(32'hbb8a5459),
	.w7(32'hbadb2872),
	.w8(32'h3b642a24),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b189d8d),
	.w1(32'h3a52ab0d),
	.w2(32'hb9043ce6),
	.w3(32'hb982146c),
	.w4(32'hba6b4e66),
	.w5(32'hb98859be),
	.w6(32'hbaa8e227),
	.w7(32'hbb25a2fc),
	.w8(32'hbabc0cc8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabccd4),
	.w1(32'h39a86c8b),
	.w2(32'hba5063b0),
	.w3(32'h3a6eb4aa),
	.w4(32'h3a7ee109),
	.w5(32'h3afa8276),
	.w6(32'hba6dad42),
	.w7(32'hbb0215f8),
	.w8(32'h3a05fcd2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae55d29),
	.w1(32'h3b1e9603),
	.w2(32'h3b3808b9),
	.w3(32'h3b545151),
	.w4(32'h3b90c26a),
	.w5(32'hba026de7),
	.w6(32'h3b3e0daf),
	.w7(32'h3b662c43),
	.w8(32'hba82262f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab69770),
	.w1(32'hbb15d3db),
	.w2(32'hbb07ea3c),
	.w3(32'hbb2e618f),
	.w4(32'hbad74f04),
	.w5(32'hba0d6fcd),
	.w6(32'hbb856f50),
	.w7(32'hbb794242),
	.w8(32'hbaf748fd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9b9d6),
	.w1(32'h3ab88a01),
	.w2(32'h3a519fd0),
	.w3(32'hb7354f86),
	.w4(32'h396bf7b6),
	.w5(32'h3b321d63),
	.w6(32'h3a9f8d46),
	.w7(32'h3aa5c609),
	.w8(32'h3b1cfa61),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060ba8),
	.w1(32'h3bd493ce),
	.w2(32'h3c05f416),
	.w3(32'h3bce2176),
	.w4(32'h3bab86a3),
	.w5(32'hba1225c3),
	.w6(32'h3bc11272),
	.w7(32'h3bf9ea64),
	.w8(32'hbaed176e),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba327be7),
	.w1(32'h38bcbe64),
	.w2(32'hba0aef73),
	.w3(32'hba8324ad),
	.w4(32'hba6d12e5),
	.w5(32'h3b0a477f),
	.w6(32'hba1d37b6),
	.w7(32'hba5ccf16),
	.w8(32'h3b2950cc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0296),
	.w1(32'h3b05b041),
	.w2(32'hba81bad3),
	.w3(32'h3a964e0b),
	.w4(32'h39d76e0a),
	.w5(32'h3baf3c2d),
	.w6(32'h39eea2a1),
	.w7(32'hbab3bd50),
	.w8(32'h3bace9c3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e6551),
	.w1(32'h3ba7aed0),
	.w2(32'h3b1bcfaf),
	.w3(32'h3b0ac776),
	.w4(32'h3ab848bd),
	.w5(32'h3b99f6a7),
	.w6(32'h3b63beb5),
	.w7(32'h3a29409a),
	.w8(32'h3b6e2713),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a8a88),
	.w1(32'h3a335bc2),
	.w2(32'h39458c3e),
	.w3(32'h3b176ac0),
	.w4(32'h3b30c657),
	.w5(32'h3a48645f),
	.w6(32'h3a42db56),
	.w7(32'h39e33c50),
	.w8(32'hb9486e95),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c0b3c),
	.w1(32'h3b0e5703),
	.w2(32'h3a829802),
	.w3(32'h3b31cd71),
	.w4(32'h3a2b632b),
	.w5(32'hba3d0b6a),
	.w6(32'h38e327f4),
	.w7(32'hb965b9ae),
	.w8(32'hb96a2eee),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab79883),
	.w1(32'hbb7d451c),
	.w2(32'hbbd0eb51),
	.w3(32'hbb659c78),
	.w4(32'hbbcf2e21),
	.w5(32'hbbf9d093),
	.w6(32'hbb83203e),
	.w7(32'hbc1d0578),
	.w8(32'hbc207bd1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840f8b),
	.w1(32'hb9f0751e),
	.w2(32'h3ac07f04),
	.w3(32'h3a254f13),
	.w4(32'h3a9584d8),
	.w5(32'h37c277a7),
	.w6(32'hb95d21a0),
	.w7(32'h3a5162c8),
	.w8(32'h3a97b54a),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962fb2),
	.w1(32'h3a027f58),
	.w2(32'hbaaf9aed),
	.w3(32'h3ad18f6d),
	.w4(32'h3b045f64),
	.w5(32'h3b1411b3),
	.w6(32'h3b29a2c3),
	.w7(32'h3a3fd2df),
	.w8(32'hbb237bdd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ab45e),
	.w1(32'h3ba5c095),
	.w2(32'h3c021397),
	.w3(32'h3ae5532a),
	.w4(32'h3ba8bebe),
	.w5(32'h3ae26799),
	.w6(32'h3a116820),
	.w7(32'h3b744d7f),
	.w8(32'h3adf9304),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25d265),
	.w1(32'h3ba89864),
	.w2(32'h3b684275),
	.w3(32'h3a375a8e),
	.w4(32'h3b24bf0f),
	.w5(32'h3b360c98),
	.w6(32'hbb4c2f84),
	.w7(32'hbac3643e),
	.w8(32'h3b6305d0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b79d5),
	.w1(32'h3aa3500a),
	.w2(32'h3b174932),
	.w3(32'h3af90dff),
	.w4(32'h3b17bfa4),
	.w5(32'h3b209c81),
	.w6(32'h3a8a03d3),
	.w7(32'h3a5b1047),
	.w8(32'hbaabb12b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a3886),
	.w1(32'h3b44248e),
	.w2(32'h3b7e36bb),
	.w3(32'h39ed3468),
	.w4(32'h3ad79d65),
	.w5(32'h3b9b4ff5),
	.w6(32'hba94d649),
	.w7(32'h3b1283f5),
	.w8(32'h3b9f6e5d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1369ca),
	.w1(32'h3a86b2af),
	.w2(32'h38f40324),
	.w3(32'h3a60ee85),
	.w4(32'hb9f503c2),
	.w5(32'h3a8d7fe2),
	.w6(32'h39caf7da),
	.w7(32'h39299926),
	.w8(32'h3ad50755),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3063c),
	.w1(32'h3bd118de),
	.w2(32'h3c087316),
	.w3(32'h3ba09f48),
	.w4(32'h3bbd4de0),
	.w5(32'hb8bc004a),
	.w6(32'h3b2b4596),
	.w7(32'h3b6a63cd),
	.w8(32'hbb6ef3df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae71fce),
	.w1(32'h39b627ad),
	.w2(32'h3abcd0b9),
	.w3(32'hbafa08c3),
	.w4(32'h3b5f78e1),
	.w5(32'h3bac9417),
	.w6(32'hbb1a0af8),
	.w7(32'h3aca41fe),
	.w8(32'h3b752d11),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39781076),
	.w1(32'hbac86b0f),
	.w2(32'hbc034f95),
	.w3(32'hbac8103a),
	.w4(32'hbacea173),
	.w5(32'hbb755fc4),
	.w6(32'hbb14f280),
	.w7(32'hbb03df3a),
	.w8(32'hbb9c8b5b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1aefbe),
	.w1(32'h3b401a1d),
	.w2(32'hba9b2d94),
	.w3(32'h3b0ccc85),
	.w4(32'hba45c460),
	.w5(32'h3a9a3ddf),
	.w6(32'hba43b68a),
	.w7(32'h3abdba09),
	.w8(32'h3ada8fbc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b23aa),
	.w1(32'h397b5755),
	.w2(32'h3bad9333),
	.w3(32'h3ad00ad2),
	.w4(32'h393604d4),
	.w5(32'h3be6a3e2),
	.w6(32'hbb31e112),
	.w7(32'h39b24ab0),
	.w8(32'h3be2aaa3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee5618),
	.w1(32'hbb47a08b),
	.w2(32'hbb9198d1),
	.w3(32'h3a251bfe),
	.w4(32'h38b114d8),
	.w5(32'h3af7e391),
	.w6(32'hbac2c228),
	.w7(32'hbb898f2a),
	.w8(32'hbbc382cb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edadbc),
	.w1(32'hba929f81),
	.w2(32'hb970cd72),
	.w3(32'h39e695d4),
	.w4(32'h3ab53d50),
	.w5(32'h3ab3262a),
	.w6(32'h393c17dd),
	.w7(32'hbad25f94),
	.w8(32'h3b0727ae),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eae926),
	.w1(32'h3b308cd3),
	.w2(32'hbaf9fa99),
	.w3(32'h3bb0a254),
	.w4(32'h3b8aaffe),
	.w5(32'hbb261677),
	.w6(32'h3b9a4d2a),
	.w7(32'h3ac85f3b),
	.w8(32'hbba6ee22),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9b817),
	.w1(32'h3b4b1ce5),
	.w2(32'h3a0aa83e),
	.w3(32'hb9b18c5c),
	.w4(32'h37b2e39f),
	.w5(32'h3bcd9e48),
	.w6(32'h3b3d47e3),
	.w7(32'h38512e7c),
	.w8(32'h3b67d361),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab2d28),
	.w1(32'h3ae70f2a),
	.w2(32'h3aa5f214),
	.w3(32'h3b351303),
	.w4(32'h3b479da3),
	.w5(32'hbb5ef557),
	.w6(32'h3b45586b),
	.w7(32'hba728790),
	.w8(32'hbb00499e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cc819),
	.w1(32'hbb438380),
	.w2(32'hbaf660e9),
	.w3(32'hbb40b0b3),
	.w4(32'hbb1ad200),
	.w5(32'hbb0bc993),
	.w6(32'hbbab38a5),
	.w7(32'hbb287f8e),
	.w8(32'hbb2a37bd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c8d3),
	.w1(32'hbb1a0f0b),
	.w2(32'h3b85c96f),
	.w3(32'hbb4a5f4e),
	.w4(32'h3ab48ee3),
	.w5(32'h3a40507b),
	.w6(32'hbba4ec9c),
	.w7(32'hbab8fca8),
	.w8(32'hba724000),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a4b1),
	.w1(32'h3b419bba),
	.w2(32'h3bd0ffc0),
	.w3(32'h3b2127a8),
	.w4(32'h3ba7b5c4),
	.w5(32'h3ba2ca93),
	.w6(32'hbab59d38),
	.w7(32'h3b5f7241),
	.w8(32'h3b99579d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa39fb4),
	.w1(32'hb9fc183b),
	.w2(32'hbb004fb1),
	.w3(32'h3981c538),
	.w4(32'hba48acfe),
	.w5(32'hba09d5c3),
	.w6(32'hbb26da47),
	.w7(32'hbb807730),
	.w8(32'hbb1b299a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38c1e7),
	.w1(32'h3aa87989),
	.w2(32'h3b924f96),
	.w3(32'h3a47e47e),
	.w4(32'h3b0d1051),
	.w5(32'hbb00a9c2),
	.w6(32'hbadb7af5),
	.w7(32'h3b2a0ed0),
	.w8(32'hbb6745d4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a5e73),
	.w1(32'hb9bb94ce),
	.w2(32'h39d38a14),
	.w3(32'hba300e0f),
	.w4(32'h3aa53d4c),
	.w5(32'hb9c28344),
	.w6(32'hbb18982a),
	.w7(32'h3b2f7c8b),
	.w8(32'hb924df86),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945aaa),
	.w1(32'hbbcd1236),
	.w2(32'hbbaf1b02),
	.w3(32'h3b03fc81),
	.w4(32'h39b90340),
	.w5(32'h3b56b717),
	.w6(32'hb9e98b57),
	.w7(32'hbab303da),
	.w8(32'hba1368d5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf69a2),
	.w1(32'h3a9c618d),
	.w2(32'h3b203a54),
	.w3(32'hba57e123),
	.w4(32'h3a960588),
	.w5(32'hb90a16f2),
	.w6(32'h3a910009),
	.w7(32'hbac6422e),
	.w8(32'hba9db185),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb179ba2),
	.w1(32'hbb14ae85),
	.w2(32'hb8da71ed),
	.w3(32'hbb0efb53),
	.w4(32'hba21876e),
	.w5(32'hbb093ef1),
	.w6(32'hbb26c03f),
	.w7(32'hbaa8a75b),
	.w8(32'hb96857f2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99565e2),
	.w1(32'hba117a40),
	.w2(32'hb9f51789),
	.w3(32'hbb09611f),
	.w4(32'hbafc2645),
	.w5(32'hbaf2e4ee),
	.w6(32'hbac0ad5e),
	.w7(32'hbada4b74),
	.w8(32'hbb3e3d2f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f0c2),
	.w1(32'hbb608f12),
	.w2(32'h3aa55a68),
	.w3(32'hb88a5486),
	.w4(32'h3b0ab795),
	.w5(32'hbb1b9a34),
	.w6(32'h3a6d1c79),
	.w7(32'h39f327c4),
	.w8(32'h39aa3768),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2ed14),
	.w1(32'hbb2a6027),
	.w2(32'hbaca4ada),
	.w3(32'hbb21f372),
	.w4(32'hbad7f3ce),
	.w5(32'hbb8ae5da),
	.w6(32'hbb0c55b7),
	.w7(32'hba4e5cb7),
	.w8(32'hbbcaa45b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c346),
	.w1(32'hbbbac1dd),
	.w2(32'hbad3ae31),
	.w3(32'hbbc40173),
	.w4(32'hba1d1b23),
	.w5(32'h3b06e938),
	.w6(32'hbbd14df5),
	.w7(32'hbb0a37ca),
	.w8(32'h3a93d844),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6f5c),
	.w1(32'hbaa2c3ef),
	.w2(32'h3a4e026a),
	.w3(32'hb7dbe56a),
	.w4(32'hba228ff1),
	.w5(32'h3b6b9aee),
	.w6(32'hbb303cc4),
	.w7(32'hb988b950),
	.w8(32'h3b7d9b2c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e2a0a),
	.w1(32'h3936ce9f),
	.w2(32'h3b92060a),
	.w3(32'h3a13e48e),
	.w4(32'h3b3bbe14),
	.w5(32'h3b6ded08),
	.w6(32'hb88b9e38),
	.w7(32'h3b0089d9),
	.w8(32'hbb3ceb7a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bdc84),
	.w1(32'h3b882a1f),
	.w2(32'h3b23ffac),
	.w3(32'h3ae06219),
	.w4(32'h3ba679a3),
	.w5(32'hbb1f16ec),
	.w6(32'h3b16f42a),
	.w7(32'h3be0074e),
	.w8(32'hb96f3dfd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399837fe),
	.w1(32'hbace1276),
	.w2(32'hb9b97ce0),
	.w3(32'hbbb818d5),
	.w4(32'hbb1bfa1f),
	.w5(32'h3b97f4df),
	.w6(32'hbb9bf068),
	.w7(32'hbb4e8b79),
	.w8(32'h3b8e10f3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa07ba),
	.w1(32'h3b63254e),
	.w2(32'h3b9ecbfe),
	.w3(32'h3b799958),
	.w4(32'h3b6899de),
	.w5(32'hbaaac21d),
	.w6(32'h3b836f86),
	.w7(32'h3bafa591),
	.w8(32'hbb18af45),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60bc10),
	.w1(32'hbb9290f1),
	.w2(32'hb92a5159),
	.w3(32'h3b08a45f),
	.w4(32'h3b8e8dbe),
	.w5(32'hbaf79af2),
	.w6(32'hbae37111),
	.w7(32'h3b5a9db3),
	.w8(32'h3aa23cdf),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00ebc8),
	.w1(32'hba60a241),
	.w2(32'h3a33a1ab),
	.w3(32'hbad8ef69),
	.w4(32'h38aba62b),
	.w5(32'h39c63198),
	.w6(32'hbabfe99c),
	.w7(32'h3ac4e470),
	.w8(32'hb7575906),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135c47),
	.w1(32'hbb120058),
	.w2(32'h39fdb63d),
	.w3(32'h3ad386ea),
	.w4(32'h3b531fa2),
	.w5(32'hbadf00b0),
	.w6(32'h3b297d29),
	.w7(32'h3b80e53e),
	.w8(32'hbb3728da),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919c0d6),
	.w1(32'h3852c766),
	.w2(32'h3ae38e2f),
	.w3(32'h3ad28619),
	.w4(32'h3a070df8),
	.w5(32'h3b1ef0a0),
	.w6(32'hb99d0d97),
	.w7(32'hbac4084f),
	.w8(32'hb88ae7bf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7557a8),
	.w1(32'h3a7d99ca),
	.w2(32'h39e7880e),
	.w3(32'hba240083),
	.w4(32'hba8cba2a),
	.w5(32'hbba7f421),
	.w6(32'h3ae8d388),
	.w7(32'h3a227a13),
	.w8(32'hbaca5890),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57b5b3),
	.w1(32'hbb29b062),
	.w2(32'hbb7517cf),
	.w3(32'hbbb6a671),
	.w4(32'hbb9cb27b),
	.w5(32'h3b1097eb),
	.w6(32'h3b25ce84),
	.w7(32'hbb64b372),
	.w8(32'h3abce6c7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1d785),
	.w1(32'h3b0fbd89),
	.w2(32'h3b5ddda2),
	.w3(32'h3add59d1),
	.w4(32'h3b8c7685),
	.w5(32'hb959804f),
	.w6(32'hbb87d90b),
	.w7(32'h3b11fa1d),
	.w8(32'hbacb501d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079b0f),
	.w1(32'hbb493274),
	.w2(32'hb9bed73c),
	.w3(32'hbb010161),
	.w4(32'hbb063cdd),
	.w5(32'h3a8e02bd),
	.w6(32'hbb8b1c77),
	.w7(32'hbb494538),
	.w8(32'h3a97f6e6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae91987),
	.w1(32'h3a86a0f6),
	.w2(32'h3b071ec5),
	.w3(32'h3a79e608),
	.w4(32'h3b5c58e6),
	.w5(32'h3b44e8cc),
	.w6(32'hbaf7f217),
	.w7(32'h3b06c8b1),
	.w8(32'h3bdb51e2),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1a25e),
	.w1(32'h3b1e0320),
	.w2(32'h3b3908d8),
	.w3(32'h3af9d986),
	.w4(32'h3ad4a1b5),
	.w5(32'hbb493673),
	.w6(32'h3b5e61ce),
	.w7(32'h3abf94a9),
	.w8(32'hbbcbfbc5),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae00687),
	.w1(32'hba7f91b0),
	.w2(32'h3b511890),
	.w3(32'h39d2839b),
	.w4(32'h3a04f9bf),
	.w5(32'hb9d1b54d),
	.w6(32'hbb538a0b),
	.w7(32'h3a071885),
	.w8(32'h39cca8ab),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e9d2f),
	.w1(32'hbb2c443b),
	.w2(32'hba2c78c4),
	.w3(32'hbad2aac6),
	.w4(32'hbb06caee),
	.w5(32'h3ae889c0),
	.w6(32'hbbaa0258),
	.w7(32'hbb18df01),
	.w8(32'h3acc5022),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba29c77),
	.w1(32'h3acb2f5c),
	.w2(32'h3922623c),
	.w3(32'h3a326d6a),
	.w4(32'h3b09bdcf),
	.w5(32'h3b2be3b8),
	.w6(32'hbac93809),
	.w7(32'h3961b07a),
	.w8(32'h3ae70452),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20c637),
	.w1(32'h3ac4afac),
	.w2(32'h3b7c250b),
	.w3(32'h3b8bd803),
	.w4(32'h3ba56ef1),
	.w5(32'h3b8f2fd1),
	.w6(32'hb9d607bb),
	.w7(32'h3bae8300),
	.w8(32'h3b9ccc8c),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bab73),
	.w1(32'h3ae2d325),
	.w2(32'h3a20507e),
	.w3(32'h3bbf8d16),
	.w4(32'h3b49c1b3),
	.w5(32'hba5b2bc1),
	.w6(32'h3bb0947f),
	.w7(32'hbb373d5c),
	.w8(32'hbbbb47a6),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a46e2),
	.w1(32'hbaef4d91),
	.w2(32'hbb5fc84d),
	.w3(32'hbad52c43),
	.w4(32'hbb15c0d4),
	.w5(32'h3b09b80e),
	.w6(32'hbb7811c4),
	.w7(32'hbb8d3435),
	.w8(32'hba89009b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39269d33),
	.w1(32'h3b6ff8df),
	.w2(32'h3c08fef4),
	.w3(32'h3ba988a6),
	.w4(32'h3bcdd7e0),
	.w5(32'h3c01f486),
	.w6(32'h3b2fb9e0),
	.w7(32'h3b9f194a),
	.w8(32'h3c0e9752),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce7c70),
	.w1(32'h3b4813df),
	.w2(32'h3aab5c1e),
	.w3(32'h3b2af0fe),
	.w4(32'h3b0e50ac),
	.w5(32'hba80a83c),
	.w6(32'hba709551),
	.w7(32'h367894a7),
	.w8(32'hbb8ecedd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64f18c),
	.w1(32'hbaaf76eb),
	.w2(32'hbb16f37e),
	.w3(32'h3a8cfbc3),
	.w4(32'h3b32a3d9),
	.w5(32'h39963361),
	.w6(32'hbb61926d),
	.w7(32'hbaf5f733),
	.w8(32'h3aa30928),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0be4a),
	.w1(32'h3a874c31),
	.w2(32'h3aa22ddf),
	.w3(32'hb9cf8256),
	.w4(32'h3a67a4b6),
	.w5(32'hba19c296),
	.w6(32'hba1b0977),
	.w7(32'h3aeabd79),
	.w8(32'hb9d4dbae),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b8c8),
	.w1(32'hbadd3ecb),
	.w2(32'hbaab2223),
	.w3(32'hbb5b7daa),
	.w4(32'hbaa5e919),
	.w5(32'h3abe633b),
	.w6(32'hba0c8680),
	.w7(32'hbab3990d),
	.w8(32'hb91aea59),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f59aba),
	.w1(32'hbb0fc0f3),
	.w2(32'hba8fae81),
	.w3(32'hbabebd43),
	.w4(32'h3a9b19bd),
	.w5(32'hb9478063),
	.w6(32'hbb79a278),
	.w7(32'hba9b5c5f),
	.w8(32'hbb2b0a6f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee31b),
	.w1(32'hbb2524e8),
	.w2(32'h3aa54727),
	.w3(32'h3a8f0b3a),
	.w4(32'h3bd02e7e),
	.w5(32'hbb0da0d5),
	.w6(32'hbb0f666e),
	.w7(32'h3b798709),
	.w8(32'hbb1148fe),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1194be),
	.w1(32'hbb125da1),
	.w2(32'hbb4848f4),
	.w3(32'h3a837fab),
	.w4(32'h3a851dce),
	.w5(32'h38609ce3),
	.w6(32'hbb341e3e),
	.w7(32'hbb4cf2a5),
	.w8(32'h3ad8a9f9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7638e),
	.w1(32'h3b976066),
	.w2(32'h3baa121e),
	.w3(32'h3a8fb572),
	.w4(32'h3b06c93f),
	.w5(32'h3b8564b0),
	.w6(32'h3767e286),
	.w7(32'h3ac9071d),
	.w8(32'h3b72514b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace64d1),
	.w1(32'hbb3f3ea7),
	.w2(32'hba5591c5),
	.w3(32'h3b03fe78),
	.w4(32'h3a523a41),
	.w5(32'h3bf92685),
	.w6(32'h3ab86ad2),
	.w7(32'hba8971f5),
	.w8(32'h3be54201),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b369af4),
	.w1(32'h3a70cea6),
	.w2(32'h3a365a2e),
	.w3(32'h3bd05abe),
	.w4(32'h3b6dd7d0),
	.w5(32'hbae3af1c),
	.w6(32'h3b0f966b),
	.w7(32'h396a32e0),
	.w8(32'hb9f574c6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add54e5),
	.w1(32'h3ad26383),
	.w2(32'h3ba64355),
	.w3(32'h3a078996),
	.w4(32'h39fe806c),
	.w5(32'hb9c946dc),
	.w6(32'h3aa3be8d),
	.w7(32'h3a43940b),
	.w8(32'h3ac91d26),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08f491),
	.w1(32'hba1a7e9a),
	.w2(32'hbab92dcc),
	.w3(32'hba667570),
	.w4(32'h394a2b91),
	.w5(32'hbad3109f),
	.w6(32'hbb72075f),
	.w7(32'hb9d0894a),
	.w8(32'hbabebb7a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac648c),
	.w1(32'hbafe3806),
	.w2(32'hba1b2fef),
	.w3(32'hbb2c2a54),
	.w4(32'h37a3ee7b),
	.w5(32'hbb548887),
	.w6(32'hbbae1623),
	.w7(32'hba8b7de4),
	.w8(32'hbb22f943),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b79610),
	.w1(32'hba77348e),
	.w2(32'h3a880cae),
	.w3(32'h39438540),
	.w4(32'h3ac2fee8),
	.w5(32'h3b25a065),
	.w6(32'hba802082),
	.w7(32'h3afe99b9),
	.w8(32'h3bc2c68c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8532b3),
	.w1(32'h3b5ea3f3),
	.w2(32'h3b9897a7),
	.w3(32'h39eaa055),
	.w4(32'h3afdb7c0),
	.w5(32'hba879173),
	.w6(32'h3b2e843a),
	.w7(32'h3bac3e3c),
	.w8(32'hbaca3d2c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5470b7),
	.w1(32'h3a313e05),
	.w2(32'h3b122c7b),
	.w3(32'hba9a40b8),
	.w4(32'h3ae05e34),
	.w5(32'h3bbaad94),
	.w6(32'h3a3bad2f),
	.w7(32'h3a830357),
	.w8(32'h3b999352),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd029),
	.w1(32'h3b3e8a82),
	.w2(32'h3b8c9c34),
	.w3(32'h3b924b91),
	.w4(32'h3b3175fd),
	.w5(32'h3b9ddce4),
	.w6(32'h3ba1caaa),
	.w7(32'h3b875d3d),
	.w8(32'h3b942b8c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0d377),
	.w1(32'hba2769b6),
	.w2(32'h3ac95f83),
	.w3(32'h397328c4),
	.w4(32'h3b07d36f),
	.w5(32'h3a817102),
	.w6(32'h3bc0c746),
	.w7(32'h3ae4fb81),
	.w8(32'h3a68e515),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eeb25),
	.w1(32'h3b074cdf),
	.w2(32'h3b1126d1),
	.w3(32'h3a43cedd),
	.w4(32'hb9d6582b),
	.w5(32'hbb221894),
	.w6(32'h3b401440),
	.w7(32'h3a20b4c6),
	.w8(32'hbb5c9f5b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3176a3),
	.w1(32'hbb6a50a4),
	.w2(32'hbb8d1290),
	.w3(32'hbb3dcbf9),
	.w4(32'hbb91b0f4),
	.w5(32'hbac437e5),
	.w6(32'hb7c19777),
	.w7(32'hbb5f7048),
	.w8(32'hba7960cc),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2813ac),
	.w1(32'h3a9f4e79),
	.w2(32'h3aa227cd),
	.w3(32'hbb026cf1),
	.w4(32'hb85945fc),
	.w5(32'h3a92a5ca),
	.w6(32'hbb951276),
	.w7(32'hbb0b43cb),
	.w8(32'h3b04311e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3727f),
	.w1(32'h3a4191df),
	.w2(32'hbb2e939d),
	.w3(32'h3aef61b1),
	.w4(32'hba4ea51a),
	.w5(32'hbafa16a1),
	.w6(32'h3b3ca20a),
	.w7(32'hbb28e097),
	.w8(32'hb8ad4bfc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7be78),
	.w1(32'h39e27e78),
	.w2(32'h3b202a51),
	.w3(32'hbb538d4a),
	.w4(32'hbab53f79),
	.w5(32'hbb22dcda),
	.w6(32'h3b58370d),
	.w7(32'h3adfef23),
	.w8(32'hbb2051ec),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac95bda),
	.w1(32'h3b66e04b),
	.w2(32'h3b6b8f23),
	.w3(32'h3b3296c7),
	.w4(32'h3b6bb2a6),
	.w5(32'hbb0ebace),
	.w6(32'hb9218041),
	.w7(32'h3b4aa539),
	.w8(32'h3b116fff),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0156b9),
	.w1(32'h3a4d8ecd),
	.w2(32'h3a51a9fb),
	.w3(32'hbb1a1bcc),
	.w4(32'hbac08147),
	.w5(32'h3b4599d6),
	.w6(32'hb8acfd62),
	.w7(32'h3a85655b),
	.w8(32'h3b606adf),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e7611),
	.w1(32'h3bafb1db),
	.w2(32'h3baa5642),
	.w3(32'h3bdb5a0c),
	.w4(32'h3baee27a),
	.w5(32'h3bc22395),
	.w6(32'h3ba44338),
	.w7(32'h3aba7f82),
	.w8(32'h3b8eec0b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f10e8),
	.w1(32'h3b2ccfcd),
	.w2(32'hb8d08ca0),
	.w3(32'h3bbd9840),
	.w4(32'h3a4f7ed2),
	.w5(32'hbb842638),
	.w6(32'h39d9b158),
	.w7(32'hbb41a1d1),
	.w8(32'hbb52d9a0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0fe43),
	.w1(32'hbb328da4),
	.w2(32'hbb1ec1e4),
	.w3(32'hbb8a0be2),
	.w4(32'hbb1f5e67),
	.w5(32'h3990e4a8),
	.w6(32'hbb9791bc),
	.w7(32'hba8beee6),
	.w8(32'hbb6e1420),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaa267),
	.w1(32'hb9581aca),
	.w2(32'h3b10684c),
	.w3(32'h3b38a58c),
	.w4(32'h3acdfcff),
	.w5(32'h3c8122c4),
	.w6(32'hbb424dfb),
	.w7(32'hbb8b8b2e),
	.w8(32'h3c744a38),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c182165),
	.w1(32'h3be9d992),
	.w2(32'h3ba7774a),
	.w3(32'h3c2c4220),
	.w4(32'h3bf5c672),
	.w5(32'hbb89391a),
	.w6(32'h3c0c5620),
	.w7(32'h3b7edd27),
	.w8(32'hbba13f87),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c3e77),
	.w1(32'hbaee9501),
	.w2(32'h398a2a72),
	.w3(32'hbb633a33),
	.w4(32'hb9ef92c7),
	.w5(32'hbac8246a),
	.w6(32'hbba9ad68),
	.w7(32'hbb792677),
	.w8(32'h3a302b47),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09faf3),
	.w1(32'hba295fdf),
	.w2(32'hbab94bb9),
	.w3(32'hbaa59fd7),
	.w4(32'hbb11836c),
	.w5(32'hbab8c1b6),
	.w6(32'hba488ba5),
	.w7(32'hbae93577),
	.w8(32'hba78b928),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9864d2),
	.w1(32'hbb86100b),
	.w2(32'hbae41675),
	.w3(32'hbb51533b),
	.w4(32'hbb62f871),
	.w5(32'hba1f9739),
	.w6(32'hbbb0c694),
	.w7(32'hbbe5d6bd),
	.w8(32'hbb0a9273),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211fb8),
	.w1(32'h3a03543e),
	.w2(32'h3ae91650),
	.w3(32'hbb231487),
	.w4(32'hbaeb84bd),
	.w5(32'h3a713f4a),
	.w6(32'hbbb116d1),
	.w7(32'hba88c8cd),
	.w8(32'hba90b983),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f4370),
	.w1(32'hba76ab8b),
	.w2(32'hbac8b54e),
	.w3(32'h3ac79b39),
	.w4(32'hb9e1d7bc),
	.w5(32'h3599501c),
	.w6(32'hba39ac01),
	.w7(32'hbb0cbbdb),
	.w8(32'h3acfb6e9),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a4864),
	.w1(32'h3b2e23b7),
	.w2(32'h3b06f4d7),
	.w3(32'hba0cba4e),
	.w4(32'h396de0ac),
	.w5(32'hbacaa8ed),
	.w6(32'hbae719e4),
	.w7(32'h3aafbf6e),
	.w8(32'hbb97fe30),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb583bcc),
	.w1(32'hbae76913),
	.w2(32'hbaa9df24),
	.w3(32'hbaf02155),
	.w4(32'hb9df0181),
	.w5(32'h39c2d946),
	.w6(32'hbb79e0d3),
	.w7(32'h38bba0f3),
	.w8(32'hb7e013b9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c39853),
	.w1(32'hba857d74),
	.w2(32'h3a0abc89),
	.w3(32'h39304f33),
	.w4(32'h3aa98866),
	.w5(32'h3c1d6d48),
	.w6(32'h3a3a540b),
	.w7(32'hb99f806f),
	.w8(32'h3bf1564e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90c18),
	.w1(32'hb9c72162),
	.w2(32'h397b6ac9),
	.w3(32'h3bf44c8d),
	.w4(32'h3b649001),
	.w5(32'h3b82afac),
	.w6(32'hbb0c158b),
	.w7(32'hba4c8ec0),
	.w8(32'h3bc47445),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b695aee),
	.w1(32'h3bb405b8),
	.w2(32'h3b927065),
	.w3(32'h3be36ef0),
	.w4(32'h3b8dd755),
	.w5(32'h3a9bff6e),
	.w6(32'h3c09b1a2),
	.w7(32'h3b9e5508),
	.w8(32'hbaca7d92),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7274e8),
	.w1(32'hb9e42035),
	.w2(32'hb9052e4f),
	.w3(32'h397b137f),
	.w4(32'h3a6601c5),
	.w5(32'h3b466d6f),
	.w6(32'hb8407763),
	.w7(32'hb964e329),
	.w8(32'h3b1552d9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a435c15),
	.w1(32'h3a0791d4),
	.w2(32'h38f25e30),
	.w3(32'h39a5d3f1),
	.w4(32'h3996e7cb),
	.w5(32'hbab58df3),
	.w6(32'h3afd8cda),
	.w7(32'h3a53bda0),
	.w8(32'h3a88c238),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab800b),
	.w1(32'h3a968f79),
	.w2(32'hbb2bf474),
	.w3(32'hba9a3f38),
	.w4(32'hba880236),
	.w5(32'h3b86026a),
	.w6(32'h38d1a60b),
	.w7(32'hbb53eb3a),
	.w8(32'h3b210407),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a224908),
	.w1(32'h3b347142),
	.w2(32'h3a027ac2),
	.w3(32'h3b8d9b77),
	.w4(32'h3b6d295c),
	.w5(32'h3a6c7c27),
	.w6(32'h3b690690),
	.w7(32'h3ac16f9d),
	.w8(32'h3b510b36),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38cf57),
	.w1(32'h3a9f4ca3),
	.w2(32'h3a903fed),
	.w3(32'hbae0ea93),
	.w4(32'hba224f82),
	.w5(32'hbb9aeac1),
	.w6(32'hbb00e3dc),
	.w7(32'h3a8ee90e),
	.w8(32'hbb79483e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d04b37),
	.w1(32'hb9a8cbf5),
	.w2(32'h3b5f4c5a),
	.w3(32'hbb57de77),
	.w4(32'h3b0044cd),
	.w5(32'h3bd426ae),
	.w6(32'hbbc6bb85),
	.w7(32'hba21c13b),
	.w8(32'h3b7803d8),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa3d0),
	.w1(32'h3b254a30),
	.w2(32'h3baff669),
	.w3(32'h3b077de5),
	.w4(32'h3b48caee),
	.w5(32'h3b569c47),
	.w6(32'hb9e80a0a),
	.w7(32'h3b097810),
	.w8(32'h3b33ba44),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47c1b0),
	.w1(32'hbac2f193),
	.w2(32'hba921516),
	.w3(32'hbb3c0e0c),
	.w4(32'hba709829),
	.w5(32'hbad014a5),
	.w6(32'hbad5120e),
	.w7(32'h3a6e5e6a),
	.w8(32'hbadc1c49),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949db43),
	.w1(32'h3a8c1f50),
	.w2(32'h3b022dc8),
	.w3(32'hbb95bff9),
	.w4(32'hbb8542b0),
	.w5(32'hba0c8802),
	.w6(32'hbb88e3a5),
	.w7(32'hbb10c9d1),
	.w8(32'h3ab261c6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae1a2e),
	.w1(32'hba08785e),
	.w2(32'hbb15e38f),
	.w3(32'hba94d790),
	.w4(32'h390280a1),
	.w5(32'h399b0b1c),
	.w6(32'hba9ffbd4),
	.w7(32'hbad7894a),
	.w8(32'h3a0bb91d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b159e80),
	.w1(32'h3a2f69c4),
	.w2(32'h3a99647a),
	.w3(32'h3a561f0d),
	.w4(32'h3b0a1eee),
	.w5(32'h3ba008a5),
	.w6(32'h38205b8e),
	.w7(32'h3a78662b),
	.w8(32'h3ac1f4fb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f2eab),
	.w1(32'h3ac7596e),
	.w2(32'h39fcae30),
	.w3(32'h3b99ba84),
	.w4(32'h3acd5432),
	.w5(32'h3b3aaa5c),
	.w6(32'h3a074827),
	.w7(32'h37bc6e72),
	.w8(32'hb877e96a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39176d56),
	.w1(32'hbb05789b),
	.w2(32'hbab8abe4),
	.w3(32'h3b33f229),
	.w4(32'h3b2f36ff),
	.w5(32'h3b00c393),
	.w6(32'hbb3b6ece),
	.w7(32'h392a484a),
	.w8(32'h39ba2197),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae78e4),
	.w1(32'h3b875513),
	.w2(32'h3be141c7),
	.w3(32'h3b752302),
	.w4(32'h3bdef4e6),
	.w5(32'h3b4a8f22),
	.w6(32'hbaff6b9f),
	.w7(32'h3b780468),
	.w8(32'h3a9b4030),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f9fa8),
	.w1(32'h3ae5132b),
	.w2(32'h3ba0d62d),
	.w3(32'h3a1bcbbd),
	.w4(32'h3ad5047c),
	.w5(32'hba9597b3),
	.w6(32'h3a9f98e2),
	.w7(32'h3b1be374),
	.w8(32'hba521058),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba607419),
	.w1(32'hbb4e35e9),
	.w2(32'hbb3d5bf9),
	.w3(32'hbb008628),
	.w4(32'hbb543c5b),
	.w5(32'hba5a702c),
	.w6(32'hbb27a577),
	.w7(32'hbbddc71f),
	.w8(32'hbb4109a7),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9066160),
	.w1(32'hbaefe74b),
	.w2(32'h39e5377c),
	.w3(32'hbb20a926),
	.w4(32'hba270ded),
	.w5(32'h3b11d3fb),
	.w6(32'hbba527da),
	.w7(32'hba243342),
	.w8(32'h3b44f6e4),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bd743),
	.w1(32'h3ad841cf),
	.w2(32'h392b4aa8),
	.w3(32'h3ba9e6fc),
	.w4(32'h3b6ab5dd),
	.w5(32'h3a0abd67),
	.w6(32'h39e4d718),
	.w7(32'h3ae8a8ac),
	.w8(32'h3989043c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51414e),
	.w1(32'h398e8373),
	.w2(32'hb7cb7f54),
	.w3(32'hba641a42),
	.w4(32'hbb643aee),
	.w5(32'hbb80bb63),
	.w6(32'hbacf24c7),
	.w7(32'hbaed986c),
	.w8(32'hbb6a4e22),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eeec0),
	.w1(32'hbaacba94),
	.w2(32'hbb0a0c06),
	.w3(32'hbb15b0d6),
	.w4(32'hbb2e8d7b),
	.w5(32'h3b6afd5c),
	.w6(32'h3abaf5d2),
	.w7(32'hbb4ccfc0),
	.w8(32'h3abea9d3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a928dc0),
	.w1(32'h3ae46369),
	.w2(32'h3af6a8d3),
	.w3(32'h3b4fd6ab),
	.w4(32'h3b6a348d),
	.w5(32'hbad250d6),
	.w6(32'hba0e1256),
	.w7(32'h3a5d207d),
	.w8(32'hbb66b50c),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb883f93),
	.w1(32'hba17fb34),
	.w2(32'hba1898bd),
	.w3(32'hb9ab732c),
	.w4(32'hba722f83),
	.w5(32'h3bd2242d),
	.w6(32'h3a1995fb),
	.w7(32'hba86cde3),
	.w8(32'h3bbd20ce),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0aa1a),
	.w1(32'hb9292f21),
	.w2(32'hb85a1d96),
	.w3(32'h3bba0e64),
	.w4(32'h3b64beca),
	.w5(32'h3b240fe6),
	.w6(32'h38e51c21),
	.w7(32'h392bfb5e),
	.w8(32'h3b1633b8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20d90),
	.w1(32'hbb5e8bb6),
	.w2(32'hbab5a5aa),
	.w3(32'hba9e2bbf),
	.w4(32'hba6ea33a),
	.w5(32'h3a3e8cc4),
	.w6(32'hba7f9aa1),
	.w7(32'hbb18ceb7),
	.w8(32'hba9a6bfe),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c93d0),
	.w1(32'hbaad5b0c),
	.w2(32'h3b8b3922),
	.w3(32'h3a86450e),
	.w4(32'h3b3ea90e),
	.w5(32'h3b4df769),
	.w6(32'hbb4cb0eb),
	.w7(32'h3aa4fa00),
	.w8(32'h3b8b2cc5),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68e4be),
	.w1(32'h3a10278a),
	.w2(32'h3ad94ee7),
	.w3(32'h3aca1241),
	.w4(32'h3acd9fe8),
	.w5(32'h3a39edb2),
	.w6(32'hbaf7e127),
	.w7(32'h3a8972ce),
	.w8(32'hbbb8e0ec),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc93594),
	.w1(32'hba583da9),
	.w2(32'h3acbe9a0),
	.w3(32'hb9f17fcb),
	.w4(32'h3b31df12),
	.w5(32'h3b6013e2),
	.w6(32'hbbbe0714),
	.w7(32'hbadee2fb),
	.w8(32'h3a8c42af),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b08a),
	.w1(32'hbaf5fd22),
	.w2(32'hbaecabb9),
	.w3(32'hba8054c7),
	.w4(32'hb9c46927),
	.w5(32'h3b5d8292),
	.w6(32'hb977d6d3),
	.w7(32'hbaa0f559),
	.w8(32'h3afe520c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21fc6f),
	.w1(32'hba0362cc),
	.w2(32'hba37d415),
	.w3(32'h3ab74806),
	.w4(32'h384c2ae6),
	.w5(32'h3c59de7e),
	.w6(32'hb83d623a),
	.w7(32'hbb0bee95),
	.w8(32'h3c3429b2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b4ae7),
	.w1(32'h3c4ade69),
	.w2(32'h3c85c829),
	.w3(32'h3c534b45),
	.w4(32'h3c8a52ce),
	.w5(32'h3b6b0932),
	.w6(32'h3bfe412f),
	.w7(32'h3c85932b),
	.w8(32'h3b86726e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94459f4),
	.w1(32'hbade9d4f),
	.w2(32'hbb3de4f7),
	.w3(32'h3b88f7f0),
	.w4(32'hba9a2929),
	.w5(32'h39b4edbc),
	.w6(32'h3ae7e4a3),
	.w7(32'hbb5e9139),
	.w8(32'hbb389e1f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15c02a),
	.w1(32'h3a49bf32),
	.w2(32'h3ae8697c),
	.w3(32'h3ad5a4a9),
	.w4(32'h3a3ad52d),
	.w5(32'h3a31f107),
	.w6(32'hba63ae2b),
	.w7(32'h3a7d4b9f),
	.w8(32'h3b380eae),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab93d23),
	.w1(32'h3a30f8ac),
	.w2(32'h3a8bac82),
	.w3(32'h3ac71177),
	.w4(32'h3b6da342),
	.w5(32'h3b43635f),
	.w6(32'h3b762578),
	.w7(32'h3a7d28d5),
	.w8(32'hbb35e63f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f58cd),
	.w1(32'hbb970c2f),
	.w2(32'hbb44462b),
	.w3(32'h3b1a78f5),
	.w4(32'h3b39eb1e),
	.w5(32'h3ae49f4e),
	.w6(32'hbadaa881),
	.w7(32'h3a910901),
	.w8(32'h3b862eb1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25337f),
	.w1(32'h3adc2cb7),
	.w2(32'h3a86b4ab),
	.w3(32'h3a3cdeb8),
	.w4(32'h3a9dd554),
	.w5(32'hbb8c57b1),
	.w6(32'h3a8769d8),
	.w7(32'h3b54e490),
	.w8(32'hbc087cbb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7afb45),
	.w1(32'hb93483bb),
	.w2(32'hbb1a035d),
	.w3(32'hbb8e458c),
	.w4(32'h3abc7d94),
	.w5(32'h3b77337d),
	.w6(32'hbba1b6ed),
	.w7(32'h39d16c7e),
	.w8(32'h3b920f2f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89913a),
	.w1(32'hbb16d97c),
	.w2(32'hbaa26d93),
	.w3(32'h3b0cfbcd),
	.w4(32'h3b094363),
	.w5(32'h39cf5a49),
	.w6(32'hbb1b2325),
	.w7(32'hbb71082a),
	.w8(32'hbbcca067),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba800643),
	.w1(32'hb8e85ac7),
	.w2(32'hbb7e7216),
	.w3(32'hbaeeb30b),
	.w4(32'hba884406),
	.w5(32'h3bea10e5),
	.w6(32'hbb487d24),
	.w7(32'hbb4c4c69),
	.w8(32'h3bbeef4d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2a70a),
	.w1(32'h3b43dda0),
	.w2(32'h3b92d862),
	.w3(32'hb8fc38d6),
	.w4(32'h3afe7b9b),
	.w5(32'h39ad08f5),
	.w6(32'h3ba5e0d4),
	.w7(32'h3b972b38),
	.w8(32'h3af8e9a4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4e517),
	.w1(32'h391e54cc),
	.w2(32'hb9c116d2),
	.w3(32'h39edaeeb),
	.w4(32'h396c81f1),
	.w5(32'h3a0e138f),
	.w6(32'hb945b434),
	.w7(32'hba3962fe),
	.w8(32'hba315703),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990e413),
	.w1(32'h394cdb41),
	.w2(32'h3a1d00e8),
	.w3(32'h3ae67b8c),
	.w4(32'h3ab0fc5e),
	.w5(32'h3b1bf4dc),
	.w6(32'hba4c4a46),
	.w7(32'h3a6a516e),
	.w8(32'h3a4d7d47),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ddc17),
	.w1(32'h3ab62f01),
	.w2(32'hb9585670),
	.w3(32'h3aa6cfa0),
	.w4(32'h3b167048),
	.w5(32'h3aa717da),
	.w6(32'h3aa08d16),
	.w7(32'hbae99db0),
	.w8(32'hba8b7d13),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c59d7),
	.w1(32'hba17de41),
	.w2(32'h3ac182b3),
	.w3(32'h3ae935e5),
	.w4(32'h3b9dccb6),
	.w5(32'h3a45cd63),
	.w6(32'hbb174f68),
	.w7(32'hb634b2f0),
	.w8(32'h3aa5f7e7),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa47158),
	.w1(32'h3a765b51),
	.w2(32'h3a575def),
	.w3(32'hba1e4ec3),
	.w4(32'hba964131),
	.w5(32'hb7948cfb),
	.w6(32'hbaaaab40),
	.w7(32'hbb0d9ac4),
	.w8(32'hb7dbb112),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2fa79),
	.w1(32'h39384ac0),
	.w2(32'hb9b6f0f7),
	.w3(32'h39b3a3a7),
	.w4(32'h3967e776),
	.w5(32'hb98c38f4),
	.w6(32'h3a32b6a2),
	.w7(32'h39e66693),
	.w8(32'h388d9650),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaa914),
	.w1(32'hb95b00cc),
	.w2(32'hb9fd17d3),
	.w3(32'h3b1204b4),
	.w4(32'h3901b62e),
	.w5(32'hba4d4e63),
	.w6(32'h38fbd126),
	.w7(32'hbad5ec90),
	.w8(32'hbad7bf40),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21103a),
	.w1(32'h3a3efb4c),
	.w2(32'h3b395813),
	.w3(32'h3a9a820c),
	.w4(32'h3a8e24b8),
	.w5(32'h3b0de1d2),
	.w6(32'h3974dd9f),
	.w7(32'h394ac1de),
	.w8(32'h3ac04de2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5cd2b04),
	.w1(32'hb79e8d36),
	.w2(32'hb82b23d2),
	.w3(32'h37996d6b),
	.w4(32'hb6e857f0),
	.w5(32'hb8459b12),
	.w6(32'hb7c21e17),
	.w7(32'hb7efc7ba),
	.w8(32'hb7bc4cea),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4d4e3),
	.w1(32'hba4edcfc),
	.w2(32'hbb4c08a3),
	.w3(32'hb9bb5549),
	.w4(32'hb7a7a4dc),
	.w5(32'hbab16499),
	.w6(32'h38fdd807),
	.w7(32'hbaaaae7d),
	.w8(32'hbb806e07),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5ee98),
	.w1(32'h38fbbbcb),
	.w2(32'h3961157a),
	.w3(32'h3903c6c2),
	.w4(32'h386b3c82),
	.w5(32'hb96676b5),
	.w6(32'hb9123cf5),
	.w7(32'hba8a8685),
	.w8(32'hbabed067),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a53b44),
	.w1(32'hb8fbadb2),
	.w2(32'hb9171dd8),
	.w3(32'h3780fad9),
	.w4(32'hb96d4f9f),
	.w5(32'hb94ba029),
	.w6(32'hb817e9ee),
	.w7(32'hb6e7b2cc),
	.w8(32'hb6bd7525),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ac98c),
	.w1(32'hba702e96),
	.w2(32'hba95658b),
	.w3(32'hb9d41429),
	.w4(32'hb9960935),
	.w5(32'hba53d366),
	.w6(32'hb9bd306b),
	.w7(32'hba6d9992),
	.w8(32'hbaca1bb7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c52dbc),
	.w1(32'h385e1383),
	.w2(32'h38b31a75),
	.w3(32'h389c041e),
	.w4(32'h38b14449),
	.w5(32'h391128ad),
	.w6(32'hb7aeecf7),
	.w7(32'hb7c2819b),
	.w8(32'h388f03a4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b0525),
	.w1(32'hba3ebf08),
	.w2(32'hb907199f),
	.w3(32'hb9dcd5d3),
	.w4(32'hba0ec35b),
	.w5(32'hb8d0afab),
	.w6(32'hb956f329),
	.w7(32'hb9254347),
	.w8(32'h3802cb4a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79752e6),
	.w1(32'hb65de418),
	.w2(32'hb7369476),
	.w3(32'hb51036bd),
	.w4(32'hb7af6cd5),
	.w5(32'hb6dcda4f),
	.w6(32'hb71aad3b),
	.w7(32'hb7b401c7),
	.w8(32'h375aa7ee),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369b0ebc),
	.w1(32'h373eebc5),
	.w2(32'hb5c074b6),
	.w3(32'h36e9d4c9),
	.w4(32'h37bf4206),
	.w5(32'h3590198e),
	.w6(32'h37025b01),
	.w7(32'hb69fed5a),
	.w8(32'hb800ba00),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4a3f7),
	.w1(32'h3aba710d),
	.w2(32'h3a6a634e),
	.w3(32'h3abef71a),
	.w4(32'h3a6e8398),
	.w5(32'h396988e2),
	.w6(32'h3abe5cd1),
	.w7(32'h3aa87267),
	.w8(32'h3a7aae72),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2726),
	.w1(32'h3a9c228c),
	.w2(32'h3adfa387),
	.w3(32'h3ae93b0a),
	.w4(32'h3aeee0a6),
	.w5(32'h3b1ac882),
	.w6(32'hb98f41b8),
	.w7(32'hba30b468),
	.w8(32'h36b53542),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cf7c0),
	.w1(32'h3b077fbf),
	.w2(32'h3a88c438),
	.w3(32'h3b0162a0),
	.w4(32'h3a0e452f),
	.w5(32'hba13eaf3),
	.w6(32'h39d3666c),
	.w7(32'hbac674ae),
	.w8(32'hbb009cee),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5af0e),
	.w1(32'hb92c640a),
	.w2(32'h3aa49acc),
	.w3(32'h3a6e965a),
	.w4(32'h3a0eab90),
	.w5(32'h3af35024),
	.w6(32'hb9e476ed),
	.w7(32'hba934c53),
	.w8(32'h36d29f1f),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80a82e6),
	.w1(32'hb942b928),
	.w2(32'hb9a3a2de),
	.w3(32'h36efca8e),
	.w4(32'hb9343e9e),
	.w5(32'hb9acd447),
	.w6(32'h39253ff5),
	.w7(32'h3707a80c),
	.w8(32'hb963aa6e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd55e7),
	.w1(32'hb9bd523c),
	.w2(32'hb99e1922),
	.w3(32'hb925d5a0),
	.w4(32'hb8f6a6ee),
	.w5(32'hb89e4a2f),
	.w6(32'h38d9be5f),
	.w7(32'hb88d7886),
	.w8(32'hb8cdec0e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59e95e2),
	.w1(32'h368f6bd0),
	.w2(32'h36dfceea),
	.w3(32'hb4a7e635),
	.w4(32'hb6aef7e7),
	.w5(32'h3711a2dd),
	.w6(32'hb69a09a8),
	.w7(32'hb6d91f69),
	.w8(32'hb7258851),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da9e30),
	.w1(32'h376dabb9),
	.w2(32'h381ff0ec),
	.w3(32'hb84a28c5),
	.w4(32'hb873d70d),
	.w5(32'hb83a3293),
	.w6(32'hb86ab711),
	.w7(32'hb84fcae9),
	.w8(32'hb7c4d717),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868e914),
	.w1(32'hba28ab22),
	.w2(32'hba86e727),
	.w3(32'hb80962f8),
	.w4(32'hb9d56e79),
	.w5(32'hbac4ba86),
	.w6(32'hb9e251ba),
	.w7(32'hbad207f4),
	.w8(32'hbb1b5ce8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bcae9b),
	.w1(32'h39c22608),
	.w2(32'h39ce4e1b),
	.w3(32'h39b046d0),
	.w4(32'h39d2cae8),
	.w5(32'h39b138a4),
	.w6(32'h39aa1f78),
	.w7(32'h39d10314),
	.w8(32'h396db076),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ecbba),
	.w1(32'hb9eed02c),
	.w2(32'hba0bbd28),
	.w3(32'hba425fc1),
	.w4(32'hb9c7f145),
	.w5(32'hba86e6cc),
	.w6(32'hb9ff2542),
	.w7(32'h372bade5),
	.w8(32'hba3817e1),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f3541),
	.w1(32'hba30332c),
	.w2(32'hb9ec5b02),
	.w3(32'hb9c5db29),
	.w4(32'hb9bc69b9),
	.w5(32'hb9a5dbc0),
	.w6(32'hb9fbacc3),
	.w7(32'hb8dfbd58),
	.w8(32'h391fd39f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78befe4),
	.w1(32'hb7802041),
	.w2(32'h36f3e0a0),
	.w3(32'hb789e3f8),
	.w4(32'hb79363e9),
	.w5(32'hb701be4a),
	.w6(32'hb7d22735),
	.w7(32'hb73bb88f),
	.w8(32'hb75356b9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c1883),
	.w1(32'hb96222aa),
	.w2(32'h3899b4cb),
	.w3(32'hb96953c8),
	.w4(32'h38cfa519),
	.w5(32'h393ded76),
	.w6(32'hb9b3e55c),
	.w7(32'hb9ae3066),
	.w8(32'hb94eec48),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d45991),
	.w1(32'hb8c1d70c),
	.w2(32'hb98b42bb),
	.w3(32'hb91a6ef2),
	.w4(32'hb8aff63b),
	.w5(32'hb949cdd6),
	.w6(32'h3858f4cc),
	.w7(32'h3814bb8b),
	.w8(32'hb912d507),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f02a0),
	.w1(32'hbb1aa23d),
	.w2(32'hbae99c88),
	.w3(32'h3a43d531),
	.w4(32'hb8a85c16),
	.w5(32'hbaf489b5),
	.w6(32'hbaf560b8),
	.w7(32'hbb495cbe),
	.w8(32'hbb94c967),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb756785e),
	.w1(32'hb8e5d021),
	.w2(32'hb8b855f3),
	.w3(32'hb4567c50),
	.w4(32'hb8a6aeb0),
	.w5(32'hb87a9e3a),
	.w6(32'hb76f3b0e),
	.w7(32'hb85ef5f2),
	.w8(32'hb7571912),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d0ba9),
	.w1(32'h3b76049c),
	.w2(32'h3b59a5aa),
	.w3(32'h3adf1266),
	.w4(32'h3a39f12c),
	.w5(32'h38cf5ebe),
	.w6(32'hb9c9ea52),
	.w7(32'hba0db012),
	.w8(32'hb9a9b059),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule