module layer_8_featuremap_45(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae236b2),
	.w1(32'hbaf7e069),
	.w2(32'hbabd2fcc),
	.w3(32'hba8679e3),
	.w4(32'hbac22cc6),
	.w5(32'hbb09a7c0),
	.w6(32'h3b378bfe),
	.w7(32'h3b57327d),
	.w8(32'h3899f800),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeade47),
	.w1(32'hbb227688),
	.w2(32'hbae774c1),
	.w3(32'hbaaf7951),
	.w4(32'hbaf05d49),
	.w5(32'hbaf1d98f),
	.w6(32'h35dda742),
	.w7(32'hbad1afca),
	.w8(32'hbaafc872),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8419f),
	.w1(32'hbb202ddd),
	.w2(32'h3a0a8b08),
	.w3(32'hbbdbb896),
	.w4(32'hbb829cdf),
	.w5(32'hbb42b785),
	.w6(32'hbbddbf5b),
	.w7(32'hbbaad214),
	.w8(32'hbb140298),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820b20),
	.w1(32'hba05e50f),
	.w2(32'h397a50b7),
	.w3(32'hb9a29ff0),
	.w4(32'h38800612),
	.w5(32'h3a095643),
	.w6(32'h3bbaf7cc),
	.w7(32'h3b662d27),
	.w8(32'h3a1be51b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca090),
	.w1(32'hbb9eabf1),
	.w2(32'hbac6b30b),
	.w3(32'hbb9f6508),
	.w4(32'hbbb962bd),
	.w5(32'hbb621173),
	.w6(32'h39f79bc9),
	.w7(32'hba9e944b),
	.w8(32'hba762d05),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc67ea6),
	.w1(32'h3bccba68),
	.w2(32'h3ba85c79),
	.w3(32'h3b21d912),
	.w4(32'h3af5f6e2),
	.w5(32'h384878e4),
	.w6(32'h390cba18),
	.w7(32'h3a7d0c9a),
	.w8(32'h3b22aab2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc66f),
	.w1(32'hba904da5),
	.w2(32'hba3d5176),
	.w3(32'hb9f630fe),
	.w4(32'hba554b63),
	.w5(32'hba0406fd),
	.w6(32'hba466a56),
	.w7(32'hba001b9f),
	.w8(32'hb99b2cd3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072752),
	.w1(32'hbb1dbd33),
	.w2(32'h39fb5076),
	.w3(32'hbc0ba4ca),
	.w4(32'hbc0874c0),
	.w5(32'hbb917e6c),
	.w6(32'hbb9c8bbe),
	.w7(32'hbba7f71a),
	.w8(32'hbbaa51c6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2deddb),
	.w1(32'hbbecdae0),
	.w2(32'hba73346f),
	.w3(32'hbbf9fd76),
	.w4(32'hbc04806f),
	.w5(32'hbb5809e6),
	.w6(32'hbbe1adea),
	.w7(32'hbbaa3c52),
	.w8(32'h3a5f83e0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ce9ac),
	.w1(32'h3a2be8a7),
	.w2(32'h3ac585ef),
	.w3(32'hba215f75),
	.w4(32'h3a6c2b57),
	.w5(32'hba25d447),
	.w6(32'hbadceca0),
	.w7(32'h39fd00fa),
	.w8(32'h3ab68ae5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290ec9),
	.w1(32'hbc048440),
	.w2(32'hbbcff707),
	.w3(32'hbba8df6e),
	.w4(32'hbbfa115c),
	.w5(32'hbba0c379),
	.w6(32'h3b526e33),
	.w7(32'h3b1033a8),
	.w8(32'hbaf5fec7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9af2b63),
	.w1(32'hbb05f5d7),
	.w2(32'hbb01e089),
	.w3(32'hba75152c),
	.w4(32'hbaa69d3d),
	.w5(32'hbb212502),
	.w6(32'hb997dae0),
	.w7(32'h3a1bba86),
	.w8(32'hba8c9dc7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121801),
	.w1(32'h3a204343),
	.w2(32'h3b823ee5),
	.w3(32'hbb966964),
	.w4(32'hbb1aac9a),
	.w5(32'h3a29ed74),
	.w6(32'hbb95fbc4),
	.w7(32'hbb87b202),
	.w8(32'h390dbe7d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba895a20),
	.w1(32'hbacf5731),
	.w2(32'hbad423d9),
	.w3(32'hbac125c1),
	.w4(32'hbaff4c53),
	.w5(32'hbae70b5e),
	.w6(32'hbad5c424),
	.w7(32'hbacdae7e),
	.w8(32'hba5aec32),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3808be),
	.w1(32'hba54f902),
	.w2(32'hba75c647),
	.w3(32'hba68de00),
	.w4(32'hba8a824c),
	.w5(32'hba7d2efe),
	.w6(32'hba78c750),
	.w7(32'hba8c77c8),
	.w8(32'hb9b5e717),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5b3d6),
	.w1(32'hbac661d4),
	.w2(32'hba74db2f),
	.w3(32'hbb0831ce),
	.w4(32'hbaf5d469),
	.w5(32'hba973f43),
	.w6(32'hbb18db64),
	.w7(32'hbac473b5),
	.w8(32'hba6fef88),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2976d8),
	.w1(32'h38bcbf32),
	.w2(32'hba80e0d9),
	.w3(32'hbaf46bb7),
	.w4(32'hbacfb499),
	.w5(32'hbafa5b9c),
	.w6(32'hbb1f064e),
	.w7(32'hb9e6fc87),
	.w8(32'hba289ccd),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb522f0d),
	.w1(32'hba29b442),
	.w2(32'h3a909bca),
	.w3(32'hbbc52c91),
	.w4(32'hbba5d779),
	.w5(32'hbb8b4e60),
	.w6(32'hbb8121eb),
	.w7(32'hbb6e1226),
	.w8(32'h3acd3a75),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80d834),
	.w1(32'hbcd5dbee),
	.w2(32'hbc54b8b4),
	.w3(32'hbbc1aeb6),
	.w4(32'hbc132853),
	.w5(32'hbb61b5da),
	.w6(32'h3c206b98),
	.w7(32'h3ba9d550),
	.w8(32'hbb0fe259),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1e0e9),
	.w1(32'hbb7efed8),
	.w2(32'h3a61f144),
	.w3(32'hbc252f1d),
	.w4(32'hbc367934),
	.w5(32'hbbad402a),
	.w6(32'h3bc0fc46),
	.w7(32'h3a2f5344),
	.w8(32'h3b1649e4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8caff9),
	.w1(32'h3ac549c0),
	.w2(32'hbb469b72),
	.w3(32'h3b817808),
	.w4(32'h3b5bd8d5),
	.w5(32'h3a591aeb),
	.w6(32'h3b45744c),
	.w7(32'h3bee597a),
	.w8(32'h3bc2dfd5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e3b1),
	.w1(32'h3b8c6f90),
	.w2(32'h3b641b6b),
	.w3(32'hbb71a57b),
	.w4(32'h3b18da50),
	.w5(32'h3ab239f5),
	.w6(32'hba6d7c2f),
	.w7(32'h3a7dfa00),
	.w8(32'h3b824502),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9570cc4),
	.w1(32'hbc6f1223),
	.w2(32'hbbdccde0),
	.w3(32'hbc013245),
	.w4(32'hbc952c84),
	.w5(32'hbc58be7f),
	.w6(32'h3c5a4b6a),
	.w7(32'h3c2be258),
	.w8(32'hba1addae),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70a953),
	.w1(32'h3ac5b212),
	.w2(32'h3b0a99fd),
	.w3(32'hb9b0e7a0),
	.w4(32'hbb64bb9c),
	.w5(32'hbb226dcf),
	.w6(32'hb9c41637),
	.w7(32'hbb6dcf15),
	.w8(32'hbac4c3a6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba355eea),
	.w1(32'hbb37927b),
	.w2(32'hbb7e3071),
	.w3(32'hba0242ed),
	.w4(32'hbb0af25c),
	.w5(32'hbb93f50c),
	.w6(32'hbb0ed0a3),
	.w7(32'hbaa196f2),
	.w8(32'hbad46e63),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9063bf),
	.w1(32'hbb57f572),
	.w2(32'h374eab29),
	.w3(32'h3aa7408b),
	.w4(32'hbbb51b4f),
	.w5(32'hbb0250f2),
	.w6(32'h3c423b64),
	.w7(32'h3be48d06),
	.w8(32'h3bb75a47),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b532149),
	.w1(32'h3b06f2f9),
	.w2(32'h3afd6d0d),
	.w3(32'h3b7c2b1b),
	.w4(32'h3b14452a),
	.w5(32'h3b049229),
	.w6(32'h3b6ca055),
	.w7(32'h3b2af96e),
	.w8(32'h3a08eb2b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba27b85),
	.w1(32'hbd212509),
	.w2(32'hbd5d72fc),
	.w3(32'hbc6cd12f),
	.w4(32'hbd5e93d5),
	.w5(32'hbcc440f8),
	.w6(32'h3ca35b52),
	.w7(32'h3dd6568f),
	.w8(32'h3d4584f1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e526f),
	.w1(32'hbb7b4dc9),
	.w2(32'hbab2d092),
	.w3(32'hbb01f170),
	.w4(32'hbb9cc8df),
	.w5(32'hbb37e2aa),
	.w6(32'h3b49b5d7),
	.w7(32'h3b236bfc),
	.w8(32'h3aa525f5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955634b),
	.w1(32'h38f0b381),
	.w2(32'h39afbf25),
	.w3(32'hba80bc1c),
	.w4(32'hba12ac54),
	.w5(32'hba5574b4),
	.w6(32'hbad6355f),
	.w7(32'hbab89d9b),
	.w8(32'hbaf4b431),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb84732),
	.w1(32'h3bd21b2f),
	.w2(32'h3b4edfe6),
	.w3(32'h3bfabbac),
	.w4(32'h3bede1b5),
	.w5(32'h3b83d363),
	.w6(32'h3bd7731d),
	.w7(32'h3bcc60ba),
	.w8(32'h3b1fdde3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1422c7),
	.w1(32'hbacf125e),
	.w2(32'hbaabf9e1),
	.w3(32'hba8ffdbf),
	.w4(32'hbae21bff),
	.w5(32'hb9dfec14),
	.w6(32'h3b01cd7b),
	.w7(32'h3a1addc7),
	.w8(32'h3b1bfa17),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f971e1),
	.w1(32'hb7b47946),
	.w2(32'hb9f5e653),
	.w3(32'hb98b5915),
	.w4(32'hb94284e3),
	.w5(32'hb98a8d33),
	.w6(32'hba1acff3),
	.w7(32'hba145365),
	.w8(32'hba38f4e5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984c58a),
	.w1(32'hba191997),
	.w2(32'hba098c93),
	.w3(32'hb9f80fa1),
	.w4(32'hb9f635a3),
	.w5(32'hb9dd6cf9),
	.w6(32'hb91e2959),
	.w7(32'hba534b79),
	.w8(32'hba0659e0),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba97670),
	.w1(32'h3bbf7443),
	.w2(32'h3b7bd96a),
	.w3(32'h3b4a7b73),
	.w4(32'h3b2399c8),
	.w5(32'h3a1399a9),
	.w6(32'h3a5d16bd),
	.w7(32'hb9983b0d),
	.w8(32'h3aab5938),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39478927),
	.w1(32'hbbfef462),
	.w2(32'hbbfbd97c),
	.w3(32'h3aea680c),
	.w4(32'hbae3a6da),
	.w5(32'hbb21b929),
	.w6(32'h3ba634bb),
	.w7(32'h3b1d13d3),
	.w8(32'h3a002aaf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925bf33),
	.w1(32'hb9c0c596),
	.w2(32'h394782e9),
	.w3(32'h398fdb3f),
	.w4(32'h39242e84),
	.w5(32'h3996d6a7),
	.w6(32'hb8484a52),
	.w7(32'h392efb91),
	.w8(32'hb9909268),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5976b0),
	.w1(32'hbac796be),
	.w2(32'hbaaf6d13),
	.w3(32'hba7f1940),
	.w4(32'h3a9c43a5),
	.w5(32'h39f19caf),
	.w6(32'h3b2d8b06),
	.w7(32'h3b72a1ce),
	.w8(32'h3aab500f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4acd9),
	.w1(32'hbac5cf46),
	.w2(32'hbade59e2),
	.w3(32'hbad1acae),
	.w4(32'hbb026f3b),
	.w5(32'hbadeafcc),
	.w6(32'hbad9ed76),
	.w7(32'hbaf8158b),
	.w8(32'hba871edb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45fc72),
	.w1(32'hba8c3d33),
	.w2(32'h392fa2d3),
	.w3(32'hb88093de),
	.w4(32'hb915761c),
	.w5(32'h3a0a1a31),
	.w6(32'hb940cb2f),
	.w7(32'h3a8b2702),
	.w8(32'h3aeb1802),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0332bf),
	.w1(32'hba944589),
	.w2(32'h3b155c74),
	.w3(32'h3b00aa9d),
	.w4(32'hbbbd9b11),
	.w5(32'hbbd2403b),
	.w6(32'h3c492210),
	.w7(32'h3bacb3a5),
	.w8(32'hbb14c230),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae506de),
	.w1(32'hbaa8c766),
	.w2(32'h3ab9c525),
	.w3(32'hba970e5b),
	.w4(32'hbae69bc2),
	.w5(32'h3939b2a9),
	.w6(32'h3a3ce723),
	.w7(32'h3a8dc271),
	.w8(32'h3bee3fe3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac13081),
	.w1(32'h3a010ef4),
	.w2(32'h3a67de3e),
	.w3(32'h3b4cdc3a),
	.w4(32'hbaa63323),
	.w5(32'hba7ea1f6),
	.w6(32'h3aa51e7f),
	.w7(32'h3ab5f3b3),
	.w8(32'hbae715e4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac761ab),
	.w1(32'hbb897593),
	.w2(32'hbb3a4841),
	.w3(32'hbba6fdfc),
	.w4(32'hbbcf1436),
	.w5(32'hbbdf5ca6),
	.w6(32'hba3f93c1),
	.w7(32'hb9b26b8b),
	.w8(32'hbb425ac2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb232ef1),
	.w1(32'hbbaa8692),
	.w2(32'h3b122b55),
	.w3(32'hbc163f09),
	.w4(32'hbc025d3a),
	.w5(32'hbb072c8f),
	.w6(32'h3b9610ad),
	.w7(32'h3ba84139),
	.w8(32'h3a3f31a5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c0e42),
	.w1(32'hbb839af3),
	.w2(32'hba3178c2),
	.w3(32'hba821943),
	.w4(32'h3a2ebbd5),
	.w5(32'h3b280bed),
	.w6(32'hba2c9cfa),
	.w7(32'h3a69f08a),
	.w8(32'h3c17ed31),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29b0a5),
	.w1(32'hbbd53481),
	.w2(32'hbc01bfeb),
	.w3(32'hbb19bcae),
	.w4(32'hbc039177),
	.w5(32'hbbb9c8cc),
	.w6(32'h3a622cd4),
	.w7(32'hbaee0fab),
	.w8(32'hbb3e3814),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153a06),
	.w1(32'hbc798708),
	.w2(32'hbb9c6bf6),
	.w3(32'hbc53acb1),
	.w4(32'hbc6b08e2),
	.w5(32'hbbbb1bcd),
	.w6(32'hbb3dede3),
	.w7(32'h3ad19303),
	.w8(32'h3ba056f9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb2606),
	.w1(32'h392906f8),
	.w2(32'h3b2504ca),
	.w3(32'h3a1c0e20),
	.w4(32'h378bdfd9),
	.w5(32'h3ab9d320),
	.w6(32'h3a9e9c5e),
	.w7(32'h3b0bc8a4),
	.w8(32'hbb193032),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19b88a),
	.w1(32'hbb599008),
	.w2(32'h39d7dcab),
	.w3(32'h390b33f7),
	.w4(32'hbaeb0504),
	.w5(32'h3abf194a),
	.w6(32'h3bc97978),
	.w7(32'h3b5d72e1),
	.w8(32'h3a34e491),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba16ad8c),
	.w1(32'h3bd9b716),
	.w2(32'h3ba3ed07),
	.w3(32'h3ab7d617),
	.w4(32'h3c07effb),
	.w5(32'h3bdadf6f),
	.w6(32'h3b49152d),
	.w7(32'h3c0343a2),
	.w8(32'h3bc00a62),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd53361),
	.w1(32'hbc8e0ba0),
	.w2(32'hbbfde7e7),
	.w3(32'hbce4cbdb),
	.w4(32'hbd1b6d5a),
	.w5(32'hbcc45bd5),
	.w6(32'hbb21e605),
	.w7(32'hbbbcbd34),
	.w8(32'hbb2e9ac5),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becc0ea),
	.w1(32'h3b365b21),
	.w2(32'hbb85fada),
	.w3(32'hbbceb9c7),
	.w4(32'hbc1d8715),
	.w5(32'hbc21c1d5),
	.w6(32'h3bd699e2),
	.w7(32'hbb549854),
	.w8(32'h3b64d883),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39661ccd),
	.w1(32'h3a9c21b1),
	.w2(32'h3a577518),
	.w3(32'hbaf44e9b),
	.w4(32'h395e89c1),
	.w5(32'h3aeecc57),
	.w6(32'hb9312e5a),
	.w7(32'hbab829fd),
	.w8(32'h3b25d9fd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1a391),
	.w1(32'hbbaf26eb),
	.w2(32'hbbc8b202),
	.w3(32'h378fa48b),
	.w4(32'hbba9b404),
	.w5(32'hbb9bc45e),
	.w6(32'hbaf23ee0),
	.w7(32'hbaff77fd),
	.w8(32'h3ac76ac2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d92e4),
	.w1(32'hbc131031),
	.w2(32'hbb483b26),
	.w3(32'hbb3cb89a),
	.w4(32'hba41842f),
	.w5(32'hba2d7846),
	.w6(32'h3ab99430),
	.w7(32'h3bd9b0c9),
	.w8(32'hbb46b2c7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f910),
	.w1(32'h3ad3daa1),
	.w2(32'h3b9bc1d2),
	.w3(32'hbafb5f35),
	.w4(32'h3b007721),
	.w5(32'h3b6b7026),
	.w6(32'hbb821c65),
	.w7(32'h3b061f7b),
	.w8(32'h3b99e383),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8143e4),
	.w1(32'hbb9dc046),
	.w2(32'hb8961c69),
	.w3(32'hbb004245),
	.w4(32'hbc013fc7),
	.w5(32'hbbb8d6d7),
	.w6(32'h3a707845),
	.w7(32'hb95f0458),
	.w8(32'h3a515a27),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab892d1),
	.w1(32'hbbadaa62),
	.w2(32'hbac67323),
	.w3(32'hbb6e2c68),
	.w4(32'hbba79a38),
	.w5(32'hbae2f5e8),
	.w6(32'hba4eb843),
	.w7(32'h3b92a724),
	.w8(32'hb9de0b67),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8938f3),
	.w1(32'h3bbea0d9),
	.w2(32'h3aea1437),
	.w3(32'hb911a3e6),
	.w4(32'h3878f6f1),
	.w5(32'h39d3fd61),
	.w6(32'h3b2946ab),
	.w7(32'h3abac8f0),
	.w8(32'h3b0b8333),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bc7ba),
	.w1(32'hbbe12354),
	.w2(32'hbb03673d),
	.w3(32'h39963ede),
	.w4(32'h3a738d92),
	.w5(32'h3a728491),
	.w6(32'hbbd5fc58),
	.w7(32'hbb430282),
	.w8(32'hbbab3de5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc30dd9),
	.w1(32'hbbd92d02),
	.w2(32'hbb69ade6),
	.w3(32'hbb66e69f),
	.w4(32'hbb60eccb),
	.w5(32'hbadc7394),
	.w6(32'hbb9cf247),
	.w7(32'hbb377c62),
	.w8(32'hba6b9f27),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba244007),
	.w1(32'hbba7a186),
	.w2(32'hbb46c327),
	.w3(32'hba8b5fe0),
	.w4(32'hbba72465),
	.w5(32'hbbbe94e4),
	.w6(32'h3b1d3ab5),
	.w7(32'h395e344d),
	.w8(32'h3ae05a79),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd44f92),
	.w1(32'hbbed598c),
	.w2(32'hbadd9d89),
	.w3(32'hbc2f6103),
	.w4(32'hbc5d188c),
	.w5(32'hbb3eb939),
	.w6(32'hbb81a5ae),
	.w7(32'hbad9b955),
	.w8(32'hbba0b7d6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a377443),
	.w1(32'h39d134d2),
	.w2(32'h39f052d5),
	.w3(32'h3936f9c7),
	.w4(32'hbaa7fa7b),
	.w5(32'hbaa8703d),
	.w6(32'h39fa54e7),
	.w7(32'hb90c4d99),
	.w8(32'hb83423d5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8052b1),
	.w1(32'hbb1c8c66),
	.w2(32'hbaa72a32),
	.w3(32'hbb3967f5),
	.w4(32'hbb7ba72b),
	.w5(32'hbb68938b),
	.w6(32'hb9e152c5),
	.w7(32'hba96643e),
	.w8(32'hbb30bf3a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc15614),
	.w1(32'hbbbe6c92),
	.w2(32'hbb5d6e81),
	.w3(32'hbbfad64d),
	.w4(32'hbbf0a9de),
	.w5(32'hbbf7388b),
	.w6(32'hbbe7cd3c),
	.w7(32'hbbb16180),
	.w8(32'hbb7d1a49),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa81c4b),
	.w1(32'hbb1a8ab4),
	.w2(32'h38a7e330),
	.w3(32'h3b882773),
	.w4(32'h3b896ace),
	.w5(32'h3bb74a07),
	.w6(32'h3b08b358),
	.w7(32'h3b19da73),
	.w8(32'h3b205f1c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb136f35),
	.w1(32'hbafa5d6c),
	.w2(32'hba21b89d),
	.w3(32'hbb1b49e9),
	.w4(32'hbb0c555d),
	.w5(32'hba291db5),
	.w6(32'hba8effd6),
	.w7(32'hba9115ce),
	.w8(32'h3a9f96e5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be305ee),
	.w1(32'hbc263f27),
	.w2(32'hbbfd966d),
	.w3(32'hbbede4c2),
	.w4(32'hbc7ab036),
	.w5(32'hbc0ea817),
	.w6(32'h3be2d145),
	.w7(32'h3c80dd9f),
	.w8(32'h3bad2846),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab3dda),
	.w1(32'h3a3fba8c),
	.w2(32'h397d1fa3),
	.w3(32'hb7f425e5),
	.w4(32'h38f9fe72),
	.w5(32'hba282d1f),
	.w6(32'h3a0d090d),
	.w7(32'h39947981),
	.w8(32'hb9ea2698),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb446238),
	.w1(32'hbba8a210),
	.w2(32'hba92fca9),
	.w3(32'hbbd4a23b),
	.w4(32'hbbfdb089),
	.w5(32'hbb3dd7a4),
	.w6(32'hba8ecfac),
	.w7(32'hba71b3df),
	.w8(32'h399e8911),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8787df8),
	.w1(32'h3a9fd9b6),
	.w2(32'h3a1b7510),
	.w3(32'hbab30378),
	.w4(32'hba08755d),
	.w5(32'hba37373a),
	.w6(32'hb8f37db8),
	.w7(32'hba1910ea),
	.w8(32'hb9d9af8c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0066c6),
	.w1(32'hbbde0173),
	.w2(32'hbbba8dd4),
	.w3(32'hbc19261d),
	.w4(32'hbbede0a0),
	.w5(32'hbbe49186),
	.w6(32'hbb15b5e1),
	.w7(32'h3b960308),
	.w8(32'hbb194acd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7afc16),
	.w1(32'hbb7fcf6f),
	.w2(32'hbb5af33c),
	.w3(32'hbb658fcf),
	.w4(32'hbb691f78),
	.w5(32'hbb3ecf9a),
	.w6(32'hbb505b63),
	.w7(32'hbb2d48c5),
	.w8(32'hbaf8fea9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb652ca3),
	.w1(32'hbbd045dd),
	.w2(32'hbb94229c),
	.w3(32'hbb511111),
	.w4(32'hbb92e387),
	.w5(32'hbb9c695d),
	.w6(32'h3a9855d1),
	.w7(32'h3a1d5692),
	.w8(32'hbabca79c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0370c4),
	.w1(32'hbae25977),
	.w2(32'hbab00c80),
	.w3(32'hbb02939c),
	.w4(32'hbb01eb2b),
	.w5(32'hbad3d92a),
	.w6(32'hbadaad41),
	.w7(32'hbabfc6d9),
	.w8(32'h38d52021),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a6f8d),
	.w1(32'hbc787a3c),
	.w2(32'hbc02b9d4),
	.w3(32'hbb599f76),
	.w4(32'hbc154d38),
	.w5(32'hbbad605c),
	.w6(32'h3b862fce),
	.w7(32'h3b909794),
	.w8(32'hbb11289c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3c0d1),
	.w1(32'hbb912fdf),
	.w2(32'hbb1b6443),
	.w3(32'hbaf3e565),
	.w4(32'hbabf91f8),
	.w5(32'hbb29c448),
	.w6(32'hbb5d249c),
	.w7(32'hba063ea6),
	.w8(32'h39d96db5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b75a3),
	.w1(32'hbb0f610e),
	.w2(32'hbb07ecba),
	.w3(32'hbb7ba04f),
	.w4(32'hbb5f02a8),
	.w5(32'hbb2d4eed),
	.w6(32'hbaeab54b),
	.w7(32'hbab91fa8),
	.w8(32'hbbfe69ed),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5a6a),
	.w1(32'hbbece148),
	.w2(32'hbba47e2c),
	.w3(32'hbb63ac23),
	.w4(32'hbb08b02f),
	.w5(32'hbae2c4d2),
	.w6(32'hbbca7815),
	.w7(32'hbb689202),
	.w8(32'hbb168cb1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbedd1),
	.w1(32'hbaf65a51),
	.w2(32'h3a9c1be5),
	.w3(32'hbc02c7b5),
	.w4(32'hbc0491c6),
	.w5(32'hbb8c3cbf),
	.w6(32'hbb931a83),
	.w7(32'hbab7f3fd),
	.w8(32'hb9e031bb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f0c58),
	.w1(32'hbb92abb9),
	.w2(32'h3b3022bb),
	.w3(32'hbbe293c9),
	.w4(32'hbbc0b179),
	.w5(32'hba00f3c6),
	.w6(32'h3b811814),
	.w7(32'h3bc0547f),
	.w8(32'h3b13c004),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc2f3),
	.w1(32'h3b81b309),
	.w2(32'hba72e206),
	.w3(32'h3af5703e),
	.w4(32'hbbbcef1e),
	.w5(32'h396f2819),
	.w6(32'h3c547440),
	.w7(32'h3c232586),
	.w8(32'h3bed8d91),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98d8fa),
	.w1(32'hbbc22971),
	.w2(32'h3bba192e),
	.w3(32'hbbdf3a03),
	.w4(32'hbc0973ba),
	.w5(32'hb8def86a),
	.w6(32'h3c4401f1),
	.w7(32'h3c07462d),
	.w8(32'h3b59a279),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafa823),
	.w1(32'hbbb526d6),
	.w2(32'hbbaf4d91),
	.w3(32'hbb89ede0),
	.w4(32'hbc4fd72e),
	.w5(32'hbc29e144),
	.w6(32'h3b8a7395),
	.w7(32'hb9c8f55b),
	.w8(32'h3ba05d04),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c48e9),
	.w1(32'h3ae0860f),
	.w2(32'h3b769cfe),
	.w3(32'h3baf3ef7),
	.w4(32'h3b6926e6),
	.w5(32'h3bb06142),
	.w6(32'h3b8581c1),
	.w7(32'h3b8dc404),
	.w8(32'hbaf8252c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a5cef),
	.w1(32'hbb481913),
	.w2(32'hb92f8622),
	.w3(32'hbb78974e),
	.w4(32'hbb6df5ac),
	.w5(32'hba13a5ec),
	.w6(32'hbb0e6cb1),
	.w7(32'hb982e6f8),
	.w8(32'hbb26996b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881c2e5),
	.w1(32'h3b4d94e4),
	.w2(32'h3ab0b1f8),
	.w3(32'hb897f92e),
	.w4(32'h3aaf6c6a),
	.w5(32'h3ac4113c),
	.w6(32'hba774cff),
	.w7(32'hbb366787),
	.w8(32'h3ba680ae),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcea01f),
	.w1(32'h3936159b),
	.w2(32'h3a80069a),
	.w3(32'h3bb240fa),
	.w4(32'hb73e8059),
	.w5(32'h3b02e792),
	.w6(32'h3bdf5d4f),
	.w7(32'h3b9bbced),
	.w8(32'h3b84dfa4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95da48),
	.w1(32'h3b15621e),
	.w2(32'h3b9d55e7),
	.w3(32'h3b53c9a9),
	.w4(32'hb945b284),
	.w5(32'h3b1060ab),
	.w6(32'h3b14c2b2),
	.w7(32'h3b806e6c),
	.w8(32'h3abfef6c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fde11),
	.w1(32'h3a9aaa2c),
	.w2(32'hba264c14),
	.w3(32'h3abba2d5),
	.w4(32'h3a2647cf),
	.w5(32'hba505589),
	.w6(32'h3997a0c6),
	.w7(32'hba952900),
	.w8(32'hbbe09041),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaeb360),
	.w1(32'hbb35f5fe),
	.w2(32'h3bb6faeb),
	.w3(32'hbc3458ba),
	.w4(32'hbc3d12bd),
	.w5(32'hbb9b0699),
	.w6(32'h39998d1e),
	.w7(32'h3bbdbfce),
	.w8(32'h3b72029f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba882c21),
	.w1(32'hbb3a2dc7),
	.w2(32'h3b0fa3e4),
	.w3(32'hbb91cab6),
	.w4(32'hbbb172d8),
	.w5(32'hbb150a2b),
	.w6(32'hbaf566b6),
	.w7(32'hbb243e10),
	.w8(32'hbbcc1b2e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d8f2),
	.w1(32'hbb6e9c42),
	.w2(32'h3b07d3d0),
	.w3(32'h3aafb078),
	.w4(32'h3b58b405),
	.w5(32'h3bf0cb93),
	.w6(32'hbbdc0c04),
	.w7(32'hbbbb0f8a),
	.w8(32'h3bdf2ab7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf69774),
	.w1(32'h3c1126b2),
	.w2(32'h3c070f14),
	.w3(32'h3bfc6010),
	.w4(32'h3c0ada61),
	.w5(32'h3c128299),
	.w6(32'h3c3ed1a1),
	.w7(32'h3c33c8e0),
	.w8(32'h3bcc5f08),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a4c00),
	.w1(32'hbc795f68),
	.w2(32'hbbb68e89),
	.w3(32'hbc162c8a),
	.w4(32'hbc3c66ca),
	.w5(32'hbb5f9fac),
	.w6(32'h3bf53b66),
	.w7(32'h3b40a9be),
	.w8(32'h3bf2288c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6eae4a),
	.w1(32'h3abb926c),
	.w2(32'h39e3af8a),
	.w3(32'hba00b794),
	.w4(32'hbb81cbda),
	.w5(32'hbb145606),
	.w6(32'h3ac6126e),
	.w7(32'hbb0fc217),
	.w8(32'h37c9bef1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdde7a),
	.w1(32'hbb45ff98),
	.w2(32'hba18719c),
	.w3(32'h37dd7e7e),
	.w4(32'hbac21626),
	.w5(32'hb8dc7438),
	.w6(32'hbafe7c55),
	.w7(32'h3a3b36ab),
	.w8(32'hbad6b9a5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e9f27),
	.w1(32'hba6dcabd),
	.w2(32'h39556b82),
	.w3(32'hbb1f4f26),
	.w4(32'hbac64ef2),
	.w5(32'hba13453e),
	.w6(32'hba8694d5),
	.w7(32'hb753c411),
	.w8(32'hbabcf115),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb175567),
	.w1(32'hbb01455a),
	.w2(32'hba9a2295),
	.w3(32'hbacc0962),
	.w4(32'hbabe677b),
	.w5(32'hb9c203db),
	.w6(32'hbaefd9a9),
	.w7(32'hbb0294d7),
	.w8(32'hbb70b742),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb45f0e),
	.w1(32'hbbbf2c45),
	.w2(32'hbbcb532e),
	.w3(32'hbbaa2c23),
	.w4(32'hbbabf003),
	.w5(32'hbbc79961),
	.w6(32'hbac31ea6),
	.w7(32'hbab167b3),
	.w8(32'hbacc829f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad49cf),
	.w1(32'hbbb01814),
	.w2(32'hbb85ccd7),
	.w3(32'hbb7738ea),
	.w4(32'hbb8154c7),
	.w5(32'hbb682bd5),
	.w6(32'hbb9225d6),
	.w7(32'hbae6e1c8),
	.w8(32'h3ba5f993),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c112f44),
	.w1(32'h3c378d2e),
	.w2(32'h3c1fe545),
	.w3(32'h3a35f7fe),
	.w4(32'h3b3fb11c),
	.w5(32'h3b62f637),
	.w6(32'h3acdc4b7),
	.w7(32'h3b32e241),
	.w8(32'h3bcb32cf),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add15bb),
	.w1(32'h3aeab664),
	.w2(32'h3af71037),
	.w3(32'h3ac3857d),
	.w4(32'h3a7fc465),
	.w5(32'h3adff790),
	.w6(32'h39eefd07),
	.w7(32'h39d79b62),
	.w8(32'hb9030dd1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8610),
	.w1(32'hbb8bbb70),
	.w2(32'hba139150),
	.w3(32'hbc2164f7),
	.w4(32'hbc59bec5),
	.w5(32'hbbeabc73),
	.w6(32'hb92a9b37),
	.w7(32'h3abd66b2),
	.w8(32'h3a83a21b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6ac8b),
	.w1(32'hbb3ba5f5),
	.w2(32'hbad53c4f),
	.w3(32'h3b1b9f63),
	.w4(32'hbae7920e),
	.w5(32'hbad01f8f),
	.w6(32'h3bd12012),
	.w7(32'h3b431edc),
	.w8(32'h39d99384),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9329e7f),
	.w1(32'hb7f85d6d),
	.w2(32'h3a495073),
	.w3(32'hbb877ada),
	.w4(32'hbb56b151),
	.w5(32'hbb1614a4),
	.w6(32'hbb1a0427),
	.w7(32'hbb127c76),
	.w8(32'hb9897e44),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1041bc),
	.w1(32'h3b3d4578),
	.w2(32'h3ac7147f),
	.w3(32'h3b3427fe),
	.w4(32'h3b3ba7df),
	.w5(32'h3b11a1be),
	.w6(32'h3afa312b),
	.w7(32'h3ae45eff),
	.w8(32'h3b078e87),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01068e),
	.w1(32'hbc0761ba),
	.w2(32'hbb74f908),
	.w3(32'hbb933a7f),
	.w4(32'hbb8f507c),
	.w5(32'hbb01574d),
	.w6(32'h397ffe37),
	.w7(32'h3a0cd257),
	.w8(32'h3a4a69b8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034dda),
	.w1(32'h3ab3e327),
	.w2(32'h3b3d4faf),
	.w3(32'h3b2c55a4),
	.w4(32'h3b832c0a),
	.w5(32'h3b8d3274),
	.w6(32'h3b6ab3ca),
	.w7(32'h3b877666),
	.w8(32'h3bccb7db),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb551e2),
	.w1(32'hbb06c065),
	.w2(32'hba7d9e61),
	.w3(32'hbb1d4b72),
	.w4(32'h3a6e6e13),
	.w5(32'hb89146b2),
	.w6(32'h3940a9cc),
	.w7(32'h3b088865),
	.w8(32'h39cc6dd6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d46858),
	.w1(32'h3b6b3a65),
	.w2(32'h3af9c9d8),
	.w3(32'h3a9a330f),
	.w4(32'h3b5eb703),
	.w5(32'h39ff5371),
	.w6(32'hba9fccad),
	.w7(32'h3ac607b8),
	.w8(32'hb774eb2c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3874373b),
	.w1(32'hb9f83f53),
	.w2(32'hb936c9fa),
	.w3(32'h392ee8c1),
	.w4(32'hb9fb4b43),
	.w5(32'hb945b51d),
	.w6(32'hb883d9d5),
	.w7(32'hba3a76df),
	.w8(32'hba064c84),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba164b94),
	.w1(32'hba36399a),
	.w2(32'hba62c96a),
	.w3(32'hba28adfd),
	.w4(32'hbb0fcc54),
	.w5(32'hba909037),
	.w6(32'hb9cfd98e),
	.w7(32'hba38def8),
	.w8(32'hb9b97646),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba561cf4),
	.w1(32'hbaadb938),
	.w2(32'hbae6a0fa),
	.w3(32'hbacd4502),
	.w4(32'hbaa7f6e1),
	.w5(32'hbaac93a3),
	.w6(32'h3a051e36),
	.w7(32'h3935a70f),
	.w8(32'hb8762399),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4b4e0),
	.w1(32'h3adaeb5a),
	.w2(32'h3a6e5004),
	.w3(32'h3a2b44f9),
	.w4(32'h3a402123),
	.w5(32'h39981e46),
	.w6(32'h3ae406b0),
	.w7(32'h3b3236cd),
	.w8(32'h3b2c87d9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6737bc),
	.w1(32'hba9da133),
	.w2(32'h3808d7e2),
	.w3(32'hbb233910),
	.w4(32'hbb08832b),
	.w5(32'hba86be53),
	.w6(32'h390b6936),
	.w7(32'h3b0b2147),
	.w8(32'h3a220945),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f27fa4),
	.w1(32'hb2456b46),
	.w2(32'h37504d67),
	.w3(32'h37c08b3a),
	.w4(32'h36b2df42),
	.w5(32'h38134394),
	.w6(32'hb697ec54),
	.w7(32'hb69fe036),
	.w8(32'h37da8cdc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5d9ff),
	.w1(32'h389922f0),
	.w2(32'hb8bc8ca9),
	.w3(32'hb656e887),
	.w4(32'h39970382),
	.w5(32'h396962df),
	.w6(32'hb839333b),
	.w7(32'hb87b6477),
	.w8(32'hb94a7961),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba949ee),
	.w1(32'h3bb5ebc4),
	.w2(32'h3b855e68),
	.w3(32'hbb515da2),
	.w4(32'hbb99977b),
	.w5(32'hbb5ee8c5),
	.w6(32'hbb3186db),
	.w7(32'hb9c82194),
	.w8(32'h3a59fc90),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07f896),
	.w1(32'hbc083ad0),
	.w2(32'hbc0f479d),
	.w3(32'h3b19bfa7),
	.w4(32'hbb2eb047),
	.w5(32'hbb8d797f),
	.w6(32'h3bd5e11e),
	.w7(32'h3b0df717),
	.w8(32'hbb1f94b9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3334),
	.w1(32'hba82727f),
	.w2(32'hba81ef02),
	.w3(32'hba822f2d),
	.w4(32'hb563d22f),
	.w5(32'hba28ca4d),
	.w6(32'hb922eef5),
	.w7(32'h3970b824),
	.w8(32'hb7244a17),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d2bb),
	.w1(32'h3b5c772e),
	.w2(32'hba012093),
	.w3(32'h3b4bc680),
	.w4(32'h3b78eeb2),
	.w5(32'h39a6785a),
	.w6(32'h3960c080),
	.w7(32'h39f0a31a),
	.w8(32'hbaee8da1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ad8aa),
	.w1(32'hbaa4191c),
	.w2(32'hba03bc8d),
	.w3(32'hbb670708),
	.w4(32'hba4768e9),
	.w5(32'hb95414f6),
	.w6(32'hba13fc8c),
	.w7(32'h3a23855d),
	.w8(32'h3a70f324),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ee397),
	.w1(32'hb982a410),
	.w2(32'h3a7cb964),
	.w3(32'hbacf98fd),
	.w4(32'h3a3acd48),
	.w5(32'h3ac546c9),
	.w6(32'h3ac3f10f),
	.w7(32'h3aaa9f3b),
	.w8(32'h3aba028e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb144175),
	.w1(32'hbb2945e8),
	.w2(32'hbb3424bf),
	.w3(32'hb9c80ea2),
	.w4(32'h3a86695a),
	.w5(32'hba9a580d),
	.w6(32'h3ad0ef21),
	.w7(32'h3b0f9246),
	.w8(32'h3a69cba3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec3f74),
	.w1(32'hba37c1bf),
	.w2(32'hbab40d5a),
	.w3(32'hba472827),
	.w4(32'h3a9d163e),
	.w5(32'h3a620d8f),
	.w6(32'h3a6ec856),
	.w7(32'h3b844ad5),
	.w8(32'h3b1e3375),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule