module layer_6_featuremap_36(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56a665),
	.w1(32'h3986f845),
	.w2(32'h3af746ee),
	.w3(32'hbb96087a),
	.w4(32'hba432267),
	.w5(32'h3b03ad8a),
	.w6(32'hbac498ad),
	.w7(32'h3b9b53e4),
	.w8(32'h3b36bae2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a579e17),
	.w1(32'h3af9c6d8),
	.w2(32'h3b9c2e7d),
	.w3(32'h3b8cf01a),
	.w4(32'h3b4521e6),
	.w5(32'hbad0c111),
	.w6(32'h3c211ae7),
	.w7(32'h3be25b19),
	.w8(32'h3bbee45c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93cc9a),
	.w1(32'h3c74090b),
	.w2(32'h3ce5d5cc),
	.w3(32'hbcff094c),
	.w4(32'h3ba81fb5),
	.w5(32'h3a98d764),
	.w6(32'hbcd22302),
	.w7(32'h3d44063b),
	.w8(32'hbcc750db),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28927d),
	.w1(32'h3b65d876),
	.w2(32'hbac5a534),
	.w3(32'hb9b9b616),
	.w4(32'hbb173711),
	.w5(32'hbaaa88c8),
	.w6(32'h3b8709a6),
	.w7(32'hb8b8e7d8),
	.w8(32'hbb21e5f0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6661a),
	.w1(32'h3b4f6b49),
	.w2(32'hba14edeb),
	.w3(32'hbc540f24),
	.w4(32'h3c91af39),
	.w5(32'hbb24c770),
	.w6(32'h3b1dcf27),
	.w7(32'h3c8a5464),
	.w8(32'hbc989778),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca26747),
	.w1(32'hbb93c952),
	.w2(32'h39a6f501),
	.w3(32'hbba01ded),
	.w4(32'hbbf766d9),
	.w5(32'hba0eaab1),
	.w6(32'hbc286fd5),
	.w7(32'hbb57ab69),
	.w8(32'h3b1e543b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b350dc9),
	.w1(32'hbaf48381),
	.w2(32'hbbbb6512),
	.w3(32'h3b9e5cd5),
	.w4(32'h3a33fad8),
	.w5(32'h3ade7650),
	.w6(32'h3c124ff9),
	.w7(32'hbb486630),
	.w8(32'h3a9391bb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c997f3),
	.w1(32'hbccb502d),
	.w2(32'hbc9fbafc),
	.w3(32'h3cfdb1a9),
	.w4(32'hbc32b0c9),
	.w5(32'hbc45eb52),
	.w6(32'h3c089663),
	.w7(32'hbd684d65),
	.w8(32'hbc3e302d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29b3cb),
	.w1(32'h3c3eba1c),
	.w2(32'hbc6e932b),
	.w3(32'h3a0592d2),
	.w4(32'h3af41ca7),
	.w5(32'hbb1bd64f),
	.w6(32'h3c2ec0eb),
	.w7(32'h3c5efc8f),
	.w8(32'hbb893e87),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b0167),
	.w1(32'h3b281183),
	.w2(32'h3b13a725),
	.w3(32'hbba00d5f),
	.w4(32'hbb15cda1),
	.w5(32'hba117852),
	.w6(32'hbb27af2d),
	.w7(32'h3b815fad),
	.w8(32'hb8978ec0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab65c1f),
	.w1(32'h3c57583f),
	.w2(32'h3c694606),
	.w3(32'hbca49549),
	.w4(32'h3ce93d0c),
	.w5(32'hbaa3a9da),
	.w6(32'hba7c575a),
	.w7(32'h3d21cf33),
	.w8(32'hbcdf812e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0323f),
	.w1(32'h3aa64f77),
	.w2(32'h3b716964),
	.w3(32'hbc2a78b0),
	.w4(32'h3c05678e),
	.w5(32'hbc0df699),
	.w6(32'hba8c2a4a),
	.w7(32'h3af4c635),
	.w8(32'hbbc44e43),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35d7d0),
	.w1(32'hbc0c1807),
	.w2(32'h3c3c7239),
	.w3(32'hbbb8422e),
	.w4(32'h3c1325f2),
	.w5(32'hbbc460db),
	.w6(32'hbbfd97ff),
	.w7(32'h3c1f9a52),
	.w8(32'hbae2e521),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6fbc4),
	.w1(32'h3b46bcac),
	.w2(32'h3c16e2f6),
	.w3(32'hbc17a5c9),
	.w4(32'hbb8f31f8),
	.w5(32'h3a6cd6c3),
	.w6(32'hbbc0464b),
	.w7(32'h3bd683d6),
	.w8(32'h3be26e6f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ed851),
	.w1(32'hbbb1ce75),
	.w2(32'hbb9e3ca4),
	.w3(32'h3b3873e9),
	.w4(32'hb9772b39),
	.w5(32'hbc3037bb),
	.w6(32'hbb08856b),
	.w7(32'hbbf72a9d),
	.w8(32'hbc616ef3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe9ee1),
	.w1(32'hbb2a2abf),
	.w2(32'h3a1d5eb2),
	.w3(32'hbb1a8c3a),
	.w4(32'hbb90ac97),
	.w5(32'h3b3017fd),
	.w6(32'hbc0185f5),
	.w7(32'hbab63d57),
	.w8(32'h3afae9f0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39247832),
	.w1(32'h3c8a339d),
	.w2(32'hbab719ef),
	.w3(32'hbb029bd7),
	.w4(32'h3cad3e6a),
	.w5(32'hbcd545b5),
	.w6(32'h3bf89b51),
	.w7(32'h3cb77154),
	.w8(32'hbd106888),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82eef4),
	.w1(32'hbac82798),
	.w2(32'h3b9e5034),
	.w3(32'hbb99e32c),
	.w4(32'h3a9dba18),
	.w5(32'h3b85303a),
	.w6(32'hbad7a041),
	.w7(32'h3bd11416),
	.w8(32'h3b8b5524),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95a7b2),
	.w1(32'h3a809a67),
	.w2(32'h3a075382),
	.w3(32'h3b643387),
	.w4(32'hbb8a90ed),
	.w5(32'hbb271c10),
	.w6(32'hba7c9477),
	.w7(32'hbb4001fa),
	.w8(32'hba643523),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d02499),
	.w1(32'hb9d73639),
	.w2(32'hbca4aa12),
	.w3(32'hbb001d8b),
	.w4(32'hbca348b0),
	.w5(32'hbc80d281),
	.w6(32'hbbcce900),
	.w7(32'hbcbbcb16),
	.w8(32'hbb84afa5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cd72a),
	.w1(32'h3a094350),
	.w2(32'hbbb8e80f),
	.w3(32'hb9aa0a0d),
	.w4(32'hbb1a1d6b),
	.w5(32'hbb074b6c),
	.w6(32'h39d4856a),
	.w7(32'hbba5c52e),
	.w8(32'hbb1b9a04),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5a69f),
	.w1(32'h3c74e5c4),
	.w2(32'hbb9b088a),
	.w3(32'hbb229fd0),
	.w4(32'h3bb65f19),
	.w5(32'h3b56dac2),
	.w6(32'h3c8ad2d9),
	.w7(32'h3c313d1e),
	.w8(32'hbbb1088a),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097150),
	.w1(32'h3cc3cfea),
	.w2(32'hbb541b5f),
	.w3(32'h39f7638c),
	.w4(32'h3cca1977),
	.w5(32'hbc140907),
	.w6(32'h3d0c6c9b),
	.w7(32'h3d0146c5),
	.w8(32'hbd1b9cbb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd127ef3),
	.w1(32'hbc0e71b5),
	.w2(32'hbc9e0dbf),
	.w3(32'h3d1869e0),
	.w4(32'hbccc6013),
	.w5(32'hbc8e3395),
	.w6(32'h3c7404bb),
	.w7(32'hbd229d04),
	.w8(32'hbbcc84f4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81223a),
	.w1(32'h3ac65d9c),
	.w2(32'hbb4dc4a7),
	.w3(32'hbc33a5bc),
	.w4(32'hbbb34464),
	.w5(32'h3b29ec69),
	.w6(32'h3a8fbb7f),
	.w7(32'h3bb7acbf),
	.w8(32'h3c011f91),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b66b5),
	.w1(32'hbbe55b58),
	.w2(32'hbc3a7d03),
	.w3(32'hbbcc9e95),
	.w4(32'h3aef4f8b),
	.w5(32'hbcb31f93),
	.w6(32'h3b6e7478),
	.w7(32'hbb6a3345),
	.w8(32'hbcb83b0d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4ef4b),
	.w1(32'h3c363e37),
	.w2(32'h3b6c98c7),
	.w3(32'hbc564cc8),
	.w4(32'hbb65a7fd),
	.w5(32'h3bbb9952),
	.w6(32'hbab66a58),
	.w7(32'h3c83f2c9),
	.w8(32'hba2ab7d9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07d955),
	.w1(32'hb9c8370c),
	.w2(32'h3aac3e76),
	.w3(32'h3c21b5b7),
	.w4(32'h3a4c9040),
	.w5(32'h3b36e840),
	.w6(32'h3b66b17f),
	.w7(32'hbbada857),
	.w8(32'h3bb0dd2b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a5b6f),
	.w1(32'h3b430a01),
	.w2(32'h39a46839),
	.w3(32'h3b85cb73),
	.w4(32'h3b14aba1),
	.w5(32'hbaa71152),
	.w6(32'h3b8c055d),
	.w7(32'hb8faf02a),
	.w8(32'hbafb8df6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c8e5),
	.w1(32'h3c5b32a1),
	.w2(32'h3b457de7),
	.w3(32'hbc2b9efe),
	.w4(32'hbbb9ad5a),
	.w5(32'h388c8cb4),
	.w6(32'h3bc35963),
	.w7(32'h3bb1bd57),
	.w8(32'h3b1cc182),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01aa7c),
	.w1(32'hbc861e4a),
	.w2(32'hbc42dfb4),
	.w3(32'h39b86d5b),
	.w4(32'hbc1e7c0c),
	.w5(32'h3b6999f9),
	.w6(32'hbc1dd45c),
	.w7(32'hbcd6454e),
	.w8(32'hba99a089),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a137b),
	.w1(32'hbc299f65),
	.w2(32'h3cd8ecc5),
	.w3(32'hbc378f0a),
	.w4(32'hbc413d1b),
	.w5(32'h39d68ae7),
	.w6(32'hbce51783),
	.w7(32'h3bccaa38),
	.w8(32'h3cd45334),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8e71d),
	.w1(32'h3cc157cd),
	.w2(32'hbbcdd6a3),
	.w3(32'h3bc6b066),
	.w4(32'h3d378186),
	.w5(32'hbc0ac20d),
	.w6(32'h3ce5b0cc),
	.w7(32'h3bf511dc),
	.w8(32'hbccf0d04),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce92c6f),
	.w1(32'h3b878609),
	.w2(32'h3c7b85f6),
	.w3(32'h3b1bb5b3),
	.w4(32'h3bdcef0f),
	.w5(32'h3afad9ed),
	.w6(32'h3b81460b),
	.w7(32'h3caaa80b),
	.w8(32'h3b820770),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90689b),
	.w1(32'h3a5b1aef),
	.w2(32'hbba25cf1),
	.w3(32'h3a3c1733),
	.w4(32'h39951a51),
	.w5(32'hbbb93bb5),
	.w6(32'h3baf5ac2),
	.w7(32'hbb00853d),
	.w8(32'hbbf7ef44),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0217a8),
	.w1(32'h3b4c368b),
	.w2(32'h3b8de302),
	.w3(32'hbc59324d),
	.w4(32'h3b740a95),
	.w5(32'h3b282061),
	.w6(32'hbb6480bb),
	.w7(32'h3c207374),
	.w8(32'h3bac938e),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afc3e5),
	.w1(32'h3a317a03),
	.w2(32'h3bbdb4a9),
	.w3(32'hbbbbab90),
	.w4(32'h3ad9e13d),
	.w5(32'hbac7ff4f),
	.w6(32'hbb0f909e),
	.w7(32'h3bb0b935),
	.w8(32'h3b9000e4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bbb21),
	.w1(32'h3ba7f2d6),
	.w2(32'h3b4b2d6d),
	.w3(32'h3bc186de),
	.w4(32'h3a9d9d99),
	.w5(32'hbab81419),
	.w6(32'h3bd5489a),
	.w7(32'h39943914),
	.w8(32'hb8db8358),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0170ca),
	.w1(32'h3c1a950d),
	.w2(32'hbb11251d),
	.w3(32'hbaea3388),
	.w4(32'h3c5f0cc7),
	.w5(32'h3bcb0b0f),
	.w6(32'h3c1eb389),
	.w7(32'h3cae9a38),
	.w8(32'hbc1cc85d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3c036),
	.w1(32'h3bdd5a56),
	.w2(32'h3cea9873),
	.w3(32'hbc98aa74),
	.w4(32'h3b407831),
	.w5(32'h3c6e6fe2),
	.w6(32'hbc9f084d),
	.w7(32'h3d14d298),
	.w8(32'h3c8dd258),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b2c88),
	.w1(32'hbb10c502),
	.w2(32'hbd1515ff),
	.w3(32'h3d01f938),
	.w4(32'h3c64fa87),
	.w5(32'hbc8bd627),
	.w6(32'h3d088990),
	.w7(32'hbd2837d6),
	.w8(32'hbc8188d5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c990968),
	.w1(32'h3b91360c),
	.w2(32'hbb14e3cd),
	.w3(32'h3afeb2d2),
	.w4(32'hbb1181ee),
	.w5(32'hbb212d33),
	.w6(32'h3baefe8f),
	.w7(32'hbae05d76),
	.w8(32'hbb1b6d03),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c90ddf),
	.w1(32'h3b9f2f8b),
	.w2(32'h3b0e767b),
	.w3(32'hb956a5cd),
	.w4(32'h3be3f5d7),
	.w5(32'h3b2c4556),
	.w6(32'h3bc40997),
	.w7(32'h3c3ac5d5),
	.w8(32'h39aefd0b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e207c0),
	.w1(32'hbc360f8d),
	.w2(32'hbc1d7399),
	.w3(32'h3b80941a),
	.w4(32'hba631e55),
	.w5(32'hbb8a04fe),
	.w6(32'hbba34598),
	.w7(32'hbc0a43a7),
	.w8(32'hbc150b5d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e323f),
	.w1(32'h3ac154a8),
	.w2(32'h3ba91d38),
	.w3(32'hbbb280b3),
	.w4(32'hbb8ff197),
	.w5(32'hbb51dae4),
	.w6(32'hbb4d2ec8),
	.w7(32'hba1d9fa9),
	.w8(32'h3b5290ef),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a14a),
	.w1(32'h3cd14750),
	.w2(32'hbd1bdf49),
	.w3(32'hbc81c1ec),
	.w4(32'h3cb12d5d),
	.w5(32'h3b032152),
	.w6(32'h3d17aa90),
	.w7(32'h3d07ca6a),
	.w8(32'hbd5ce73a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd779e44),
	.w1(32'hbae37cfa),
	.w2(32'hbb944858),
	.w3(32'h3c273430),
	.w4(32'hbb3365ab),
	.w5(32'hbb4c6412),
	.w6(32'h3c3c17cf),
	.w7(32'hbc06b1af),
	.w8(32'h3aff87f8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139255),
	.w1(32'h3be734d1),
	.w2(32'hbcea844b),
	.w3(32'hbc99b97f),
	.w4(32'h3c936b67),
	.w5(32'hbca44f40),
	.w6(32'hbba9af11),
	.w7(32'h3cead941),
	.w8(32'hbd38a3d8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd38628e),
	.w1(32'hbbd9482b),
	.w2(32'hba96a655),
	.w3(32'hbbfa7145),
	.w4(32'hbbdf6d27),
	.w5(32'hbb95318e),
	.w6(32'hbba79016),
	.w7(32'hbba83456),
	.w8(32'h3ae8a2e3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b795729),
	.w1(32'h3c2c117f),
	.w2(32'hbb267411),
	.w3(32'hbcca6dd7),
	.w4(32'hbba71505),
	.w5(32'h3cc286bf),
	.w6(32'hbc511402),
	.w7(32'h3d1f74e7),
	.w8(32'h3c5e8b31),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dbb34),
	.w1(32'hba09f20b),
	.w2(32'hbbb465ce),
	.w3(32'hbb963bf8),
	.w4(32'hbb9b0712),
	.w5(32'hbb8c44f8),
	.w6(32'h39c7a211),
	.w7(32'hbb8dce1b),
	.w8(32'hbbaec5a3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba32cb6),
	.w1(32'hbb283013),
	.w2(32'hbca4feae),
	.w3(32'h3bd457d4),
	.w4(32'hbc72674a),
	.w5(32'hbca54bae),
	.w6(32'h3bd6ca4a),
	.w7(32'hbcaad1af),
	.w8(32'hbc9cd2ef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e616),
	.w1(32'h3b0fba3a),
	.w2(32'hbb8e3fef),
	.w3(32'hba0f11fb),
	.w4(32'hbbf6105c),
	.w5(32'hbb484b91),
	.w6(32'h3a0278be),
	.w7(32'hbbe216f5),
	.w8(32'hbaa5788d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19756f),
	.w1(32'h3c01a852),
	.w2(32'hbb4cfb07),
	.w3(32'h3c272103),
	.w4(32'h3b1919ac),
	.w5(32'hb8fee757),
	.w6(32'h3c36b3a5),
	.w7(32'hbb653aab),
	.w8(32'hbb69abb2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac3aec),
	.w1(32'h3b196729),
	.w2(32'hbaf90f76),
	.w3(32'hbb05a225),
	.w4(32'hbbc54575),
	.w5(32'hbad707cc),
	.w6(32'h3b1e8bf8),
	.w7(32'hbb781847),
	.w8(32'hbb27e554),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87bbe4),
	.w1(32'h3910551a),
	.w2(32'h3ba18199),
	.w3(32'h3ba3e04a),
	.w4(32'h3bcf4b83),
	.w5(32'h3bb3b942),
	.w6(32'h3bd8bf27),
	.w7(32'h3c011d4e),
	.w8(32'h3ba07f75),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d608d),
	.w1(32'h3bde8cce),
	.w2(32'h3bd08920),
	.w3(32'hb9aadee3),
	.w4(32'hba8000ef),
	.w5(32'h3b954edd),
	.w6(32'h3a0f8736),
	.w7(32'hbaf8ccf6),
	.w8(32'h3ba8556f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0474c6),
	.w1(32'hbb7dfef0),
	.w2(32'hbbc735f4),
	.w3(32'hbbe067fb),
	.w4(32'h3b782da4),
	.w5(32'hb8988ed4),
	.w6(32'hbb407d68),
	.w7(32'hbb5b30c4),
	.w8(32'h3b10f635),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba438f1d),
	.w1(32'h3a76ea82),
	.w2(32'h3c2e5004),
	.w3(32'hba13bb92),
	.w4(32'h3be3845e),
	.w5(32'h3bb7b2e1),
	.w6(32'h3b1a2e10),
	.w7(32'h3c5856ee),
	.w8(32'h3c31b07b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8afdd),
	.w1(32'hbbaba0e4),
	.w2(32'h3a98afdb),
	.w3(32'hbba7440e),
	.w4(32'hbb955bd6),
	.w5(32'hbbbebc3c),
	.w6(32'hbc3f71f2),
	.w7(32'hbbe2c0e4),
	.w8(32'hbb492340),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba237ce),
	.w1(32'h3a61f2b9),
	.w2(32'h3aa1fb54),
	.w3(32'h3a00efe1),
	.w4(32'h3afd9807),
	.w5(32'h3a0201eb),
	.w6(32'h3ab82eb9),
	.w7(32'h3b32dcb7),
	.w8(32'h3ae65dbd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacf997),
	.w1(32'h3c954ed5),
	.w2(32'h3bf360fe),
	.w3(32'h3c42e962),
	.w4(32'h3c256848),
	.w5(32'h3c864142),
	.w6(32'h3c584696),
	.w7(32'h3c1bdc3a),
	.w8(32'h3c514aca),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247b99),
	.w1(32'hbc1a8e20),
	.w2(32'hbb5d2b78),
	.w3(32'hbb7e1ccf),
	.w4(32'h3a52ace4),
	.w5(32'h3c0686f3),
	.w6(32'hbc9a3a61),
	.w7(32'h3affc19b),
	.w8(32'h3bd60960),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa24c45),
	.w1(32'hbbddfb9d),
	.w2(32'hbbbb9256),
	.w3(32'hbc973b10),
	.w4(32'hbc53c889),
	.w5(32'hbbf9bfbb),
	.w6(32'hbc76306b),
	.w7(32'hbc59bd1d),
	.w8(32'hbbada100),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule