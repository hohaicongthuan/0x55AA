module layer_10_featuremap_290(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c8540),
	.w1(32'h3bdc5c21),
	.w2(32'h3c83d8bc),
	.w3(32'hbc1290c4),
	.w4(32'h3c2adab5),
	.w5(32'hbc93b3c0),
	.w6(32'hbc78c8fe),
	.w7(32'h3b403b14),
	.w8(32'hba8ec96d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c824fe2),
	.w1(32'hba9aca7c),
	.w2(32'hbc5f27d1),
	.w3(32'hbbec8de2),
	.w4(32'h3bc5f3f8),
	.w5(32'h39dd7c02),
	.w6(32'hbcf2d23a),
	.w7(32'h3ac26c45),
	.w8(32'h3adc4756),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16fd75),
	.w1(32'hbb89a21b),
	.w2(32'hbbb43447),
	.w3(32'h39c58d9a),
	.w4(32'h3bb729cc),
	.w5(32'h3b4b0366),
	.w6(32'hbc440c0e),
	.w7(32'h3a0f742e),
	.w8(32'h3acbc9b5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b29f9),
	.w1(32'h3ad9476d),
	.w2(32'h3a3f64ed),
	.w3(32'h3be425c0),
	.w4(32'h3b5f87ae),
	.w5(32'hbb88b859),
	.w6(32'hbbfc04e2),
	.w7(32'h3aa1fd33),
	.w8(32'h3b5c0b53),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbf75e),
	.w1(32'hbb945908),
	.w2(32'hbbbea0fc),
	.w3(32'h3b561512),
	.w4(32'hbb219903),
	.w5(32'h3c525be1),
	.w6(32'h3c780d71),
	.w7(32'h3bc05d73),
	.w8(32'hbba55885),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42ece5),
	.w1(32'hbab6e867),
	.w2(32'h3c499435),
	.w3(32'h3bd45514),
	.w4(32'h3c8eccbe),
	.w5(32'h3bcacff6),
	.w6(32'hbce5ac8b),
	.w7(32'h3b264f36),
	.w8(32'h3bee39dd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab03a1),
	.w1(32'hb659986e),
	.w2(32'h3b5220ad),
	.w3(32'hba33e958),
	.w4(32'h3c4029b2),
	.w5(32'h3c8e69d5),
	.w6(32'hbd237f78),
	.w7(32'hbbaecc67),
	.w8(32'h3c447704),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e6904),
	.w1(32'h3ae116b6),
	.w2(32'h3bef8526),
	.w3(32'h3a7a88cf),
	.w4(32'hbb306607),
	.w5(32'h3c844aa9),
	.w6(32'hbc471f8d),
	.w7(32'hbb4af39e),
	.w8(32'h3c1f27d5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27cd5a),
	.w1(32'h3a4d33cf),
	.w2(32'h3bb5d322),
	.w3(32'h3c1fae99),
	.w4(32'h3bf5c718),
	.w5(32'h3c10460b),
	.w6(32'hbbb96554),
	.w7(32'h396d4d8f),
	.w8(32'hbc3a6c6d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb57049),
	.w1(32'hbbef0760),
	.w2(32'h3c12b3cf),
	.w3(32'h3b4b719e),
	.w4(32'h3c96e8eb),
	.w5(32'h3ba84934),
	.w6(32'hbced8ff6),
	.w7(32'h38257cf6),
	.w8(32'hbc2e7178),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c6d09),
	.w1(32'hbadbd91a),
	.w2(32'h3c1612df),
	.w3(32'h3a51d5ea),
	.w4(32'h3c5187bf),
	.w5(32'hbbf92e13),
	.w6(32'hbd05ed9c),
	.w7(32'hbb52e4be),
	.w8(32'h3c2a4e8e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbccee0),
	.w1(32'hb9d8908d),
	.w2(32'hbaee0c33),
	.w3(32'hbbbb39e3),
	.w4(32'hbb486660),
	.w5(32'h3aefbdbd),
	.w6(32'hbc60e83a),
	.w7(32'h3b9e9335),
	.w8(32'h3bb59baa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cd501),
	.w1(32'h3bfabdc0),
	.w2(32'h3c3d65cb),
	.w3(32'h3ae70b58),
	.w4(32'hbbd31e39),
	.w5(32'h3b8af8e1),
	.w6(32'h3c21e1ee),
	.w7(32'h3c51d99d),
	.w8(32'hba16e43b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2034f3),
	.w1(32'h3c1f8d96),
	.w2(32'h3bac61cb),
	.w3(32'h3bb233ac),
	.w4(32'h3b8bd2a0),
	.w5(32'h3b86378d),
	.w6(32'h3bfb9980),
	.w7(32'h3b31c508),
	.w8(32'hbbae8c35),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15b248),
	.w1(32'hbc133f50),
	.w2(32'h3b4b37b3),
	.w3(32'hbc325406),
	.w4(32'hbc19f395),
	.w5(32'h3b21f35b),
	.w6(32'hbcde7e6b),
	.w7(32'hbacaa06d),
	.w8(32'hb99dbc6e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adff014),
	.w1(32'h3b9badfa),
	.w2(32'h3aaaadea),
	.w3(32'h3b8b03e0),
	.w4(32'h3c11bee1),
	.w5(32'h3bf68c98),
	.w6(32'hbc038bf5),
	.w7(32'h3ba666a1),
	.w8(32'h3c327d37),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc799cf),
	.w1(32'h3c5a8f4e),
	.w2(32'h3c398d3e),
	.w3(32'hbb9fbcc5),
	.w4(32'h3c279039),
	.w5(32'h3a1a04cb),
	.w6(32'hbd002baa),
	.w7(32'h3c122224),
	.w8(32'hba19a718),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af77d0e),
	.w1(32'hbc11559c),
	.w2(32'hbadd03ce),
	.w3(32'hbbda6614),
	.w4(32'h3b32078b),
	.w5(32'h3b366cce),
	.w6(32'hbc56d844),
	.w7(32'hba46728f),
	.w8(32'h3ae074a6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3859963b),
	.w1(32'h3adb5afb),
	.w2(32'h3ba4eb12),
	.w3(32'hbba0223b),
	.w4(32'hbb5b8b9a),
	.w5(32'h3b983da2),
	.w6(32'hb74475dc),
	.w7(32'hba5751a2),
	.w8(32'h3a669f52),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd5174),
	.w1(32'hba42a70d),
	.w2(32'h3bb060fd),
	.w3(32'hbb6ea6e0),
	.w4(32'h3afe7acd),
	.w5(32'h3ab58ef0),
	.w6(32'h39f95c8d),
	.w7(32'h3b723ad9),
	.w8(32'h3bd250e1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2347ac),
	.w1(32'h3bd8b85a),
	.w2(32'h38d14738),
	.w3(32'hba29ec4e),
	.w4(32'h3ba23b37),
	.w5(32'h3c1b5955),
	.w6(32'h3b714df0),
	.w7(32'hbba69032),
	.w8(32'h3be93f38),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13c5d5),
	.w1(32'hbae1df48),
	.w2(32'hbb625a33),
	.w3(32'h3c274eb5),
	.w4(32'h3b36cef8),
	.w5(32'h3a91a272),
	.w6(32'h3c15fe37),
	.w7(32'h3b01f732),
	.w8(32'h39f247dc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c0190),
	.w1(32'hbbc20300),
	.w2(32'hbb7c1cfe),
	.w3(32'hbb4d3e6a),
	.w4(32'hbac0bb92),
	.w5(32'hbbde0fbc),
	.w6(32'hbc4e7a25),
	.w7(32'h3a1a5984),
	.w8(32'h3b45ec7d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d892c),
	.w1(32'h3bc28c1b),
	.w2(32'h3bf45a59),
	.w3(32'hbb930125),
	.w4(32'hbbad9852),
	.w5(32'hbba5e578),
	.w6(32'hba81c10b),
	.w7(32'hbc2e6526),
	.w8(32'h3ab17f82),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57774d),
	.w1(32'hbbdbc911),
	.w2(32'hbadad77b),
	.w3(32'hbb6d75d9),
	.w4(32'hbaccc4e8),
	.w5(32'h3c44efd2),
	.w6(32'hbafde25a),
	.w7(32'h3ba29f7c),
	.w8(32'hbb2eda61),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d290),
	.w1(32'hbc29252c),
	.w2(32'h3c060d0a),
	.w3(32'hbb95b23b),
	.w4(32'h3c0654ec),
	.w5(32'hbac1f1a0),
	.w6(32'hbd364782),
	.w7(32'hbb8cba05),
	.w8(32'hb9a40985),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b7c6),
	.w1(32'h3c17f114),
	.w2(32'h3bf9598b),
	.w3(32'h3c5a4c87),
	.w4(32'h3bdb19f8),
	.w5(32'h3c7ee43d),
	.w6(32'hbb43a761),
	.w7(32'h3c2bbb96),
	.w8(32'h3adfca5c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dfc66),
	.w1(32'h3ac21657),
	.w2(32'h3c0829c3),
	.w3(32'h3c3055dd),
	.w4(32'h3c2ec816),
	.w5(32'h3b4ae19d),
	.w6(32'h3b80b501),
	.w7(32'h3b69cbc5),
	.w8(32'h3b55767a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873e35),
	.w1(32'hbab422f7),
	.w2(32'h3abb9954),
	.w3(32'hba34b123),
	.w4(32'h3a22a8c5),
	.w5(32'h3b948f6c),
	.w6(32'h3b484d88),
	.w7(32'hba8094e8),
	.w8(32'hba143c6b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd80be),
	.w1(32'h3b79d492),
	.w2(32'h3ae3add1),
	.w3(32'h3bb847bd),
	.w4(32'h3b961e12),
	.w5(32'h3b9b12e6),
	.w6(32'h3c4cb94e),
	.w7(32'h3c05c204),
	.w8(32'h3b0f0e33),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fb43f),
	.w1(32'hbc80b96f),
	.w2(32'hbbd3794d),
	.w3(32'hbb300c44),
	.w4(32'h39e213f7),
	.w5(32'h3aecac73),
	.w6(32'hbbc80259),
	.w7(32'hb9ac0d43),
	.w8(32'h3bc3f361),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be63ea2),
	.w1(32'h3b74111f),
	.w2(32'h3bb3321b),
	.w3(32'hbc6cccd5),
	.w4(32'hbc111cac),
	.w5(32'h3b2ab3f5),
	.w6(32'hbaba38d5),
	.w7(32'h3bd4f1fb),
	.w8(32'hbb7e71c2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45cefe),
	.w1(32'h3ba450a0),
	.w2(32'hbb8aab05),
	.w3(32'hbbfc259d),
	.w4(32'hbb7d8e77),
	.w5(32'h3b56d748),
	.w6(32'hbc07ae37),
	.w7(32'hba30f846),
	.w8(32'h3c0e947b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c005fbb),
	.w1(32'hbc145445),
	.w2(32'hba83d906),
	.w3(32'hbc02903d),
	.w4(32'h3abf86cc),
	.w5(32'h3a1cf368),
	.w6(32'hbc8b57a3),
	.w7(32'h3b712a20),
	.w8(32'hbb42fee7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35f0f7),
	.w1(32'h3b27df69),
	.w2(32'h3af202b2),
	.w3(32'h39729c89),
	.w4(32'hba993992),
	.w5(32'h3b6ba493),
	.w6(32'hba50f888),
	.w7(32'h3b38719b),
	.w8(32'hbb63b26b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae15707),
	.w1(32'hbad57915),
	.w2(32'h3c62355a),
	.w3(32'h3a79d688),
	.w4(32'h3bfc54f5),
	.w5(32'hbac34ed5),
	.w6(32'hbc33d939),
	.w7(32'h3b2bcdb9),
	.w8(32'h3c0006c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3dc1b),
	.w1(32'hbbb6a188),
	.w2(32'h3b0f8f6f),
	.w3(32'hbc4d9304),
	.w4(32'h3a0c4608),
	.w5(32'h3b5973fa),
	.w6(32'h3a81d190),
	.w7(32'h3c4d8eab),
	.w8(32'hbc501fa4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3219f5),
	.w1(32'h3af77421),
	.w2(32'h3c31b123),
	.w3(32'h3bc7097e),
	.w4(32'h3c845e63),
	.w5(32'hbc0736da),
	.w6(32'hbcfaa823),
	.w7(32'h3bcf40ba),
	.w8(32'h3b5a68b4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e7a2),
	.w1(32'h3bb3c157),
	.w2(32'hb72ec91b),
	.w3(32'hbb770efd),
	.w4(32'hbbaf64d3),
	.w5(32'hbbf7a952),
	.w6(32'hbc63217d),
	.w7(32'hbb5ac756),
	.w8(32'hbc287247),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf754a9),
	.w1(32'hbb9b2066),
	.w2(32'hba8a06ac),
	.w3(32'hbbf32b79),
	.w4(32'h3c88b3eb),
	.w5(32'hb96c37bf),
	.w6(32'h3c44c4ce),
	.w7(32'hbb4cdadf),
	.w8(32'hb9f23a32),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea7a38),
	.w1(32'h3a87d4d6),
	.w2(32'hbb818e79),
	.w3(32'h3a75d30b),
	.w4(32'hbb90dcde),
	.w5(32'h3b515e56),
	.w6(32'h38a80154),
	.w7(32'hbc16691b),
	.w8(32'hbbfd86d7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc1b5a),
	.w1(32'hbbe76802),
	.w2(32'h3c026967),
	.w3(32'hbb2a447f),
	.w4(32'h3c1a0388),
	.w5(32'h3b828c6a),
	.w6(32'hbd359727),
	.w7(32'h3b201064),
	.w8(32'hbb512716),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b989f9d),
	.w1(32'h3c2f9f6e),
	.w2(32'h3b0dff61),
	.w3(32'h3b08b9c1),
	.w4(32'h3b34ca75),
	.w5(32'h3bed77f8),
	.w6(32'h3b726703),
	.w7(32'hbbc9ff25),
	.w8(32'h3be7b3f0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c981fe8),
	.w1(32'h3c2c58a5),
	.w2(32'h3bd0734f),
	.w3(32'h3c9edc06),
	.w4(32'h3c102487),
	.w5(32'h3c2ae6be),
	.w6(32'hbd03721b),
	.w7(32'h3af61393),
	.w8(32'h3aee7399),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5aeda),
	.w1(32'h3bfa771d),
	.w2(32'h3c0bd653),
	.w3(32'h3c1c4827),
	.w4(32'h3c108cc4),
	.w5(32'h3c157cf4),
	.w6(32'h3c4acf6c),
	.w7(32'h3bbfc0b4),
	.w8(32'h3b3e6ca8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bddbb88),
	.w1(32'h3ba9b650),
	.w2(32'h3bf1ffe2),
	.w3(32'h3c5ff8fe),
	.w4(32'h3c437636),
	.w5(32'hbba508bb),
	.w6(32'hbbadcb1f),
	.w7(32'hbb9137ad),
	.w8(32'hbbafe729),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e2b3),
	.w1(32'hbb16bffb),
	.w2(32'hbbb69e2a),
	.w3(32'h3addd485),
	.w4(32'h3aafdf45),
	.w5(32'h3b9c636e),
	.w6(32'h3b8c8166),
	.w7(32'hba50ba95),
	.w8(32'h3bbdaf0b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8c11f),
	.w1(32'h3bd4d7ee),
	.w2(32'hbb8aacfd),
	.w3(32'h3b540777),
	.w4(32'hbb6405d6),
	.w5(32'h3b9e4a71),
	.w6(32'hba621b3c),
	.w7(32'h3aca6540),
	.w8(32'hbbc4ae20),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f83aa),
	.w1(32'h3b963dec),
	.w2(32'h3c18e158),
	.w3(32'h3b3408d1),
	.w4(32'hbb38c57d),
	.w5(32'h3b648d7c),
	.w6(32'hbbbef3cb),
	.w7(32'h3b3836b9),
	.w8(32'hbc01069f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdf292),
	.w1(32'hbba9b262),
	.w2(32'hbafb0b52),
	.w3(32'h3b6df1e0),
	.w4(32'h3a722624),
	.w5(32'h3b07f92b),
	.w6(32'hbca1439d),
	.w7(32'h3b51e170),
	.w8(32'h3a0d8c89),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14fb78),
	.w1(32'hbbaca2ab),
	.w2(32'hbc470fc0),
	.w3(32'hbb9da6cb),
	.w4(32'hbbad6a16),
	.w5(32'hbc0e4b6a),
	.w6(32'h3ac0a1a8),
	.w7(32'hbc1ed6b2),
	.w8(32'hbac60a23),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf613d8),
	.w1(32'hbb51000c),
	.w2(32'h39511aae),
	.w3(32'h3b949a42),
	.w4(32'hb9f3b0dd),
	.w5(32'h3b3d8c88),
	.w6(32'hbbf6b9dc),
	.w7(32'h3b0637a3),
	.w8(32'hbc0c0578),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93cff0),
	.w1(32'h3ad09a3c),
	.w2(32'hba76054b),
	.w3(32'hbb0de78c),
	.w4(32'h3aa8fb2c),
	.w5(32'h3c30f1f0),
	.w6(32'hbc0ad7ab),
	.w7(32'hbc0ef7a6),
	.w8(32'h3c01cfcb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1171d3),
	.w1(32'h3ac9545b),
	.w2(32'hba703c0c),
	.w3(32'h3b9279f6),
	.w4(32'hbb956b59),
	.w5(32'h3bc7d8ac),
	.w6(32'hbc923527),
	.w7(32'hbb3bc212),
	.w8(32'h3ab6314f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb589ce3),
	.w1(32'hbb9107cc),
	.w2(32'h3ba67102),
	.w3(32'hbad1ec56),
	.w4(32'h3b748730),
	.w5(32'h3bc8d73d),
	.w6(32'hbaa5e7c7),
	.w7(32'h3b2354f7),
	.w8(32'hbaa577e1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e40ab),
	.w1(32'hbb7b0d04),
	.w2(32'hba48623c),
	.w3(32'h3bc3f3ae),
	.w4(32'h3b8ec274),
	.w5(32'h3b794d74),
	.w6(32'hbb799580),
	.w7(32'h3abe9fa3),
	.w8(32'h3bea0abe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929e33),
	.w1(32'h3b9fc47a),
	.w2(32'hbb0cc3c0),
	.w3(32'h3bf794e2),
	.w4(32'hbbc0dade),
	.w5(32'h3c21479c),
	.w6(32'h3c80aa05),
	.w7(32'hbb9a50fc),
	.w8(32'hbb5d0d03),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39452b8c),
	.w1(32'h3c14f560),
	.w2(32'h3c2911f0),
	.w3(32'h3bf52617),
	.w4(32'h3bdf8fd9),
	.w5(32'h3c14f20f),
	.w6(32'hb99d728e),
	.w7(32'hbaaa50d9),
	.w8(32'hb7046f55),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2c30c),
	.w1(32'hb995c6b2),
	.w2(32'h3b820c23),
	.w3(32'hba8acdb3),
	.w4(32'h3ac04fd1),
	.w5(32'hbb5fa3e7),
	.w6(32'hbcff3e53),
	.w7(32'hbba22786),
	.w8(32'hbb9adaa9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a462f0d),
	.w1(32'h3c88cc0c),
	.w2(32'hbc590d42),
	.w3(32'h3c4f94b1),
	.w4(32'hbc26e399),
	.w5(32'h3b051b95),
	.w6(32'h3cb63550),
	.w7(32'hbc1c3abc),
	.w8(32'hbb9d9987),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd744d0),
	.w1(32'hbb1c722a),
	.w2(32'h3bf07e92),
	.w3(32'hbbf12794),
	.w4(32'hbbaa45ad),
	.w5(32'h3bd2c2e2),
	.w6(32'hbc5758cf),
	.w7(32'hb92ca7b0),
	.w8(32'hba71197e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43404b),
	.w1(32'hbaef33fe),
	.w2(32'h3c3d69c2),
	.w3(32'h3b4ab178),
	.w4(32'h3c206b64),
	.w5(32'hbafd52f8),
	.w6(32'hbd0ef670),
	.w7(32'h3b735968),
	.w8(32'hbb21163a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b3dcd),
	.w1(32'hbb01cd40),
	.w2(32'hba7395a3),
	.w3(32'hbaca6343),
	.w4(32'hb9872e56),
	.w5(32'h3b7e8b63),
	.w6(32'hbb2bbec5),
	.w7(32'hba8d61a7),
	.w8(32'h3acacb31),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7828ce),
	.w1(32'hb95541c5),
	.w2(32'hb9891ecb),
	.w3(32'hbac2fb56),
	.w4(32'h3aa5e2ba),
	.w5(32'h399fb7ca),
	.w6(32'hb9e8806f),
	.w7(32'h3ad3e34d),
	.w8(32'h3b57870d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7186df),
	.w1(32'h3b04b153),
	.w2(32'hbaf0d838),
	.w3(32'h3b93ae10),
	.w4(32'h3b8ce7ed),
	.w5(32'h3b5c2de5),
	.w6(32'h3bca97a2),
	.w7(32'h39d73b14),
	.w8(32'h3b6a8ab8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7b19d),
	.w1(32'hbbb0893e),
	.w2(32'hbb1b3b38),
	.w3(32'hbb6db0db),
	.w4(32'h3b4d2d15),
	.w5(32'h3b6398e3),
	.w6(32'hbc0a86fd),
	.w7(32'h3baa619b),
	.w8(32'hbc11f6d2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bb9f9),
	.w1(32'hbc0ecdaa),
	.w2(32'h3c51bf64),
	.w3(32'h3a9a5cdc),
	.w4(32'h3bb59b66),
	.w5(32'h3bc76b05),
	.w6(32'hbcbd8c40),
	.w7(32'h3c7fc022),
	.w8(32'h3c3fd474),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52d69d),
	.w1(32'h3c899534),
	.w2(32'hbb6a8e8a),
	.w3(32'h3c45603b),
	.w4(32'hba0dac66),
	.w5(32'h3bc66df7),
	.w6(32'h3bd4b168),
	.w7(32'hbb2b2731),
	.w8(32'hbbd5a1c9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f643),
	.w1(32'h3b8b56db),
	.w2(32'h34c55700),
	.w3(32'h3b8b823e),
	.w4(32'h3b4344b7),
	.w5(32'h3b8cc30e),
	.w6(32'h3b63ff74),
	.w7(32'hbbfc32ea),
	.w8(32'hbb4feaa8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e141),
	.w1(32'hbba57c48),
	.w2(32'h3c1dfc1c),
	.w3(32'h3b2e43ee),
	.w4(32'hbacfeb29),
	.w5(32'h3b481322),
	.w6(32'hbcf3ea92),
	.w7(32'h3bab169f),
	.w8(32'h3c08453e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa5d0b),
	.w1(32'h3bd89773),
	.w2(32'h3b8dabfd),
	.w3(32'hb8f083db),
	.w4(32'h39f6195a),
	.w5(32'hba093ad8),
	.w6(32'h3b5a8fd7),
	.w7(32'h3b91e496),
	.w8(32'h3bea080c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9faa6a),
	.w1(32'hbaf2febd),
	.w2(32'h3a9b1c80),
	.w3(32'hbc03e856),
	.w4(32'hbac1bd83),
	.w5(32'hbbcde5b4),
	.w6(32'hbaecaa04),
	.w7(32'hbb67ae9b),
	.w8(32'hbc2b5a3f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba24f4e),
	.w1(32'hbab18121),
	.w2(32'h3b45d9e1),
	.w3(32'hbae71902),
	.w4(32'hbc020ec6),
	.w5(32'hbb5cd532),
	.w6(32'hbc9c08e7),
	.w7(32'hbc588349),
	.w8(32'h3acc3de2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf31faf),
	.w1(32'h3b17fea3),
	.w2(32'hbc0f8024),
	.w3(32'hbbd4b83b),
	.w4(32'hba346df6),
	.w5(32'hbaa7a3d9),
	.w6(32'hbc6c8380),
	.w7(32'h38f48682),
	.w8(32'hbc78ab07),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd328ae),
	.w1(32'h3c2074ee),
	.w2(32'h3c3361bb),
	.w3(32'h3a9febed),
	.w4(32'h3c108fd0),
	.w5(32'h3a4a466b),
	.w6(32'hbc883a04),
	.w7(32'h3bba20dd),
	.w8(32'h3b10b104),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a12d77),
	.w1(32'h3b9c5d58),
	.w2(32'h3a76c30e),
	.w3(32'h3a0b4ea2),
	.w4(32'hbbb8555d),
	.w5(32'hb9a21bbe),
	.w6(32'h3c151a33),
	.w7(32'hb99f5187),
	.w8(32'h3b553e62),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba166640),
	.w1(32'hb92c243c),
	.w2(32'hba36f38e),
	.w3(32'hbbbb4bef),
	.w4(32'hbb1529f5),
	.w5(32'hbb98d29c),
	.w6(32'hbbee6b03),
	.w7(32'hbb5fc1ce),
	.w8(32'hbb289902),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd58f6),
	.w1(32'hbc09d428),
	.w2(32'hbc0ce4ce),
	.w3(32'hbbd704da),
	.w4(32'hbb6fadb8),
	.w5(32'h39daf2c4),
	.w6(32'h3a4609c1),
	.w7(32'hbbc82523),
	.w8(32'hbb72f50b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b308a),
	.w1(32'hbb99ac72),
	.w2(32'h3af7b409),
	.w3(32'hbbebedea),
	.w4(32'hbb7bbf75),
	.w5(32'h3c05ac63),
	.w6(32'h3b0a6e93),
	.w7(32'h3a9e024f),
	.w8(32'h3c125f73),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cabe5),
	.w1(32'hbbafce9e),
	.w2(32'h3bbb44d3),
	.w3(32'h3aa581c3),
	.w4(32'h3c158891),
	.w5(32'h38361e56),
	.w6(32'hbcd3eb0a),
	.w7(32'h3c5218e0),
	.w8(32'h3c4368cf),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54f5b3),
	.w1(32'h3c178a35),
	.w2(32'hbb3b6e56),
	.w3(32'h3bdf94b6),
	.w4(32'hbc7c2f7c),
	.w5(32'h3b57bca5),
	.w6(32'h3d010bc9),
	.w7(32'hbb6e45e6),
	.w8(32'hbb9408bf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17d723),
	.w1(32'h3a8291a6),
	.w2(32'h3baf01fe),
	.w3(32'hba1ee4e9),
	.w4(32'hba87dd10),
	.w5(32'h3b11573d),
	.w6(32'hbb7b5a17),
	.w7(32'h3a66eaf6),
	.w8(32'h3b0e25d6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59b2aa),
	.w1(32'h39bec597),
	.w2(32'h3b02fd26),
	.w3(32'hba42234b),
	.w4(32'hba89c7cd),
	.w5(32'h3acddb41),
	.w6(32'h3ae59122),
	.w7(32'hbb714c9f),
	.w8(32'hbb54ecae),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be16545),
	.w1(32'hba2fceb7),
	.w2(32'hba5b967a),
	.w3(32'hbb560751),
	.w4(32'h3b847c1e),
	.w5(32'hbab90694),
	.w6(32'hbc0b0098),
	.w7(32'hbb17bfa8),
	.w8(32'h392dd752),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64bb3b),
	.w1(32'hbbee1a48),
	.w2(32'hbb10614f),
	.w3(32'hba158d0c),
	.w4(32'h3a81207b),
	.w5(32'h3bfee720),
	.w6(32'hbbbf0786),
	.w7(32'hba683253),
	.w8(32'h3a20db18),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f3039),
	.w1(32'hbab65dfb),
	.w2(32'h3bd694cf),
	.w3(32'hbb0964ea),
	.w4(32'h3be0a3e1),
	.w5(32'h3b837445),
	.w6(32'hbcc764ca),
	.w7(32'hbc6fbeaf),
	.w8(32'hbb9db5dd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ce8d),
	.w1(32'h3b8d7684),
	.w2(32'h3b3f331f),
	.w3(32'h3c1aafb1),
	.w4(32'h3b82aa83),
	.w5(32'hba373b55),
	.w6(32'hbca4c00f),
	.w7(32'hba77abd3),
	.w8(32'h3b0b7241),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8705dc),
	.w1(32'hb77ca162),
	.w2(32'h3ba51ce4),
	.w3(32'hbc0a6afd),
	.w4(32'hbb38b5ed),
	.w5(32'h3bcf54a5),
	.w6(32'hbaf00b3a),
	.w7(32'h3c0766c7),
	.w8(32'h3be2e8fd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ba511),
	.w1(32'h3b9d6ac0),
	.w2(32'h3c285da5),
	.w3(32'hbafb9d28),
	.w4(32'h3c392504),
	.w5(32'h3acd5581),
	.w6(32'hbcdb3ee7),
	.w7(32'h3c2ad864),
	.w8(32'hbbcba237),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d05701),
	.w1(32'hbb1d0e98),
	.w2(32'hba9b5550),
	.w3(32'h3b769878),
	.w4(32'h3c138189),
	.w5(32'hbb952db2),
	.w6(32'hbbd69e0d),
	.w7(32'h3b469e36),
	.w8(32'h3c00886b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad34314),
	.w1(32'hbc030eec),
	.w2(32'hbbd0eb89),
	.w3(32'hbbc59fd8),
	.w4(32'h3b8037b5),
	.w5(32'h3b8935ff),
	.w6(32'h3a23c10c),
	.w7(32'hbb03c928),
	.w8(32'h3b57f46f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9932),
	.w1(32'hbb3f12bd),
	.w2(32'hbb02fff8),
	.w3(32'h3ad805b9),
	.w4(32'h3b862e02),
	.w5(32'h3bdbd5d0),
	.w6(32'h3996dcdd),
	.w7(32'h3b18c1f7),
	.w8(32'h3b65f0f5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17f86c),
	.w1(32'h3c24b9e3),
	.w2(32'h3ab2a3f4),
	.w3(32'h3c20f57f),
	.w4(32'hbabe0f4d),
	.w5(32'h3a2d59a4),
	.w6(32'hbc56085a),
	.w7(32'h3abb0b9a),
	.w8(32'h3b199f67),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb090ab7),
	.w1(32'hbb2eee4b),
	.w2(32'hbc40aca0),
	.w3(32'hbb8eea62),
	.w4(32'hbbe4f75a),
	.w5(32'h3c177452),
	.w6(32'hbbc9edba),
	.w7(32'hbbfeed80),
	.w8(32'hbb357a6e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0390d2),
	.w1(32'hbc5c8f1b),
	.w2(32'h3b7b814e),
	.w3(32'hbad10abd),
	.w4(32'h3c52460d),
	.w5(32'h3b1f5e49),
	.w6(32'hbc9f8f62),
	.w7(32'h3bab9798),
	.w8(32'h3b7d0ca0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf638e3),
	.w1(32'h3b880175),
	.w2(32'h3ba88917),
	.w3(32'hbb928ea9),
	.w4(32'h3b2e39d0),
	.w5(32'hbc704c45),
	.w6(32'hba9ee08d),
	.w7(32'h3b157c4f),
	.w8(32'hbc157fbb),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbca879),
	.w1(32'hbb1b01c4),
	.w2(32'hbc9f9f84),
	.w3(32'hb9d9508c),
	.w4(32'hbb0f8d96),
	.w5(32'hbb687ff9),
	.w6(32'h3c96daf6),
	.w7(32'hbc68f27f),
	.w8(32'h3a6654dd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04c861),
	.w1(32'h3a44caa1),
	.w2(32'hbc61dec8),
	.w3(32'hbb1a3300),
	.w4(32'hbb1f2547),
	.w5(32'h3b41e085),
	.w6(32'hbc4d6d58),
	.w7(32'hbcb36145),
	.w8(32'hbaff861e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6d952),
	.w1(32'hb89ec222),
	.w2(32'hbb00b253),
	.w3(32'hb9e27de0),
	.w4(32'hba6078b0),
	.w5(32'h3b388cf7),
	.w6(32'hbbe2a526),
	.w7(32'hbb9f00e2),
	.w8(32'hbc0c0486),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72849e),
	.w1(32'hbc948ce9),
	.w2(32'h3c085669),
	.w3(32'hbbd769ef),
	.w4(32'h3caf1841),
	.w5(32'h3bad52e1),
	.w6(32'hbcf80ba3),
	.w7(32'h3d030c87),
	.w8(32'hbb921cb3),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe450cb),
	.w1(32'hbbcb5ecc),
	.w2(32'hbb6c432b),
	.w3(32'h3ae09358),
	.w4(32'h3bba750e),
	.w5(32'hbb4fbc32),
	.w6(32'h3b5ed1d7),
	.w7(32'h3c20e7d4),
	.w8(32'hbb806fae),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2241fc),
	.w1(32'hbac2fadc),
	.w2(32'hbb680eab),
	.w3(32'hba8bbd64),
	.w4(32'hba0d9b70),
	.w5(32'h3b95dd05),
	.w6(32'h3b1424ab),
	.w7(32'hbb50a669),
	.w8(32'hba6045b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3922b3),
	.w1(32'h3b782533),
	.w2(32'hbb5d3d7f),
	.w3(32'hbb7ffeda),
	.w4(32'h3920ac8e),
	.w5(32'h3b41fbf2),
	.w6(32'hbb88a658),
	.w7(32'hbb02fa3c),
	.w8(32'h3cacbc37),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4df5),
	.w1(32'h3c1b7752),
	.w2(32'hbb1c8693),
	.w3(32'hbb9186de),
	.w4(32'hbc30dde0),
	.w5(32'hbbb1efba),
	.w6(32'h3c12449e),
	.w7(32'hbcb06bc1),
	.w8(32'hbc8a5849),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cbe0f),
	.w1(32'hbba4f8c1),
	.w2(32'h3b08f48c),
	.w3(32'hb9c56f81),
	.w4(32'h3c02c880),
	.w5(32'hbb8bb96b),
	.w6(32'hbc55c1d7),
	.w7(32'h3c9d263d),
	.w8(32'hbca427a9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62e343),
	.w1(32'hbca7d6ce),
	.w2(32'hba2416b3),
	.w3(32'h3afd0712),
	.w4(32'h3c559022),
	.w5(32'h398cad5c),
	.w6(32'hbc800fa1),
	.w7(32'h3d098574),
	.w8(32'hbc33371c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb004e0),
	.w1(32'hbc852fc9),
	.w2(32'h3c528da0),
	.w3(32'hbaebb18d),
	.w4(32'h3c6bac86),
	.w5(32'hba3899e3),
	.w6(32'hbcbdeef5),
	.w7(32'h3cb058c6),
	.w8(32'h3986cb78),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab706d8),
	.w1(32'hbb94be22),
	.w2(32'h3aa4f81b),
	.w3(32'hbbac5d8e),
	.w4(32'h3a584bb0),
	.w5(32'h3b8634bd),
	.w6(32'hbbcfec70),
	.w7(32'h3adc6842),
	.w8(32'h3af1ea11),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85e2f5d),
	.w1(32'hbb274c08),
	.w2(32'hbb0873fc),
	.w3(32'hbb873af8),
	.w4(32'hbb831c4d),
	.w5(32'h3b1c2940),
	.w6(32'hbc0313b9),
	.w7(32'hbc2c5121),
	.w8(32'h3b594c82),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b919b50),
	.w1(32'hbb67e240),
	.w2(32'hbbfd482d),
	.w3(32'h39e94d6e),
	.w4(32'hbc134e88),
	.w5(32'hbbb785d3),
	.w6(32'hbad1490b),
	.w7(32'hbc10ac59),
	.w8(32'hbc06194e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9fe33),
	.w1(32'hbacc615f),
	.w2(32'h3bb4d2ab),
	.w3(32'hbb93b203),
	.w4(32'h3b3c86e9),
	.w5(32'h3a4eba80),
	.w6(32'hbb83d9e2),
	.w7(32'h3c0a465a),
	.w8(32'hbbadd0fb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857fee),
	.w1(32'hbb5521f7),
	.w2(32'hbba17987),
	.w3(32'h3bdd2191),
	.w4(32'h3ba18400),
	.w5(32'h3baeb9bc),
	.w6(32'h3980ab22),
	.w7(32'hbbe1451a),
	.w8(32'h3bb47cb4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6de669),
	.w1(32'h3b591cdb),
	.w2(32'hbbc60714),
	.w3(32'hbb6b34a3),
	.w4(32'hbbfeca4e),
	.w5(32'hbac4dc45),
	.w6(32'hb788e0c7),
	.w7(32'hbbd24af9),
	.w8(32'hbbab9533),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc10020),
	.w1(32'hbb28f1f7),
	.w2(32'h3bd97857),
	.w3(32'h3b237d18),
	.w4(32'h3bf602e4),
	.w5(32'h397ff30e),
	.w6(32'h3b52c3c6),
	.w7(32'h3c337c32),
	.w8(32'hbc0ba02a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1baef6),
	.w1(32'hbccd2aa2),
	.w2(32'h3c3148d6),
	.w3(32'h3c78e3dc),
	.w4(32'h39ac8a18),
	.w5(32'h3a46152c),
	.w6(32'h3b4c2d60),
	.w7(32'h3cd1d94c),
	.w8(32'hbbc68b1c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2491),
	.w1(32'hbb7b93be),
	.w2(32'hbb32d362),
	.w3(32'hb88495c1),
	.w4(32'h3c5f3a1b),
	.w5(32'h3b953fc8),
	.w6(32'hbc0ac82e),
	.w7(32'hbadd637e),
	.w8(32'h3abf8dd0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8c813),
	.w1(32'h3a3840b0),
	.w2(32'hbb414e33),
	.w3(32'h3bb0a247),
	.w4(32'hbba835ae),
	.w5(32'hbc484bce),
	.w6(32'h3b8a98b4),
	.w7(32'hbb95797e),
	.w8(32'hbb5973b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8053a),
	.w1(32'hbc071fc0),
	.w2(32'hbb5aaabe),
	.w3(32'hbbeac3f9),
	.w4(32'h3c15e57d),
	.w5(32'h3c1f19a8),
	.w6(32'hbc2f54bf),
	.w7(32'h3cad2f6f),
	.w8(32'h3b02eccd),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcff60b),
	.w1(32'h3acd2021),
	.w2(32'hbaa474cc),
	.w3(32'hbab4245b),
	.w4(32'h3a818701),
	.w5(32'h3a417f6b),
	.w6(32'hbc2ee2ca),
	.w7(32'hbaea2a73),
	.w8(32'hbaf0f371),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670210),
	.w1(32'hbb47e7c4),
	.w2(32'hb9104768),
	.w3(32'hbad425d8),
	.w4(32'hb99e5301),
	.w5(32'h3a4f7461),
	.w6(32'hbbdbf3a6),
	.w7(32'hbc10d9e8),
	.w8(32'hbb1ba1c6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c1cbf),
	.w1(32'hbae1caf4),
	.w2(32'hbb4d897d),
	.w3(32'h3b83a355),
	.w4(32'h3c364602),
	.w5(32'h3b6e4279),
	.w6(32'hbb5c68f7),
	.w7(32'h3b83743b),
	.w8(32'h3984020e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b659e4d),
	.w1(32'h3aad0a92),
	.w2(32'hb91be072),
	.w3(32'hbb6d72e3),
	.w4(32'hbb086734),
	.w5(32'h3ba26da7),
	.w6(32'h3a022a12),
	.w7(32'hbb0794be),
	.w8(32'h3a54f61a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5b7f8),
	.w1(32'h3a0b7a6f),
	.w2(32'h3b5c978e),
	.w3(32'h3bf87b73),
	.w4(32'h3b983fb4),
	.w5(32'hbaaefe07),
	.w6(32'h3b267ee7),
	.w7(32'h3a00d251),
	.w8(32'h3b5d1c56),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b9709),
	.w1(32'h3a4282ed),
	.w2(32'h3aa2f01f),
	.w3(32'hbb60e1fc),
	.w4(32'hbb387b56),
	.w5(32'h3b849ea9),
	.w6(32'h3b31b422),
	.w7(32'h3b558e87),
	.w8(32'h3a41c14d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b290cf3),
	.w1(32'hbb8c39d8),
	.w2(32'hbb6411dc),
	.w3(32'hba2e8691),
	.w4(32'hbbda2b63),
	.w5(32'hbbb394f1),
	.w6(32'h3be0e84d),
	.w7(32'h3b1b0912),
	.w8(32'hbbe40b0e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb039c),
	.w1(32'hbbfa8cd6),
	.w2(32'hbb057cb1),
	.w3(32'hbb1eafa7),
	.w4(32'hbab55cb2),
	.w5(32'h39513298),
	.w6(32'h3c3bc707),
	.w7(32'h3b0ba910),
	.w8(32'h3b451f30),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa99efa),
	.w1(32'hbb1cf568),
	.w2(32'h3a12817b),
	.w3(32'h3b11469b),
	.w4(32'hbaec54d9),
	.w5(32'hbb251262),
	.w6(32'h39fd7f4c),
	.w7(32'h3bc1a9c5),
	.w8(32'hbc76f3b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa00da),
	.w1(32'hbc4fc743),
	.w2(32'h3acbb620),
	.w3(32'h3c20411c),
	.w4(32'hbb6752fa),
	.w5(32'hbb0ad4b4),
	.w6(32'h3ca6dd9f),
	.w7(32'hbac589b0),
	.w8(32'hbab1f478),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6faba5),
	.w1(32'hbb91b366),
	.w2(32'hbc1a66ab),
	.w3(32'hbbb3f34c),
	.w4(32'hbbd11e7a),
	.w5(32'hb8e4cb05),
	.w6(32'hbb9950e0),
	.w7(32'hbc4a5879),
	.w8(32'hb77246bf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3785f2ac),
	.w1(32'hbbd28d01),
	.w2(32'hb827bf88),
	.w3(32'hb98c30ae),
	.w4(32'h3a6c8682),
	.w5(32'h3b4cdd6a),
	.w6(32'hbb08823b),
	.w7(32'h3c49151f),
	.w8(32'h39d04b7e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf604f5),
	.w1(32'hbc24e4d9),
	.w2(32'h3ba099c3),
	.w3(32'h3b0ad09e),
	.w4(32'h3b36dc86),
	.w5(32'hbb2459ad),
	.w6(32'h3bf354f4),
	.w7(32'h3c701f02),
	.w8(32'h3bc29085),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc78527),
	.w1(32'h3b94eab0),
	.w2(32'hb9aca23c),
	.w3(32'h3a898b4a),
	.w4(32'hbb661976),
	.w5(32'hbb870560),
	.w6(32'h3bb8452e),
	.w7(32'hbb8b3574),
	.w8(32'h3af43216),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b667ca8),
	.w1(32'hbb84aff2),
	.w2(32'hbb8b3af5),
	.w3(32'hbbf1983b),
	.w4(32'hbbed985b),
	.w5(32'h3b971d11),
	.w6(32'hbbc9166a),
	.w7(32'h3bd9bc82),
	.w8(32'h3b694b68),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43018),
	.w1(32'h3a503670),
	.w2(32'h39c370b3),
	.w3(32'h3b32ac74),
	.w4(32'hbb420d3c),
	.w5(32'h3bd2ed19),
	.w6(32'h3af28a55),
	.w7(32'h3a9a2ecc),
	.w8(32'h3b89169b),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb27ae),
	.w1(32'hba7ec16f),
	.w2(32'h39c6030c),
	.w3(32'h3ba44876),
	.w4(32'h3ab6ac26),
	.w5(32'h3b675509),
	.w6(32'hba291e55),
	.w7(32'h3bde3bf6),
	.w8(32'h3b48e89c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6cb85),
	.w1(32'h3b781783),
	.w2(32'hbc1da854),
	.w3(32'h3ba36927),
	.w4(32'h3b44c8d0),
	.w5(32'h3bc0f018),
	.w6(32'hbb11e770),
	.w7(32'hbb766f83),
	.w8(32'h3c0bbcff),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ff434),
	.w1(32'h3b910999),
	.w2(32'h39b421c5),
	.w3(32'h3b058bf0),
	.w4(32'hbb85e952),
	.w5(32'h3b0794b2),
	.w6(32'h3b865951),
	.w7(32'hbada27bf),
	.w8(32'h3b935560),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bbdcb),
	.w1(32'h39973f0a),
	.w2(32'hb8ea498b),
	.w3(32'hbacc27e5),
	.w4(32'hbb977c90),
	.w5(32'h3a22c9f9),
	.w6(32'hbb427164),
	.w7(32'hbb36c7f5),
	.w8(32'h3ac3e6dc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b0d5),
	.w1(32'h3acf1832),
	.w2(32'h3a8c08a3),
	.w3(32'hbacc4d62),
	.w4(32'hbb280e53),
	.w5(32'hbb58829e),
	.w6(32'h3accd0b9),
	.w7(32'h3ab3aeaf),
	.w8(32'hbc6088fd),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14b3fd),
	.w1(32'hbc2d8e00),
	.w2(32'h3c0cc12d),
	.w3(32'h3a9f3acf),
	.w4(32'h3c266784),
	.w5(32'hbb6ab4c4),
	.w6(32'hbc26ab29),
	.w7(32'h3cb645cc),
	.w8(32'hbbba2fd4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc112b67),
	.w1(32'hbb29654b),
	.w2(32'h3b806a19),
	.w3(32'hbb80d279),
	.w4(32'h3b79b774),
	.w5(32'hbb83804c),
	.w6(32'hbb495d36),
	.w7(32'h3c136d44),
	.w8(32'hbb66b820),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb393e1e),
	.w1(32'hbbb4fbc1),
	.w2(32'h3b33ff30),
	.w3(32'hbb78e672),
	.w4(32'hbaa23c51),
	.w5(32'hbb80eff3),
	.w6(32'h3c8896be),
	.w7(32'hb941603e),
	.w8(32'hbba30ca2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac33100),
	.w1(32'h3bce1a13),
	.w2(32'h3bb74a95),
	.w3(32'hbb55a1e1),
	.w4(32'h39cf4952),
	.w5(32'h3ae06b35),
	.w6(32'h3b0759ef),
	.w7(32'h3bb4d00e),
	.w8(32'hb9fd4d23),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0407b),
	.w1(32'h38b3b4e8),
	.w2(32'hba663158),
	.w3(32'hbbfc2bab),
	.w4(32'hbb1cefa5),
	.w5(32'hbacded6b),
	.w6(32'hbb67cd79),
	.w7(32'hba6276ec),
	.w8(32'hbbb02db1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c78fe),
	.w1(32'hbb0b038a),
	.w2(32'h3bf442a4),
	.w3(32'hbb18a087),
	.w4(32'h3a4b493f),
	.w5(32'hbb4ce467),
	.w6(32'hbbc7eb9e),
	.w7(32'h3bfa2e90),
	.w8(32'hbc11d639),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954d88),
	.w1(32'hbbd4be32),
	.w2(32'h3acf3763),
	.w3(32'h3a691e75),
	.w4(32'h3bda2aa6),
	.w5(32'hbb536de1),
	.w6(32'h39bd0a46),
	.w7(32'h3c4de842),
	.w8(32'hbb537b71),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97fa5e),
	.w1(32'h3c84fbd7),
	.w2(32'h3bcd8e79),
	.w3(32'hbaca6527),
	.w4(32'h3b81ce7b),
	.w5(32'hbb12c790),
	.w6(32'hbbdba942),
	.w7(32'h3c13c4d7),
	.w8(32'hbbb9eb44),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6813c9),
	.w1(32'hbb50a5a1),
	.w2(32'hb974026e),
	.w3(32'h3b437f36),
	.w4(32'hbb75c98f),
	.w5(32'h3bee5bee),
	.w6(32'h3c1b5108),
	.w7(32'h3c16fd35),
	.w8(32'h3be3d6a9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18390),
	.w1(32'h3b4f62e6),
	.w2(32'h3b537537),
	.w3(32'hbb8462d2),
	.w4(32'h3bf44369),
	.w5(32'h3b8a46ae),
	.w6(32'hbba5abd4),
	.w7(32'h3bb25925),
	.w8(32'h3b63f3dd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a979993),
	.w1(32'h3aea7792),
	.w2(32'hbb881add),
	.w3(32'h3a8c0f8f),
	.w4(32'hbc316f40),
	.w5(32'h3b3aea8c),
	.w6(32'hba5e7f5c),
	.w7(32'hbc5b788b),
	.w8(32'h3b835037),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5410d),
	.w1(32'h39a2557b),
	.w2(32'h3a96c646),
	.w3(32'hbb68009e),
	.w4(32'hbb11e16b),
	.w5(32'hbbba7359),
	.w6(32'hbb13739b),
	.w7(32'h3956847f),
	.w8(32'h3b85963b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fdf53),
	.w1(32'h3bc28a8e),
	.w2(32'h3b75c91b),
	.w3(32'hbbfaaded),
	.w4(32'h3bdd4ff2),
	.w5(32'hba3a4598),
	.w6(32'hbb880942),
	.w7(32'h3c400ef2),
	.w8(32'hbb55ed23),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac30824),
	.w1(32'hbba47ce6),
	.w2(32'hbb03d96c),
	.w3(32'h3b8b214d),
	.w4(32'h3b0b62a8),
	.w5(32'h3b1b1048),
	.w6(32'h3bbeed7a),
	.w7(32'h3b84526f),
	.w8(32'hba814dfc),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab14132),
	.w1(32'hb9ecbaa1),
	.w2(32'hba3a5db5),
	.w3(32'hba480008),
	.w4(32'h392c32c5),
	.w5(32'hbb8d6a91),
	.w6(32'h3b096d8b),
	.w7(32'hba1ee183),
	.w8(32'hbc6665b8),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b64a9),
	.w1(32'hbc2a8c8e),
	.w2(32'hbba9bb28),
	.w3(32'hba0bee5e),
	.w4(32'h3c30e706),
	.w5(32'h3ad49789),
	.w6(32'hbc2b3d1a),
	.w7(32'h3ba09269),
	.w8(32'h3b8f3ea6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f2745),
	.w1(32'hbb7aef8c),
	.w2(32'hbbf117d9),
	.w3(32'hbba571f6),
	.w4(32'hbc1ea958),
	.w5(32'hbbbc3c1a),
	.w6(32'hbb90752b),
	.w7(32'hbc0a8a43),
	.w8(32'hbbc845e1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ec1ef),
	.w1(32'hbc157271),
	.w2(32'h3bb5564a),
	.w3(32'hbb05827a),
	.w4(32'hbc109515),
	.w5(32'hbb6433b7),
	.w6(32'h3c53d5e2),
	.w7(32'h3bfcf9f0),
	.w8(32'hbb98a4ec),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc8ade),
	.w1(32'hb9826f4c),
	.w2(32'h3aa01945),
	.w3(32'h3b65e308),
	.w4(32'hba432774),
	.w5(32'hbc0a89ec),
	.w6(32'h3a1f434a),
	.w7(32'h3b7e6ef1),
	.w8(32'hbbd72b53),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66d285),
	.w1(32'hbbe0fd12),
	.w2(32'hbbd09dca),
	.w3(32'hbac42e10),
	.w4(32'h3cc0dcfd),
	.w5(32'hb9aa1123),
	.w6(32'hbc63c71a),
	.w7(32'h3cc8e19f),
	.w8(32'hbc81edb2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72f969),
	.w1(32'hbc3de1fc),
	.w2(32'h3c22f20d),
	.w3(32'h3abd3448),
	.w4(32'hbb76c2af),
	.w5(32'hbb0cfea0),
	.w6(32'h3c8b6f5b),
	.w7(32'h3ca37332),
	.w8(32'hbc1abf9a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ef9c9),
	.w1(32'hbb22b006),
	.w2(32'hbc259b9f),
	.w3(32'h3bdda124),
	.w4(32'h3ca13849),
	.w5(32'hbb3eee09),
	.w6(32'hbba2c0c8),
	.w7(32'hba633041),
	.w8(32'hbc5aa421),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6b99),
	.w1(32'hbcaa59fe),
	.w2(32'hbbdc7d69),
	.w3(32'hbc6252e0),
	.w4(32'h3b37a106),
	.w5(32'hb8885146),
	.w6(32'hbcb836e2),
	.w7(32'h3c78b3ac),
	.w8(32'h3ad59fcd),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa66a),
	.w1(32'hbbb36719),
	.w2(32'hbc0a915a),
	.w3(32'h3b89470d),
	.w4(32'hbae311cb),
	.w5(32'hbbeb56b7),
	.w6(32'h3bd52aaa),
	.w7(32'h38223e9f),
	.w8(32'hbc82ea81),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeeb85b),
	.w1(32'hbbe8bc8b),
	.w2(32'h3afec67e),
	.w3(32'hba87939a),
	.w4(32'h3c8baba7),
	.w5(32'hbbd3c7d2),
	.w6(32'hbb8dd0b7),
	.w7(32'h3d1a5495),
	.w8(32'hbc05e907),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca1697),
	.w1(32'hbb1211a7),
	.w2(32'hbb29e59c),
	.w3(32'hbb5efa41),
	.w4(32'h3cae1e3e),
	.w5(32'h3b4e8ab1),
	.w6(32'hbba9ae05),
	.w7(32'h3c7f3a9d),
	.w8(32'hbb2535e0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63767f),
	.w1(32'h3b79b780),
	.w2(32'hbbdf4f1a),
	.w3(32'h3b6d484a),
	.w4(32'h3a65ea65),
	.w5(32'hb8df4f96),
	.w6(32'h3b0d45ab),
	.w7(32'h3ba3fab9),
	.w8(32'h3ba0b8f6),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb940b5),
	.w1(32'h3bef2d0f),
	.w2(32'h3a094008),
	.w3(32'hbb5d7dcf),
	.w4(32'hbbf7b10e),
	.w5(32'h3b218862),
	.w6(32'h3b986c7c),
	.w7(32'hbb1fba41),
	.w8(32'h3c6c3554),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a33ec),
	.w1(32'h3c4f4480),
	.w2(32'h3b5158d0),
	.w3(32'hba9f94a5),
	.w4(32'hbc9b97d2),
	.w5(32'h3adb49d6),
	.w6(32'h3bb7a8fb),
	.w7(32'hbd01fcd5),
	.w8(32'hbba0d8a8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb815aaa),
	.w1(32'hba9965fd),
	.w2(32'h3ba61528),
	.w3(32'h3ba4e770),
	.w4(32'h3c3d2fc3),
	.w5(32'hbaf3963d),
	.w6(32'hba41109a),
	.w7(32'h3bbd3b1c),
	.w8(32'hbbe27e06),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb626c30),
	.w1(32'hbb5a69df),
	.w2(32'hba5f4b9c),
	.w3(32'h3b0400ad),
	.w4(32'hbb1e3f45),
	.w5(32'hbb61bb2e),
	.w6(32'h39767add),
	.w7(32'h3b6a0a08),
	.w8(32'hbc1b2014),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba51a1a),
	.w1(32'h3a6112dd),
	.w2(32'h38a66fff),
	.w3(32'h3c09550c),
	.w4(32'h3c2c85ed),
	.w5(32'hbc14c537),
	.w6(32'h3b3ff49e),
	.w7(32'h3c892db4),
	.w8(32'hbcdb8a16),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b79f0),
	.w1(32'hbcbd8149),
	.w2(32'h3c1e4c41),
	.w3(32'hbc267bce),
	.w4(32'h3b691497),
	.w5(32'h3a8478b2),
	.w6(32'hbcf0d841),
	.w7(32'h3d28f4ad),
	.w8(32'hba3962e6),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b261df9),
	.w1(32'h3a25ec2a),
	.w2(32'hbafa0cee),
	.w3(32'h3ab3749e),
	.w4(32'hbb6077ac),
	.w5(32'hbbb3b70e),
	.w6(32'hbbea38c5),
	.w7(32'hbc2028f6),
	.w8(32'hb9112738),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb1b4),
	.w1(32'hbbf47bef),
	.w2(32'h3bd206b6),
	.w3(32'hbbd0916e),
	.w4(32'h3c7ca8a1),
	.w5(32'hbb698766),
	.w6(32'hbc01902e),
	.w7(32'h3c5ae68d),
	.w8(32'hbb3499d3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3a978),
	.w1(32'hbc15da4a),
	.w2(32'h3bfc636b),
	.w3(32'hbb8a96b0),
	.w4(32'h3c2542e7),
	.w5(32'h3be0b439),
	.w6(32'hbc4429bf),
	.w7(32'h3c15876d),
	.w8(32'h3c442ecd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee1014),
	.w1(32'h3c38a54f),
	.w2(32'hbc00db9e),
	.w3(32'h3a8edc26),
	.w4(32'hbc8138e0),
	.w5(32'hbb4cd5d3),
	.w6(32'h3c1517aa),
	.w7(32'hbcad1bbd),
	.w8(32'hbb168aba),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc42c7e),
	.w1(32'hbb125371),
	.w2(32'h39fa8a21),
	.w3(32'hbbbb7d7b),
	.w4(32'hb980d6ce),
	.w5(32'h3bb56cb7),
	.w6(32'h3a1f688f),
	.w7(32'h3bab4e1f),
	.w8(32'h3b5db2dd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba353e3),
	.w1(32'h3b984ba8),
	.w2(32'hbb5c6903),
	.w3(32'h3b978a92),
	.w4(32'hbc2f5ab8),
	.w5(32'hbb3b4865),
	.w6(32'h3c1c7585),
	.w7(32'hbc0bed8a),
	.w8(32'h39a56a04),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812fa0),
	.w1(32'hbc74700e),
	.w2(32'hba5370c6),
	.w3(32'hba7686af),
	.w4(32'h3c6f61f5),
	.w5(32'hbc19a533),
	.w6(32'hbca2bbf9),
	.w7(32'h3c8b9265),
	.w8(32'hbc6a725c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b054cb3),
	.w1(32'hbc1e2ec0),
	.w2(32'h39e2c07c),
	.w3(32'h3b8b8f3b),
	.w4(32'h3c1f7b20),
	.w5(32'hbb592acd),
	.w6(32'hbc1b7adb),
	.w7(32'h3d06880a),
	.w8(32'hbb0f964a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce8692),
	.w1(32'h3a9819fa),
	.w2(32'hbba392ec),
	.w3(32'hbc0a42e1),
	.w4(32'h39316ee9),
	.w5(32'hbc0f94c6),
	.w6(32'hbae4d1c5),
	.w7(32'hbbdc14a6),
	.w8(32'hbc3e6ab7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa6057),
	.w1(32'hba48d0f0),
	.w2(32'hba8ce194),
	.w3(32'hbb246117),
	.w4(32'h3bc70347),
	.w5(32'h3a9e7233),
	.w6(32'hbb46124b),
	.w7(32'h3c39d69a),
	.w8(32'hbb7183dd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec978),
	.w1(32'hbbc52b1a),
	.w2(32'h3bba48d3),
	.w3(32'h3bd0a76b),
	.w4(32'h3b104290),
	.w5(32'hbb671ec1),
	.w6(32'h3b5c5b4c),
	.w7(32'h3c993842),
	.w8(32'hbc21068d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad354b7),
	.w1(32'hbc6a7676),
	.w2(32'hbb1ce0f2),
	.w3(32'h3ad81387),
	.w4(32'hbbdfe084),
	.w5(32'h3a13a27d),
	.w6(32'hbaff0ef1),
	.w7(32'h3c206a19),
	.w8(32'hbb864057),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03cf91),
	.w1(32'hbb175803),
	.w2(32'hba6d8c45),
	.w3(32'h3b860705),
	.w4(32'h3b392b94),
	.w5(32'hbb8e3397),
	.w6(32'h3bb44bd3),
	.w7(32'h3be857de),
	.w8(32'hbc15f069),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d584b),
	.w1(32'hbb8e082b),
	.w2(32'hbb16b60d),
	.w3(32'hbb84c390),
	.w4(32'hbba98d39),
	.w5(32'h3b25e73b),
	.w6(32'hbb82fa7b),
	.w7(32'hbb27d578),
	.w8(32'hb9174b6e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993958d),
	.w1(32'h3a3261c6),
	.w2(32'hbbcd202c),
	.w3(32'h3b25cb84),
	.w4(32'hbbbfa83f),
	.w5(32'h3b817579),
	.w6(32'h3becedb5),
	.w7(32'hbb5c3f5f),
	.w8(32'h3ba7feb0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba382a8),
	.w1(32'h3b86b663),
	.w2(32'hbabf1c59),
	.w3(32'hbc1190d0),
	.w4(32'hbc743bc2),
	.w5(32'hbb4cf987),
	.w6(32'h3a3f0c6b),
	.w7(32'hbc901427),
	.w8(32'h3b33d479),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be47fcf),
	.w1(32'h3bcae6cc),
	.w2(32'hb8e4f18b),
	.w3(32'h3a64e698),
	.w4(32'hbbeeb8e4),
	.w5(32'hbbffb40a),
	.w6(32'h3b8b67bd),
	.w7(32'hbb272342),
	.w8(32'hbb2e36cd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a6025),
	.w1(32'h3b8e1ca9),
	.w2(32'h3b05843e),
	.w3(32'hbb925c53),
	.w4(32'h3aebe372),
	.w5(32'hbbbd2620),
	.w6(32'hbb293e1f),
	.w7(32'h3b7dc59c),
	.w8(32'h3bb0befe),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb6d22),
	.w1(32'h39bb91fa),
	.w2(32'hbbb34e2a),
	.w3(32'h39b20e6b),
	.w4(32'h3a8202d7),
	.w5(32'h3a87c997),
	.w6(32'h3c3be051),
	.w7(32'h3b645d52),
	.w8(32'hbb7f7228),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae97195),
	.w1(32'hbb8425b0),
	.w2(32'h389d9122),
	.w3(32'h3ba6e0f9),
	.w4(32'h3b664bf0),
	.w5(32'h3a10abe6),
	.w6(32'h3b409f8f),
	.w7(32'h3c008ac1),
	.w8(32'hbbacbf18),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2e0d2),
	.w1(32'hbbacb695),
	.w2(32'h3b51c175),
	.w3(32'h3b1698c3),
	.w4(32'hbc006a4e),
	.w5(32'hbad3dc18),
	.w6(32'h3bb3e537),
	.w7(32'h3c07df63),
	.w8(32'hba84b02c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58b4b0),
	.w1(32'hbb9702a6),
	.w2(32'h3b14b2fe),
	.w3(32'h3b86dc65),
	.w4(32'hbb6174c5),
	.w5(32'h3906cb99),
	.w6(32'h3bb930f3),
	.w7(32'h3c1d0965),
	.w8(32'hbb07ca42),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4b305),
	.w1(32'h3b660b4b),
	.w2(32'hbb7dccec),
	.w3(32'h3ada7d2e),
	.w4(32'hbbb1a8b0),
	.w5(32'hbb0a2591),
	.w6(32'h3b8eb65b),
	.w7(32'hbc14f53e),
	.w8(32'h3a9b4181),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbe5d9),
	.w1(32'hb9331fe8),
	.w2(32'hb8a94007),
	.w3(32'hbbaf4f99),
	.w4(32'hbb9a60e5),
	.w5(32'hbbdac8ee),
	.w6(32'hba85dee8),
	.w7(32'hbc25d54d),
	.w8(32'hbbfb3e7e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf52c52),
	.w1(32'hbc6a1810),
	.w2(32'hbb57523a),
	.w3(32'hbb14ce75),
	.w4(32'h3b9dc893),
	.w5(32'hbbe8776e),
	.w6(32'hbba6c494),
	.w7(32'h3bf6ffc2),
	.w8(32'hbcf368ab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc375923),
	.w1(32'hbcb57c3e),
	.w2(32'h3baccccb),
	.w3(32'h3b33da43),
	.w4(32'h3cab7f83),
	.w5(32'hbb042ea7),
	.w6(32'hbcdbd93e),
	.w7(32'h3d6aecfe),
	.w8(32'hbbe7f859),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ab49),
	.w1(32'h3b2a66b4),
	.w2(32'hbbad9a04),
	.w3(32'h3c0b66f4),
	.w4(32'h3c27daf2),
	.w5(32'h3b919ea6),
	.w6(32'hbaa2f957),
	.w7(32'h3b44b59e),
	.w8(32'h3bcf0727),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b719576),
	.w1(32'hbb41409f),
	.w2(32'h3a0c690f),
	.w3(32'hbb4c47a3),
	.w4(32'hbb99d9d1),
	.w5(32'h3a7230d9),
	.w6(32'hbbd3a1ca),
	.w7(32'hbb909681),
	.w8(32'h3bf47d26),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8f9f6),
	.w1(32'h3bc6d750),
	.w2(32'h3a30177e),
	.w3(32'hba64199c),
	.w4(32'hbbfa24a1),
	.w5(32'hbb7e7668),
	.w6(32'h3c0f54d7),
	.w7(32'h3b50c227),
	.w8(32'hbc15aa52),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb82a2f),
	.w1(32'hbc4e7c90),
	.w2(32'hbb830d27),
	.w3(32'hbc2e8967),
	.w4(32'h3c5466cd),
	.w5(32'h3ae1e84d),
	.w6(32'hbc9d36f7),
	.w7(32'h3c8eb43a),
	.w8(32'hb9e6a3bd),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacfa96),
	.w1(32'hbae3a974),
	.w2(32'hbbb46136),
	.w3(32'hbad5f2ab),
	.w4(32'hbbd4ed72),
	.w5(32'hba1196fc),
	.w6(32'h39c28442),
	.w7(32'hbba1251f),
	.w8(32'h3b2aa3e6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a078b),
	.w1(32'hbaedf065),
	.w2(32'h3bb9ccc5),
	.w3(32'h3aed20e4),
	.w4(32'h3c54914a),
	.w5(32'h3b872d01),
	.w6(32'h3bb87d2e),
	.w7(32'h3c8a4c0b),
	.w8(32'h3a8e2af9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94bea73),
	.w1(32'h3ab57db5),
	.w2(32'h396ee8ab),
	.w3(32'hbae91534),
	.w4(32'h3b8de738),
	.w5(32'hbb61501b),
	.w6(32'hbb404f68),
	.w7(32'hb9221fd7),
	.w8(32'hbc2993d6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab879e6),
	.w1(32'hbc86d6cd),
	.w2(32'hbbcb1728),
	.w3(32'hbb521a2e),
	.w4(32'h3baae2b3),
	.w5(32'h3af758be),
	.w6(32'hbc5d9a73),
	.w7(32'h3cb4710d),
	.w8(32'h3ca5cb8e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c540fe3),
	.w1(32'h3c3b0e2e),
	.w2(32'hbaedfcdc),
	.w3(32'hbc6dcd04),
	.w4(32'hbcd8cd43),
	.w5(32'h3b54b78f),
	.w6(32'hbb45a71d),
	.w7(32'hbcc4715e),
	.w8(32'h3b5d7a0e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d13c9),
	.w1(32'h3b59d84d),
	.w2(32'h3baa05c6),
	.w3(32'h3b603dac),
	.w4(32'h39954fbe),
	.w5(32'h3b5703d5),
	.w6(32'h3b19ac15),
	.w7(32'h3bb20697),
	.w8(32'h3c108ee2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bdc50),
	.w1(32'h3c71f68c),
	.w2(32'hbb82e2c7),
	.w3(32'hbb15ea79),
	.w4(32'hbc8b16d4),
	.w5(32'hbad15932),
	.w6(32'h3b819e54),
	.w7(32'hbc9da0af),
	.w8(32'hbc4287ae),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb697a9),
	.w1(32'hbb37a5bd),
	.w2(32'hbb5f668b),
	.w3(32'h3ac795f0),
	.w4(32'h3c36e2f6),
	.w5(32'hbab1e93e),
	.w6(32'hbc078aaf),
	.w7(32'h3c7ac05f),
	.w8(32'hba0a31c4),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074e96),
	.w1(32'hbb6df414),
	.w2(32'hb9ec8d7b),
	.w3(32'hbbfa0254),
	.w4(32'h3b884ee7),
	.w5(32'h3b6531d7),
	.w6(32'h39d0107f),
	.w7(32'h3ac56072),
	.w8(32'h3c3c82e6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd68a6),
	.w1(32'h3bcda8ea),
	.w2(32'h37a522c2),
	.w3(32'hbc09e01a),
	.w4(32'hbc463b46),
	.w5(32'hbb5602ce),
	.w6(32'h3c09872c),
	.w7(32'hbc877d2d),
	.w8(32'hbb1c04be),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e147),
	.w1(32'hbbf71e94),
	.w2(32'hb9c0ed6f),
	.w3(32'hbb58b6b0),
	.w4(32'h3aac583e),
	.w5(32'h3aab9928),
	.w6(32'hbabe790d),
	.w7(32'h3b105766),
	.w8(32'h3ba57084),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf7224),
	.w1(32'h3b9aa5b9),
	.w2(32'h3b43b4b6),
	.w3(32'hbb258f44),
	.w4(32'hbaf04ce2),
	.w5(32'hbbb399cb),
	.w6(32'h3b802532),
	.w7(32'h3a0b220b),
	.w8(32'hbc74611b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11bf6d),
	.w1(32'hbc10226a),
	.w2(32'hba80ec2f),
	.w3(32'hb88a8f41),
	.w4(32'h3bf428cf),
	.w5(32'hbb8d111f),
	.w6(32'hbba11d41),
	.w7(32'h3ca9c419),
	.w8(32'hbb2be23c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdf465),
	.w1(32'hbb86e567),
	.w2(32'hbbbcc71d),
	.w3(32'h3a566a1f),
	.w4(32'h3b1ee645),
	.w5(32'h3b940c68),
	.w6(32'h3b8f57ee),
	.w7(32'h3b97268a),
	.w8(32'h3a38ea4d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e4173),
	.w1(32'h3b0ade63),
	.w2(32'h3b984d17),
	.w3(32'h3a280d55),
	.w4(32'h3b474b7b),
	.w5(32'hb8b5facf),
	.w6(32'hba7e1dc8),
	.w7(32'h3c0444fc),
	.w8(32'h3bc32064),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84be85),
	.w1(32'h3bbf8150),
	.w2(32'h3c2b2e56),
	.w3(32'h3b6856d6),
	.w4(32'hba888455),
	.w5(32'h3bdcb766),
	.w6(32'h3bb42537),
	.w7(32'h3aa24b04),
	.w8(32'h3c24889c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12e85a),
	.w1(32'hbab5be80),
	.w2(32'h3aa1411c),
	.w3(32'hba5d2e87),
	.w4(32'hbb0b3376),
	.w5(32'hbaf85b59),
	.w6(32'h3ba7554a),
	.w7(32'hbb8d2402),
	.w8(32'hbba216cb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb910f14),
	.w1(32'hbb18dba7),
	.w2(32'hbb7f50a1),
	.w3(32'h3b810e2b),
	.w4(32'hbc2d1025),
	.w5(32'hbc57fee1),
	.w6(32'hbbe043c4),
	.w7(32'hbc52447c),
	.w8(32'hbcccfc0a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12500d),
	.w1(32'hbd05a285),
	.w2(32'h3a8186dc),
	.w3(32'hbb6cfb08),
	.w4(32'h3be73012),
	.w5(32'h3b962dc5),
	.w6(32'hbc902f76),
	.w7(32'h3c49c160),
	.w8(32'h3b3320e0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd63ece),
	.w1(32'h3b71ade1),
	.w2(32'h3b95e3de),
	.w3(32'h3bb47271),
	.w4(32'hbb9b7085),
	.w5(32'h3bc8dd74),
	.w6(32'hbb2c93a7),
	.w7(32'hbbb3bf8d),
	.w8(32'h3c3934ec),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55820),
	.w1(32'h3aa08a6f),
	.w2(32'hbc202d4d),
	.w3(32'h3b6069fe),
	.w4(32'hbb0a1b61),
	.w5(32'hbb3fc672),
	.w6(32'h3ad2cbe0),
	.w7(32'hbc2ab686),
	.w8(32'hbc74426c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf56781),
	.w1(32'hbc174f5c),
	.w2(32'h3ac9e6d2),
	.w3(32'h3b3f3083),
	.w4(32'h3b9d998f),
	.w5(32'h3c0ca513),
	.w6(32'hbbfff5a5),
	.w7(32'h3cf229c2),
	.w8(32'h3ce901c3),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9907b7),
	.w1(32'h3ca527e4),
	.w2(32'hbb44470c),
	.w3(32'hbc71b3b3),
	.w4(32'hbd075814),
	.w5(32'h3a32ab22),
	.w6(32'h3c3eb4c6),
	.w7(32'hbd303673),
	.w8(32'hbb959327),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c0b5a),
	.w1(32'hbc103a64),
	.w2(32'h3a61bc26),
	.w3(32'h3a9e8f37),
	.w4(32'h3c45262a),
	.w5(32'h37722605),
	.w6(32'hbbfc3380),
	.w7(32'h3c0d3ade),
	.w8(32'hb8959d06),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb869f469),
	.w1(32'hba23dfd8),
	.w2(32'hbacb0193),
	.w3(32'hb9bc32c6),
	.w4(32'hba231985),
	.w5(32'hba2be390),
	.w6(32'hba783ab1),
	.w7(32'hba9226ba),
	.w8(32'hba628189),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0d487),
	.w1(32'hba2543ca),
	.w2(32'hba5b88cf),
	.w3(32'hbadd640f),
	.w4(32'hba50e67f),
	.w5(32'hb91a92fc),
	.w6(32'hb9326a3a),
	.w7(32'hb99ae44f),
	.w8(32'hba082529),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba004812),
	.w1(32'hb9c75264),
	.w2(32'hb973cf16),
	.w3(32'h3a2832bd),
	.w4(32'h3946c40f),
	.w5(32'h3b8a1de6),
	.w6(32'h3a8eae1c),
	.w7(32'h39d5b47b),
	.w8(32'h3b5cd876),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cce4e),
	.w1(32'h3b4d4e21),
	.w2(32'h3b3409f0),
	.w3(32'h3baf38df),
	.w4(32'h3ba65e71),
	.w5(32'h3a2cc6e3),
	.w6(32'h3ba8dd6a),
	.w7(32'h3b8c3d5a),
	.w8(32'hb98714b0),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ef9da),
	.w1(32'hbacb0c1c),
	.w2(32'hb9b7b77d),
	.w3(32'hbb5a33e6),
	.w4(32'hb986d306),
	.w5(32'hbaeeae3f),
	.w6(32'hbbaba836),
	.w7(32'hbaee0772),
	.w8(32'hbaaf0eee),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34751e),
	.w1(32'hb99fa4f7),
	.w2(32'hb8c86b8f),
	.w3(32'hbad081d8),
	.w4(32'hba82cfb0),
	.w5(32'hba623ee3),
	.w6(32'hbae4d7d1),
	.w7(32'hba3caffc),
	.w8(32'hbaa74191),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad7184),
	.w1(32'hbafea854),
	.w2(32'hbb09e748),
	.w3(32'hbacd256a),
	.w4(32'hbb267001),
	.w5(32'hba8e8364),
	.w6(32'hbada58bf),
	.w7(32'hbb29270c),
	.w8(32'hba748f50),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6c588),
	.w1(32'hba117466),
	.w2(32'hbb2ac57d),
	.w3(32'hbaf83137),
	.w4(32'hbb2c27a4),
	.w5(32'hba3292b9),
	.w6(32'hbabf0842),
	.w7(32'hbb0d9120),
	.w8(32'hb9606b18),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07dc48),
	.w1(32'h3a19b2fa),
	.w2(32'h3a303c3f),
	.w3(32'hb89319fc),
	.w4(32'hb9b2b9f1),
	.w5(32'hb8cafb76),
	.w6(32'h39ad8c1a),
	.w7(32'hb898a972),
	.w8(32'hb9e39c8b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b680b),
	.w1(32'hba083ba2),
	.w2(32'h38ab36d4),
	.w3(32'h39cdcb19),
	.w4(32'h3a40ef11),
	.w5(32'hb9714970),
	.w6(32'h39890208),
	.w7(32'h39be9472),
	.w8(32'hb938c451),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba268b88),
	.w1(32'hb91b8352),
	.w2(32'hba474d17),
	.w3(32'h38a1113d),
	.w4(32'hb951cf22),
	.w5(32'h39adbe58),
	.w6(32'hb8e8e2a3),
	.w7(32'hb9d6c6fc),
	.w8(32'hb8a11fbb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae238a),
	.w1(32'h38da6f9b),
	.w2(32'h37bc6773),
	.w3(32'h39d8ae19),
	.w4(32'h39e59cc8),
	.w5(32'hba8ef761),
	.w6(32'hb98827dc),
	.w7(32'hb906c041),
	.w8(32'hba84fafc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b38cac),
	.w1(32'hba9361d6),
	.w2(32'hbaeb41d4),
	.w3(32'hba94987e),
	.w4(32'hbaaec570),
	.w5(32'h39b613cf),
	.w6(32'hbabe8e5a),
	.w7(32'hbaff89b5),
	.w8(32'h39db7a1f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c1f3e),
	.w1(32'hbacc5d9a),
	.w2(32'hb8840dc2),
	.w3(32'h3adb9e25),
	.w4(32'hb81472fe),
	.w5(32'h39cab87f),
	.w6(32'hba5c39a0),
	.w7(32'h39cf3cb0),
	.w8(32'h3ac6cb88),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb832cf97),
	.w1(32'h39732924),
	.w2(32'h3a8fc2c1),
	.w3(32'h39ca0482),
	.w4(32'h3a21f356),
	.w5(32'h3af57cac),
	.w6(32'hb98a28d7),
	.w7(32'h39ee8639),
	.w8(32'h3ae208f8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47419),
	.w1(32'h3a8d9332),
	.w2(32'h3b14a891),
	.w3(32'h3ab03a8a),
	.w4(32'h3af19f2d),
	.w5(32'h395cc988),
	.w6(32'h3a6636bb),
	.w7(32'h3b070aff),
	.w8(32'h3921f54c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d27f5c),
	.w1(32'h3a305c91),
	.w2(32'hb9945494),
	.w3(32'hb856ea00),
	.w4(32'hba0b2990),
	.w5(32'h3ae836b1),
	.w6(32'h399239a3),
	.w7(32'hb9c600d5),
	.w8(32'h3aeffba1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0b4eb),
	.w1(32'h3ac9de1e),
	.w2(32'h3911b2d4),
	.w3(32'h3ab167e0),
	.w4(32'h3a81b834),
	.w5(32'h3b23d024),
	.w6(32'h3addff59),
	.w7(32'h3a49561e),
	.w8(32'h3b25f02b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afab72e),
	.w1(32'h3b0eb6ce),
	.w2(32'h3b18b618),
	.w3(32'h3b25c9cc),
	.w4(32'h3b1ad036),
	.w5(32'hb9b2ec45),
	.w6(32'h3b2636cf),
	.w7(32'h3b2a5d95),
	.w8(32'hba7240ce),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf74aac),
	.w1(32'hba966a35),
	.w2(32'hba043097),
	.w3(32'h38db547f),
	.w4(32'h3a767904),
	.w5(32'hb99e2dd0),
	.w6(32'hb98555de),
	.w7(32'hb9df7971),
	.w8(32'hba04dfec),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b271d),
	.w1(32'hba2ff79d),
	.w2(32'h39b59fdd),
	.w3(32'hba2d0bf7),
	.w4(32'hb9986738),
	.w5(32'hbaa14952),
	.w6(32'hb9f8ce71),
	.w7(32'hb84efdbd),
	.w8(32'hbaa513c9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d4d06),
	.w1(32'hbb33710f),
	.w2(32'hbb2bfbd1),
	.w3(32'hbae1db3a),
	.w4(32'hbac25114),
	.w5(32'hba8aaf95),
	.w6(32'hbb128317),
	.w7(32'hbaf52129),
	.w8(32'hba5f0af5),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a264c35),
	.w1(32'h3a50a6db),
	.w2(32'h3a77d108),
	.w3(32'h390fbf5f),
	.w4(32'h3aa8a58a),
	.w5(32'hb9128aab),
	.w6(32'h3a14e2e5),
	.w7(32'h3af44d5c),
	.w8(32'hb98a3898),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9583be4),
	.w1(32'hbaba42b5),
	.w2(32'hb91bd46d),
	.w3(32'hbaa3b186),
	.w4(32'hb9533df9),
	.w5(32'hb9989bd7),
	.w6(32'hbabdec36),
	.w7(32'hb9a6a330),
	.w8(32'hba190b8c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3859fd),
	.w1(32'hb98d45bf),
	.w2(32'hb9d2fc27),
	.w3(32'hbaa09ebf),
	.w4(32'hbad158ac),
	.w5(32'hba54691b),
	.w6(32'hba6a8cd5),
	.w7(32'hbaa9f036),
	.w8(32'hbac82114),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba583d74),
	.w1(32'hbad862a8),
	.w2(32'hba8a424c),
	.w3(32'hba22eaff),
	.w4(32'hb9aa8164),
	.w5(32'hba45e154),
	.w6(32'hbac8e812),
	.w7(32'hba14379e),
	.w8(32'hbad11866),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b446c2),
	.w1(32'h3813997c),
	.w2(32'hba09a0f3),
	.w3(32'hba9389ae),
	.w4(32'hba8c0117),
	.w5(32'h3b18e4db),
	.w6(32'hbad06070),
	.w7(32'hbb00be80),
	.w8(32'h3a8a9cd5),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33d6f3),
	.w1(32'hba8e7f0c),
	.w2(32'h3b22d1d1),
	.w3(32'h3b6e4836),
	.w4(32'h3b443e53),
	.w5(32'h39312bd4),
	.w6(32'h3a3a1bef),
	.w7(32'h3b6438f2),
	.w8(32'h3b3d462c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c7027),
	.w1(32'h39670fb5),
	.w2(32'hb9391e8e),
	.w3(32'h3987979d),
	.w4(32'h37949b9b),
	.w5(32'hb78c05e2),
	.w6(32'h39810ef3),
	.w7(32'hb82cda4c),
	.w8(32'h3a20de1c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac122f),
	.w1(32'h382455aa),
	.w2(32'hba61e5dd),
	.w3(32'hba9ac37e),
	.w4(32'hbafdde4b),
	.w5(32'h3a84f0dc),
	.w6(32'h3aa336ab),
	.w7(32'hba188122),
	.w8(32'hba8d18c4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule