module layer_10_featuremap_180(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ea84f),
	.w1(32'hbcdde444),
	.w2(32'h3d013200),
	.w3(32'h3bff1b97),
	.w4(32'hbc387b98),
	.w5(32'hbbda95f0),
	.w6(32'hbbc91889),
	.w7(32'hbbcb797f),
	.w8(32'hbb4ddbd1),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f057),
	.w1(32'hbbb4fa4e),
	.w2(32'h3bd7b8a9),
	.w3(32'h3ab1f2b5),
	.w4(32'hb8d160a5),
	.w5(32'h3bab333c),
	.w6(32'hbb0b9f3a),
	.w7(32'h3aaf9b88),
	.w8(32'h3b6ef6d0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4f07),
	.w1(32'h3bbe2302),
	.w2(32'hbb61e8fa),
	.w3(32'h3a5b5176),
	.w4(32'h3b0f4dfb),
	.w5(32'h3934d423),
	.w6(32'hb8f89c37),
	.w7(32'hbbae227b),
	.w8(32'hbba76dc5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73d82),
	.w1(32'hbcb51e72),
	.w2(32'h3a11d256),
	.w3(32'hbad60400),
	.w4(32'hbb8e9ce3),
	.w5(32'h39ca895e),
	.w6(32'hbc04bc78),
	.w7(32'hbb217fba),
	.w8(32'h3bdc0dd3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d7a2c),
	.w1(32'hbb251449),
	.w2(32'hbcdaddb9),
	.w3(32'h3b967e31),
	.w4(32'hbbe37f69),
	.w5(32'h3af2703a),
	.w6(32'hbc1b764b),
	.w7(32'h3b7cb269),
	.w8(32'h3c039be9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c774893),
	.w1(32'hbced41c8),
	.w2(32'hbc1aac37),
	.w3(32'h3c15d2f7),
	.w4(32'hbc60ab42),
	.w5(32'h3b106ac2),
	.w6(32'hbca25233),
	.w7(32'hbc07b7d9),
	.w8(32'h3b95b06c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c78d798),
	.w1(32'hbb828bbd),
	.w2(32'hbc9bc9f3),
	.w3(32'h3c23541d),
	.w4(32'hbbda00fa),
	.w5(32'hbb7eb64a),
	.w6(32'hbbf9e824),
	.w7(32'hbc05a4c7),
	.w8(32'hbbd7f77f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce351a),
	.w1(32'h3a673032),
	.w2(32'h3aada2a4),
	.w3(32'hbb656a35),
	.w4(32'h3b817201),
	.w5(32'h3b882db6),
	.w6(32'hbb3d0bff),
	.w7(32'hbb7a5e7d),
	.w8(32'hba2d0aff),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b71a9),
	.w1(32'hbbaa0f3b),
	.w2(32'hbb5a456c),
	.w3(32'h3b91b071),
	.w4(32'hbb67072d),
	.w5(32'hbb8df189),
	.w6(32'hbb123c55),
	.w7(32'hbbdd8edd),
	.w8(32'hbb2a9c9c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3243bc),
	.w1(32'h3bb583aa),
	.w2(32'hbb9221c5),
	.w3(32'h3923cf02),
	.w4(32'h3b347548),
	.w5(32'hbc38c827),
	.w6(32'h3bc05749),
	.w7(32'hbb5be70b),
	.w8(32'hbb88e00b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bbe49),
	.w1(32'h3be6c076),
	.w2(32'h3bba562b),
	.w3(32'hbb002c89),
	.w4(32'hba93982b),
	.w5(32'h3b2222a2),
	.w6(32'hbb9f10a1),
	.w7(32'hba5bf912),
	.w8(32'h3aa5da8b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea03d1),
	.w1(32'h3b8d5419),
	.w2(32'hbbf84af0),
	.w3(32'h3c22a55e),
	.w4(32'h3b985b31),
	.w5(32'h391146a0),
	.w6(32'hbbb155e0),
	.w7(32'hbabd14f3),
	.w8(32'hbbe8d556),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22f19a),
	.w1(32'h3b05df06),
	.w2(32'hbb2c6bf6),
	.w3(32'hbb83ab4b),
	.w4(32'h395cee40),
	.w5(32'hbb4cb3ed),
	.w6(32'hba913eaf),
	.w7(32'hbb103a2f),
	.w8(32'hbba3f466),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917a3d1),
	.w1(32'h3cd2bf13),
	.w2(32'hba4c9a65),
	.w3(32'h3a1b885b),
	.w4(32'h3b5ac0ea),
	.w5(32'hbc835104),
	.w6(32'h3c17b6cc),
	.w7(32'hbbd9ac74),
	.w8(32'hbc861de0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1026c0),
	.w1(32'h3c185d46),
	.w2(32'h3b6baa1b),
	.w3(32'hbc9eddbc),
	.w4(32'h3c638af8),
	.w5(32'h3b16415a),
	.w6(32'hbc25c016),
	.w7(32'h3bc78cca),
	.w8(32'h3bfb1924),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13d8f7),
	.w1(32'hbbbebe98),
	.w2(32'h3b7eae3a),
	.w3(32'hbb03fa75),
	.w4(32'h3aa3f1a2),
	.w5(32'hbac3cc7c),
	.w6(32'hbb6099e5),
	.w7(32'hbb8fe14a),
	.w8(32'hba15e1b2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bbd86),
	.w1(32'hbb6441c5),
	.w2(32'h39787fbf),
	.w3(32'h3a84ca7f),
	.w4(32'h3b17f8cc),
	.w5(32'h3bde93f1),
	.w6(32'hbbbc7de1),
	.w7(32'h3bd7e07c),
	.w8(32'hbab3dc94),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d55ec),
	.w1(32'h3b2dd9e6),
	.w2(32'hbb1c2465),
	.w3(32'hbc04652f),
	.w4(32'h3a28c1a4),
	.w5(32'hbbb7b776),
	.w6(32'h3a16319b),
	.w7(32'hbb67c0a3),
	.w8(32'hbbecfcdf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba1db0),
	.w1(32'hb969f3f2),
	.w2(32'hb9deec6a),
	.w3(32'hbb5cd1a4),
	.w4(32'hb9883d56),
	.w5(32'hbaa7dace),
	.w6(32'hbb325c84),
	.w7(32'hb928ead0),
	.w8(32'hbbd46119),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca1894),
	.w1(32'hbb8c172d),
	.w2(32'hbbb55ae8),
	.w3(32'h3ab9d13b),
	.w4(32'hbb71ebe0),
	.w5(32'hbbaac92d),
	.w6(32'hbb60df32),
	.w7(32'hbbf5239b),
	.w8(32'hbb898e20),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac4854),
	.w1(32'h3ac80873),
	.w2(32'h3b13df9b),
	.w3(32'hbb4051cb),
	.w4(32'h3a68023b),
	.w5(32'h3ad009f1),
	.w6(32'hbb4a9995),
	.w7(32'hbaf3d2db),
	.w8(32'hba8dc711),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a1536),
	.w1(32'h3d361375),
	.w2(32'hb9caa9b2),
	.w3(32'h3a1988f9),
	.w4(32'h3a79dd45),
	.w5(32'h3b306ac7),
	.w6(32'h3c103364),
	.w7(32'hba7433ef),
	.w8(32'hbbda059f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c7b1f),
	.w1(32'h3b997bce),
	.w2(32'hbb7e0c64),
	.w3(32'hbc10b4db),
	.w4(32'h3b0aaed2),
	.w5(32'hbbbd3978),
	.w6(32'h3b5bee2d),
	.w7(32'h39a65fa5),
	.w8(32'hb7c09ae8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacd160),
	.w1(32'hbb481745),
	.w2(32'hba3901e9),
	.w3(32'hbb36083d),
	.w4(32'hba772a5f),
	.w5(32'hbb1198de),
	.w6(32'hbb2f43a7),
	.w7(32'hba5fd5d5),
	.w8(32'h3a2ef900),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39803aa3),
	.w1(32'hbc273dde),
	.w2(32'h39e9dc8d),
	.w3(32'h3a8cb47f),
	.w4(32'hbb27ccc2),
	.w5(32'hbc07679d),
	.w6(32'hbbb73000),
	.w7(32'hbb5e3228),
	.w8(32'h3bc96b97),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb96e8),
	.w1(32'h3b70b991),
	.w2(32'h368f65a0),
	.w3(32'hbb8f52df),
	.w4(32'hbbb9913b),
	.w5(32'hbb97808a),
	.w6(32'h3c0f0fc7),
	.w7(32'h3bc440a7),
	.w8(32'h3b537491),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e3e6),
	.w1(32'hbb77dfac),
	.w2(32'hbb807d78),
	.w3(32'h39e98576),
	.w4(32'hba943b4f),
	.w5(32'hbb039e58),
	.w6(32'hbb05319a),
	.w7(32'hbb6d2d39),
	.w8(32'hbadbb3df),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b5d3),
	.w1(32'hbbeb1431),
	.w2(32'hbafc5ff0),
	.w3(32'h3b139a37),
	.w4(32'hbbe08930),
	.w5(32'hbbaaa984),
	.w6(32'h3b96ae2f),
	.w7(32'h3b34f483),
	.w8(32'h3bc881a3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97ab2c),
	.w1(32'hba90f80a),
	.w2(32'hbbe250da),
	.w3(32'h3be6f806),
	.w4(32'h3a6e7542),
	.w5(32'hbad71465),
	.w6(32'hbadae134),
	.w7(32'hbb14e115),
	.w8(32'h3abd247c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b65b7),
	.w1(32'hba1c720d),
	.w2(32'hbb6ac4c7),
	.w3(32'h3aa86fd1),
	.w4(32'h3a6fcc10),
	.w5(32'hbb89c9b4),
	.w6(32'h3b02f913),
	.w7(32'h3ad8cf7b),
	.w8(32'hbadafc5e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba07a5f),
	.w1(32'hbadee7af),
	.w2(32'hbaaddbcd),
	.w3(32'hbbce602c),
	.w4(32'hbab8999c),
	.w5(32'hb907dd8e),
	.w6(32'hbb257b74),
	.w7(32'hbb176030),
	.w8(32'hba2af886),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf84052),
	.w1(32'hbb96096e),
	.w2(32'hbb0d5bf6),
	.w3(32'hba04dc4c),
	.w4(32'hbaadbff4),
	.w5(32'h389649e7),
	.w6(32'hbb7f1343),
	.w7(32'hbb2f0318),
	.w8(32'h38b7ee91),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93974b3),
	.w1(32'hbbd66b9f),
	.w2(32'hbd0152ad),
	.w3(32'h3a76c732),
	.w4(32'hbc1b4e18),
	.w5(32'hbcced610),
	.w6(32'hbb96af34),
	.w7(32'hbcf192db),
	.w8(32'hbca1a89a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fdb58),
	.w1(32'h3ae0697b),
	.w2(32'h3be49cbf),
	.w3(32'hbc4284bd),
	.w4(32'h3c3e3466),
	.w5(32'h3c6c735f),
	.w6(32'h3c005a2a),
	.w7(32'h3c6162ca),
	.w8(32'h3c0943ac),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0609),
	.w1(32'hbc57d842),
	.w2(32'h3bb7ccf0),
	.w3(32'h3bd80da2),
	.w4(32'hbba5740f),
	.w5(32'hbab12020),
	.w6(32'hbc0ea283),
	.w7(32'hb8edc4a3),
	.w8(32'h3c0f99b5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70c3bc),
	.w1(32'hbba66595),
	.w2(32'hbbcf3fc9),
	.w3(32'h3ba55365),
	.w4(32'hbb002b75),
	.w5(32'hbbb3a4d3),
	.w6(32'hbbb74a6c),
	.w7(32'hbb78909e),
	.w8(32'hbb6f371c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88ad9b),
	.w1(32'hbc3d5a5d),
	.w2(32'hbbb5fc5b),
	.w3(32'hbb57d95a),
	.w4(32'h3acb08a5),
	.w5(32'h3b011cce),
	.w6(32'hbc1dbba3),
	.w7(32'h3b8e8d74),
	.w8(32'h3c30bd80),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94e1f0),
	.w1(32'h3a8a6b34),
	.w2(32'hbb833ef8),
	.w3(32'h3b8a969f),
	.w4(32'h3abc15e7),
	.w5(32'h3b576fd7),
	.w6(32'h3afcc8d1),
	.w7(32'h3ae71e25),
	.w8(32'h3a7b4a69),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1e60f),
	.w1(32'hbbc43198),
	.w2(32'h3a9082c5),
	.w3(32'h3a09be00),
	.w4(32'hba9804a5),
	.w5(32'h3b76e206),
	.w6(32'h39b04ece),
	.w7(32'h3b892f52),
	.w8(32'h3c3f5b0b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac05a4),
	.w1(32'hbb52db23),
	.w2(32'hbbbfb3bb),
	.w3(32'h3b989e4c),
	.w4(32'hbafe19cf),
	.w5(32'hba01d37a),
	.w6(32'hbb686b4e),
	.w7(32'hb95723db),
	.w8(32'hbb039ee9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeaa63),
	.w1(32'hbb17428c),
	.w2(32'hbb71171d),
	.w3(32'hbab2b541),
	.w4(32'h39d4fdf1),
	.w5(32'hbb2bf0e6),
	.w6(32'hba1dc730),
	.w7(32'h3a0f9fd6),
	.w8(32'hba18ea81),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77390d),
	.w1(32'h38081f41),
	.w2(32'hba9fef37),
	.w3(32'hbb9eb189),
	.w4(32'h3a8f4053),
	.w5(32'hba231cff),
	.w6(32'hbabedeb0),
	.w7(32'h3b1deec0),
	.w8(32'h3a367fd9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70197f),
	.w1(32'h39ce5383),
	.w2(32'hbaaa5c87),
	.w3(32'hbaa9bed5),
	.w4(32'h3a921cd5),
	.w5(32'hb961cc89),
	.w6(32'hb949a985),
	.w7(32'h3a956945),
	.w8(32'h3a8ba686),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc2f3d),
	.w1(32'h3c5bf53c),
	.w2(32'hbbda651c),
	.w3(32'h39788a1b),
	.w4(32'h3b689e7d),
	.w5(32'hbc31bf47),
	.w6(32'h3c4a4785),
	.w7(32'hb9ac60cd),
	.w8(32'hbbb5385e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accb808),
	.w1(32'h3d21fa64),
	.w2(32'h3c4701b6),
	.w3(32'hba45b412),
	.w4(32'h3c3f72d6),
	.w5(32'hbc405ca9),
	.w6(32'h3d0462a3),
	.w7(32'h3bd8c550),
	.w8(32'hbc51c4ca),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd428b7),
	.w1(32'h3cc7013f),
	.w2(32'hbcc14473),
	.w3(32'hbc8130b7),
	.w4(32'hbac2fda5),
	.w5(32'hbc314fbf),
	.w6(32'h3c1c92d5),
	.w7(32'hb957963c),
	.w8(32'hbc6afa26),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3e76d),
	.w1(32'hbb5a8e11),
	.w2(32'hb9bd3067),
	.w3(32'hbc23ccb3),
	.w4(32'h3b3d3ad4),
	.w5(32'h3c13fbd5),
	.w6(32'hbb865cf8),
	.w7(32'h3bf06526),
	.w8(32'h3a54647b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c677396),
	.w1(32'hbbc01090),
	.w2(32'hbbb9ffcf),
	.w3(32'h3886135c),
	.w4(32'hba831bff),
	.w5(32'hbb383781),
	.w6(32'hbba8bdbd),
	.w7(32'hbb803d67),
	.w8(32'hbc5377f5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12662b),
	.w1(32'hbb8a0c4a),
	.w2(32'hbbc50cc5),
	.w3(32'hbaea4577),
	.w4(32'hbacbe280),
	.w5(32'hbb2c4618),
	.w6(32'hbb32458a),
	.w7(32'hbb20ebb2),
	.w8(32'hb82c9f31),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21912b),
	.w1(32'h3c180d7e),
	.w2(32'h3a0345fb),
	.w3(32'hbae71bd2),
	.w4(32'h3b22eaba),
	.w5(32'hba021fa6),
	.w6(32'h3b90ac12),
	.w7(32'h3a94327c),
	.w8(32'hb9464f1a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c2e30),
	.w1(32'h3d2c014b),
	.w2(32'hbc56b75b),
	.w3(32'hba5a0524),
	.w4(32'h3cab776c),
	.w5(32'hbbf3dc92),
	.w6(32'h3c96ef66),
	.w7(32'h3aa3615b),
	.w8(32'hbc9ccf38),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf362e6),
	.w1(32'hbced9640),
	.w2(32'h3d2827eb),
	.w3(32'hbca938d8),
	.w4(32'hbc99c49d),
	.w5(32'hbc9025da),
	.w6(32'hbcc13df2),
	.w7(32'hbcd02664),
	.w8(32'hbbb83255),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dfc24),
	.w1(32'hbc8d8cfe),
	.w2(32'h3bd5109a),
	.w3(32'hbba24a2b),
	.w4(32'hbb0948f1),
	.w5(32'h3b728103),
	.w6(32'hbc3ceac8),
	.w7(32'hbbbf3946),
	.w8(32'hbb846698),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be22e5b),
	.w1(32'hbc56ac7c),
	.w2(32'hbca6d73e),
	.w3(32'hba9e16f7),
	.w4(32'hbc1a3fa3),
	.w5(32'hb9c2ef65),
	.w6(32'hbc9f61a2),
	.w7(32'hbc379a33),
	.w8(32'hb97c0706),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81aa80),
	.w1(32'hbc0eb50e),
	.w2(32'h3bbd2311),
	.w3(32'h3bb93ebd),
	.w4(32'h3a7060e0),
	.w5(32'h3bc6b5ee),
	.w6(32'hbbacf5bb),
	.w7(32'h39519869),
	.w8(32'hbaa2466f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b536563),
	.w1(32'hba03d8ec),
	.w2(32'hba840c29),
	.w3(32'h3a91faee),
	.w4(32'h3ad53773),
	.w5(32'h3b16bdb1),
	.w6(32'h3b85383e),
	.w7(32'hbb6f466a),
	.w8(32'hbab722a3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a7835),
	.w1(32'h3ceaf6f7),
	.w2(32'hbb36bc45),
	.w3(32'hbb01628a),
	.w4(32'h3bf5c17d),
	.w5(32'hbbec288c),
	.w6(32'h3c849f55),
	.w7(32'h3b2b9061),
	.w8(32'hbc970899),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07b8e4),
	.w1(32'hbc651d0e),
	.w2(32'hbccac8c8),
	.w3(32'hbcb1b667),
	.w4(32'hbc96614f),
	.w5(32'hbbd37e76),
	.w6(32'hbccc3503),
	.w7(32'hb703db91),
	.w8(32'hbc6eb3b0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d65c7),
	.w1(32'hbbbc0b57),
	.w2(32'h3b1a203c),
	.w3(32'hbc78f6c3),
	.w4(32'hba71c2cf),
	.w5(32'h3a88f30c),
	.w6(32'hbb23eb84),
	.w7(32'hbbcc46cf),
	.w8(32'hba701c54),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cc2f2),
	.w1(32'hbc0cb3b6),
	.w2(32'h3af4a8a9),
	.w3(32'h3b3cae05),
	.w4(32'hbb915679),
	.w5(32'hba091eaa),
	.w6(32'hbbadcade),
	.w7(32'hbb1bf8a5),
	.w8(32'h3b2515fd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45c8e8),
	.w1(32'h3969db72),
	.w2(32'h3ad007f4),
	.w3(32'h3b82a2b7),
	.w4(32'h3b1ebc8c),
	.w5(32'h3aca84db),
	.w6(32'hbaa88b0a),
	.w7(32'h3b804474),
	.w8(32'hbaf8cda8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bb7ae),
	.w1(32'hb897a3cc),
	.w2(32'h3ae45ab7),
	.w3(32'h3aca64d1),
	.w4(32'hbb8f5e64),
	.w5(32'hbabd4b19),
	.w6(32'hbaebd42d),
	.w7(32'hbacdf91b),
	.w8(32'h3a8cc046),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a9650),
	.w1(32'hbc60abe7),
	.w2(32'hbc9615a1),
	.w3(32'h3a6dfc61),
	.w4(32'hbbe7ba15),
	.w5(32'hbcb83fc3),
	.w6(32'hbc098853),
	.w7(32'hbc70471e),
	.w8(32'hbb7d5776),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0123b1),
	.w1(32'h3bc495fa),
	.w2(32'hbaea680f),
	.w3(32'hbbc020c7),
	.w4(32'h3b49c894),
	.w5(32'hbb45f4d8),
	.w6(32'h3bd6867c),
	.w7(32'h3af92ac2),
	.w8(32'h3b957007),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba916d2),
	.w1(32'hbae40978),
	.w2(32'hb91acd52),
	.w3(32'h3aec6536),
	.w4(32'h3abe918f),
	.w5(32'h3ae72eb4),
	.w6(32'hba9c5423),
	.w7(32'hbb3d944a),
	.w8(32'h3a6232d1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b000eff),
	.w1(32'h3c083453),
	.w2(32'hbc3fb16a),
	.w3(32'h3b18f1d0),
	.w4(32'h3b93114c),
	.w5(32'h3bedffb8),
	.w6(32'hbbb8c778),
	.w7(32'h3bf9cd64),
	.w8(32'hbb866846),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14f1fe),
	.w1(32'hbbd7f9ce),
	.w2(32'hbb360d94),
	.w3(32'h3a970237),
	.w4(32'hbb571016),
	.w5(32'hbb4362bb),
	.w6(32'hbb9900eb),
	.w7(32'hbb5a8c2e),
	.w8(32'hbb8d991b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd60e3),
	.w1(32'h36b07048),
	.w2(32'hbbe42362),
	.w3(32'hbc542261),
	.w4(32'hba8b9c9c),
	.w5(32'hbbce70bc),
	.w6(32'hbb144115),
	.w7(32'hbb046c2e),
	.w8(32'hbbe49539),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002154),
	.w1(32'hbbb3bf66),
	.w2(32'h3b1a167a),
	.w3(32'hbb2b55ef),
	.w4(32'hb7833b18),
	.w5(32'hba13d69c),
	.w6(32'hbb976df7),
	.w7(32'hbaf2835e),
	.w8(32'hbb1df52d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58adbf),
	.w1(32'h3d6ca76d),
	.w2(32'hbd18b47d),
	.w3(32'hbbade5c8),
	.w4(32'h3c792675),
	.w5(32'hbc664fee),
	.w6(32'h3cc94bbd),
	.w7(32'h3ba52d2e),
	.w8(32'hbcaa33e1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20b2d0),
	.w1(32'hbbce00b0),
	.w2(32'h3b4768c6),
	.w3(32'hbce2e81a),
	.w4(32'hbabc6d15),
	.w5(32'hba3da2e0),
	.w6(32'hbb6ea22b),
	.w7(32'hbb3ec7f1),
	.w8(32'h3a993c42),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7de0e2),
	.w1(32'hbbaf7ce4),
	.w2(32'hbb1f808e),
	.w3(32'hbac5f5e9),
	.w4(32'hbb478944),
	.w5(32'h3b7d4c90),
	.w6(32'hbba72f9e),
	.w7(32'h3a3a157a),
	.w8(32'h3b7a49bf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e589a),
	.w1(32'hbc15e6e3),
	.w2(32'h3b043575),
	.w3(32'h3b43366e),
	.w4(32'hbb3db383),
	.w5(32'h3a233a50),
	.w6(32'hbbe2f144),
	.w7(32'hbb328380),
	.w8(32'h3b4eef86),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ee15),
	.w1(32'hbba76e03),
	.w2(32'hbb89c445),
	.w3(32'h3b9ffd99),
	.w4(32'hba35d61a),
	.w5(32'hbb106c97),
	.w6(32'hbbb5d0b8),
	.w7(32'hbb9c9ba4),
	.w8(32'hbb39c7de),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dc7bf),
	.w1(32'hbbc62038),
	.w2(32'h3c27b286),
	.w3(32'hbaf9aa96),
	.w4(32'h3b3f265b),
	.w5(32'hba84cd3b),
	.w6(32'hbb8916de),
	.w7(32'hba6df1b3),
	.w8(32'h3a8fe0ee),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6b6e3),
	.w1(32'hbba6118d),
	.w2(32'hbc810871),
	.w3(32'h3b697eb5),
	.w4(32'hbbcf75ab),
	.w5(32'hbc74c4e1),
	.w6(32'h3c0ae186),
	.w7(32'hbc426f33),
	.w8(32'hbc9f7c87),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccbda71),
	.w1(32'h3c0f869f),
	.w2(32'hbb9534e8),
	.w3(32'hbc2676de),
	.w4(32'h3af8fc71),
	.w5(32'hbb10d59b),
	.w6(32'h3b62b77a),
	.w7(32'hbb16a220),
	.w8(32'hba0d5db8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4e02),
	.w1(32'h3b5d41d4),
	.w2(32'hbb338a81),
	.w3(32'h3b4fd2d9),
	.w4(32'h3b8d3c99),
	.w5(32'hbbc2b27e),
	.w6(32'h3c11f8f5),
	.w7(32'hbb514612),
	.w8(32'h3b8e920f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b675979),
	.w1(32'hbbe11464),
	.w2(32'h3b4a2511),
	.w3(32'h3b7b200d),
	.w4(32'h3b023aa1),
	.w5(32'h3b5ed495),
	.w6(32'hbb6de8b6),
	.w7(32'h3b95e350),
	.w8(32'hbb12816d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde4f26),
	.w1(32'hbbba5485),
	.w2(32'hbb3b1cf7),
	.w3(32'hbb09a35f),
	.w4(32'hbb48e867),
	.w5(32'hbabe0276),
	.w6(32'hbbb21c97),
	.w7(32'hbb3d48af),
	.w8(32'h39c55e99),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f0026),
	.w1(32'hbb13d311),
	.w2(32'hbad68b29),
	.w3(32'hb9ab1831),
	.w4(32'hba955091),
	.w5(32'h3a6a04cd),
	.w6(32'h3a4a2266),
	.w7(32'h3ad99263),
	.w8(32'hb90207a3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb264b8f),
	.w1(32'hbb423bf2),
	.w2(32'h3a7e4194),
	.w3(32'hbb0a59f6),
	.w4(32'hba982cb4),
	.w5(32'h39648eaf),
	.w6(32'hbb2afb78),
	.w7(32'hb9c84a4d),
	.w8(32'hbbdef828),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad85c4),
	.w1(32'hbb87801c),
	.w2(32'hb9b103ef),
	.w3(32'hbba13d7e),
	.w4(32'h36ca7ca1),
	.w5(32'hbbca71fe),
	.w6(32'hba70b19d),
	.w7(32'hba681148),
	.w8(32'h3a9854d7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3e3b5),
	.w1(32'hbb4dc1ae),
	.w2(32'h3bb8ac18),
	.w3(32'hbba1eb0c),
	.w4(32'hbab13d73),
	.w5(32'h3b5995f8),
	.w6(32'h3ad0fddf),
	.w7(32'h3ab37ae8),
	.w8(32'hbb867e67),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81cb89),
	.w1(32'hbc287860),
	.w2(32'hbb557104),
	.w3(32'h3aaba804),
	.w4(32'hbb9f5c25),
	.w5(32'h3aa48c7a),
	.w6(32'h3b0e8fba),
	.w7(32'h3c1c2111),
	.w8(32'h3b580daf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36be2d),
	.w1(32'h3b934d51),
	.w2(32'hbb06ce06),
	.w3(32'h3b9f4327),
	.w4(32'h39dddd6f),
	.w5(32'hb9231cac),
	.w6(32'h3b4074dd),
	.w7(32'hb9de49d1),
	.w8(32'hbc305e96),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc602f75),
	.w1(32'h3cc1e83a),
	.w2(32'h3bffc11d),
	.w3(32'hbc03e441),
	.w4(32'h3c588405),
	.w5(32'h3b0499b4),
	.w6(32'h3caefe6c),
	.w7(32'h3bdf70d4),
	.w8(32'hbbfef6f6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f6d59),
	.w1(32'hbaeb2c6f),
	.w2(32'hba44271d),
	.w3(32'hbac4fb19),
	.w4(32'hb9bda815),
	.w5(32'h392d4250),
	.w6(32'hbb2f988a),
	.w7(32'hbae99277),
	.w8(32'hba090f9f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa610b9),
	.w1(32'hbc5831ae),
	.w2(32'h3abdcfdf),
	.w3(32'hbb3debaf),
	.w4(32'hbba65c28),
	.w5(32'h3a9a5053),
	.w6(32'hbc26cd62),
	.w7(32'hbb468d2d),
	.w8(32'hba580002),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd07b8a),
	.w1(32'hbb0eea5f),
	.w2(32'hba8a0706),
	.w3(32'hb749beac),
	.w4(32'hbaed2016),
	.w5(32'h395d772d),
	.w6(32'hbbb37b9a),
	.w7(32'hbb9b414e),
	.w8(32'hbb671a94),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed8bf8),
	.w1(32'hba896c84),
	.w2(32'hb942a89f),
	.w3(32'h3b044a7f),
	.w4(32'h3a625140),
	.w5(32'h3a8f7be8),
	.w6(32'h3a67933f),
	.w7(32'h3a76a9fc),
	.w8(32'h3b343124),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb769943),
	.w1(32'h3c9245fe),
	.w2(32'hbc3c3824),
	.w3(32'h3b22ccdb),
	.w4(32'h3beb465a),
	.w5(32'hbc14c4ea),
	.w6(32'h3c137933),
	.w7(32'h3a5ee2ec),
	.w8(32'hbc44a794),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc812219),
	.w1(32'hbc76d3d5),
	.w2(32'h3c46f371),
	.w3(32'hbc7ba484),
	.w4(32'hbbafd3cc),
	.w5(32'h3c128169),
	.w6(32'hbbf3bdda),
	.w7(32'hbaa38aa2),
	.w8(32'h3bdef2c7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4898a3),
	.w1(32'hbb46b824),
	.w2(32'hbb981961),
	.w3(32'h3ad73152),
	.w4(32'hba9afc40),
	.w5(32'hbac2c17f),
	.w6(32'hbb9dfd9d),
	.w7(32'hbbcc81a5),
	.w8(32'hbb7d03b9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63cf03),
	.w1(32'hba27c2b5),
	.w2(32'hba9e0b20),
	.w3(32'h39d27180),
	.w4(32'hba9a1de7),
	.w5(32'hba7c82eb),
	.w6(32'h3a49c7c0),
	.w7(32'h3ae9ad16),
	.w8(32'h3ba2ac7a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81cca1),
	.w1(32'hbc693691),
	.w2(32'hbc3d1fd0),
	.w3(32'h3a617f12),
	.w4(32'hbc3921e1),
	.w5(32'h3c270c62),
	.w6(32'hbb4b9c37),
	.w7(32'hbb04dbff),
	.w8(32'h3b57c3ea),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b3b9d),
	.w1(32'hb98cdd27),
	.w2(32'hba8acbcd),
	.w3(32'h3c7b7b91),
	.w4(32'h3b613cce),
	.w5(32'hbbb4b33b),
	.w6(32'h3aaf5b81),
	.w7(32'hbb80fdf6),
	.w8(32'hbbfbd0cd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ffdf),
	.w1(32'hbc3bac44),
	.w2(32'hbc336ef0),
	.w3(32'hbb585070),
	.w4(32'hbc26f580),
	.w5(32'hbc8b8e4e),
	.w6(32'hbc41c101),
	.w7(32'hbcc166e5),
	.w8(32'h3a178588),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd4b80),
	.w1(32'hbc00a718),
	.w2(32'hba8ea994),
	.w3(32'h3c7dec78),
	.w4(32'h39d14dbc),
	.w5(32'h3b25a3ec),
	.w6(32'hbb0dd872),
	.w7(32'h3b260ea9),
	.w8(32'hba52f826),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f1f31),
	.w1(32'hbc15f266),
	.w2(32'h3c674b32),
	.w3(32'hbb8835ac),
	.w4(32'h3ba12d29),
	.w5(32'h3bf876ca),
	.w6(32'hbc3b22aa),
	.w7(32'h3a900a69),
	.w8(32'h3c24e7dd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c542625),
	.w1(32'h3ba5eec9),
	.w2(32'hbc5748f4),
	.w3(32'h3ac9a901),
	.w4(32'hbc4561a5),
	.w5(32'h3c1c2fc6),
	.w6(32'hbc472d43),
	.w7(32'h3c588c88),
	.w8(32'hbb7b9270),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b98cc),
	.w1(32'hbb7b3ba3),
	.w2(32'hbd0f7b0c),
	.w3(32'hbc852cb2),
	.w4(32'hbc858017),
	.w5(32'h3bee51b9),
	.w6(32'h3b1efadc),
	.w7(32'h3beab1f2),
	.w8(32'h3ac4d1b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd65a3),
	.w1(32'h3c54ceae),
	.w2(32'hbc091e9b),
	.w3(32'h3b8a0e09),
	.w4(32'h3b280b0e),
	.w5(32'hbb642b8e),
	.w6(32'h3bb44720),
	.w7(32'hba2b365e),
	.w8(32'h3b0aabd4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c5be2),
	.w1(32'hbbf058be),
	.w2(32'hbb829a7d),
	.w3(32'h3bd3769d),
	.w4(32'hbb86b0fc),
	.w5(32'h3b74c6c8),
	.w6(32'hbbad7656),
	.w7(32'h3783f243),
	.w8(32'h3b27e76b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f02ff),
	.w1(32'h3c0848db),
	.w2(32'h3b36f46a),
	.w3(32'h3873a9ce),
	.w4(32'h3c0640b4),
	.w5(32'h3b413799),
	.w6(32'hbb7a2b61),
	.w7(32'hbb0ee9f5),
	.w8(32'h3c1ba47d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d76c1),
	.w1(32'hbbc2bd19),
	.w2(32'hbc35820c),
	.w3(32'h3bbdf45d),
	.w4(32'hbbaf3437),
	.w5(32'hbc0191af),
	.w6(32'hbb6bcf38),
	.w7(32'hbbedbdac),
	.w8(32'hbbdf0f38),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f049c),
	.w1(32'h3b605b44),
	.w2(32'h3b7427a7),
	.w3(32'hbabdd54f),
	.w4(32'h3b64d151),
	.w5(32'h3b8e695f),
	.w6(32'h3a15c10a),
	.w7(32'hbac25d45),
	.w8(32'hbb2318ff),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a9e6),
	.w1(32'h39056196),
	.w2(32'h3af65c03),
	.w3(32'hba84e01b),
	.w4(32'h39b8e4c6),
	.w5(32'h3aea5d70),
	.w6(32'hbb287798),
	.w7(32'hba9351b3),
	.w8(32'hb892474e),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5dc388),
	.w1(32'h3be83945),
	.w2(32'hbbdd503c),
	.w3(32'h3a81a06c),
	.w4(32'hba97fa0a),
	.w5(32'hbb9b070d),
	.w6(32'h3b5cc14b),
	.w7(32'hbb257883),
	.w8(32'hbb781536),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f21b2),
	.w1(32'h3ceccbc6),
	.w2(32'h3c483961),
	.w3(32'h3b1d66a1),
	.w4(32'h3c4172be),
	.w5(32'hbbcab370),
	.w6(32'h3cb2eeac),
	.w7(32'hb9c3d713),
	.w8(32'hbc821f5b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0d247),
	.w1(32'hbc2b25e0),
	.w2(32'h3bc51ee5),
	.w3(32'hbc174ba3),
	.w4(32'hbb2eaf98),
	.w5(32'h3a8b0239),
	.w6(32'hbbcb71fe),
	.w7(32'hbbdd556a),
	.w8(32'h3bb33de2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b489805),
	.w1(32'hbc35d458),
	.w2(32'h3d12f626),
	.w3(32'h3b160626),
	.w4(32'hbbe5ae49),
	.w5(32'hbccd38a2),
	.w6(32'hbbce50e4),
	.w7(32'hbc85beeb),
	.w8(32'h3b29e30a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26ec99),
	.w1(32'hbc491a3e),
	.w2(32'h3ab58028),
	.w3(32'hbbcd191c),
	.w4(32'hbb634f0e),
	.w5(32'hbaad81b8),
	.w6(32'hbc4a3373),
	.w7(32'hbbefc122),
	.w8(32'hba12b8a2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4654c),
	.w1(32'h3bde5b24),
	.w2(32'h39e3e605),
	.w3(32'h3b8746cc),
	.w4(32'h3b979797),
	.w5(32'hba808173),
	.w6(32'hb9be2372),
	.w7(32'h3b088bde),
	.w8(32'h3bb718b2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb056),
	.w1(32'h3c926f01),
	.w2(32'hbb1d005d),
	.w3(32'hbabdc93b),
	.w4(32'h3b5c8553),
	.w5(32'hbc652b4a),
	.w6(32'h3be64a09),
	.w7(32'hbab79912),
	.w8(32'hbbe074ff),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc352ef6),
	.w1(32'h3c0e1123),
	.w2(32'hbbb75aa3),
	.w3(32'hbba89e2a),
	.w4(32'hb89356ed),
	.w5(32'hbb088f52),
	.w6(32'h3b964c66),
	.w7(32'hba128988),
	.w8(32'h3b0876e7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22eb4b),
	.w1(32'hbba2169e),
	.w2(32'hbb32cd84),
	.w3(32'h3b97e9cd),
	.w4(32'hbad48e5a),
	.w5(32'h3a200ded),
	.w6(32'hbba74248),
	.w7(32'hba3d26e9),
	.w8(32'h3b5ec72d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b340feb),
	.w1(32'hbc15519b),
	.w2(32'hbb0d02ef),
	.w3(32'h3b7ddb24),
	.w4(32'hbb84e7df),
	.w5(32'h3ab360de),
	.w6(32'hbbfb7cd6),
	.w7(32'hbb1bca6b),
	.w8(32'h3ba24045),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d719),
	.w1(32'h3c40799f),
	.w2(32'h3b27ff3b),
	.w3(32'h3bf9e70d),
	.w4(32'hbadd14bf),
	.w5(32'hbb8a4b15),
	.w6(32'hb942d9e6),
	.w7(32'hbb2840da),
	.w8(32'hba2fdc73),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94d905),
	.w1(32'h3b7e652a),
	.w2(32'hbc47677e),
	.w3(32'hbb4791c5),
	.w4(32'hba48cc56),
	.w5(32'hbb2c6203),
	.w6(32'hbbfd5761),
	.w7(32'hb8e442ee),
	.w8(32'hbbdb06b9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf14cc6),
	.w1(32'hbbff5a76),
	.w2(32'hba9bfdfa),
	.w3(32'hbb12e86f),
	.w4(32'hbc02986e),
	.w5(32'h39e6cb14),
	.w6(32'hbbd09a30),
	.w7(32'hbade2ea5),
	.w8(32'h3aff5265),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c249c10),
	.w1(32'hbc216736),
	.w2(32'h3991ac15),
	.w3(32'h3b62d293),
	.w4(32'hbb454fb9),
	.w5(32'hbb399a87),
	.w6(32'hbc0867dd),
	.w7(32'hbc4f44e4),
	.w8(32'hbba845d4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70b843),
	.w1(32'hbb8cc82c),
	.w2(32'h3ad71102),
	.w3(32'hbbab06a4),
	.w4(32'hbb28f0ed),
	.w5(32'h3adce503),
	.w6(32'hbae116a8),
	.w7(32'h3aa23d18),
	.w8(32'h3bcdbc22),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab59e4d),
	.w1(32'hbc6bae2e),
	.w2(32'hbcce079f),
	.w3(32'h3b8ac15c),
	.w4(32'hbc87aceb),
	.w5(32'h3a5c005a),
	.w6(32'h3b910151),
	.w7(32'h3bde33a7),
	.w8(32'hbb028e9b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1040a8),
	.w1(32'hbce58b10),
	.w2(32'hba74373e),
	.w3(32'h3bac79d3),
	.w4(32'hbc045534),
	.w5(32'h3c55473b),
	.w6(32'hbc87e18f),
	.w7(32'hbc0b40a2),
	.w8(32'h369305b4),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5319f),
	.w1(32'hbba1a2e5),
	.w2(32'hbb4330ad),
	.w3(32'h3bcc0a13),
	.w4(32'hbabef3b4),
	.w5(32'hbaf27bfd),
	.w6(32'hbb9cf125),
	.w7(32'hbb821370),
	.w8(32'hba4e37a4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c568),
	.w1(32'h3a810961),
	.w2(32'h3bd25c97),
	.w3(32'hbac75dd5),
	.w4(32'hbacb9a63),
	.w5(32'h3b980219),
	.w6(32'hbb73e2ef),
	.w7(32'h3add6fbf),
	.w8(32'hbb043a59),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0427da),
	.w1(32'hbabc70d9),
	.w2(32'hbb300ebb),
	.w3(32'hbb3f395a),
	.w4(32'hbbe0f3ec),
	.w5(32'hbaaaf84e),
	.w6(32'hbc1fe448),
	.w7(32'hbbfc3d2e),
	.w8(32'hbc4da1fb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e050bf),
	.w1(32'h3a615219),
	.w2(32'h3bb67cb4),
	.w3(32'hbb1da60e),
	.w4(32'hbb11de5c),
	.w5(32'hbb566e81),
	.w6(32'hb966e956),
	.w7(32'h3a6551e4),
	.w8(32'hbb394f5f),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be17fd1),
	.w1(32'hbbd12ab3),
	.w2(32'hbbb6a63b),
	.w3(32'hbb99f534),
	.w4(32'hbbb323f1),
	.w5(32'hbbb54e34),
	.w6(32'hbba55ae8),
	.w7(32'hbbd6730e),
	.w8(32'hbbbf3055),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09ede4),
	.w1(32'hbb4793f1),
	.w2(32'hbadb9008),
	.w3(32'hbbd6770b),
	.w4(32'hba866c14),
	.w5(32'hbad122d7),
	.w6(32'hbb44a913),
	.w7(32'hbb4ca8e2),
	.w8(32'hbbb1aed9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fd9d0),
	.w1(32'h3b6cf7de),
	.w2(32'h3bb97bb8),
	.w3(32'hbb28c925),
	.w4(32'h3c595b9b),
	.w5(32'h3c5faca3),
	.w6(32'h3acd54e9),
	.w7(32'h3ba6ef1c),
	.w8(32'h3b7c8a17),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd61c67),
	.w1(32'h3b93d783),
	.w2(32'h3b1509ff),
	.w3(32'h3c438ed9),
	.w4(32'h3be02726),
	.w5(32'h3bad7def),
	.w6(32'hbb6af992),
	.w7(32'hba09f9cf),
	.w8(32'hbb1c6f5b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8073f0),
	.w1(32'hbaad68d4),
	.w2(32'h3c0114a6),
	.w3(32'h3b3e898c),
	.w4(32'hbb45ec88),
	.w5(32'h3b91799c),
	.w6(32'hbb3c6861),
	.w7(32'h3bb8e0f9),
	.w8(32'hba228009),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08624),
	.w1(32'hbc0f9f1c),
	.w2(32'hbc7bb046),
	.w3(32'h3b3da054),
	.w4(32'hbbd13eea),
	.w5(32'hbc612883),
	.w6(32'hbbd355a4),
	.w7(32'hbc4f4a28),
	.w8(32'hbc47efd1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53a0bc),
	.w1(32'hbacaa8c4),
	.w2(32'h38d5fc28),
	.w3(32'hbc268305),
	.w4(32'hbb1357c9),
	.w5(32'h3a219954),
	.w6(32'hbbaf3a77),
	.w7(32'hbac2c810),
	.w8(32'hbbb0df15),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21a5fe),
	.w1(32'h3b7d8068),
	.w2(32'h3ba5ad2c),
	.w3(32'hbb6513bc),
	.w4(32'h3b523f5d),
	.w5(32'h3b7f89a9),
	.w6(32'h39d25b70),
	.w7(32'h3b632306),
	.w8(32'hba997515),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4145e),
	.w1(32'hbba69c83),
	.w2(32'hbbfb0a58),
	.w3(32'h39ff2e75),
	.w4(32'h3ab8dca0),
	.w5(32'hbb48437f),
	.w6(32'hb9ed61e8),
	.w7(32'hbbd3d783),
	.w8(32'hbb868dbc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7172a),
	.w1(32'h3baf39c3),
	.w2(32'h3c0439e4),
	.w3(32'hbb3dd31d),
	.w4(32'hbba88f1f),
	.w5(32'hbb839d3a),
	.w6(32'h3b7c9395),
	.w7(32'h3bc57176),
	.w8(32'h3b378a68),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2cbe9),
	.w1(32'h3a679f42),
	.w2(32'hba95d108),
	.w3(32'hbbcde740),
	.w4(32'h3c0fd6e9),
	.w5(32'h3c7f42a2),
	.w6(32'hbb954b23),
	.w7(32'hbba862d5),
	.w8(32'hbc0a63ed),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8439ba),
	.w1(32'h3ac691ae),
	.w2(32'h3badb5af),
	.w3(32'h3c49995b),
	.w4(32'hbb7be367),
	.w5(32'hbb330c16),
	.w6(32'hb95942ab),
	.w7(32'h3b78561d),
	.w8(32'hb9b282b3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd4b4c),
	.w1(32'h3c1ee96d),
	.w2(32'h3c85cc14),
	.w3(32'hba27b969),
	.w4(32'h3bda6de9),
	.w5(32'h3c7e6079),
	.w6(32'h3c1cbc07),
	.w7(32'h3c2affe8),
	.w8(32'h3c0cf3db),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c929d7c),
	.w1(32'h3b87235c),
	.w2(32'h3b9e8771),
	.w3(32'h3c30f9e1),
	.w4(32'h3c55d49b),
	.w5(32'h3c96514a),
	.w6(32'hbb9442e7),
	.w7(32'h3ada6941),
	.w8(32'hbbd3ac18),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a033dc4),
	.w1(32'h3b6aef10),
	.w2(32'h3ba90af4),
	.w3(32'h3ba5dddc),
	.w4(32'h3a8fd075),
	.w5(32'h3b60be2f),
	.w6(32'h3a4cd5c5),
	.w7(32'h3b5ad93c),
	.w8(32'hbb1980d2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c52ad1),
	.w1(32'h3c055c70),
	.w2(32'h3bb8e653),
	.w3(32'hbb045de6),
	.w4(32'h3b52c8da),
	.w5(32'hba819157),
	.w6(32'h3c01d80b),
	.w7(32'h3bb33560),
	.w8(32'h3b86f537),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0b7d4),
	.w1(32'hbbb17ab5),
	.w2(32'hbbfa2a02),
	.w3(32'h3a33eaf2),
	.w4(32'hba87276b),
	.w5(32'hbba508ac),
	.w6(32'h3a9c4055),
	.w7(32'hbb84c60b),
	.w8(32'hbab4c168),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd3961),
	.w1(32'hbb0a57fe),
	.w2(32'hbb2f5690),
	.w3(32'hbb8e50ed),
	.w4(32'hba46d2aa),
	.w5(32'hbb011481),
	.w6(32'h3a842b1e),
	.w7(32'hb9bffaa5),
	.w8(32'hbaa236f1),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65354c),
	.w1(32'hb8d67362),
	.w2(32'h38d3a432),
	.w3(32'hbb378105),
	.w4(32'hbb09ed9a),
	.w5(32'hbb15e610),
	.w6(32'hba982b85),
	.w7(32'hbadd71ff),
	.w8(32'hbbe1c4af),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3120c5),
	.w1(32'h3adc2546),
	.w2(32'h3be98c2e),
	.w3(32'hbb165082),
	.w4(32'hba87a164),
	.w5(32'h3baf461d),
	.w6(32'hbad30cae),
	.w7(32'h3b8bbb2c),
	.w8(32'h3b16bc87),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0614a),
	.w1(32'h3bfe39a1),
	.w2(32'h3c838f57),
	.w3(32'h3be5f67c),
	.w4(32'hbb447644),
	.w5(32'h3b0d5ca4),
	.w6(32'hbb3570b9),
	.w7(32'h3b4846c8),
	.w8(32'hbbb5d9c0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38f1b6),
	.w1(32'h3b19aaa5),
	.w2(32'hbb2a43a6),
	.w3(32'h3b89bf5c),
	.w4(32'h3b2ca613),
	.w5(32'hbb2f5879),
	.w6(32'h3b9ac961),
	.w7(32'h3a16b3af),
	.w8(32'h3af4bc7d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e66c),
	.w1(32'hbb8da838),
	.w2(32'hbb1df306),
	.w3(32'h3b5cdc65),
	.w4(32'hbb96dc90),
	.w5(32'hbba3c43c),
	.w6(32'hbc332abf),
	.w7(32'hbbeb86ea),
	.w8(32'hbc118748),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77d4cd),
	.w1(32'hba8b05e0),
	.w2(32'hbb850e81),
	.w3(32'hbb845a94),
	.w4(32'hbbb06b0e),
	.w5(32'hbba13cee),
	.w6(32'h3bae7e2c),
	.w7(32'h3ae09ed9),
	.w8(32'hbb61f7e5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd0d57),
	.w1(32'h3a9fd092),
	.w2(32'hb9f0c022),
	.w3(32'hbbc6bf21),
	.w4(32'h3b26e361),
	.w5(32'h3a6c0d39),
	.w6(32'h3abdd265),
	.w7(32'hbaa908bf),
	.w8(32'hbaed0d5b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9232d57),
	.w1(32'h3aa2ebbe),
	.w2(32'h3b54b854),
	.w3(32'h38a6b27a),
	.w4(32'h395a0640),
	.w5(32'h3b378b6f),
	.w6(32'hba666c69),
	.w7(32'h3a69fb62),
	.w8(32'hbab4c9d2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a241c),
	.w1(32'hbbbec72d),
	.w2(32'hbbd33928),
	.w3(32'hbabefd2b),
	.w4(32'hbbbaa79f),
	.w5(32'hbb8ae576),
	.w6(32'hbbb5f929),
	.w7(32'hbb9d0f93),
	.w8(32'hbc1f030b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18597c),
	.w1(32'hbbf21047),
	.w2(32'hbbf0717d),
	.w3(32'hbbd24f6a),
	.w4(32'hbb9ad584),
	.w5(32'hbbb6bb9c),
	.w6(32'hbb2e4897),
	.w7(32'hbb68997f),
	.w8(32'h3b44389a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba000f4e),
	.w1(32'h3b6b2a5b),
	.w2(32'h3abea7a8),
	.w3(32'h3aa5b9af),
	.w4(32'h3bb16c8a),
	.w5(32'h3b859f3c),
	.w6(32'h3b5c47fc),
	.w7(32'h3b51076a),
	.w8(32'h3b743afd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d4d10),
	.w1(32'h3b72c42f),
	.w2(32'h3c0219a6),
	.w3(32'h3b69a383),
	.w4(32'h3aa11e30),
	.w5(32'h3b8489e5),
	.w6(32'h3a67eaa2),
	.w7(32'h3b9a9ebe),
	.w8(32'h3b456f6d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8e757),
	.w1(32'hbb023f90),
	.w2(32'h3ae20bf6),
	.w3(32'h3af3beab),
	.w4(32'hbac9a8c9),
	.w5(32'h3ab63283),
	.w6(32'hbb6cc4af),
	.w7(32'hb9b76987),
	.w8(32'hb8e25fe4),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af479cc),
	.w1(32'hba8bc346),
	.w2(32'h3baa1664),
	.w3(32'h3a3ee7dd),
	.w4(32'hbb1b5932),
	.w5(32'h3a77fdd1),
	.w6(32'hbb21f201),
	.w7(32'h3980f862),
	.w8(32'hbb02e70e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866170),
	.w1(32'hbb0e3d24),
	.w2(32'hbb223aa1),
	.w3(32'h3b027817),
	.w4(32'hba52913f),
	.w5(32'hba863cab),
	.w6(32'h38125966),
	.w7(32'hbb9eed9a),
	.w8(32'hbc0492de),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9adca),
	.w1(32'hbc336f4e),
	.w2(32'hbc60f241),
	.w3(32'hbbca8141),
	.w4(32'hbc1b5f1b),
	.w5(32'hbc396c80),
	.w6(32'hbbbd1840),
	.w7(32'hbc1bf706),
	.w8(32'hbc286646),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6efa79),
	.w1(32'h3a0b0e95),
	.w2(32'h3adac4a8),
	.w3(32'hbc33a6ae),
	.w4(32'hbb80c874),
	.w5(32'hbab2517d),
	.w6(32'hbab323e1),
	.w7(32'h3ac0e156),
	.w8(32'hba77705e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fef60),
	.w1(32'hbc147743),
	.w2(32'hbbea476c),
	.w3(32'hbae86765),
	.w4(32'hbc0c6cb6),
	.w5(32'hbc0ef4bc),
	.w6(32'hbbbd28ef),
	.w7(32'hbbb46928),
	.w8(32'hbb6e0279),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb658765),
	.w1(32'hbbce4f48),
	.w2(32'hbc1c1a88),
	.w3(32'hbbabd64c),
	.w4(32'hbb92d1fd),
	.w5(32'hbc0ab39e),
	.w6(32'hbb2caaac),
	.w7(32'hbc00b4c1),
	.w8(32'hbbdc8fdf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e1811),
	.w1(32'hbb61c8e5),
	.w2(32'hbb02941a),
	.w3(32'hbbfd18ee),
	.w4(32'hbb98ba46),
	.w5(32'hbb2fae31),
	.w6(32'hbbd1f66a),
	.w7(32'hbb8052ba),
	.w8(32'hbbe605c4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3987),
	.w1(32'hbb8c238c),
	.w2(32'hbb983a73),
	.w3(32'hbbd816fa),
	.w4(32'hbb405ff0),
	.w5(32'hbba0b082),
	.w6(32'hba94a237),
	.w7(32'hbb4be79a),
	.w8(32'hbb1ce8a6),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b4249),
	.w1(32'h3aaf27d7),
	.w2(32'hbbb62960),
	.w3(32'hbb879319),
	.w4(32'h3af02a1e),
	.w5(32'hbaa39bf6),
	.w6(32'h3ac47197),
	.w7(32'hbb1e56d1),
	.w8(32'hbbb7284a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a956e),
	.w1(32'hbbeaf61e),
	.w2(32'hbb343cf8),
	.w3(32'h3ad891b6),
	.w4(32'hbc410ae3),
	.w5(32'hbc211a85),
	.w6(32'hbbf4b64c),
	.w7(32'hbb3d1835),
	.w8(32'hbbdf06dc),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf97791),
	.w1(32'hbbaaf2a8),
	.w2(32'hba9448e9),
	.w3(32'hbc750e8b),
	.w4(32'hbba0575a),
	.w5(32'hbb48880b),
	.w6(32'hbaf3b4dc),
	.w7(32'h3a07a043),
	.w8(32'h389ebd60),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55abc9),
	.w1(32'h3bb5e20c),
	.w2(32'hbb180c34),
	.w3(32'h3acfd7cc),
	.w4(32'h3c26eef0),
	.w5(32'h3b1e19f3),
	.w6(32'h3c79b19e),
	.w7(32'h3b9920e2),
	.w8(32'h3bd85b46),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f7e71),
	.w1(32'hbb069611),
	.w2(32'h3bed2855),
	.w3(32'h3b2847ef),
	.w4(32'hbc39e6bd),
	.w5(32'hbc3bad7a),
	.w6(32'h3b4025a3),
	.w7(32'h3c1d8c7e),
	.w8(32'h3c19f6ac),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4160),
	.w1(32'h3b70f874),
	.w2(32'h396f3cdc),
	.w3(32'hbb93eb9b),
	.w4(32'hbb8f5f07),
	.w5(32'hbc2cf8a3),
	.w6(32'h3babcf72),
	.w7(32'h3b68a48d),
	.w8(32'hbb1ae4f7),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd27ab4),
	.w1(32'h39b3de7d),
	.w2(32'hbb21687d),
	.w3(32'hbc5b2399),
	.w4(32'h3c6901a8),
	.w5(32'h3c54dec8),
	.w6(32'hbbff0b0f),
	.w7(32'hbc30fb49),
	.w8(32'hbc54a65b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b958698),
	.w1(32'h39ea11f7),
	.w2(32'hb80b0611),
	.w3(32'h3c7de5f7),
	.w4(32'h3aa93200),
	.w5(32'h39c6e8a2),
	.w6(32'h3b93b67e),
	.w7(32'h3b66a96c),
	.w8(32'h3b904ccf),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c7798),
	.w1(32'hbbc8970e),
	.w2(32'hbb06e409),
	.w3(32'h3b5bcd8b),
	.w4(32'hbb7e898f),
	.w5(32'hbae8295d),
	.w6(32'hbb7da315),
	.w7(32'hbb1b80ad),
	.w8(32'hbb0e19cb),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7153b9f),
	.w1(32'h3af7b99a),
	.w2(32'h3b907d17),
	.w3(32'hb9d1a3d7),
	.w4(32'hb9a33ef3),
	.w5(32'h3b1d283e),
	.w6(32'hbb6f3a11),
	.w7(32'hb98034ed),
	.w8(32'hbb3feaf7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b419c40),
	.w1(32'h3c162373),
	.w2(32'h3bd95d09),
	.w3(32'hba68d81a),
	.w4(32'h3c2a712e),
	.w5(32'h3be9f76b),
	.w6(32'h3b855e72),
	.w7(32'h3a95b01c),
	.w8(32'hbb9b63a7),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20bad1),
	.w1(32'h3a8a5d8a),
	.w2(32'h394fb482),
	.w3(32'hbb2f83ea),
	.w4(32'h3b32846c),
	.w5(32'h3c14f469),
	.w6(32'h3b6273f5),
	.w7(32'h3a2a81ea),
	.w8(32'hbba6a6eb),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89ea6),
	.w1(32'h3c031565),
	.w2(32'h3c84a225),
	.w3(32'h3c151447),
	.w4(32'h3b55a92c),
	.w5(32'h3c1e2f6c),
	.w6(32'h3af4abd1),
	.w7(32'h3c240461),
	.w8(32'h3b06fbc8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a6228),
	.w1(32'hbc1c0e4e),
	.w2(32'hbbeba67f),
	.w3(32'h3b1d0d10),
	.w4(32'hbc128b1b),
	.w5(32'hbbd0c3e3),
	.w6(32'hbc076aac),
	.w7(32'hbbce01a3),
	.w8(32'hbb767bae),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b302d),
	.w1(32'h3b04ceaf),
	.w2(32'hbaaa417a),
	.w3(32'hbb7a6a83),
	.w4(32'h3a89aed6),
	.w5(32'hba79e930),
	.w6(32'h3b33de21),
	.w7(32'hba367d66),
	.w8(32'hb9d8cbaf),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9b4c3),
	.w1(32'hbb5e453c),
	.w2(32'hbbdccf28),
	.w3(32'hb9e97e24),
	.w4(32'hbb4250d1),
	.w5(32'hbb6102fd),
	.w6(32'hbb8163f4),
	.w7(32'hbba0cc80),
	.w8(32'hbb0129f7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16bfb4),
	.w1(32'h3b81e7ed),
	.w2(32'h3c29f174),
	.w3(32'hbb2c8f0c),
	.w4(32'hbbc0658f),
	.w5(32'hbb3a8259),
	.w6(32'hba46a2c5),
	.w7(32'h3add1c91),
	.w8(32'hbb97cb79),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba158a9e),
	.w1(32'h3c6df29c),
	.w2(32'h3c6bec47),
	.w3(32'hbbe81952),
	.w4(32'h3c92e8d8),
	.w5(32'h3ca96463),
	.w6(32'h3aa08ed0),
	.w7(32'h3bfc51ba),
	.w8(32'hbb2613f9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c4273),
	.w1(32'hbc0905ce),
	.w2(32'hbc23bcb6),
	.w3(32'h3b209634),
	.w4(32'hbbd2a7ee),
	.w5(32'hbc01887a),
	.w6(32'hbbade85e),
	.w7(32'hbbf964e8),
	.w8(32'hbbf69aed),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2a66),
	.w1(32'hbbb05d3c),
	.w2(32'hbbf956d6),
	.w3(32'hbc31c09c),
	.w4(32'hbc215da2),
	.w5(32'hbc34074b),
	.w6(32'hbc45dee4),
	.w7(32'hbc3fdf42),
	.w8(32'hbc9309bd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a490),
	.w1(32'hbba32285),
	.w2(32'hbbc0491a),
	.w3(32'hbb8c36b2),
	.w4(32'hbb24e32d),
	.w5(32'hbb9f4daa),
	.w6(32'h3b874819),
	.w7(32'h3a15d4f7),
	.w8(32'hba12d2a9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcc4d3),
	.w1(32'hbb5c59e1),
	.w2(32'h3b02b1d2),
	.w3(32'hbb88b753),
	.w4(32'hbbf18260),
	.w5(32'hbbef2c3a),
	.w6(32'hbb80feb9),
	.w7(32'h386defdb),
	.w8(32'hb9fd0332),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b879484),
	.w1(32'h3b7f5cad),
	.w2(32'h3c3168c2),
	.w3(32'hbbadcc9a),
	.w4(32'h3b40572f),
	.w5(32'h3be9c3fd),
	.w6(32'h3ad645c0),
	.w7(32'h3b9dc6e8),
	.w8(32'h3ae95a5c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8d577),
	.w1(32'h3ab25d34),
	.w2(32'hbb4b8ecb),
	.w3(32'h3b201556),
	.w4(32'h3bb14409),
	.w5(32'h3a506bda),
	.w6(32'h3bf6cbd8),
	.w7(32'h3a7efad7),
	.w8(32'h3b393811),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e422),
	.w1(32'hbb7e09a3),
	.w2(32'hbb971f1e),
	.w3(32'h3ac45d5d),
	.w4(32'hbb4baf7a),
	.w5(32'hbb6de6a5),
	.w6(32'hbb35006e),
	.w7(32'hbb878eb1),
	.w8(32'hbba60acd),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb162b),
	.w1(32'h3c651edd),
	.w2(32'h3c381bba),
	.w3(32'hbbb858fb),
	.w4(32'h3c0fabbe),
	.w5(32'h3c14b475),
	.w6(32'h3bde9e9d),
	.w7(32'h3c01d053),
	.w8(32'hbb88731c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe49a98),
	.w1(32'h3b8ff685),
	.w2(32'h3b4159ce),
	.w3(32'hbb70a5fb),
	.w4(32'h3b42106c),
	.w5(32'h3b0e571e),
	.w6(32'h3b96c6fc),
	.w7(32'h3b4e4a0f),
	.w8(32'h3ac59736),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac38b25),
	.w1(32'hbadd94fa),
	.w2(32'hbc01066a),
	.w3(32'hba385352),
	.w4(32'h3b30fbb6),
	.w5(32'hbb6e5ec2),
	.w6(32'h3b72533e),
	.w7(32'hba69c670),
	.w8(32'h3a5cb5ee),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ee9d2),
	.w1(32'h3bb78562),
	.w2(32'h3c02b6b0),
	.w3(32'h3adfcbe0),
	.w4(32'h39488ba9),
	.w5(32'h3b7e17d6),
	.w6(32'h3b0ae9d0),
	.w7(32'h3bb78fed),
	.w8(32'h3aa592f0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87aa52),
	.w1(32'h3c2cebc0),
	.w2(32'h3b4da623),
	.w3(32'hbabcf9f7),
	.w4(32'h3c18553d),
	.w5(32'h399fa9c1),
	.w6(32'h39bf1e25),
	.w7(32'hbb2cfbe5),
	.w8(32'hbc769839),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fbd1f),
	.w1(32'hbbd8932a),
	.w2(32'hbc241b73),
	.w3(32'hbc5e0e82),
	.w4(32'hbbacd318),
	.w5(32'hbc08bbd5),
	.w6(32'hbb239545),
	.w7(32'hbbd3b8aa),
	.w8(32'hbbe561d0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a565),
	.w1(32'hb98acc52),
	.w2(32'h3adfd616),
	.w3(32'hbc039125),
	.w4(32'hbb7a1a91),
	.w5(32'hb9dc3e85),
	.w6(32'hbb9139b4),
	.w7(32'hba6fedef),
	.w8(32'hbb3eb60f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb549220),
	.w1(32'hbb0d0b31),
	.w2(32'hb9c5e2ee),
	.w3(32'hbb993f7e),
	.w4(32'hbb54dd47),
	.w5(32'hbb332317),
	.w6(32'hbbf9aecb),
	.w7(32'hbb6921e9),
	.w8(32'hbbad7136),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d68e9),
	.w1(32'hba163ef5),
	.w2(32'h3b2d322e),
	.w3(32'hbbaef3bd),
	.w4(32'hbb058e32),
	.w5(32'h3aa5c2f2),
	.w6(32'hbab90843),
	.w7(32'h3b0b0330),
	.w8(32'h3ac25292),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57fcb9),
	.w1(32'hbbab432f),
	.w2(32'hbbdc6307),
	.w3(32'h39ea4cff),
	.w4(32'hbbbabc24),
	.w5(32'hbbdb03b0),
	.w6(32'hbb8a40a6),
	.w7(32'hbbac67a4),
	.w8(32'hbbe0397a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0072a3),
	.w1(32'hbb0a0ee6),
	.w2(32'hba0cee54),
	.w3(32'hbbdec902),
	.w4(32'h3b1c595f),
	.w5(32'h3c9153eb),
	.w6(32'hbb2b69ba),
	.w7(32'hbb6f02df),
	.w8(32'hbb7d36de),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b46e4),
	.w1(32'h3b2a2fab),
	.w2(32'h3b80ddd9),
	.w3(32'h3c8b4b0a),
	.w4(32'h3a35fcc7),
	.w5(32'h3b31ed03),
	.w6(32'hbb0e4146),
	.w7(32'h3ae92f2e),
	.w8(32'hbb216c49),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84b9cc),
	.w1(32'hbba824bc),
	.w2(32'hbb6f12c6),
	.w3(32'h3ab1ac74),
	.w4(32'hbb90c7f6),
	.w5(32'hbb860dd7),
	.w6(32'hbb8e321d),
	.w7(32'hbb9d339e),
	.w8(32'hbbbc2ece),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc236ed1),
	.w1(32'hbb53ecc8),
	.w2(32'hbc10bf3f),
	.w3(32'hbbfcc761),
	.w4(32'hbb97f71e),
	.w5(32'hbbdaff69),
	.w6(32'h3b4d9796),
	.w7(32'hbb3523cd),
	.w8(32'hbb1bdab6),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa166e),
	.w1(32'h3b7b13e9),
	.w2(32'h3c1e738e),
	.w3(32'hbb0134df),
	.w4(32'h39c868fa),
	.w5(32'h3bc72b3f),
	.w6(32'hbab12aca),
	.w7(32'h3b84a0f1),
	.w8(32'hba793da0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7fc9),
	.w1(32'hba773af5),
	.w2(32'hbc013df2),
	.w3(32'h39e9c371),
	.w4(32'h39dde87e),
	.w5(32'hbbaff976),
	.w6(32'h3b3883b0),
	.w7(32'hbb45dd55),
	.w8(32'hbb3d99c2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42217e),
	.w1(32'hbbdfc967),
	.w2(32'hbb1a9941),
	.w3(32'h38bf1005),
	.w4(32'hbc0d2069),
	.w5(32'hbbba6953),
	.w6(32'hbbe9dd81),
	.w7(32'hbbad55e7),
	.w8(32'hbbf5c4b1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf897),
	.w1(32'h3aa512d6),
	.w2(32'h3a39f605),
	.w3(32'hbc105b50),
	.w4(32'hbb151f6c),
	.w5(32'hbb2bd005),
	.w6(32'h3ad173a9),
	.w7(32'h3ace823e),
	.w8(32'hbb0916b8),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265edc),
	.w1(32'hbbcc8f8f),
	.w2(32'hbc38b467),
	.w3(32'hbc06dd58),
	.w4(32'hbbd30b66),
	.w5(32'hbc161144),
	.w6(32'hbbc2572f),
	.w7(32'hbc1a7fd3),
	.w8(32'hbc38956c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e11d9),
	.w1(32'h3bde9822),
	.w2(32'hba652555),
	.w3(32'hbc0b365f),
	.w4(32'h3b27346e),
	.w5(32'hbb919a8d),
	.w6(32'h3c0c26af),
	.w7(32'h3b85d58c),
	.w8(32'hb989fde0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabad227),
	.w1(32'h3b9444b0),
	.w2(32'h3b980003),
	.w3(32'hbb818438),
	.w4(32'h3aa7590e),
	.w5(32'h3aa0e425),
	.w6(32'h3ba3fe07),
	.w7(32'h3ba6c79a),
	.w8(32'h3adfbc06),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9bcd9),
	.w1(32'hbbff5770),
	.w2(32'h3ba530d3),
	.w3(32'h3b732f49),
	.w4(32'hbb93f9fb),
	.w5(32'h3c2d1c64),
	.w6(32'hbc17a40f),
	.w7(32'hbb5a0707),
	.w8(32'h3b3e23fb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3227b9),
	.w1(32'h3b413778),
	.w2(32'h3bce6822),
	.w3(32'h3c4b1559),
	.w4(32'hb7d9d4f5),
	.w5(32'h3b5948cd),
	.w6(32'h3a62d26c),
	.w7(32'h3bab9598),
	.w8(32'h3b465f07),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2aeed),
	.w1(32'hba3a2454),
	.w2(32'hbb04be1e),
	.w3(32'h3aa2b577),
	.w4(32'hbad4f997),
	.w5(32'hbb25f0e6),
	.w6(32'hbaf2ea8f),
	.w7(32'hbb5dc13b),
	.w8(32'hbb2bbc23),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1635ed),
	.w1(32'h3af78d86),
	.w2(32'h399adc75),
	.w3(32'hbac42ab3),
	.w4(32'h39975438),
	.w5(32'h3b252520),
	.w6(32'hbb0ad4d6),
	.w7(32'h3b7ee984),
	.w8(32'hbb2d8c86),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babaec7),
	.w1(32'h3ad242a5),
	.w2(32'h3b5d2c0c),
	.w3(32'h39feb2f6),
	.w4(32'hbb18848f),
	.w5(32'hba321214),
	.w6(32'hbb901ef5),
	.w7(32'hbb19bd87),
	.w8(32'hbb4b1926),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083547),
	.w1(32'h3bf826a2),
	.w2(32'h3b4c6da4),
	.w3(32'h3b7d5c71),
	.w4(32'h3c02a980),
	.w5(32'h3a9fefb0),
	.w6(32'h3c1efeb8),
	.w7(32'h3b8910f7),
	.w8(32'h3ba2eff9),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81824a2),
	.w1(32'hbab3f6b6),
	.w2(32'h3b2ab8d5),
	.w3(32'h3a9a7fa9),
	.w4(32'hbadee1a2),
	.w5(32'h3b10632f),
	.w6(32'hba83b619),
	.w7(32'hba0609aa),
	.w8(32'hbb242ffd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf6626),
	.w1(32'hbba15775),
	.w2(32'hbc29312b),
	.w3(32'hbb936ef4),
	.w4(32'hbb0e599a),
	.w5(32'hbbb83a38),
	.w6(32'hb9b9a284),
	.w7(32'hbb90d58f),
	.w8(32'h3b0e1c01),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb630055),
	.w1(32'hbb8a3fd8),
	.w2(32'hbb5272e0),
	.w3(32'h39a4631a),
	.w4(32'hba89c896),
	.w5(32'hb9bba407),
	.w6(32'hbb030519),
	.w7(32'hbb185d9e),
	.w8(32'hbb2ccb30),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80957b),
	.w1(32'hbb25a56c),
	.w2(32'h3c15c5a1),
	.w3(32'hb9fd3a76),
	.w4(32'hbb978656),
	.w5(32'h3c0a0c4c),
	.w6(32'hbba51b09),
	.w7(32'h3b05fe8e),
	.w8(32'hba2cbe0a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b979c83),
	.w1(32'h3b83d3be),
	.w2(32'h3a543de1),
	.w3(32'h3b9a2fe0),
	.w4(32'h3b9653a6),
	.w5(32'h39fac67a),
	.w6(32'h3b65f862),
	.w7(32'h3a0aed8f),
	.w8(32'hba490f5d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219c29),
	.w1(32'h3ac0c577),
	.w2(32'h3b865221),
	.w3(32'hb9a3285b),
	.w4(32'h3b5b361a),
	.w5(32'h3bd73eb0),
	.w6(32'h3b695e30),
	.w7(32'h3b11cbb4),
	.w8(32'hbab7615a),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1faae2),
	.w1(32'hbba185e6),
	.w2(32'hbb4b38b2),
	.w3(32'h3b20dc48),
	.w4(32'hbbb79355),
	.w5(32'hbb9b8382),
	.w6(32'hbb924af1),
	.w7(32'hbbcdb265),
	.w8(32'hbbe4c7ed),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde6396),
	.w1(32'h3bc93faf),
	.w2(32'h3c1628c5),
	.w3(32'hbbf67212),
	.w4(32'hba8458bb),
	.w5(32'h3b88be30),
	.w6(32'hba4447b8),
	.w7(32'h3b835003),
	.w8(32'hbb2e5997),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ead91),
	.w1(32'h3bf694f5),
	.w2(32'h3bf8da6f),
	.w3(32'hbad44433),
	.w4(32'h3b96d489),
	.w5(32'h3bfdf432),
	.w6(32'h39a5de31),
	.w7(32'h3bb6be91),
	.w8(32'hbb6645ba),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b3911),
	.w1(32'h3ca76d22),
	.w2(32'h3c89fab0),
	.w3(32'hbb005903),
	.w4(32'h3bbc747e),
	.w5(32'h3a96c2a2),
	.w6(32'h3c93d11c),
	.w7(32'h3ca16a4f),
	.w8(32'h3c2d9fca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9beaa0b),
	.w1(32'h3bb05566),
	.w2(32'h3c21cbc7),
	.w3(32'hbc407ae8),
	.w4(32'h3b1f5ae6),
	.w5(32'h3bd83fa9),
	.w6(32'hbbebc1cd),
	.w7(32'hba1eff45),
	.w8(32'hbbc1f4f5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be60503),
	.w1(32'hba7d48cb),
	.w2(32'h3b4f498d),
	.w3(32'h3b03421e),
	.w4(32'hbb600490),
	.w5(32'h3af2735c),
	.w6(32'hbbc8989e),
	.w7(32'hbabdfcc0),
	.w8(32'hbb77c856),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988d78b),
	.w1(32'h3af5fb9b),
	.w2(32'h3b6cba92),
	.w3(32'hbaae390d),
	.w4(32'h38c01f3f),
	.w5(32'h3b19f6f7),
	.w6(32'hbb2c8d1b),
	.w7(32'h39fefd49),
	.w8(32'hbae8b072),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b387720),
	.w1(32'hb9425d0b),
	.w2(32'h3a67a32b),
	.w3(32'h3a33c0b2),
	.w4(32'hbb274676),
	.w5(32'h3937c74a),
	.w6(32'hbb203e9a),
	.w7(32'hbad86f85),
	.w8(32'hbb968205),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bac3f),
	.w1(32'hbbc39629),
	.w2(32'hbb7ca915),
	.w3(32'h390b9b18),
	.w4(32'hbb8b0cd4),
	.w5(32'hbb40944c),
	.w6(32'hbb9bc03b),
	.w7(32'hbb8ca9ab),
	.w8(32'hbb8dc40d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe79dd6),
	.w1(32'h3b90cfb9),
	.w2(32'h3c1dacdf),
	.w3(32'hbbb57023),
	.w4(32'h39c798b4),
	.w5(32'h3b7f24a8),
	.w6(32'h3a9aebc5),
	.w7(32'h3bc4e23d),
	.w8(32'h3b88d235),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cfb00),
	.w1(32'h3b59eb20),
	.w2(32'h3bab51fc),
	.w3(32'h3b997b0d),
	.w4(32'h3aaa0488),
	.w5(32'h3b6ad5fc),
	.w6(32'hbae03052),
	.w7(32'h3ae052dd),
	.w8(32'hba6d09f4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e00aa),
	.w1(32'hbc32b144),
	.w2(32'hba6bdc85),
	.w3(32'h3a7cb9d8),
	.w4(32'hbc278862),
	.w5(32'hbb92f1c5),
	.w6(32'hbbfc79e5),
	.w7(32'hbb61965d),
	.w8(32'h3b87acff),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ae22a),
	.w1(32'h380f29c7),
	.w2(32'hba410404),
	.w3(32'hbb06c546),
	.w4(32'h38dfd4dc),
	.w5(32'h3ab3f2da),
	.w6(32'hbaf55521),
	.w7(32'hb927652f),
	.w8(32'hbba30dbd),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39dab),
	.w1(32'hbbbed3d8),
	.w2(32'hb91e0c9f),
	.w3(32'h39e256dc),
	.w4(32'hbbccb94d),
	.w5(32'hbb6eaa56),
	.w6(32'h39b73ee0),
	.w7(32'h3b4739d5),
	.w8(32'h3be0ad1a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadc896),
	.w1(32'h3a8320c6),
	.w2(32'h3b23adc6),
	.w3(32'h3c279789),
	.w4(32'hbb608344),
	.w5(32'hba0c8d9f),
	.w6(32'hbb62ca18),
	.w7(32'hb9a48da0),
	.w8(32'hbbed9748),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba769bbb),
	.w1(32'hbc2d6e67),
	.w2(32'hbc3cd4c0),
	.w3(32'hbb6e0f28),
	.w4(32'hbc2146b4),
	.w5(32'hbc388921),
	.w6(32'hbc27da42),
	.w7(32'hbc4f6210),
	.w8(32'hbc7523f4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fcaad),
	.w1(32'hbbadd9dd),
	.w2(32'h3c495e60),
	.w3(32'hbc182269),
	.w4(32'hbc261b45),
	.w5(32'h3ac9dd4a),
	.w6(32'hbc0f86e6),
	.w7(32'h3ad5a553),
	.w8(32'h3b2ba645),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81bf36),
	.w1(32'h3b7c68a7),
	.w2(32'h3bd70bd1),
	.w3(32'h3b94e826),
	.w4(32'h3ab1c0d3),
	.w5(32'h3b98f212),
	.w6(32'hbb55cdad),
	.w7(32'h3ac33d94),
	.w8(32'hbb1125e5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89b7e8),
	.w1(32'hbaaea3f0),
	.w2(32'h3ab1daa1),
	.w3(32'h3a8bdf6f),
	.w4(32'hbbae6c49),
	.w5(32'hbb034b96),
	.w6(32'hbb90842f),
	.w7(32'hb9b9f844),
	.w8(32'hbb467dad),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99516ad),
	.w1(32'hba9d5892),
	.w2(32'h3b20d8de),
	.w3(32'hbb7a51b2),
	.w4(32'hbba0c524),
	.w5(32'hb9a8f3ca),
	.w6(32'hbba4067a),
	.w7(32'hb8d4d7c5),
	.w8(32'hbb77ae69),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71b3c9),
	.w1(32'h3b91ea66),
	.w2(32'h3c898adf),
	.w3(32'hbb566f8a),
	.w4(32'hbbdb1566),
	.w5(32'hbba70f12),
	.w6(32'hb86854d0),
	.w7(32'h3c1bb130),
	.w8(32'h3c391879),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a9a18),
	.w1(32'h398953e6),
	.w2(32'hbb7e1d66),
	.w3(32'hbb2acd78),
	.w4(32'hba136430),
	.w5(32'hbb61cbce),
	.w6(32'h3b203300),
	.w7(32'hbb15afd3),
	.w8(32'hbb57ae41),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2c3ac),
	.w1(32'hba8e3d43),
	.w2(32'h3c1f9e02),
	.w3(32'h38589fcb),
	.w4(32'hbb5cdfb5),
	.w5(32'h3beee4b4),
	.w6(32'hbbbc8782),
	.w7(32'h3b42cded),
	.w8(32'hb8c852a9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bfac4),
	.w1(32'h3b4fb612),
	.w2(32'h3bfe26b7),
	.w3(32'h3a866532),
	.w4(32'h39714c9e),
	.w5(32'h3b91c36c),
	.w6(32'hbb9081a7),
	.w7(32'h3a865d94),
	.w8(32'hbc0e411b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40064e),
	.w1(32'hbb836afd),
	.w2(32'hbaf4c04f),
	.w3(32'hbb8e59ef),
	.w4(32'hbbd00800),
	.w5(32'hbb85ca92),
	.w6(32'hbc01f986),
	.w7(32'hbb9a8620),
	.w8(32'hbc0034bf),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb647ee5),
	.w1(32'h3b98cce9),
	.w2(32'h3c039f68),
	.w3(32'hbbde251c),
	.w4(32'hbb9b2974),
	.w5(32'hbb3e95e8),
	.w6(32'h3c16a593),
	.w7(32'h3c77ffae),
	.w8(32'h3c41c08f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5342),
	.w1(32'h3bab7c38),
	.w2(32'h3cb0108d),
	.w3(32'hbba7350e),
	.w4(32'h3a307824),
	.w5(32'h3c790f93),
	.w6(32'hbabf39b1),
	.w7(32'h3c264096),
	.w8(32'h3b170690),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c472936),
	.w1(32'h3bcdfe41),
	.w2(32'h3c351a4c),
	.w3(32'h3c5548f7),
	.w4(32'h3b989469),
	.w5(32'h3bc88f7e),
	.w6(32'h3af5ffe6),
	.w7(32'h3bd9ccb1),
	.w8(32'h3b46d1f1),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bea30),
	.w1(32'hb8ac680c),
	.w2(32'h364bf987),
	.w3(32'h39a2edb0),
	.w4(32'hb8721530),
	.w5(32'h3895555e),
	.w6(32'hb8125fb6),
	.w7(32'hb8f7f249),
	.w8(32'hb886b24e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c690b2),
	.w1(32'hba36d1d3),
	.w2(32'hbb1f96d7),
	.w3(32'hbae792b8),
	.w4(32'h395ccf34),
	.w5(32'h38964586),
	.w6(32'h3ab12a7b),
	.w7(32'h3a7abbc2),
	.w8(32'hb9c3a7f8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule