module layer_10_featuremap_112(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93ae0e),
	.w1(32'h39f66408),
	.w2(32'h3a64ed2a),
	.w3(32'hba20a192),
	.w4(32'h390158d4),
	.w5(32'h3a6db790),
	.w6(32'hbacad5ce),
	.w7(32'hba78712e),
	.w8(32'hbb38d39c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f1c123),
	.w1(32'hbac5895b),
	.w2(32'hbafeafaa),
	.w3(32'hbb51281d),
	.w4(32'hbb0467be),
	.w5(32'hbb1e0f69),
	.w6(32'hba94599a),
	.w7(32'hba9b3500),
	.w8(32'hbad93a10),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c3c6),
	.w1(32'hbae11850),
	.w2(32'hbb6f6dc6),
	.w3(32'hbb1b6295),
	.w4(32'hba2ee3bd),
	.w5(32'hba8b0717),
	.w6(32'h3a2ce4d5),
	.w7(32'hb967d4e4),
	.w8(32'hb9a6749f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c68df),
	.w1(32'hbb5c10a8),
	.w2(32'hbb7c1b44),
	.w3(32'h39251972),
	.w4(32'h3ab43b24),
	.w5(32'hbad11a1f),
	.w6(32'hbb3306de),
	.w7(32'hbb3d95b3),
	.w8(32'hbb0641c4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6906f),
	.w1(32'h3b0d50ba),
	.w2(32'h3a1f368b),
	.w3(32'h3b0fc4f6),
	.w4(32'h3a129530),
	.w5(32'h38e820d8),
	.w6(32'h3a962ae5),
	.w7(32'h3a04ce8e),
	.w8(32'hb964ffff),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa73812),
	.w1(32'hb995c87f),
	.w2(32'hba4953b9),
	.w3(32'h3a437711),
	.w4(32'hb9fb1dc5),
	.w5(32'hbaa60049),
	.w6(32'h3a2e59af),
	.w7(32'hb6e976c9),
	.w8(32'hba0f5228),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec50b8),
	.w1(32'hbb268ca8),
	.w2(32'hbb641d06),
	.w3(32'hbaa9c682),
	.w4(32'hbb019f1e),
	.w5(32'hbb2a5078),
	.w6(32'hbb13b95e),
	.w7(32'hbb5ee1b7),
	.w8(32'hbadb52b2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7002),
	.w1(32'h39d16e02),
	.w2(32'h38315246),
	.w3(32'hbadb9403),
	.w4(32'h39f49a5f),
	.w5(32'h3a1d76fa),
	.w6(32'h39cf0f3e),
	.w7(32'h39a1014d),
	.w8(32'h390981a9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9745f11),
	.w1(32'hba63af0a),
	.w2(32'hbac0f9ec),
	.w3(32'h39983287),
	.w4(32'hba230465),
	.w5(32'hba4f0706),
	.w6(32'hba3ba6b7),
	.w7(32'hba9578b0),
	.w8(32'hb98e582b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e54787),
	.w1(32'hba7ec06b),
	.w2(32'hbacb113c),
	.w3(32'hba29a05b),
	.w4(32'hbb0e69d7),
	.w5(32'hbb427c02),
	.w6(32'hbaf745f3),
	.w7(32'hba5741de),
	.w8(32'hbafb6df0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4422e1),
	.w1(32'hbb2141d3),
	.w2(32'hbb8d94c2),
	.w3(32'hbb3e7518),
	.w4(32'hb9a3b863),
	.w5(32'hbaae2280),
	.w6(32'h39d37dcc),
	.w7(32'hba3ec05f),
	.w8(32'hbb648060),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed889),
	.w1(32'h3b4229cc),
	.w2(32'h3b117ba3),
	.w3(32'hbadbb67e),
	.w4(32'h3acafead),
	.w5(32'h3aa701e3),
	.w6(32'hba16d61d),
	.w7(32'h386f529f),
	.w8(32'hbadfd94c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4a138),
	.w1(32'hb9d3f2ad),
	.w2(32'hbacd17c1),
	.w3(32'h39d4724a),
	.w4(32'hba6dd23a),
	.w5(32'hbad38cac),
	.w6(32'h38f9693b),
	.w7(32'h38d6d409),
	.w8(32'h380c5e95),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b73a67),
	.w1(32'hb9b613b9),
	.w2(32'hba6eb725),
	.w3(32'hba8726e1),
	.w4(32'hba3c8201),
	.w5(32'hba3783fd),
	.w6(32'hb8403de5),
	.w7(32'hb9ab65d5),
	.w8(32'hba3a36c6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b93f),
	.w1(32'h3b84249e),
	.w2(32'h3b5cfcb3),
	.w3(32'hba5bf587),
	.w4(32'h3ad40645),
	.w5(32'h3a99d6f6),
	.w6(32'hbb077fbc),
	.w7(32'hbafdd374),
	.w8(32'hbb809e4e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a119f29),
	.w1(32'hba816499),
	.w2(32'hba8889c2),
	.w3(32'hba023147),
	.w4(32'hba82be44),
	.w5(32'hba9222b9),
	.w6(32'hba3f2f97),
	.w7(32'hba20fce7),
	.w8(32'hb9d9a33f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9942cf5),
	.w1(32'hbb060c6a),
	.w2(32'hbb94a600),
	.w3(32'hba4ad9c6),
	.w4(32'hbac2aca8),
	.w5(32'hbb6644c1),
	.w6(32'h3825a78f),
	.w7(32'hbb2d1622),
	.w8(32'hbabfc8da),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb020861),
	.w1(32'hbb12cc24),
	.w2(32'hbb7b6fee),
	.w3(32'hbb0605f3),
	.w4(32'hbb189bf1),
	.w5(32'hbb4dc56f),
	.w6(32'hbb014d73),
	.w7(32'hbb3e115e),
	.w8(32'hbaf12679),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567d27),
	.w1(32'hba26c112),
	.w2(32'hbb0d2802),
	.w3(32'hbb3d4fcd),
	.w4(32'hba65eea3),
	.w5(32'hba75a88d),
	.w6(32'hba92e9cb),
	.w7(32'hbae69633),
	.w8(32'hba19ff0b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c77f9),
	.w1(32'hb9ab509c),
	.w2(32'hbac8b1ea),
	.w3(32'hba1ebee4),
	.w4(32'hb9f36288),
	.w5(32'hba8e7387),
	.w6(32'hb9487d13),
	.w7(32'hba5f27fc),
	.w8(32'hba1fc8a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0071ad),
	.w1(32'hbb1bbfdb),
	.w2(32'hba880087),
	.w3(32'hba7d049c),
	.w4(32'hba3a886a),
	.w5(32'hb9cc2d9a),
	.w6(32'hbb03f2fc),
	.w7(32'hba905f05),
	.w8(32'h3a4b6e33),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e2535),
	.w1(32'hbb537d48),
	.w2(32'hbbca531e),
	.w3(32'h3a949578),
	.w4(32'hba0d0d68),
	.w5(32'h39e45764),
	.w6(32'hb93dce07),
	.w7(32'hbb5f29a9),
	.w8(32'hbb779160),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676fd4),
	.w1(32'hbb815e13),
	.w2(32'hbbebc543),
	.w3(32'hbb1123bc),
	.w4(32'hb9e222eb),
	.w5(32'hbbafb7a7),
	.w6(32'hbafbeab3),
	.w7(32'hbbc67bf6),
	.w8(32'hbaa32dfc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7881),
	.w1(32'hb9a82048),
	.w2(32'hba30ebf0),
	.w3(32'hb9b5a16c),
	.w4(32'h382d7778),
	.w5(32'hb9328775),
	.w6(32'h386aba88),
	.w7(32'hb7a41fb0),
	.w8(32'hb76b5c9a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d0a75),
	.w1(32'hba8a6b11),
	.w2(32'hbaf7b09d),
	.w3(32'h3a066ec8),
	.w4(32'hbac5baac),
	.w5(32'hbb60c75f),
	.w6(32'hb99acc1a),
	.w7(32'hba1be57d),
	.w8(32'hbac33986),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb431f2c),
	.w1(32'hbb80258e),
	.w2(32'hbbb56a8b),
	.w3(32'hbb478363),
	.w4(32'hbaa525c0),
	.w5(32'hbafc4ca8),
	.w6(32'hbaeac5ff),
	.w7(32'hbb037f5e),
	.w8(32'hbb1cf2ef),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2896),
	.w1(32'hba7bf245),
	.w2(32'hbabc766d),
	.w3(32'hbb2829a1),
	.w4(32'hba2d9a7a),
	.w5(32'hba808724),
	.w6(32'hba51894d),
	.w7(32'hba5ecba9),
	.w8(32'hba55f3e6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a3456),
	.w1(32'h3959f40f),
	.w2(32'hbac49a29),
	.w3(32'hba4d69b1),
	.w4(32'hba62accf),
	.w5(32'hbb1d4fff),
	.w6(32'h3ace2aa0),
	.w7(32'h3a239cee),
	.w8(32'hb9aec771),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f5aeb),
	.w1(32'h3b0a6f68),
	.w2(32'hbba8b3ba),
	.w3(32'hba711f56),
	.w4(32'h3b283af3),
	.w5(32'hbb9adb2d),
	.w6(32'h3b881051),
	.w7(32'hbb24c0f9),
	.w8(32'hba585029),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93c837),
	.w1(32'hbb3891d7),
	.w2(32'hbb9b193a),
	.w3(32'hbb3034b4),
	.w4(32'hbaa5f5c3),
	.w5(32'hbb72a669),
	.w6(32'hbb15083e),
	.w7(32'hbb65e5b5),
	.w8(32'hba926196),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67742b),
	.w1(32'hba90b3f3),
	.w2(32'hba2a3e8e),
	.w3(32'hbb405547),
	.w4(32'hba8cda91),
	.w5(32'hba288d94),
	.w6(32'hba800ca6),
	.w7(32'hb9e6631e),
	.w8(32'h39c2ae9d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37747de9),
	.w1(32'hba792de5),
	.w2(32'hbaaa53c7),
	.w3(32'h3933d4a0),
	.w4(32'hba1df585),
	.w5(32'hba30fa01),
	.w6(32'hba0dc532),
	.w7(32'hb9732838),
	.w8(32'h39173a59),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ea368a),
	.w1(32'h39dfca7b),
	.w2(32'hbb1e91d3),
	.w3(32'h385244c6),
	.w4(32'hb9960266),
	.w5(32'hba0fe26c),
	.w6(32'h3a06a49e),
	.w7(32'hbab685ed),
	.w8(32'hbac272ab),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a247c),
	.w1(32'hbb480206),
	.w2(32'hbb332257),
	.w3(32'hbb11dfda),
	.w4(32'hbad4bfde),
	.w5(32'hbac675f7),
	.w6(32'hbb3908c4),
	.w7(32'h39c87b63),
	.w8(32'h3b3c80c2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d60c5),
	.w1(32'h3a187101),
	.w2(32'h3a09b005),
	.w3(32'hbb099ee5),
	.w4(32'hbaaad4e1),
	.w5(32'hbabde766),
	.w6(32'hb982c8dd),
	.w7(32'h3977a353),
	.w8(32'h396ef39c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba699a1f),
	.w1(32'hba12f8e2),
	.w2(32'hbaa3b913),
	.w3(32'hbb114e1e),
	.w4(32'hba1550c2),
	.w5(32'hba2364fa),
	.w6(32'hb9831a75),
	.w7(32'hba42268f),
	.w8(32'hb9fd5491),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89fd24),
	.w1(32'hba998075),
	.w2(32'hbb0f16db),
	.w3(32'hb92509be),
	.w4(32'hbb1f20ce),
	.w5(32'hbb391e9b),
	.w6(32'hba79c876),
	.w7(32'h3898c74b),
	.w8(32'hb9a63198),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb0226),
	.w1(32'hbb40f132),
	.w2(32'hbb8d3e75),
	.w3(32'hbb22e8d8),
	.w4(32'hbb241fd7),
	.w5(32'hbb69e0d5),
	.w6(32'hbb04f281),
	.w7(32'hbb206428),
	.w8(32'hbae3024d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05a1b5),
	.w1(32'hba6a8540),
	.w2(32'hbb0550ee),
	.w3(32'hbaf68b70),
	.w4(32'hba7c4a55),
	.w5(32'hbae1ce13),
	.w6(32'hb80708ab),
	.w7(32'hbaa7f8c1),
	.w8(32'hbabc712e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a796),
	.w1(32'hbac39477),
	.w2(32'hba9bb9c8),
	.w3(32'hba2f3e95),
	.w4(32'hbad8cef2),
	.w5(32'hbacb91df),
	.w6(32'hbac36086),
	.w7(32'hba315afe),
	.w8(32'hb95f4e2e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ede0b9),
	.w1(32'hbb491ad9),
	.w2(32'hbbaec3f7),
	.w3(32'hbac5a405),
	.w4(32'hbac23dd4),
	.w5(32'hbba0980b),
	.w6(32'hbb2564e4),
	.w7(32'hbba567b7),
	.w8(32'hbb029cd7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b007d),
	.w1(32'hb980a873),
	.w2(32'hba9ab54a),
	.w3(32'hbb43642c),
	.w4(32'hba2daef6),
	.w5(32'hba472887),
	.w6(32'h3996ca63),
	.w7(32'h395470c0),
	.w8(32'hba128b47),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8645),
	.w1(32'hbaee6000),
	.w2(32'hbb14a2e0),
	.w3(32'hbac21ae7),
	.w4(32'hbabede68),
	.w5(32'hbb09e787),
	.w6(32'hba1793e4),
	.w7(32'hba0d34cf),
	.w8(32'h39029408),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba496658),
	.w1(32'hbb3738be),
	.w2(32'hbaa6aa19),
	.w3(32'hba3608ee),
	.w4(32'hbb20b1ae),
	.w5(32'hbad0135c),
	.w6(32'hbaf6f844),
	.w7(32'hba6b04be),
	.w8(32'hbaacfdbe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e193),
	.w1(32'hbae5c704),
	.w2(32'h35098f45),
	.w3(32'hbb839a11),
	.w4(32'hbb138e40),
	.w5(32'hb982651c),
	.w6(32'hbad04790),
	.w7(32'hb90cb8fb),
	.w8(32'h3a90c19f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f2242),
	.w1(32'hba54fa7d),
	.w2(32'hbb3f1d4c),
	.w3(32'hb995ca82),
	.w4(32'hbabf6f4f),
	.w5(32'hbae02022),
	.w6(32'hba3777cd),
	.w7(32'hbaf82cc9),
	.w8(32'hbac126b5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb219dde),
	.w1(32'h3b193238),
	.w2(32'h3b5f95f4),
	.w3(32'hbb34f4f5),
	.w4(32'h3a00482c),
	.w5(32'h3af335cd),
	.w6(32'hbadde3d0),
	.w7(32'hbab4359a),
	.w8(32'hbb1cc8ea),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087220),
	.w1(32'hbb090eeb),
	.w2(32'hbba61d4a),
	.w3(32'h3a8a0516),
	.w4(32'hbabc9f49),
	.w5(32'hbb8ef01c),
	.w6(32'hb9f29acd),
	.w7(32'hbb4dc568),
	.w8(32'hbb0ccfb1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb992646),
	.w1(32'hbab24c4f),
	.w2(32'hbb256499),
	.w3(32'hbb26bf71),
	.w4(32'hba6891e2),
	.w5(32'hbacffd2b),
	.w6(32'hb9d69970),
	.w7(32'hba2a14d8),
	.w8(32'hb90dbd49),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba668710),
	.w1(32'hb945c799),
	.w2(32'hb9ac29ee),
	.w3(32'hba61bb06),
	.w4(32'hb746551b),
	.w5(32'hb9f27e0b),
	.w6(32'h36bab64d),
	.w7(32'hb92555b3),
	.w8(32'hba4ace01),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9968367),
	.w1(32'hbaf1454d),
	.w2(32'hbb33af1c),
	.w3(32'h383be030),
	.w4(32'hba7475ae),
	.w5(32'hbaf97c2e),
	.w6(32'hba2d92e1),
	.w7(32'hbabcb725),
	.w8(32'hbad6f39d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59fb5),
	.w1(32'hba30a188),
	.w2(32'hbb0b5a24),
	.w3(32'hba997ed6),
	.w4(32'hba884bb7),
	.w5(32'hbb2a63c8),
	.w6(32'hbaef9253),
	.w7(32'hbb259823),
	.w8(32'hbb800678),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11375b),
	.w1(32'hbb4f46f7),
	.w2(32'hbb418f22),
	.w3(32'hbb0c3c3d),
	.w4(32'hbb234d2d),
	.w5(32'hbb287845),
	.w6(32'hbacdb691),
	.w7(32'hba205aec),
	.w8(32'hbab68c60),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48fd25),
	.w1(32'hbb449a6d),
	.w2(32'hbb1c17cf),
	.w3(32'hbb2c11f7),
	.w4(32'hbb915063),
	.w5(32'hbb3f13d9),
	.w6(32'hbb66cb55),
	.w7(32'hbb4c13ca),
	.w8(32'hbb0fb82e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27cd85),
	.w1(32'hbabaad66),
	.w2(32'hbab44a57),
	.w3(32'hb9bf3638),
	.w4(32'hbabe6d7d),
	.w5(32'hbad4f2db),
	.w6(32'h360708b8),
	.w7(32'h38a156c8),
	.w8(32'h3a4074d5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981fece),
	.w1(32'hbb08d6d9),
	.w2(32'hbbd45c52),
	.w3(32'hba2363db),
	.w4(32'hbb22c098),
	.w5(32'hbb951c31),
	.w6(32'hbb1231b0),
	.w7(32'hbb861db8),
	.w8(32'hbb397010),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7052bf),
	.w1(32'hbb372860),
	.w2(32'hbb650dc0),
	.w3(32'hbb2664aa),
	.w4(32'hbaff1a47),
	.w5(32'hbb20fa2a),
	.w6(32'hba986f0b),
	.w7(32'hbafd59ff),
	.w8(32'hbb10cdac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c384e),
	.w1(32'h3a346cb0),
	.w2(32'hba8d4ba4),
	.w3(32'hbb3a9de8),
	.w4(32'h3a76ca76),
	.w5(32'hba27729d),
	.w6(32'h39f57fa3),
	.w7(32'hb8a278cb),
	.w8(32'h3a220a50),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19633a),
	.w1(32'hbac0b620),
	.w2(32'hbac88f27),
	.w3(32'h3a9ab66c),
	.w4(32'hba92ea31),
	.w5(32'hba62621d),
	.w6(32'hbaa79496),
	.w7(32'hbacd9d71),
	.w8(32'hba0aa39f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b09c8),
	.w1(32'hba0847a4),
	.w2(32'hbaa36792),
	.w3(32'hb98658dc),
	.w4(32'hb9bfcca7),
	.w5(32'hba4d1b7c),
	.w6(32'h3916cf73),
	.w7(32'hb9f4db70),
	.w8(32'hb9c575c7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63701d),
	.w1(32'hba313bcd),
	.w2(32'hba572675),
	.w3(32'hb9c272f6),
	.w4(32'hbaab0a04),
	.w5(32'hb9ab3b40),
	.w6(32'hb950e3a5),
	.w7(32'h380a2e9c),
	.w8(32'hb9a2f407),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dabe9),
	.w1(32'hba314a19),
	.w2(32'hba4840d2),
	.w3(32'h3967cc7a),
	.w4(32'hb9d0a219),
	.w5(32'hb9b62ea4),
	.w6(32'h3911d54a),
	.w7(32'hb9bbbe56),
	.w8(32'hb92c4cb0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dada74),
	.w1(32'h39ba6b17),
	.w2(32'hbaf6392b),
	.w3(32'h38fac890),
	.w4(32'h39185eca),
	.w5(32'h39bce2fb),
	.w6(32'hb9746443),
	.w7(32'h39f834eb),
	.w8(32'h3b072611),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916db67),
	.w1(32'hbab6b3e4),
	.w2(32'hba3d5be6),
	.w3(32'h399a3f28),
	.w4(32'hbb08cff2),
	.w5(32'hbb0f5af0),
	.w6(32'hbace02fe),
	.w7(32'hba83dfc8),
	.w8(32'hbac6f77b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cfc91),
	.w1(32'h3ac31e40),
	.w2(32'hba5a7b90),
	.w3(32'hbb1b86ea),
	.w4(32'h3aaa6f90),
	.w5(32'hba45727f),
	.w6(32'h3aa8bb8f),
	.w7(32'hba99c98a),
	.w8(32'hbb131ac2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a0885),
	.w1(32'hba0a0b37),
	.w2(32'hbb818f74),
	.w3(32'hba985d66),
	.w4(32'h398fad80),
	.w5(32'hba3e177d),
	.w6(32'h3a1ca879),
	.w7(32'hbaac03ea),
	.w8(32'h3901fe4b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13fe60),
	.w1(32'hbac0ddba),
	.w2(32'hbb8d8fd2),
	.w3(32'h39f8d47c),
	.w4(32'hba6cbaf2),
	.w5(32'hbb20077d),
	.w6(32'hbada987a),
	.w7(32'hbb14d2d4),
	.w8(32'hba454b5a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fcfaf),
	.w1(32'hbba2ac89),
	.w2(32'hbbd6c09c),
	.w3(32'hbb28fc6c),
	.w4(32'hb9eeaec5),
	.w5(32'hbba2c080),
	.w6(32'hbb0a6368),
	.w7(32'hbbc3f395),
	.w8(32'hba4e04dd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab745f),
	.w1(32'hba201445),
	.w2(32'hba98838a),
	.w3(32'hba247caf),
	.w4(32'hb97cf936),
	.w5(32'hba65b9b1),
	.w6(32'hb98adfbc),
	.w7(32'hba445912),
	.w8(32'hba5cc8ed),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd2c5b),
	.w1(32'h3998e8bb),
	.w2(32'hbb4d6666),
	.w3(32'hbab60304),
	.w4(32'h37174e7b),
	.w5(32'hbb2cf7e1),
	.w6(32'hb94fdbdf),
	.w7(32'hbb01ea1b),
	.w8(32'hbb084256),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bbf84),
	.w1(32'hbb04619d),
	.w2(32'hbb3c7f99),
	.w3(32'hba4f988c),
	.w4(32'hbafe9fdf),
	.w5(32'hbb056c5b),
	.w6(32'hbb039996),
	.w7(32'hbb1ff2a1),
	.w8(32'hbaa24558),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b000b),
	.w1(32'hb9445a21),
	.w2(32'hbabc4526),
	.w3(32'hbad84504),
	.w4(32'hba063e4a),
	.w5(32'hba1b3440),
	.w6(32'h38b8be9e),
	.w7(32'hba5b8c1b),
	.w8(32'hba2d24bd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43657b),
	.w1(32'hba77091f),
	.w2(32'hbadd3607),
	.w3(32'hb95238e7),
	.w4(32'hba33e5c9),
	.w5(32'hba7e9dc8),
	.w6(32'hb9d37b34),
	.w7(32'hba7ccd9c),
	.w8(32'hba529b28),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e4a6),
	.w1(32'hbaadb30f),
	.w2(32'hbab1e5ae),
	.w3(32'hba0b12ff),
	.w4(32'hba82f410),
	.w5(32'hbaa198cf),
	.w6(32'hba297dd3),
	.w7(32'hb95f72dc),
	.w8(32'h3987a29b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4272e5),
	.w1(32'h390f3389),
	.w2(32'hb91125d1),
	.w3(32'hb90c27a8),
	.w4(32'hba0d7330),
	.w5(32'hba1c5315),
	.w6(32'hb93df395),
	.w7(32'hba28a158),
	.w8(32'hbaccfdcc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadccb12),
	.w1(32'h39a9dc23),
	.w2(32'hba44b4a0),
	.w3(32'hbabdb4bc),
	.w4(32'h39289a43),
	.w5(32'h389d0914),
	.w6(32'hbb030919),
	.w7(32'hbadbdae0),
	.w8(32'hbb96ff0e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5828a6),
	.w1(32'h395d822b),
	.w2(32'hba2936dd),
	.w3(32'hba695aa7),
	.w4(32'h3a0a522a),
	.w5(32'hb9ec561c),
	.w6(32'h3a81d25e),
	.w7(32'h38e77f87),
	.w8(32'h38f1ce9a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba692afa),
	.w1(32'h3a4fc654),
	.w2(32'hba811e36),
	.w3(32'h39c55ede),
	.w4(32'h3a3a636d),
	.w5(32'h39f190e5),
	.w6(32'h3a838471),
	.w7(32'h39cf8372),
	.w8(32'h3a4ef1ff),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c07ad),
	.w1(32'hbb2a39ce),
	.w2(32'hbb3bb663),
	.w3(32'h396def73),
	.w4(32'hba534934),
	.w5(32'hbb18eeaa),
	.w6(32'h3a6e52ba),
	.w7(32'h392c7151),
	.w8(32'h39dd0491),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98abbb3),
	.w1(32'hbab02160),
	.w2(32'hba95b359),
	.w3(32'hb9ed2224),
	.w4(32'hba7abcfa),
	.w5(32'hba538ce8),
	.w6(32'hbad5800f),
	.w7(32'hbac38473),
	.w8(32'h39c5a7d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ad9f9),
	.w1(32'hbb61e629),
	.w2(32'hbb90d316),
	.w3(32'h3a14e309),
	.w4(32'hba526caf),
	.w5(32'hbb48fef8),
	.w6(32'hbb308637),
	.w7(32'hbb6ee3ef),
	.w8(32'hba927bd7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70cc38),
	.w1(32'h3a67e414),
	.w2(32'h3ae282dd),
	.w3(32'hbac6a5bd),
	.w4(32'hb8e680f9),
	.w5(32'h3a029db0),
	.w6(32'h3a5b02f8),
	.w7(32'h3ae632c3),
	.w8(32'hb8aedded),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94fabab),
	.w1(32'hbb1aefcc),
	.w2(32'hbb76186e),
	.w3(32'hba8593f3),
	.w4(32'hbae08c1c),
	.w5(32'hbb395d90),
	.w6(32'hbabe7e4f),
	.w7(32'hbb1294e3),
	.w8(32'hbaf217de),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f8f78),
	.w1(32'h3a06f4b7),
	.w2(32'h3a8746cd),
	.w3(32'hbb3a3158),
	.w4(32'hba264047),
	.w5(32'h3a5c1ae8),
	.w6(32'hb9137b21),
	.w7(32'h39de1293),
	.w8(32'hb9ee1b18),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083f79),
	.w1(32'hb9b1b73a),
	.w2(32'hba0f36ee),
	.w3(32'hb9636992),
	.w4(32'hb96b178e),
	.w5(32'hbaad6550),
	.w6(32'hbaaa0895),
	.w7(32'h392e47d8),
	.w8(32'h39956d41),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae62591),
	.w1(32'hba464752),
	.w2(32'hbb289a16),
	.w3(32'h39238b4c),
	.w4(32'hb9fae3ee),
	.w5(32'hbac57537),
	.w6(32'hb99c839d),
	.w7(32'hba63cf6b),
	.w8(32'hba9936ef),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1d58),
	.w1(32'hba576a48),
	.w2(32'hba47e77b),
	.w3(32'hbb0d6179),
	.w4(32'hbaa90648),
	.w5(32'h393535f5),
	.w6(32'hbb2542a6),
	.w7(32'hbab55d0b),
	.w8(32'hbacc22bd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ab060),
	.w1(32'hba47eb58),
	.w2(32'hb9e1e508),
	.w3(32'hba332fb8),
	.w4(32'hba270a47),
	.w5(32'hba0be5ab),
	.w6(32'hba035d23),
	.w7(32'hb82f47db),
	.w8(32'h39ca66b9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc2512),
	.w1(32'hbb15eec3),
	.w2(32'hbb05c228),
	.w3(32'hb917ed24),
	.w4(32'hbb1357ab),
	.w5(32'hbb1746eb),
	.w6(32'hbabfb007),
	.w7(32'hba74a74d),
	.w8(32'hb9efbac2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ae6df),
	.w1(32'hbabee9db),
	.w2(32'hbaa31565),
	.w3(32'hbac9ccbf),
	.w4(32'hba734b9d),
	.w5(32'hba51974e),
	.w6(32'hbacc2db4),
	.w7(32'hbac00ca4),
	.w8(32'hb88e7df1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb1b44),
	.w1(32'hbab03058),
	.w2(32'hba909a14),
	.w3(32'h39d18723),
	.w4(32'hb9e240c9),
	.w5(32'hba127c32),
	.w6(32'hba15a02b),
	.w7(32'h383b35c7),
	.w8(32'h394a7097),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7af8de),
	.w1(32'hbad9ee2a),
	.w2(32'hbb21cb4f),
	.w3(32'hba1cb290),
	.w4(32'hba964c3b),
	.w5(32'hbad310ff),
	.w6(32'hbaf364de),
	.w7(32'hbb00c25a),
	.w8(32'hbabc8ba8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e4f86),
	.w1(32'h3a8533ba),
	.w2(32'h3a3ec2e2),
	.w3(32'hbacb27b1),
	.w4(32'h3915b60f),
	.w5(32'hb57adeab),
	.w6(32'h3886797d),
	.w7(32'hb8190081),
	.w8(32'hbaa775c5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76a18),
	.w1(32'hbb008dc4),
	.w2(32'hbbb12625),
	.w3(32'hbae6a4a6),
	.w4(32'h3a108da3),
	.w5(32'hbb755a30),
	.w6(32'hbabbd696),
	.w7(32'hbb8bc03b),
	.w8(32'hbb041fcb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb911416),
	.w1(32'hbb0c7e71),
	.w2(32'hbb5fe0b3),
	.w3(32'hbb03990f),
	.w4(32'hba991bcb),
	.w5(32'hba923262),
	.w6(32'hb9bf8d6b),
	.w7(32'hb9bd2707),
	.w8(32'hb8d087d5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcc254),
	.w1(32'hba7603d6),
	.w2(32'hbaef4cb1),
	.w3(32'hba19a26f),
	.w4(32'hbaae95b4),
	.w5(32'h39c68cff),
	.w6(32'hbb08151e),
	.w7(32'hbaffbff1),
	.w8(32'hbb048920),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e1aa),
	.w1(32'hbac08b34),
	.w2(32'hbba9713c),
	.w3(32'h3a6188ff),
	.w4(32'h3a8b9f54),
	.w5(32'hbb81d0da),
	.w6(32'h39ad3ba1),
	.w7(32'hbbb11da3),
	.w8(32'h398928f9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb067db1),
	.w1(32'hbabb7826),
	.w2(32'hbb7af8ea),
	.w3(32'hb9b33f7d),
	.w4(32'hba8538cd),
	.w5(32'hbb8efd30),
	.w6(32'hba8ef22f),
	.w7(32'hbb86c11e),
	.w8(32'h39b7122c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adce5cc),
	.w1(32'h38b33f76),
	.w2(32'h399874a2),
	.w3(32'h3a8daf4c),
	.w4(32'hb925f82f),
	.w5(32'h3a7af577),
	.w6(32'hbacc76bd),
	.w7(32'hb9d878aa),
	.w8(32'h3a004572),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ef4bda),
	.w1(32'hbab8c8e3),
	.w2(32'hbaf2fd24),
	.w3(32'h390b5b58),
	.w4(32'hbac62cd8),
	.w5(32'hbb19c1e9),
	.w6(32'hba04d2b9),
	.w7(32'hb93ff59b),
	.w8(32'hba4cd0dd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44a8b4),
	.w1(32'hba8433c8),
	.w2(32'hbbaff5f6),
	.w3(32'hbb2cf756),
	.w4(32'h3b3a4272),
	.w5(32'hbadbd2ca),
	.w6(32'hba4719e2),
	.w7(32'hbb632c22),
	.w8(32'hba79f304),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c59cd),
	.w1(32'h3ad1bc7d),
	.w2(32'h3af70a56),
	.w3(32'hbb0f08b1),
	.w4(32'h39222aa9),
	.w5(32'h3b3fe7d8),
	.w6(32'h3a99082c),
	.w7(32'hba321eb6),
	.w8(32'hbb0aa0a8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7882),
	.w1(32'h3a052d81),
	.w2(32'hba6c9c80),
	.w3(32'h3ae50d2a),
	.w4(32'h3a3b80cc),
	.w5(32'hba2c6cfd),
	.w6(32'h3adcb001),
	.w7(32'h3800633d),
	.w8(32'h39c2b8ba),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3ad36),
	.w1(32'h3a22a8f6),
	.w2(32'hba393b76),
	.w3(32'h3ad443ef),
	.w4(32'h3a930a0b),
	.w5(32'h3a70c11d),
	.w6(32'h3ab6612e),
	.w7(32'h3824bff4),
	.w8(32'h38e21a1a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b17fb),
	.w1(32'h3983905a),
	.w2(32'hba34ef64),
	.w3(32'hb7861384),
	.w4(32'h3a173c97),
	.w5(32'hba244745),
	.w6(32'h3a869aef),
	.w7(32'h399f6394),
	.w8(32'hb877e887),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0af572),
	.w1(32'hb9c19392),
	.w2(32'hbaa7cc22),
	.w3(32'h39a7f12f),
	.w4(32'hb9a4d948),
	.w5(32'hba112b0a),
	.w6(32'hb9ab0252),
	.w7(32'hba0060ee),
	.w8(32'hb996d9dd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942aca7),
	.w1(32'h37caf871),
	.w2(32'hba3ec46c),
	.w3(32'hb9e8fd24),
	.w4(32'h3a6ab88c),
	.w5(32'h3ab13fcb),
	.w6(32'h3adbbb3e),
	.w7(32'h3ab6a3d3),
	.w8(32'h3a570ae2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a66f9),
	.w1(32'hbb0a69e0),
	.w2(32'hba9efceb),
	.w3(32'h3aab59f9),
	.w4(32'hba5e0e58),
	.w5(32'hba3824f9),
	.w6(32'hba9c9dbe),
	.w7(32'hb7ba8a22),
	.w8(32'h3a4c3268),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dfb85),
	.w1(32'h3947c654),
	.w2(32'hb85d4c38),
	.w3(32'hb94398e6),
	.w4(32'h3a1c6fc7),
	.w5(32'h39e3411f),
	.w6(32'h3a0a47a9),
	.w7(32'hb94232cd),
	.w8(32'h39fcc2f1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaabdb4),
	.w1(32'hbac5265b),
	.w2(32'hba52813b),
	.w3(32'hb9acd243),
	.w4(32'hbaedb837),
	.w5(32'hba471050),
	.w6(32'hbb07ad7d),
	.w7(32'hba99fd52),
	.w8(32'hbb28b084),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50bef4),
	.w1(32'hba64add1),
	.w2(32'hbab4b0d9),
	.w3(32'hbac5be07),
	.w4(32'hb9a2be77),
	.w5(32'hbaad4e30),
	.w6(32'hba51ac55),
	.w7(32'hba27bc39),
	.w8(32'hbaa9e998),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafef4b1),
	.w1(32'h3af9e90e),
	.w2(32'h3b1d8b1e),
	.w3(32'hbaf5aa38),
	.w4(32'h3a57b021),
	.w5(32'h3a9296d9),
	.w6(32'h3a2624db),
	.w7(32'h3b160bae),
	.w8(32'h3a4def10),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38a738),
	.w1(32'hbaab12d5),
	.w2(32'hbb03eaec),
	.w3(32'h3a09af94),
	.w4(32'hbaa942e8),
	.w5(32'hbb046e72),
	.w6(32'hba010528),
	.w7(32'hba77e711),
	.w8(32'hbadbc186),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17e73e),
	.w1(32'h3a20cd6d),
	.w2(32'hba57b012),
	.w3(32'hbb052489),
	.w4(32'h3a9e3a53),
	.w5(32'h3a8b9ce7),
	.w6(32'h3a7f9bee),
	.w7(32'h39c93a88),
	.w8(32'h39be4c84),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369c2520),
	.w1(32'h38b41c44),
	.w2(32'h3a608d68),
	.w3(32'h3a27a0f7),
	.w4(32'hb9eaacfb),
	.w5(32'h39186e25),
	.w6(32'h39aed61c),
	.w7(32'h3a823195),
	.w8(32'h391e9ddc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb898c6bf),
	.w1(32'h39643fc4),
	.w2(32'hba291fbe),
	.w3(32'hb90f5437),
	.w4(32'h39f94995),
	.w5(32'hba287bde),
	.w6(32'h3a93daeb),
	.w7(32'h38364210),
	.w8(32'h39788a68),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba626582),
	.w1(32'h399caa6e),
	.w2(32'hb92eaf32),
	.w3(32'h39da1f1d),
	.w4(32'h3a147a81),
	.w5(32'hb88932b2),
	.w6(32'h3a3bf8e9),
	.w7(32'h390cd5dc),
	.w8(32'h39667cde),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385eee20),
	.w1(32'h3a579d4a),
	.w2(32'h39afa9f4),
	.w3(32'h3a184b41),
	.w4(32'h3a4e4ead),
	.w5(32'hb8c560d8),
	.w6(32'h3a94bb1e),
	.w7(32'h3a19697c),
	.w8(32'h39b4f512),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957b163),
	.w1(32'hba907eb9),
	.w2(32'hbaa2977f),
	.w3(32'h3954a06f),
	.w4(32'hba2f0aec),
	.w5(32'hb9cb1793),
	.w6(32'h3ac16951),
	.w7(32'h39ef2b16),
	.w8(32'h3992d604),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a181f9f),
	.w1(32'hbadcebec),
	.w2(32'hbb9a9b56),
	.w3(32'h3a5c0190),
	.w4(32'hba50b3f9),
	.w5(32'hbb3ec52f),
	.w6(32'hbae5936a),
	.w7(32'hbb5833aa),
	.w8(32'hb8bd1b7a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a9cb1),
	.w1(32'hba0adce5),
	.w2(32'hb9f3e2c3),
	.w3(32'hb9d70990),
	.w4(32'hba96456a),
	.w5(32'hba373dc0),
	.w6(32'hba46ba13),
	.w7(32'h3a50a1e5),
	.w8(32'hb8096a3a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c062e8),
	.w1(32'h398ab220),
	.w2(32'h37157d46),
	.w3(32'hba98b0b2),
	.w4(32'hb999c46f),
	.w5(32'h376c56d4),
	.w6(32'hb9bdbdb6),
	.w7(32'h3a30aeba),
	.w8(32'hba007d16),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a5bf7),
	.w1(32'hb9b8ccf5),
	.w2(32'hba6af9d0),
	.w3(32'hbb0bbf4b),
	.w4(32'hb9050cf8),
	.w5(32'hba390ee0),
	.w6(32'h38feffc4),
	.w7(32'hb986cb72),
	.w8(32'hb9a5b66c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba138b82),
	.w1(32'h3b1ff8fe),
	.w2(32'h3b208629),
	.w3(32'hb68b65fb),
	.w4(32'h3aab1654),
	.w5(32'h3b8d9288),
	.w6(32'h3ad2fa48),
	.w7(32'hb916c061),
	.w8(32'h399a1fd3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8400b),
	.w1(32'hbb3e97ee),
	.w2(32'hbad0db61),
	.w3(32'h3b1a1434),
	.w4(32'hbb4b21f0),
	.w5(32'hbb1cdd59),
	.w6(32'hbae9b26b),
	.w7(32'h38a4cf82),
	.w8(32'hba2f55a7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02b9da),
	.w1(32'hbac0b534),
	.w2(32'hba8a245e),
	.w3(32'hbb1d5d0d),
	.w4(32'hba90fe64),
	.w5(32'hba72bad0),
	.w6(32'hba860db6),
	.w7(32'hb9a26caf),
	.w8(32'h39fa630a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44b3d9),
	.w1(32'hb9657b47),
	.w2(32'h39d29fff),
	.w3(32'hb9ab67de),
	.w4(32'h38aa3069),
	.w5(32'h392983d4),
	.w6(32'hb827d9a9),
	.w7(32'h39b49533),
	.w8(32'hb8a7a378),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b0de3),
	.w1(32'h3a1aacc9),
	.w2(32'h3a5c6aa1),
	.w3(32'hb8f961d9),
	.w4(32'h3a3400ae),
	.w5(32'h3a42bf19),
	.w6(32'h39a68998),
	.w7(32'h3882817f),
	.w8(32'h396c666e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de6168),
	.w1(32'h3ab320cc),
	.w2(32'h3b0474d7),
	.w3(32'h3a444ebc),
	.w4(32'h3b163076),
	.w5(32'h3b0d3bbc),
	.w6(32'h3998d1e7),
	.w7(32'h3ae27d56),
	.w8(32'h3acdcf78),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34560),
	.w1(32'hba8d2c75),
	.w2(32'hba721077),
	.w3(32'h3a9bd083),
	.w4(32'hba7d7ccd),
	.w5(32'hba916a7d),
	.w6(32'hba897781),
	.w7(32'hba6d133a),
	.w8(32'hba8427ac),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba581be0),
	.w1(32'hbaaed32c),
	.w2(32'hba0305b3),
	.w3(32'hba5db448),
	.w4(32'hba8f997f),
	.w5(32'hba87a696),
	.w6(32'hba549ec2),
	.w7(32'hb9ad42a1),
	.w8(32'hba0656f0),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba207dc8),
	.w1(32'hba859ba7),
	.w2(32'hb9d6bf97),
	.w3(32'hba720644),
	.w4(32'hb90c2c63),
	.w5(32'hb71dcd16),
	.w6(32'h39c4eecf),
	.w7(32'hba2fe68c),
	.w8(32'hba6fa17f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22a442),
	.w1(32'h3af60ec0),
	.w2(32'h3a47793b),
	.w3(32'hba366226),
	.w4(32'h3b15d187),
	.w5(32'h3a2a0876),
	.w6(32'h3ae88ed0),
	.w7(32'hb9fc8e7a),
	.w8(32'h3abf1673),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b073adc),
	.w1(32'h3a67a389),
	.w2(32'h3abed5e1),
	.w3(32'h3a670d9c),
	.w4(32'h3ab0e128),
	.w5(32'h3aab297f),
	.w6(32'h3a2bf566),
	.w7(32'h39dced51),
	.w8(32'h39928220),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b7d7e),
	.w1(32'hba51b581),
	.w2(32'hba79b1b1),
	.w3(32'h3a7d675d),
	.w4(32'hba6161c6),
	.w5(32'hba56969f),
	.w6(32'hba78ec39),
	.w7(32'hba9fd9fb),
	.w8(32'hba4ae2c8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc686a),
	.w1(32'h3991b4f5),
	.w2(32'h3a0c931d),
	.w3(32'hba585be6),
	.w4(32'h39b550dc),
	.w5(32'h39d0ae78),
	.w6(32'h39cc7691),
	.w7(32'h3a247115),
	.w8(32'h3a32e39e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf640e),
	.w1(32'h39deba49),
	.w2(32'h39ad2a0f),
	.w3(32'h39406c4a),
	.w4(32'h3a56f182),
	.w5(32'h3a553521),
	.w6(32'hb9ac7271),
	.w7(32'hb887ce41),
	.w8(32'h396495d9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38046ed2),
	.w1(32'hba800cdc),
	.w2(32'hba80fccc),
	.w3(32'h39979725),
	.w4(32'hba2cd8af),
	.w5(32'hba3eceb0),
	.w6(32'hba3b24a3),
	.w7(32'hba80ab00),
	.w8(32'hba95ed3c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fecf7),
	.w1(32'hbac76e42),
	.w2(32'hba81c785),
	.w3(32'hb9cd9a83),
	.w4(32'hba9231c6),
	.w5(32'hb901b6d4),
	.w6(32'hba8f5836),
	.w7(32'hba035fc9),
	.w8(32'hba9eb9f6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa547e4),
	.w1(32'h3a70a498),
	.w2(32'h39cfd594),
	.w3(32'hbaa07801),
	.w4(32'h3a9f59ab),
	.w5(32'h3a9ba21c),
	.w6(32'h3a807bb9),
	.w7(32'h3a8cdf6b),
	.w8(32'h36a01366),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9866b2a),
	.w1(32'hb9593dea),
	.w2(32'h3770e6d3),
	.w3(32'hb9e77274),
	.w4(32'h39294760),
	.w5(32'h39e46fd7),
	.w6(32'hb9cfe0a9),
	.w7(32'hb93310ea),
	.w8(32'hb910b32a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446732),
	.w1(32'hb7ac96ac),
	.w2(32'h39a2370d),
	.w3(32'hb9827624),
	.w4(32'h3932eb72),
	.w5(32'hb96e0866),
	.w6(32'h378e8a08),
	.w7(32'h3a30f205),
	.w8(32'hb86226b7),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f910ae),
	.w1(32'hb994ee98),
	.w2(32'h3aafb75b),
	.w3(32'hb9d5f603),
	.w4(32'h3af1c500),
	.w5(32'h3acc7c0f),
	.w6(32'h3a4d43c9),
	.w7(32'h3a805289),
	.w8(32'h3a3cc35c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86fb76),
	.w1(32'h3a00456a),
	.w2(32'h398f3008),
	.w3(32'h3a2b2551),
	.w4(32'h3a41fe9c),
	.w5(32'h3a31aab3),
	.w6(32'h37f2545e),
	.w7(32'hb8c323c6),
	.w8(32'h390a061f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994b016),
	.w1(32'h391982fa),
	.w2(32'hb9840fb5),
	.w3(32'h3a2fc87c),
	.w4(32'hb9db465f),
	.w5(32'hba780268),
	.w6(32'h3971b8e1),
	.w7(32'hb9a21ae7),
	.w8(32'h34fed3b6),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba891be7),
	.w1(32'hba81a70b),
	.w2(32'hba651752),
	.w3(32'hba688f58),
	.w4(32'hba51db03),
	.w5(32'hb9d22fe1),
	.w6(32'hbaa2637e),
	.w7(32'hbaab0a5d),
	.w8(32'hbaa0819b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba902b0c),
	.w1(32'hba381c28),
	.w2(32'hb9ac6e70),
	.w3(32'hb9c4bed6),
	.w4(32'hba2ca26a),
	.w5(32'hba05d80c),
	.w6(32'hba080324),
	.w7(32'hb9943cd6),
	.w8(32'hb9dd85ab),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db307a),
	.w1(32'h39b53949),
	.w2(32'h38841bcc),
	.w3(32'hb9c8b804),
	.w4(32'h3a24b2b0),
	.w5(32'h39f2f972),
	.w6(32'hb99c444d),
	.w7(32'hb9d21c18),
	.w8(32'hb7eb9620),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9919ca5),
	.w1(32'h39bae1f4),
	.w2(32'h39802ed0),
	.w3(32'h38df2801),
	.w4(32'h3a772c09),
	.w5(32'h3a1a6de1),
	.w6(32'h39aebfd7),
	.w7(32'hb8e6910e),
	.w8(32'hb8de86de),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9df4a),
	.w1(32'hba2c3af3),
	.w2(32'hba493bc2),
	.w3(32'h3972c7c7),
	.w4(32'hb9957e96),
	.w5(32'h39f3fb42),
	.w6(32'hba7b985e),
	.w7(32'hbaa405cf),
	.w8(32'hbad90174),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba239f88),
	.w1(32'h3a2ab5db),
	.w2(32'h39b2cc62),
	.w3(32'hb9cea5dd),
	.w4(32'hba73dac2),
	.w5(32'hbaa44e27),
	.w6(32'hb89214c9),
	.w7(32'hba0ed86d),
	.w8(32'hba0078ea),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d30efc),
	.w1(32'h38a5034f),
	.w2(32'h390e7dd6),
	.w3(32'hb999c4ee),
	.w4(32'h37e32c3d),
	.w5(32'hb8ddbd41),
	.w6(32'hb918c1c1),
	.w7(32'h385045a5),
	.w8(32'h3679685d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391505dd),
	.w1(32'hb9c3516d),
	.w2(32'hba546246),
	.w3(32'h395c79b5),
	.w4(32'h385a7072),
	.w5(32'hb904c48b),
	.w6(32'hba1158f4),
	.w7(32'hb9fe676c),
	.w8(32'hba0c2ab1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8189097),
	.w1(32'h3a79d04d),
	.w2(32'h388a6ed9),
	.w3(32'h38ee4f78),
	.w4(32'h39babbf3),
	.w5(32'hb9c9cca9),
	.w6(32'h3a361f4f),
	.w7(32'h395f279b),
	.w8(32'hb9d5d101),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0ca4a),
	.w1(32'h39bbafa2),
	.w2(32'h39cdad3c),
	.w3(32'h390f9922),
	.w4(32'h3abcf29f),
	.w5(32'h3a9727ef),
	.w6(32'h3a42eb6d),
	.w7(32'h39f737cf),
	.w8(32'h3a1bf37d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac20241),
	.w1(32'hba69538c),
	.w2(32'hbaad30e4),
	.w3(32'hba871ad6),
	.w4(32'hb968ee09),
	.w5(32'hb9bacbdf),
	.w6(32'hbaf632bd),
	.w7(32'hbab80eb1),
	.w8(32'hbaadc49b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6dd2a3),
	.w1(32'hba70f1fd),
	.w2(32'h3a178e50),
	.w3(32'hba123792),
	.w4(32'hba4ecefe),
	.w5(32'h39c6125a),
	.w6(32'hba1b0aa6),
	.w7(32'hb83a7721),
	.w8(32'h39a0d064),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12fc93),
	.w1(32'hb9c8ee59),
	.w2(32'h3a2e4ed0),
	.w3(32'h3a111e5d),
	.w4(32'hba3afd0f),
	.w5(32'h39dbdc66),
	.w6(32'hb93589a9),
	.w7(32'h3a516d8e),
	.w8(32'h3a2e7411),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcea1b),
	.w1(32'h376d7435),
	.w2(32'h38d7327c),
	.w3(32'h3971842e),
	.w4(32'h39e7c6ff),
	.w5(32'h3975700e),
	.w6(32'hb8fa8fdd),
	.w7(32'hb975b673),
	.w8(32'hb939e5e8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9296cc8),
	.w1(32'h39798773),
	.w2(32'h39c7e304),
	.w3(32'h3923e4d3),
	.w4(32'h39d24cf2),
	.w5(32'h39e70628),
	.w6(32'hb9063668),
	.w7(32'hb97ceed2),
	.w8(32'hb9c942b6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c7461),
	.w1(32'h39388717),
	.w2(32'h387c8de0),
	.w3(32'h38921cbf),
	.w4(32'hb93655ee),
	.w5(32'hb80af06f),
	.w6(32'hba0214b8),
	.w7(32'hb8797629),
	.w8(32'hba1b7e31),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88643c),
	.w1(32'h39257dae),
	.w2(32'h3ac1b1cf),
	.w3(32'hbac4111d),
	.w4(32'h37aae369),
	.w5(32'h3a67cf6b),
	.w6(32'hba54eef6),
	.w7(32'h3a24e1ee),
	.w8(32'h3a49dbd9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e1433),
	.w1(32'hba3f76ab),
	.w2(32'hba8e9713),
	.w3(32'h3a3fab1b),
	.w4(32'h3676dbee),
	.w5(32'hb90e2335),
	.w6(32'hba942c2c),
	.w7(32'hba7e6b03),
	.w8(32'hbaa31340),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac424f4),
	.w1(32'h3935db08),
	.w2(32'h3998beb1),
	.w3(32'hba4415b3),
	.w4(32'h39b4b4f5),
	.w5(32'h376895c6),
	.w6(32'hb817c05c),
	.w7(32'hb9a55d8a),
	.w8(32'hba205764),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947a238),
	.w1(32'hba097542),
	.w2(32'hba142fcc),
	.w3(32'h392b00ac),
	.w4(32'hb8c18883),
	.w5(32'hb9a6a043),
	.w6(32'hba1c3848),
	.w7(32'hba95ce8e),
	.w8(32'hba96736d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba860e8b),
	.w1(32'hba6bdb97),
	.w2(32'hb9cd2490),
	.w3(32'hba104480),
	.w4(32'hba443e18),
	.w5(32'hba1d7c98),
	.w6(32'hba474b3c),
	.w7(32'hba1c3ad5),
	.w8(32'hb9fd0a1a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c70553),
	.w1(32'h39a695d2),
	.w2(32'h39b7a3af),
	.w3(32'hba1057af),
	.w4(32'h3a20e24c),
	.w5(32'h39f8ec33),
	.w6(32'h3a0b4493),
	.w7(32'h39c75098),
	.w8(32'h39ace2fb),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b58817),
	.w1(32'hba3319d4),
	.w2(32'hba0edddf),
	.w3(32'h3935a769),
	.w4(32'hba35016b),
	.w5(32'hba0002fd),
	.w6(32'hba2aff28),
	.w7(32'h3811e8ca),
	.w8(32'h3988ff2e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a974f),
	.w1(32'hba843913),
	.w2(32'h39b6c0b6),
	.w3(32'hba3b88e4),
	.w4(32'hbaa1695b),
	.w5(32'h391ed7b9),
	.w6(32'hba8c51c9),
	.w7(32'h3a235594),
	.w8(32'h3a74efc3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2c512),
	.w1(32'hbabac5b4),
	.w2(32'hba886bf0),
	.w3(32'h3a7d283d),
	.w4(32'hba9c9abb),
	.w5(32'hba512ee4),
	.w6(32'hba73c7ee),
	.w7(32'hba7d13e3),
	.w8(32'hbaa9825b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22e73e),
	.w1(32'h3a2fd32d),
	.w2(32'h3a60307d),
	.w3(32'hb9d70c3a),
	.w4(32'h3a2668fe),
	.w5(32'h3a6fae14),
	.w6(32'hb83c1b44),
	.w7(32'h396f8970),
	.w8(32'h39d42979),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920b0a9),
	.w1(32'hba8bbd0b),
	.w2(32'hbabed60c),
	.w3(32'h391244b6),
	.w4(32'hba27aad8),
	.w5(32'hb9d8407e),
	.w6(32'hba21e631),
	.w7(32'hba15d91a),
	.w8(32'hb9a5cfad),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2a5a7),
	.w1(32'hba3e67e8),
	.w2(32'hb98f4d64),
	.w3(32'hb841dfc3),
	.w4(32'h3996236a),
	.w5(32'hba2b2140),
	.w6(32'hba4913e3),
	.w7(32'hb9b240b9),
	.w8(32'hba3f43e3),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d46819),
	.w1(32'hba55c7b4),
	.w2(32'hba30cb05),
	.w3(32'hba0ebd37),
	.w4(32'hb9d859bf),
	.w5(32'hb792b1e3),
	.w6(32'hba0f60ec),
	.w7(32'hbaaa0afb),
	.w8(32'hba557c02),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3833c398),
	.w1(32'hb9504597),
	.w2(32'hb7b11646),
	.w3(32'h398ad8ac),
	.w4(32'h399c2567),
	.w5(32'h3a7d774a),
	.w6(32'h3a6e0046),
	.w7(32'h3ac9f8c2),
	.w8(32'h3a9bf071),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8c9ba),
	.w1(32'hb9a205ab),
	.w2(32'h3990ce69),
	.w3(32'h39b0456f),
	.w4(32'hb8c5c1c2),
	.w5(32'h3a3b3477),
	.w6(32'hb8aefbae),
	.w7(32'h39885b36),
	.w8(32'h38805b7b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21548b),
	.w1(32'h396af222),
	.w2(32'h39e5d9fd),
	.w3(32'hba35b533),
	.w4(32'h39d2afa4),
	.w5(32'h3a05f9f6),
	.w6(32'hb9f031df),
	.w7(32'hb654a97f),
	.w8(32'hb9202df0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944eae7),
	.w1(32'h387d7450),
	.w2(32'h3989dd45),
	.w3(32'h394e531a),
	.w4(32'h38a678a4),
	.w5(32'h38eef6a2),
	.w6(32'h39bce29f),
	.w7(32'h39ecafcb),
	.w8(32'h39eb880f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39572284),
	.w1(32'hba49e3eb),
	.w2(32'hbaace5c6),
	.w3(32'h39268e9b),
	.w4(32'hba8eb789),
	.w5(32'hba8b2a7d),
	.w6(32'hba1c3b34),
	.w7(32'hba8a18c1),
	.w8(32'hba527272),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77972d),
	.w1(32'h3a8e42f9),
	.w2(32'hba8fb1bd),
	.w3(32'hba4623bc),
	.w4(32'h3afd6512),
	.w5(32'h3ad685a9),
	.w6(32'h3a2b0fb2),
	.w7(32'h3ab71297),
	.w8(32'h3a1ddcd5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e27a2),
	.w1(32'h3815df25),
	.w2(32'hb60b07fe),
	.w3(32'h39bd4e07),
	.w4(32'h3a76eff9),
	.w5(32'h39ffe130),
	.w6(32'hba1e73a6),
	.w7(32'hba7f15eb),
	.w8(32'hb9f69131),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f8486),
	.w1(32'h3af0fc1b),
	.w2(32'h3a2a2268),
	.w3(32'h3a13acbd),
	.w4(32'h3b182bbc),
	.w5(32'h3a7636eb),
	.w6(32'h3af2e2e1),
	.w7(32'h39b49e5d),
	.w8(32'h39ec2528),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ca799),
	.w1(32'h371353ff),
	.w2(32'hb90f40b2),
	.w3(32'h3a05d302),
	.w4(32'hb9bb905f),
	.w5(32'hba486317),
	.w6(32'h399e767e),
	.w7(32'h38db588f),
	.w8(32'hb9776b55),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f880de),
	.w1(32'hba4060f0),
	.w2(32'h3a822550),
	.w3(32'hb9302bad),
	.w4(32'hb9e81ccb),
	.w5(32'h39dc5f63),
	.w6(32'hba957aa5),
	.w7(32'h39195fea),
	.w8(32'h3a5b284f),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad67e0),
	.w1(32'hba3fec9a),
	.w2(32'hb9eb3e13),
	.w3(32'h3a1d3a2a),
	.w4(32'hba4e429b),
	.w5(32'hba5a11ca),
	.w6(32'hba73ab33),
	.w7(32'hba934ec0),
	.w8(32'hba0aa944),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb42cb),
	.w1(32'h3a43ed3e),
	.w2(32'hb89192e6),
	.w3(32'h393781c6),
	.w4(32'h39b4a6b9),
	.w5(32'hb8f9dc10),
	.w6(32'h3a9b90b3),
	.w7(32'hba4fef90),
	.w8(32'hb83225f8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c2816),
	.w1(32'hba8d04be),
	.w2(32'hba63107b),
	.w3(32'h3a141dcf),
	.w4(32'hba85cd8f),
	.w5(32'hba8cb346),
	.w6(32'hba0120ed),
	.w7(32'hb8db07a5),
	.w8(32'h38686807),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e59d5),
	.w1(32'hba30f98b),
	.w2(32'hb8924ea2),
	.w3(32'hba9aa16b),
	.w4(32'h3964b44b),
	.w5(32'hb768e3aa),
	.w6(32'hba07161b),
	.w7(32'hb9c62b92),
	.w8(32'hb9c67868),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fc3a06),
	.w1(32'hbaf91167),
	.w2(32'hba654807),
	.w3(32'h392571d6),
	.w4(32'hba9308bd),
	.w5(32'hbaa17bfb),
	.w6(32'hbac6b6e5),
	.w7(32'hb98307a3),
	.w8(32'hb980a9b6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f92bb3),
	.w1(32'h393cd92e),
	.w2(32'h37c0a880),
	.w3(32'hb9ee2d87),
	.w4(32'h3a2d570c),
	.w5(32'h39cf7dd9),
	.w6(32'hb9621000),
	.w7(32'h385903bd),
	.w8(32'h387b565b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e11ba6),
	.w1(32'h3ad238eb),
	.w2(32'h3aefed1d),
	.w3(32'hb927036c),
	.w4(32'h3b09ff07),
	.w5(32'h3ac5ac13),
	.w6(32'h39d616c5),
	.w7(32'h3a9c0958),
	.w8(32'h3a6297d0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43a29d),
	.w1(32'hba88dfba),
	.w2(32'hbaa1cfd6),
	.w3(32'hb88b15fa),
	.w4(32'hba31df5e),
	.w5(32'hba0df938),
	.w6(32'hba3a85e9),
	.w7(32'hba484658),
	.w8(32'hba324bea),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933b363),
	.w1(32'hba284cac),
	.w2(32'h3932582d),
	.w3(32'h382c3baf),
	.w4(32'hba8cdb4b),
	.w5(32'hb9fdc71b),
	.w6(32'hb9cfea69),
	.w7(32'hb91b67f5),
	.w8(32'hb91313e5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9833203),
	.w1(32'hb88679c5),
	.w2(32'hba9a07cd),
	.w3(32'hb96c4655),
	.w4(32'hba053905),
	.w5(32'hb9176a62),
	.w6(32'h395367f7),
	.w7(32'hbaaae7e8),
	.w8(32'hba7e77b7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08c269),
	.w1(32'hbab76db6),
	.w2(32'hb9cdae1b),
	.w3(32'h3a42d82b),
	.w4(32'hbab9dca4),
	.w5(32'hb9d656f3),
	.w6(32'hba9a1bca),
	.w7(32'hb9f9cb50),
	.w8(32'hba615f41),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba760cb0),
	.w1(32'hba27dc97),
	.w2(32'hb6f890a0),
	.w3(32'hb9f11b32),
	.w4(32'hba896354),
	.w5(32'hb9fae93d),
	.w6(32'hba396d30),
	.w7(32'hb90d1861),
	.w8(32'h38cff63a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1407f),
	.w1(32'h39e87e9c),
	.w2(32'h39e82b71),
	.w3(32'hb932cc70),
	.w4(32'h3a87874a),
	.w5(32'h3a385ad9),
	.w6(32'h38b5018f),
	.w7(32'hb8981f9e),
	.w8(32'h39596e76),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a33c45),
	.w1(32'hbaa03274),
	.w2(32'hbab713aa),
	.w3(32'h3a08beef),
	.w4(32'hbb0540af),
	.w5(32'hba530112),
	.w6(32'hb9a0466f),
	.w7(32'hbaec9611),
	.w8(32'hbae42efd),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88fd06),
	.w1(32'hba407c80),
	.w2(32'hba1324cf),
	.w3(32'hb9da5091),
	.w4(32'hba211317),
	.w5(32'hb9ebedae),
	.w6(32'hba537a42),
	.w7(32'hba32a812),
	.w8(32'hba3e5e67),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a14f),
	.w1(32'h38426ffc),
	.w2(32'h398da45e),
	.w3(32'hba0844a7),
	.w4(32'h399d3a5c),
	.w5(32'h392c3fe2),
	.w6(32'h39496794),
	.w7(32'hb793ebf5),
	.w8(32'h38b47fef),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cb2e4c),
	.w1(32'h399a5dd6),
	.w2(32'h39fda9ce),
	.w3(32'h39da2b7c),
	.w4(32'h3a0a6a5d),
	.w5(32'h3a0c07e9),
	.w6(32'h398b67e9),
	.w7(32'h398745a0),
	.w8(32'h39c7d6fe),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991c886),
	.w1(32'h3972d849),
	.w2(32'h39f8203d),
	.w3(32'h3a02a274),
	.w4(32'h3a091b7e),
	.w5(32'h39cfa396),
	.w6(32'hb95f416f),
	.w7(32'hba045fd0),
	.w8(32'hba0b205b),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a0bb0),
	.w1(32'hba8b3cc9),
	.w2(32'hba81daf9),
	.w3(32'h38e6f4df),
	.w4(32'hba826e93),
	.w5(32'hba808361),
	.w6(32'hba092d53),
	.w7(32'hb9b06b5f),
	.w8(32'hb9aeabbe),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37a82b),
	.w1(32'hb99f2218),
	.w2(32'hbb4e839a),
	.w3(32'hba2db595),
	.w4(32'h38a3b7c4),
	.w5(32'hb9554d02),
	.w6(32'hb9a38e3d),
	.w7(32'hb945e17e),
	.w8(32'hbad9c33f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd786f),
	.w1(32'h3a0bb247),
	.w2(32'h3a05f7d2),
	.w3(32'hba773cca),
	.w4(32'h3a4bf037),
	.w5(32'h3a3664f0),
	.w6(32'h3a3b0582),
	.w7(32'h3a3cb3a7),
	.w8(32'h3a096094),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf2e89),
	.w1(32'hba73ea52),
	.w2(32'hb905e4e1),
	.w3(32'h3a0fbef1),
	.w4(32'hba4406a4),
	.w5(32'hb97c9452),
	.w6(32'hba7af3dd),
	.w7(32'hb98d80b4),
	.w8(32'h394c6860),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3651977c),
	.w1(32'h3a263419),
	.w2(32'hb98b941e),
	.w3(32'hb9362fbd),
	.w4(32'hb984aa2b),
	.w5(32'hba530030),
	.w6(32'h390350ab),
	.w7(32'h399ce442),
	.w8(32'hba0a68d8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad67486),
	.w1(32'hb941fa8b),
	.w2(32'hb7547b07),
	.w3(32'hba91402e),
	.w4(32'h39c67b43),
	.w5(32'h399793a5),
	.w6(32'hb91d8106),
	.w7(32'hb92c5949),
	.w8(32'hb98ae460),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae83eb),
	.w1(32'hb9d9a29d),
	.w2(32'h39581360),
	.w3(32'h39e3c92f),
	.w4(32'hba7f1282),
	.w5(32'hb98228bd),
	.w6(32'hba25af0f),
	.w7(32'hb85c46a9),
	.w8(32'h398c7191),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dafaa),
	.w1(32'hbaa203c3),
	.w2(32'hba88d95d),
	.w3(32'h39366778),
	.w4(32'hbabf6742),
	.w5(32'hbaa229e8),
	.w6(32'hba74c6be),
	.w7(32'hba80ce87),
	.w8(32'hba094f2c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1df982),
	.w1(32'hb96937c0),
	.w2(32'hb89ddc5a),
	.w3(32'hba83c0fe),
	.w4(32'hb91d68f5),
	.w5(32'h38e50fe8),
	.w6(32'hb9a00e7a),
	.w7(32'hb9bf22e6),
	.w8(32'hb98e5aab),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9845979),
	.w1(32'hba5838d2),
	.w2(32'hb9e28a42),
	.w3(32'hb7569b78),
	.w4(32'hba93a02b),
	.w5(32'hba97501b),
	.w6(32'hb9eb6251),
	.w7(32'hb95be66b),
	.w8(32'hb9441940),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef2932),
	.w1(32'hba159285),
	.w2(32'h3a3ea4aa),
	.w3(32'hba52225d),
	.w4(32'hba412d3f),
	.w5(32'hb9b6fdb7),
	.w6(32'hba961d88),
	.w7(32'h39cb0722),
	.w8(32'h3a07f840),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394dbf72),
	.w1(32'hbab9cb96),
	.w2(32'hba973d46),
	.w3(32'hbab0eef5),
	.w4(32'hbabb9e39),
	.w5(32'hba9a3836),
	.w6(32'hbad77532),
	.w7(32'hbaa7bd3b),
	.w8(32'hba91aad2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7aa09),
	.w1(32'h398af656),
	.w2(32'hb8f58c6d),
	.w3(32'hba16d0b1),
	.w4(32'h39ed5bec),
	.w5(32'h3a02868c),
	.w6(32'hb9f1d701),
	.w7(32'hb91d1daa),
	.w8(32'hba3526ee),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5145a7),
	.w1(32'h397214cf),
	.w2(32'h394c476e),
	.w3(32'hba090c54),
	.w4(32'h3a3350e6),
	.w5(32'h39ee0e81),
	.w6(32'h389f8cc1),
	.w7(32'hb971ae25),
	.w8(32'hb88ed070),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350b4849),
	.w1(32'hb5233e17),
	.w2(32'h392ceaed),
	.w3(32'h39b04af6),
	.w4(32'hb9905189),
	.w5(32'hb99fbe98),
	.w6(32'h3a0154c8),
	.w7(32'h39d1bd76),
	.w8(32'h3912a58d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb935011d),
	.w1(32'h3a415e4d),
	.w2(32'h3a0f89e4),
	.w3(32'h36b7101e),
	.w4(32'h3a83ecec),
	.w5(32'h39e7d9ad),
	.w6(32'h3a2d74cd),
	.w7(32'h378a6ab9),
	.w8(32'hb96fd457),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75dff91),
	.w1(32'h384ebef0),
	.w2(32'hb7ec79b4),
	.w3(32'h39a13fc1),
	.w4(32'h396ac63e),
	.w5(32'h39179be5),
	.w6(32'hb9da776b),
	.w7(32'hba183c2f),
	.w8(32'hb9c65542),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967b253),
	.w1(32'hba616223),
	.w2(32'hba0ebcb0),
	.w3(32'h37a484e7),
	.w4(32'hba8cce68),
	.w5(32'hba683f6b),
	.w6(32'hba69555b),
	.w7(32'hba8d60d6),
	.w8(32'hba9fbc53),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb4212),
	.w1(32'hb9f97fab),
	.w2(32'hba0981f2),
	.w3(32'hb9e246ff),
	.w4(32'hba173eaf),
	.w5(32'hba64e83f),
	.w6(32'hba08831c),
	.w7(32'hba05db64),
	.w8(32'hba41e720),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa4063),
	.w1(32'hba7275c3),
	.w2(32'h397c6d81),
	.w3(32'hba99bb4a),
	.w4(32'hba77b88c),
	.w5(32'hb9548f46),
	.w6(32'hba73980c),
	.w7(32'h37905164),
	.w8(32'h3a02ee0d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e6710),
	.w1(32'hba71a6f2),
	.w2(32'hb99cc513),
	.w3(32'h39df15ff),
	.w4(32'hbaa1bde0),
	.w5(32'hba8042f7),
	.w6(32'hba6d7a93),
	.w7(32'hba20fc4f),
	.w8(32'hba2c6255),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1910a4),
	.w1(32'hb748718e),
	.w2(32'hba112418),
	.w3(32'hba5c7bb1),
	.w4(32'hb8480a11),
	.w5(32'hb75bc0eb),
	.w6(32'h39d6e0a0),
	.w7(32'h38f9a988),
	.w8(32'hb9673b14),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0dfb42),
	.w1(32'h3867b5ed),
	.w2(32'h39637b5a),
	.w3(32'h39ad6974),
	.w4(32'hba79394d),
	.w5(32'hba3ca3a1),
	.w6(32'hb9d4939b),
	.w7(32'hb8a7a67e),
	.w8(32'h3a1c8f31),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a513837),
	.w1(32'h39333a3a),
	.w2(32'h3a431cbe),
	.w3(32'h39627e67),
	.w4(32'h3a5adeae),
	.w5(32'h3a5c15bf),
	.w6(32'hb9c3b3d6),
	.w7(32'h3a509d3f),
	.w8(32'hb98a9ee9),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c10e50),
	.w1(32'hbabbc7ab),
	.w2(32'hba332495),
	.w3(32'hb936f9de),
	.w4(32'hbad276b7),
	.w5(32'hbaa13467),
	.w6(32'hba38d839),
	.w7(32'hb9f0122e),
	.w8(32'hb94d8051),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c69dc),
	.w1(32'hba2239f1),
	.w2(32'hb9ca6e9a),
	.w3(32'hbaa8fb69),
	.w4(32'hb98fdcfd),
	.w5(32'hb8adc230),
	.w6(32'hbaa4da88),
	.w7(32'hba8787f7),
	.w8(32'hba39f8e5),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20b164),
	.w1(32'hb7645cc6),
	.w2(32'hb887b915),
	.w3(32'hb8d19e4e),
	.w4(32'hba3037bd),
	.w5(32'hba7fd4f5),
	.w6(32'hb9690840),
	.w7(32'hb9a08989),
	.w8(32'h3745cf38),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1009da),
	.w1(32'hb8de8828),
	.w2(32'hbb56f618),
	.w3(32'h3ab19323),
	.w4(32'hba861500),
	.w5(32'hbaf123e8),
	.w6(32'h39854af9),
	.w7(32'hbab4c825),
	.w8(32'h39aab440),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390f7aad),
	.w1(32'h3a1f65c9),
	.w2(32'h3a1c9f88),
	.w3(32'h39f004a1),
	.w4(32'h3a65abae),
	.w5(32'h3a82a18d),
	.w6(32'h3a6fd121),
	.w7(32'h3a2b4b72),
	.w8(32'h39fa4079),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398169e7),
	.w1(32'h399dc8d3),
	.w2(32'h3a0bd3ab),
	.w3(32'h3a35e8e6),
	.w4(32'h3a328a8b),
	.w5(32'h39a8db81),
	.w6(32'h399dd902),
	.w7(32'h37c8f339),
	.w8(32'hb6bc29c4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a38c4),
	.w1(32'h39cc75b8),
	.w2(32'h39dc79f9),
	.w3(32'h3a0eb612),
	.w4(32'h3a0fb8aa),
	.w5(32'h3a1945ab),
	.w6(32'h3a043561),
	.w7(32'h39e7b34b),
	.w8(32'h39bea8ea),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39652bef),
	.w1(32'h3a204d6b),
	.w2(32'h39cbc914),
	.w3(32'h39d7fe77),
	.w4(32'h3a3a0d06),
	.w5(32'h3a1064d2),
	.w6(32'h37889346),
	.w7(32'hb8885c2e),
	.w8(32'h391c9525),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943e8a0),
	.w1(32'hba96d07b),
	.w2(32'hb9fd414c),
	.w3(32'hb8891a21),
	.w4(32'hbaaea106),
	.w5(32'hbaa7524b),
	.w6(32'hba347e8b),
	.w7(32'hb9c30484),
	.w8(32'hb7bec2fa),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79fec37),
	.w1(32'h3911e187),
	.w2(32'hb8ac48a9),
	.w3(32'hba3eeb40),
	.w4(32'h3a403a48),
	.w5(32'h3a08314e),
	.w6(32'h37f4cf9e),
	.w7(32'hb98bc0cf),
	.w8(32'h38cb8405),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ff9c0f),
	.w1(32'h39a2da89),
	.w2(32'h39cb6833),
	.w3(32'h39a9cbfa),
	.w4(32'h39d1ff8e),
	.w5(32'h3a02fc40),
	.w6(32'h3a02c3fc),
	.w7(32'h39d115df),
	.w8(32'h39c4b2ee),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b788f),
	.w1(32'hb8ad6f99),
	.w2(32'h3944807e),
	.w3(32'h39d20d31),
	.w4(32'hb996f97f),
	.w5(32'hba41feb3),
	.w6(32'h3991ee64),
	.w7(32'h3a4bedd6),
	.w8(32'hb96bded3),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a058afb),
	.w1(32'h3a04e817),
	.w2(32'h39a0a380),
	.w3(32'h382a1bcb),
	.w4(32'h3a6f6c0d),
	.w5(32'h3a25de09),
	.w6(32'hb544efe9),
	.w7(32'h372f9bd4),
	.w8(32'hb78cde9a),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e723d),
	.w1(32'h3b211696),
	.w2(32'h3b036634),
	.w3(32'h393e98b3),
	.w4(32'h3b5e0468),
	.w5(32'h3ac96361),
	.w6(32'h3a6c5674),
	.w7(32'h3aeff2ac),
	.w8(32'h3b0c3672),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb9b3d),
	.w1(32'h3a1da375),
	.w2(32'h39d3b180),
	.w3(32'h39b0878a),
	.w4(32'h3aac6a41),
	.w5(32'h3a9db688),
	.w6(32'h39887c6b),
	.w7(32'h39423ba0),
	.w8(32'h399c57ed),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a41ef7),
	.w1(32'hba5eafae),
	.w2(32'hba3b0663),
	.w3(32'h39f86a37),
	.w4(32'hba964dc6),
	.w5(32'hba4eafa6),
	.w6(32'hba744aae),
	.w7(32'hb93baee4),
	.w8(32'hb82ff643),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac71d3),
	.w1(32'h399f2003),
	.w2(32'hba1d1471),
	.w3(32'hba1f06a4),
	.w4(32'h3a6a731a),
	.w5(32'hb95c4ca8),
	.w6(32'hba552554),
	.w7(32'hbabaf78b),
	.w8(32'hba81dbd4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2e21),
	.w1(32'h3a0d24eb),
	.w2(32'h3a171c64),
	.w3(32'hba89b567),
	.w4(32'h3a3cafc9),
	.w5(32'h3a4e4015),
	.w6(32'h3a442173),
	.w7(32'h3a26a0bc),
	.w8(32'h3a0cf26f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398335a1),
	.w1(32'h39a1477d),
	.w2(32'h3a420a34),
	.w3(32'h3a0ad6e0),
	.w4(32'h39a5fbda),
	.w5(32'h3a0ff6f2),
	.w6(32'h39de853b),
	.w7(32'h3a150f19),
	.w8(32'h3a3e6dd5),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e250c0),
	.w1(32'h3a00049d),
	.w2(32'h3a33626a),
	.w3(32'h3a041e35),
	.w4(32'h3a2b6970),
	.w5(32'h3a4d6408),
	.w6(32'h3a0490cd),
	.w7(32'h39f3cc33),
	.w8(32'h3a10ed1e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38239b4c),
	.w1(32'hb9b3f8fb),
	.w2(32'h3999165a),
	.w3(32'h39bbad3f),
	.w4(32'h3a998e41),
	.w5(32'h3acaf23c),
	.w6(32'hba03c084),
	.w7(32'hb9c6764c),
	.w8(32'hba3281f2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9babb11),
	.w1(32'hba5859f3),
	.w2(32'hb96e6dba),
	.w3(32'h389d3433),
	.w4(32'hba62fd1d),
	.w5(32'hb89e080e),
	.w6(32'hba121ab6),
	.w7(32'hba097629),
	.w8(32'hb981ef68),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ae558),
	.w1(32'h3905616d),
	.w2(32'hb98c43e7),
	.w3(32'h3a60a4ce),
	.w4(32'h3a9213d7),
	.w5(32'h37c8741f),
	.w6(32'hb98dc3ab),
	.w7(32'hba93c345),
	.w8(32'hba800f61),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33f01c),
	.w1(32'hb7be71da),
	.w2(32'hba2540dd),
	.w3(32'hb81d6d71),
	.w4(32'h3a04a106),
	.w5(32'h39a9653e),
	.w6(32'hba13d4a4),
	.w7(32'hba120025),
	.w8(32'hb7346b49),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb299f),
	.w1(32'h39a1b03e),
	.w2(32'h39e6668d),
	.w3(32'h3957dc81),
	.w4(32'h39cf765e),
	.w5(32'h39bd807f),
	.w6(32'h39b77110),
	.w7(32'h39f05071),
	.w8(32'h3a17a046),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c625a5),
	.w1(32'hb88c6843),
	.w2(32'hb948698c),
	.w3(32'h39b7f49a),
	.w4(32'h39f579d9),
	.w5(32'h3a6b9b02),
	.w6(32'h3a1017bd),
	.w7(32'h3a162245),
	.w8(32'h3a1d4cdc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a210c92),
	.w1(32'h3a2c68f3),
	.w2(32'h3a3b39af),
	.w3(32'h3aabd594),
	.w4(32'h3ad6aebf),
	.w5(32'h3ab4f638),
	.w6(32'h38e14650),
	.w7(32'hb9afc357),
	.w8(32'h39539098),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a5452),
	.w1(32'hb963e1ff),
	.w2(32'hb980aabf),
	.w3(32'h3ab9c7da),
	.w4(32'h3a2fb507),
	.w5(32'h39cd9ad8),
	.w6(32'hba1a27c3),
	.w7(32'hb9f28228),
	.w8(32'h39371b47),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35aa88b1),
	.w1(32'hbaa3346e),
	.w2(32'h39c30251),
	.w3(32'h39dd3e75),
	.w4(32'hba7ba4e7),
	.w5(32'h38ebd0d8),
	.w6(32'h3aa80d49),
	.w7(32'hba915cda),
	.w8(32'hba1b6db0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533eb0),
	.w1(32'hba1d7946),
	.w2(32'hb99c7637),
	.w3(32'h39cf7f5f),
	.w4(32'hba0de5fe),
	.w5(32'hba2f6b2c),
	.w6(32'h3ac817ea),
	.w7(32'h3aa3f8fe),
	.w8(32'h3ab0d1e9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule