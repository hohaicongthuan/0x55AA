module layer_10_featuremap_364(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd49d26a),
	.w1(32'h3d594358),
	.w2(32'hbdda5f3e),
	.w3(32'hbdeecefb),
	.w4(32'h3e04fa99),
	.w5(32'hbe149c74),
	.w6(32'h3d81af20),
	.w7(32'hbd8f65ba),
	.w8(32'hbed9856f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7791ba),
	.w1(32'hbcf71094),
	.w2(32'hbe4ab5b8),
	.w3(32'h3d3b34e3),
	.w4(32'h3d103d8e),
	.w5(32'hbcd0cde7),
	.w6(32'hbe23d329),
	.w7(32'hbe16bb01),
	.w8(32'hbdda7ac5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb39508),
	.w1(32'hbca88bd8),
	.w2(32'hbdc4287c),
	.w3(32'hbe0cc8e4),
	.w4(32'hbd242a05),
	.w5(32'hbd4e09f1),
	.w6(32'hbe8132bf),
	.w7(32'hbe552feb),
	.w8(32'hbe220fd1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdf9d947),
	.w1(32'hbe2f2af5),
	.w2(32'hbdad2445),
	.w3(32'hbf07c57d),
	.w4(32'hbe6cf5e4),
	.w5(32'hbec50924),
	.w6(32'hbd0bda7b),
	.w7(32'hbef311ca),
	.w8(32'h3d9cc150),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd18691),
	.w1(32'hbd15709c),
	.w2(32'h3b86f210),
	.w3(32'hbe2ba375),
	.w4(32'hbe939874),
	.w5(32'hbd0bcd3e),
	.w6(32'h3dcb9d92),
	.w7(32'h3e24860e),
	.w8(32'hbdc72d80),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec3e82d),
	.w1(32'hbd99a674),
	.w2(32'hbeecd9f8),
	.w3(32'hbe288037),
	.w4(32'hbcef1116),
	.w5(32'hbe666c03),
	.w6(32'h3dbbe8da),
	.w7(32'hbf1d7050),
	.w8(32'h3d1e502c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18b551),
	.w1(32'hbd98c3e9),
	.w2(32'hbd512636),
	.w3(32'hbe7f1b01),
	.w4(32'hbda7f0a6),
	.w5(32'hbe0da310),
	.w6(32'hbe80772c),
	.w7(32'h3cbc9b54),
	.w8(32'hbe040eee),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39c476),
	.w1(32'h3c39ac97),
	.w2(32'hbe63bfb9),
	.w3(32'hbdc81604),
	.w4(32'hbe0c5f2b),
	.w5(32'h3c897cda),
	.w6(32'hbd92f461),
	.w7(32'hbe7340bf),
	.w8(32'hbda37da1),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd96e58d),
	.w1(32'h3d9794f3),
	.w2(32'hbe05c2c1),
	.w3(32'h3b9c12f6),
	.w4(32'hbe8faed8),
	.w5(32'h3e89d1a2),
	.w6(32'hbf01733f),
	.w7(32'hbf0d57d4),
	.w8(32'h3ce161a2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dda861e),
	.w1(32'h3b21d156),
	.w2(32'hbdc26563),
	.w3(32'hbdcedaa8),
	.w4(32'hbe51661f),
	.w5(32'hbe3503d7),
	.w6(32'hbee6e85d),
	.w7(32'hbde22da7),
	.w8(32'hbd91c2ba),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda54e07),
	.w1(32'hbdd694e1),
	.w2(32'hbe007e5c),
	.w3(32'hbf1413a4),
	.w4(32'hbe24600d),
	.w5(32'h3b7040bd),
	.w6(32'hbf322d78),
	.w7(32'hbe128c53),
	.w8(32'hbef72410),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f9983),
	.w1(32'hbd6dbb92),
	.w2(32'hbdfea871),
	.w3(32'hbd157c45),
	.w4(32'hbe463c21),
	.w5(32'hbdf48a52),
	.w6(32'h3ef3a2b3),
	.w7(32'hbd943995),
	.w8(32'hbeb76925),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d835a17),
	.w1(32'h3dd2c0f5),
	.w2(32'h3d2b6330),
	.w3(32'h3be0ee90),
	.w4(32'h3ccdc395),
	.w5(32'h3d00ceb2),
	.w6(32'hbec13a49),
	.w7(32'h3cb08d7d),
	.w8(32'h3cbacec2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d121e2f),
	.w1(32'h3d995639),
	.w2(32'h3db15b56),
	.w3(32'h3cb17aeb),
	.w4(32'h3d020eb5),
	.w5(32'h3c85bee9),
	.w6(32'h3cf4d0ad),
	.w7(32'h3c9e0e66),
	.w8(32'h3ce148e0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad295c),
	.w1(32'h3d455cd3),
	.w2(32'h3cad3edf),
	.w3(32'h3ccc175c),
	.w4(32'h3d38900d),
	.w5(32'h3ca1e97c),
	.w6(32'h3cdef683),
	.w7(32'h3c89cdda),
	.w8(32'h3cf05e45),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d050cb1),
	.w1(32'h3d864c99),
	.w2(32'h3cf711c2),
	.w3(32'h3d0b428f),
	.w4(32'h3cf47e38),
	.w5(32'h3ce4b374),
	.w6(32'h3cfe8e80),
	.w7(32'h3d007c1a),
	.w8(32'h3cf1c122),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccab5c1),
	.w1(32'h3d4caef5),
	.w2(32'h3c9d387d),
	.w3(32'h3d29d1ae),
	.w4(32'h3bf0b797),
	.w5(32'h3cd9349c),
	.w6(32'h3d3ffdf8),
	.w7(32'h3c9af359),
	.w8(32'h3d4be4fa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95d5e3),
	.w1(32'h3d166a4f),
	.w2(32'h3ca368c6),
	.w3(32'h3c859fe9),
	.w4(32'h3cc8bcc8),
	.w5(32'h3d1454a4),
	.w6(32'h3cd3e774),
	.w7(32'h3c5f2a24),
	.w8(32'h3d0048b2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d789c41),
	.w1(32'h3d2c9cbf),
	.w2(32'h3cf89597),
	.w3(32'h3ca457dd),
	.w4(32'h3d12d4dd),
	.w5(32'h3d510c6c),
	.w6(32'h3cbcabbd),
	.w7(32'h3d4c7387),
	.w8(32'h3c7586e5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc39c5),
	.w1(32'h3d27630d),
	.w2(32'h3cd22fc2),
	.w3(32'h3ca3e38e),
	.w4(32'h3c6ec67c),
	.w5(32'h3d42a863),
	.w6(32'h3d3f5194),
	.w7(32'h3c96e755),
	.w8(32'h3d9987b6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce75860),
	.w1(32'h3d7c50d2),
	.w2(32'h3c5018d3),
	.w3(32'h3c1b937a),
	.w4(32'h3d141f6f),
	.w5(32'h3cacfbca),
	.w6(32'h3cab1685),
	.w7(32'h3d07cc92),
	.w8(32'h3cf440fb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8fa77),
	.w1(32'h3cd3a139),
	.w2(32'h3d097d25),
	.w3(32'h3ce1e60d),
	.w4(32'h3cab6cc3),
	.w5(32'h3d09fc27),
	.w6(32'h3cd382a4),
	.w7(32'h3cabd1d6),
	.w8(32'h3cbaa9fa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab4a42),
	.w1(32'h3cc5b596),
	.w2(32'h3c931e2a),
	.w3(32'h3cf1becd),
	.w4(32'h3d4cf5dd),
	.w5(32'h3d51778c),
	.w6(32'h3cd84dd1),
	.w7(32'h3ceb26d0),
	.w8(32'h3cb826b5),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f4a75),
	.w1(32'h3ccc4560),
	.w2(32'h3cee0060),
	.w3(32'h3d01cc87),
	.w4(32'h3d26bd85),
	.w5(32'h3cb7bc25),
	.w6(32'h3d101738),
	.w7(32'h3cc9ba5c),
	.w8(32'h3c767184),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bdb1c),
	.w1(32'h3d32da1c),
	.w2(32'h3cd00663),
	.w3(32'h3d1ca865),
	.w4(32'h3d740632),
	.w5(32'h3cbfea89),
	.w6(32'h3c94941d),
	.w7(32'h3c6114e1),
	.w8(32'h3d0bfd33),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0114cb),
	.w1(32'h3c98aaa2),
	.w2(32'h3cae443a),
	.w3(32'h3d290d52),
	.w4(32'h3cdd7f18),
	.w5(32'h3c8f9648),
	.w6(32'h3cbdb704),
	.w7(32'h3cfd8800),
	.w8(32'h3d179b18),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8deefa),
	.w1(32'h3cd3a4df),
	.w2(32'h3b2e0a22),
	.w3(32'h3cb898cf),
	.w4(32'h3cf09f1e),
	.w5(32'h398ebeab),
	.w6(32'h3cf5f791),
	.w7(32'h3cc77532),
	.w8(32'hbb4002ff),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ef68d),
	.w1(32'h3cb73823),
	.w2(32'hbc11a552),
	.w3(32'hbbc65dcf),
	.w4(32'hbc1423aa),
	.w5(32'h3b842960),
	.w6(32'hbad517b2),
	.w7(32'hbc5475c5),
	.w8(32'h3ac8e0a2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917d70),
	.w1(32'hbc348d43),
	.w2(32'hbbd2b3d8),
	.w3(32'hbbfef625),
	.w4(32'h3bbca719),
	.w5(32'hbba69360),
	.w6(32'h3c87cb65),
	.w7(32'hbb40afcd),
	.w8(32'h3c818d03),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76d64b),
	.w1(32'hbb76bce6),
	.w2(32'hbc2801a8),
	.w3(32'hbaccdadc),
	.w4(32'h3bbb363a),
	.w5(32'h398843a2),
	.w6(32'h3bc634ad),
	.w7(32'hbb44cd09),
	.w8(32'hbaa5cbac),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53c671),
	.w1(32'h3be8c045),
	.w2(32'h3b765717),
	.w3(32'hbc385955),
	.w4(32'h3bea17af),
	.w5(32'h3c536362),
	.w6(32'hbabf90b4),
	.w7(32'h3b966f8b),
	.w8(32'hbc8e1577),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ee63),
	.w1(32'h3c728a42),
	.w2(32'hbbe9235f),
	.w3(32'h3c3b4e2e),
	.w4(32'hbc144d58),
	.w5(32'h3b049e36),
	.w6(32'h3c1ef4a4),
	.w7(32'h3b28d5f8),
	.w8(32'hbc4890f5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3b9a),
	.w1(32'h3b6f7bd5),
	.w2(32'h3c8ea3dc),
	.w3(32'hbc395639),
	.w4(32'h3b856d5d),
	.w5(32'h3bd73601),
	.w6(32'hbc4ae9e7),
	.w7(32'h3c5e49c5),
	.w8(32'hbc2bbe24),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f20ed),
	.w1(32'hb84d553b),
	.w2(32'h3ba930b7),
	.w3(32'hba47b4d0),
	.w4(32'hbb8ea90c),
	.w5(32'h3ae0ca13),
	.w6(32'h3b15cb9b),
	.w7(32'h3ba1b3db),
	.w8(32'hba677425),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf5c68),
	.w1(32'h3c530bc6),
	.w2(32'h3ca88365),
	.w3(32'hbbdb3441),
	.w4(32'h3aa5de5c),
	.w5(32'hbbf6c258),
	.w6(32'h3cc4b512),
	.w7(32'hba62bfdb),
	.w8(32'hb83c77d6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e3c8),
	.w1(32'hbc610b75),
	.w2(32'hbc8e52cf),
	.w3(32'h3c5e80fd),
	.w4(32'h3a99c802),
	.w5(32'h3b40a381),
	.w6(32'hb93fdaf3),
	.w7(32'h3cc69e7e),
	.w8(32'h3b9f1e48),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1af930),
	.w1(32'h3bba6256),
	.w2(32'hb924c86d),
	.w3(32'hbae67007),
	.w4(32'h39a0df18),
	.w5(32'hbbc11923),
	.w6(32'hbb35e56c),
	.w7(32'hbb25e390),
	.w8(32'hbb786cd2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0017d7),
	.w1(32'hba226d88),
	.w2(32'h3c556108),
	.w3(32'hbc2de918),
	.w4(32'hbb8f7a3c),
	.w5(32'h3963ec3b),
	.w6(32'hbc4ee0b3),
	.w7(32'hbbf084b5),
	.w8(32'h3b831f31),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc0a0a),
	.w1(32'h3c91ba0c),
	.w2(32'hbc46a195),
	.w3(32'hbc699461),
	.w4(32'h3c9549d7),
	.w5(32'h3a94b874),
	.w6(32'h3c4f8569),
	.w7(32'hbc72d1f8),
	.w8(32'hbc93f3ad),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0af3b0),
	.w1(32'hbc63a8c1),
	.w2(32'h3b51dbb6),
	.w3(32'hb8df0e51),
	.w4(32'h3c24272c),
	.w5(32'hbb40dc6b),
	.w6(32'h3cadadd9),
	.w7(32'hbba583c3),
	.w8(32'h3b14421a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7041f),
	.w1(32'hbc69a7e8),
	.w2(32'h3b849721),
	.w3(32'hbb377cb6),
	.w4(32'hbc14b8c9),
	.w5(32'h3bb74114),
	.w6(32'h3acc4d2b),
	.w7(32'hba207c40),
	.w8(32'h3b663cb0),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62f5ca),
	.w1(32'hbc32d646),
	.w2(32'h3c9ba77f),
	.w3(32'hbc23830a),
	.w4(32'hbc4db578),
	.w5(32'h3b694594),
	.w6(32'h3c1a84db),
	.w7(32'h3b490ce1),
	.w8(32'hbb07cc42),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc701ba8),
	.w1(32'h3bec5597),
	.w2(32'hbb69d6ed),
	.w3(32'h3cb6a0b4),
	.w4(32'hbc3748bb),
	.w5(32'hbc5556fd),
	.w6(32'h3caba0ff),
	.w7(32'h3c48c791),
	.w8(32'h3b0bf022),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cb35a),
	.w1(32'h3aefd74e),
	.w2(32'hbc5c77b0),
	.w3(32'h3c07d14a),
	.w4(32'hba6c606a),
	.w5(32'h3be7eb59),
	.w6(32'hbc316d7e),
	.w7(32'hbbaebe07),
	.w8(32'hba58de6e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc3a0c),
	.w1(32'h3b0d4f39),
	.w2(32'h3b4932b6),
	.w3(32'h399993a0),
	.w4(32'h3b0e762c),
	.w5(32'hbbaec794),
	.w6(32'hbb996e42),
	.w7(32'hbb2551a5),
	.w8(32'h39a78608),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9611),
	.w1(32'hbb8efd6b),
	.w2(32'hbcd566f5),
	.w3(32'h3bb474fa),
	.w4(32'h3c238055),
	.w5(32'hbc5f6767),
	.w6(32'h3aea3a83),
	.w7(32'h3ca449d8),
	.w8(32'h3bf4460b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b549c),
	.w1(32'h3c5f98b9),
	.w2(32'h3bb03f4d),
	.w3(32'hbb53bd71),
	.w4(32'h3aef45a0),
	.w5(32'h3a53c0b7),
	.w6(32'h3b6020c7),
	.w7(32'h3bc2bf34),
	.w8(32'h3ba17850),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87d4d0),
	.w1(32'h3c06dc16),
	.w2(32'hbc5bf576),
	.w3(32'h3d0eeba4),
	.w4(32'h3b0f8e18),
	.w5(32'hb8e42cdf),
	.w6(32'h3c7cf505),
	.w7(32'h3ad0cb28),
	.w8(32'h3b3b95a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd3fcc),
	.w1(32'hbb8ca2c6),
	.w2(32'hbad6924b),
	.w3(32'h3b66260a),
	.w4(32'h3bac1e48),
	.w5(32'h3b86abfa),
	.w6(32'h3b87a332),
	.w7(32'h3c5e9633),
	.w8(32'hbbb9f7cb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bac76),
	.w1(32'hb952dc7f),
	.w2(32'hbcb87c01),
	.w3(32'hbca1f9cf),
	.w4(32'hbbb05983),
	.w5(32'h3b843a4a),
	.w6(32'hbbcc2c52),
	.w7(32'h3b1cb514),
	.w8(32'hbb43aed4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ebad53),
	.w1(32'h3b75d856),
	.w2(32'h3b20cd98),
	.w3(32'hbbad9df6),
	.w4(32'hbaf6f41a),
	.w5(32'hba53985d),
	.w6(32'hbaedd1a6),
	.w7(32'h3b5a8bfb),
	.w8(32'h3c5e8ce3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc924072),
	.w1(32'hbbe8a83e),
	.w2(32'hbc373b54),
	.w3(32'hba7e5002),
	.w4(32'h3c576e7f),
	.w5(32'h3c1a4639),
	.w6(32'h3a891f81),
	.w7(32'h3bfedc64),
	.w8(32'hbc19ac60),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6ed46),
	.w1(32'hbbf6fd4c),
	.w2(32'hbc02b4ac),
	.w3(32'hbbf8bd53),
	.w4(32'h3bad7d6a),
	.w5(32'h3be49252),
	.w6(32'hbb5cb18f),
	.w7(32'h3c130788),
	.w8(32'hbb28304a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51a50d),
	.w1(32'h3b2a7d31),
	.w2(32'hbbdb4fc6),
	.w3(32'hbbc4d574),
	.w4(32'h3bb59b51),
	.w5(32'h3b9d81c3),
	.w6(32'hb9171653),
	.w7(32'hbc0ec8c2),
	.w8(32'hbbb1ecaf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53a3a5),
	.w1(32'h3cafddab),
	.w2(32'hb99d2da9),
	.w3(32'hbc0927ef),
	.w4(32'h3caaf42f),
	.w5(32'hbc1bccf3),
	.w6(32'hbba93e30),
	.w7(32'hbb7ae540),
	.w8(32'hbb0dd11e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ca196),
	.w1(32'hbb5ece63),
	.w2(32'h3b03ce0d),
	.w3(32'h3c1662b2),
	.w4(32'hbace4e8d),
	.w5(32'hbc2dcc4e),
	.w6(32'h3bb70291),
	.w7(32'hbc69a370),
	.w8(32'h3ac73342),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e738cf),
	.w1(32'h3ac38668),
	.w2(32'hbb8caa5a),
	.w3(32'hba53988e),
	.w4(32'h3b60c59c),
	.w5(32'h3b6b54e5),
	.w6(32'hbb1447ac),
	.w7(32'hbc3f74ae),
	.w8(32'h3a9509a8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67db18),
	.w1(32'h3c944061),
	.w2(32'hbc99f930),
	.w3(32'hbc3b0287),
	.w4(32'hbb5915a4),
	.w5(32'h3a73df5e),
	.w6(32'hbbc79d68),
	.w7(32'hba60c3ff),
	.w8(32'h3c2cb2a0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5e22),
	.w1(32'h3b23a8b8),
	.w2(32'h3ab41cfb),
	.w3(32'hbbdadcb8),
	.w4(32'h3bc9cdb6),
	.w5(32'hbc07c85e),
	.w6(32'h3a31c693),
	.w7(32'hbc67410a),
	.w8(32'hbbfd7c48),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab0dde),
	.w1(32'hbc116474),
	.w2(32'hba46b587),
	.w3(32'hbc9437dd),
	.w4(32'h3bab9624),
	.w5(32'hbab4d9b8),
	.w6(32'hbc4a3e7f),
	.w7(32'hbc596545),
	.w8(32'hbc759ced),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdaf74c),
	.w1(32'hba646bd3),
	.w2(32'h3a7d0f41),
	.w3(32'h3c8b7a56),
	.w4(32'h3b43cbaf),
	.w5(32'hbba2199a),
	.w6(32'hbc8e3f82),
	.w7(32'h3add741c),
	.w8(32'hbb09f523),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c866f),
	.w1(32'hbc45406c),
	.w2(32'hbad8320d),
	.w3(32'h3c1e865b),
	.w4(32'hbb4a214a),
	.w5(32'hbc4eb5c1),
	.w6(32'h3bb55192),
	.w7(32'hbb5b0042),
	.w8(32'h3bfafc77),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efd76),
	.w1(32'h3bb93c6c),
	.w2(32'hbbc422b5),
	.w3(32'hbb81d6ea),
	.w4(32'hbc7fbc86),
	.w5(32'hbb010949),
	.w6(32'hbc19f865),
	.w7(32'hba7f3b84),
	.w8(32'h3aedb595),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca53252),
	.w1(32'h3bb6639c),
	.w2(32'hbc14e5c3),
	.w3(32'hbc374c04),
	.w4(32'h3b2039a3),
	.w5(32'hbc27fa74),
	.w6(32'h3b07c661),
	.w7(32'hbc60594b),
	.w8(32'h3bf27645),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa6eef),
	.w1(32'hba6ac8f8),
	.w2(32'h3a82ab72),
	.w3(32'h3ba23139),
	.w4(32'hbaf2c74b),
	.w5(32'h3c06cc62),
	.w6(32'h3b6783f5),
	.w7(32'h3b14b5ea),
	.w8(32'h3bb7e071),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e2ad),
	.w1(32'h3b1189bc),
	.w2(32'h3b0b44cc),
	.w3(32'h3c7f6136),
	.w4(32'h3b5f73e7),
	.w5(32'hbb897121),
	.w6(32'h3be6a478),
	.w7(32'hbc4ea57d),
	.w8(32'hbb94696e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05cc6b),
	.w1(32'h3b3afe37),
	.w2(32'hba0d34a2),
	.w3(32'h3ba9f5c0),
	.w4(32'hbac4a1f8),
	.w5(32'h3c71fa6d),
	.w6(32'hbaf9fc1b),
	.w7(32'hbce55b18),
	.w8(32'hbb8378ad),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e3227),
	.w1(32'hb9ea7a3d),
	.w2(32'hbc900a7d),
	.w3(32'hbc080e83),
	.w4(32'hbbf44d44),
	.w5(32'h3bd0833c),
	.w6(32'hbc569dfc),
	.w7(32'h3b46a398),
	.w8(32'h3c50edbc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb432dc4),
	.w1(32'h3c7a8f71),
	.w2(32'hbaca6231),
	.w3(32'h3b5e8335),
	.w4(32'hb96d2634),
	.w5(32'h39be80a6),
	.w6(32'hbb694df2),
	.w7(32'hbc94ca07),
	.w8(32'h3d0edd5c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0dc4b),
	.w1(32'h3c0b9e83),
	.w2(32'h3bfcac9f),
	.w3(32'hbc6facb4),
	.w4(32'hbaff0b77),
	.w5(32'hbbc66528),
	.w6(32'hbac99548),
	.w7(32'h3bb8317c),
	.w8(32'h3c48180d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb749d8),
	.w1(32'h3c6d10ae),
	.w2(32'hbc07913e),
	.w3(32'hbd3f768f),
	.w4(32'h3a8f579a),
	.w5(32'h3bef2cc6),
	.w6(32'hbc2a93e9),
	.w7(32'hb9123dfc),
	.w8(32'hb8c56b72),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d7543),
	.w1(32'hbc7729f3),
	.w2(32'hbba6d7ff),
	.w3(32'h3c46a46a),
	.w4(32'h3b6417ba),
	.w5(32'h3a5ebcb0),
	.w6(32'hbb95f173),
	.w7(32'h3b6a9645),
	.w8(32'h3b91aab6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8432dd),
	.w1(32'hba2e27e8),
	.w2(32'hbb06d4fa),
	.w3(32'hbc15e7a5),
	.w4(32'hbc45480c),
	.w5(32'h3b866918),
	.w6(32'hbaaed630),
	.w7(32'h3c1bf5e9),
	.w8(32'hbb62579f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809194),
	.w1(32'hb9c5578b),
	.w2(32'h3ba40cd9),
	.w3(32'hbbb2443c),
	.w4(32'hbb9320c4),
	.w5(32'h3b191de3),
	.w6(32'h3c3ad8e7),
	.w7(32'hb908d627),
	.w8(32'h3c02c5d3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37e41c),
	.w1(32'h3c5871dd),
	.w2(32'hbb4c9225),
	.w3(32'hbb7d3081),
	.w4(32'h3c498ba4),
	.w5(32'h3ba88914),
	.w6(32'h3bbd2531),
	.w7(32'h3be43d17),
	.w8(32'h3ac04e41),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2b00),
	.w1(32'hb8bd88d4),
	.w2(32'h3ccbaad5),
	.w3(32'h3badf283),
	.w4(32'h3bdb2408),
	.w5(32'hbc1e0056),
	.w6(32'h3c1d3bd4),
	.w7(32'h3ba91ed2),
	.w8(32'hbbb8e3aa),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3651a7),
	.w1(32'h3a3be2f5),
	.w2(32'h3ad46153),
	.w3(32'hba9ab36b),
	.w4(32'h3b8ff920),
	.w5(32'hbc6dbb2f),
	.w6(32'h3b4b3b06),
	.w7(32'h3aae7492),
	.w8(32'hbbd3d1dc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b1a6e),
	.w1(32'h3bf003e7),
	.w2(32'h3b924d91),
	.w3(32'h3bada788),
	.w4(32'hbb1ce3de),
	.w5(32'hbc0521ea),
	.w6(32'hbc44c0f2),
	.w7(32'hbbce97b4),
	.w8(32'h3c4b4bc3),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba88d89),
	.w1(32'hba1a9c83),
	.w2(32'hbb2b93de),
	.w3(32'hbc634633),
	.w4(32'hba11adba),
	.w5(32'h3ab41a22),
	.w6(32'hbb2b341a),
	.w7(32'hbc754560),
	.w8(32'hbb5e7513),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2b103),
	.w1(32'h3a9a0e34),
	.w2(32'hbc6e5c94),
	.w3(32'hbad4b3a7),
	.w4(32'h3ab41d4c),
	.w5(32'h3bd857c1),
	.w6(32'hb850a314),
	.w7(32'hba9a9859),
	.w8(32'hbb53f3c2),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2afc1),
	.w1(32'hbbd11059),
	.w2(32'hbb6c3fd2),
	.w3(32'hbaf2169a),
	.w4(32'hbb0a7b6b),
	.w5(32'h3a7f5937),
	.w6(32'h3b82ed2f),
	.w7(32'hba6ba419),
	.w8(32'h3b8068a1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319736),
	.w1(32'h3d0c9205),
	.w2(32'hbbb739ee),
	.w3(32'h3c2958c0),
	.w4(32'hbbc1b272),
	.w5(32'h3c7bb1e8),
	.w6(32'h3ad7cfb7),
	.w7(32'hbb8c87e7),
	.w8(32'hbab1fd69),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ddbcf),
	.w1(32'h3c0680bd),
	.w2(32'hbb9798fd),
	.w3(32'hbb560f23),
	.w4(32'hbad08905),
	.w5(32'h3af112c3),
	.w6(32'hba85f948),
	.w7(32'hbc06ea58),
	.w8(32'h3979ead1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3381b0),
	.w1(32'hbb0ac457),
	.w2(32'hbb1f193f),
	.w3(32'hbb0a40be),
	.w4(32'h3b4f868c),
	.w5(32'hbbfa6657),
	.w6(32'hbcce21d0),
	.w7(32'hbc8e3370),
	.w8(32'h3c015bca),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba70af6),
	.w1(32'hba5b0646),
	.w2(32'h3c0613a5),
	.w3(32'h3b335d73),
	.w4(32'h3b913562),
	.w5(32'hbbaf92ea),
	.w6(32'h395362b7),
	.w7(32'hbb430961),
	.w8(32'hbb956133),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab4557),
	.w1(32'hbc018fdf),
	.w2(32'hbbbeb800),
	.w3(32'hbb72e777),
	.w4(32'hbc04f209),
	.w5(32'h3b76b259),
	.w6(32'hbba41b6c),
	.w7(32'hbc00d2c8),
	.w8(32'hbbedc7da),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef6ce7),
	.w1(32'hbd3d1160),
	.w2(32'h3c244ba3),
	.w3(32'h3ca9d3e9),
	.w4(32'h3b4cdc85),
	.w5(32'h39a78ded),
	.w6(32'h3b9fdb90),
	.w7(32'hbbf3715b),
	.w8(32'hbb43e120),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169d5b),
	.w1(32'hbba40aca),
	.w2(32'h3a0274f2),
	.w3(32'hbb7858fe),
	.w4(32'h3ad1d334),
	.w5(32'h3cc510cc),
	.w6(32'hb91b5037),
	.w7(32'h3d5234b8),
	.w8(32'hb9b31557),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc33661),
	.w1(32'h3cb0f8df),
	.w2(32'h3b22f58a),
	.w3(32'h3b99ea38),
	.w4(32'h39ed4277),
	.w5(32'h3c76c4bb),
	.w6(32'hbae48699),
	.w7(32'hbb78bd01),
	.w8(32'h3c7932c1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3db62d),
	.w1(32'h3b7e4fbd),
	.w2(32'h3c15510c),
	.w3(32'h3b1e9183),
	.w4(32'hbc13a2cd),
	.w5(32'h3c287b0c),
	.w6(32'hbbed33e1),
	.w7(32'h3c4794ff),
	.w8(32'h3b89ebdd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4a271),
	.w1(32'h3be322dc),
	.w2(32'hbc31b2b4),
	.w3(32'hb8a50d21),
	.w4(32'h3b5ec54f),
	.w5(32'h3b6291c2),
	.w6(32'hbc4b55aa),
	.w7(32'hbb599098),
	.w8(32'hb8cdda15),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22acbc),
	.w1(32'hbbd221e7),
	.w2(32'h3c1327f3),
	.w3(32'h3c5c66e5),
	.w4(32'hbcd16540),
	.w5(32'h3bdd8678),
	.w6(32'h3c40b9b1),
	.w7(32'hbaf1cfe5),
	.w8(32'hbc186d3f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dd0a7),
	.w1(32'hbbabd790),
	.w2(32'hbc73a835),
	.w3(32'h3c5c1298),
	.w4(32'h3c8a3712),
	.w5(32'h39400ca7),
	.w6(32'hbc14864c),
	.w7(32'hbc691a0f),
	.w8(32'hbb637fc3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57a882),
	.w1(32'hbc417984),
	.w2(32'hbc322ecc),
	.w3(32'hbad953eb),
	.w4(32'h3b16d9c2),
	.w5(32'hbbd3954a),
	.w6(32'hbb3c5593),
	.w7(32'h35b7fc50),
	.w8(32'h3bda668b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c199a),
	.w1(32'hbd28fbce),
	.w2(32'hba6f9310),
	.w3(32'hbb33edae),
	.w4(32'hbc40fe39),
	.w5(32'hbb438ede),
	.w6(32'hbbb821d6),
	.w7(32'h3c570456),
	.w8(32'hbb2a55d0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c341947),
	.w1(32'h3ba6dd31),
	.w2(32'h3b4510b3),
	.w3(32'hbbaa0f27),
	.w4(32'hbb99fd0b),
	.w5(32'hbc99389b),
	.w6(32'h3c8531d7),
	.w7(32'h3cd09dba),
	.w8(32'h3b610ffa),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e076),
	.w1(32'h3bf1ba1e),
	.w2(32'hba81305d),
	.w3(32'h3cdc94a8),
	.w4(32'h3aac2097),
	.w5(32'hbd931901),
	.w6(32'h3bdaa66e),
	.w7(32'hbb856004),
	.w8(32'h38f8365e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd174d3a),
	.w1(32'hbcf48dba),
	.w2(32'h3bfea678),
	.w3(32'h3a959b71),
	.w4(32'hbb5cab4e),
	.w5(32'hbb6cdbac),
	.w6(32'h3bbb2bf2),
	.w7(32'h3bd9acb6),
	.w8(32'h3b29aaa0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b8a9),
	.w1(32'h3cd85ef2),
	.w2(32'hbd0d4be1),
	.w3(32'hbc5e8166),
	.w4(32'hbc3d8b2e),
	.w5(32'h3c9b9de0),
	.w6(32'hbbe811b7),
	.w7(32'h3d0c0266),
	.w8(32'h39d7abe7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc015844),
	.w1(32'h3b973ad7),
	.w2(32'hbba7c81b),
	.w3(32'hba9cd1a5),
	.w4(32'hbc1a0dc2),
	.w5(32'hbc357990),
	.w6(32'hbc346901),
	.w7(32'h3bd09227),
	.w8(32'hbacbc33b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8590a),
	.w1(32'h3b1e05bf),
	.w2(32'hba8487d3),
	.w3(32'h3b4e1f57),
	.w4(32'h3c187099),
	.w5(32'hb7dd81dd),
	.w6(32'h3b051c6a),
	.w7(32'hbb3f5766),
	.w8(32'h3abe9e7b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17f9ed),
	.w1(32'h3bae0fed),
	.w2(32'hbb2c63f5),
	.w3(32'hbadec899),
	.w4(32'hbbe2ffd5),
	.w5(32'h3a201ba0),
	.w6(32'h3c36b7d2),
	.w7(32'h3c2e5ae2),
	.w8(32'h3aea3749),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d4ac8),
	.w1(32'h3c9f5f9c),
	.w2(32'hbc253b4e),
	.w3(32'h3ad10758),
	.w4(32'hbc55526e),
	.w5(32'hba94f3bc),
	.w6(32'hbb4eb74e),
	.w7(32'h3c690f55),
	.w8(32'hbd64ea1a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05fa0d),
	.w1(32'h3c1cfc93),
	.w2(32'h3b18db89),
	.w3(32'h3b186a3d),
	.w4(32'h3c55ef62),
	.w5(32'hbbbcce2f),
	.w6(32'hbbfd493f),
	.w7(32'hbae52fde),
	.w8(32'h3b9f7e49),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b57da),
	.w1(32'h3ae66ac2),
	.w2(32'hbc0063cc),
	.w3(32'hbd2405b7),
	.w4(32'hbc0e51b4),
	.w5(32'h3cfa77dc),
	.w6(32'h3b316658),
	.w7(32'h3bbf776b),
	.w8(32'h3a5ad65e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c577841),
	.w1(32'hbaf5c01b),
	.w2(32'h3c35cf68),
	.w3(32'h3b869823),
	.w4(32'h3a8f516f),
	.w5(32'hbbe33a68),
	.w6(32'hbc51ec07),
	.w7(32'h3b335aec),
	.w8(32'hbc5c5a7c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19ca99),
	.w1(32'hbbafb284),
	.w2(32'h3d012aff),
	.w3(32'h3c406e72),
	.w4(32'h3a5769c6),
	.w5(32'h3b6ada1c),
	.w6(32'hbbd65c0e),
	.w7(32'hbc56db93),
	.w8(32'h3a474961),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8f2b3),
	.w1(32'h3b3bf3be),
	.w2(32'h3a812146),
	.w3(32'hbc112dfe),
	.w4(32'h3b70dfb1),
	.w5(32'h38714394),
	.w6(32'h39015173),
	.w7(32'h3b7f0b12),
	.w8(32'hbb5d023a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cb181),
	.w1(32'h3b85dd9f),
	.w2(32'hbb30bdb1),
	.w3(32'h3bb14f08),
	.w4(32'hbba30cbc),
	.w5(32'h3b042a9e),
	.w6(32'hbce157c6),
	.w7(32'hbbdb357d),
	.w8(32'h3a85827f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b4cf),
	.w1(32'hbc4b3ee9),
	.w2(32'h3a33bb1e),
	.w3(32'h39f44eac),
	.w4(32'hbaf42b6e),
	.w5(32'hbd3107ff),
	.w6(32'h3bdecb23),
	.w7(32'h38d320f5),
	.w8(32'hbb4a4a41),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40f449),
	.w1(32'h3a2afa10),
	.w2(32'hbc3c05fb),
	.w3(32'h3a258d7c),
	.w4(32'hbafb319b),
	.w5(32'hbbd5ebc5),
	.w6(32'hbacc315e),
	.w7(32'hbbdd5323),
	.w8(32'hbb385ac7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad57f0),
	.w1(32'hbaf9134f),
	.w2(32'hbb89be7c),
	.w3(32'hbb58bfa0),
	.w4(32'h3b4b5439),
	.w5(32'hbac18a03),
	.w6(32'h3c1a797b),
	.w7(32'hba66e1e4),
	.w8(32'hbc0dcdbc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18fbdb),
	.w1(32'h3a42a2b4),
	.w2(32'hbc0ebdc0),
	.w3(32'h39131f9a),
	.w4(32'h3c1d08a5),
	.w5(32'hbbba031d),
	.w6(32'hbbbd0ae0),
	.w7(32'h3ae3193a),
	.w8(32'h3a6af173),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc183f8),
	.w1(32'h3b3e4db1),
	.w2(32'hbba90dca),
	.w3(32'h3a124b96),
	.w4(32'hbabf5479),
	.w5(32'h3ad40c2b),
	.w6(32'hbb5de55f),
	.w7(32'h3b522aac),
	.w8(32'hbb824f71),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a805525),
	.w1(32'hbb31faf6),
	.w2(32'hbb8c4281),
	.w3(32'hba96cf87),
	.w4(32'hb98deebd),
	.w5(32'h3b039e53),
	.w6(32'hbc01c7e0),
	.w7(32'h3b10ee50),
	.w8(32'hbc08d37e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beadf9c),
	.w1(32'hbb976d4d),
	.w2(32'hbb00fcc2),
	.w3(32'hbb9a0319),
	.w4(32'h3b8c4600),
	.w5(32'h3b870362),
	.w6(32'hbc984e1c),
	.w7(32'hb689f6f4),
	.w8(32'h3c1c9461),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bfd1e),
	.w1(32'hbc21384e),
	.w2(32'hbc1475be),
	.w3(32'h3c23cad6),
	.w4(32'h3c7ff54e),
	.w5(32'h3cd5f8ed),
	.w6(32'h3b7146c3),
	.w7(32'h3b3201bc),
	.w8(32'hbc7e6c83),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf96f56),
	.w1(32'h3c74a5de),
	.w2(32'hba4ae80a),
	.w3(32'h3a07bc3c),
	.w4(32'hbbb2b573),
	.w5(32'h3bfc6ff7),
	.w6(32'hbc548552),
	.w7(32'hbbdd9a2c),
	.w8(32'hbb032510),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8fc80),
	.w1(32'hbba138be),
	.w2(32'h3c534cd5),
	.w3(32'h3b94b2e9),
	.w4(32'hbc206bb3),
	.w5(32'hbb742124),
	.w6(32'h3ccfacd7),
	.w7(32'h3b261ff9),
	.w8(32'h3bed19a2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80fea4a),
	.w1(32'hbc0eb0ac),
	.w2(32'h3cd1f841),
	.w3(32'h3d003948),
	.w4(32'hbc01a8e5),
	.w5(32'h3b94ecfd),
	.w6(32'h3b6662b0),
	.w7(32'hbbbe7000),
	.w8(32'hbc385e95),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb533f8),
	.w1(32'hbbd2e323),
	.w2(32'hbb93042f),
	.w3(32'h3c7aa8b0),
	.w4(32'h3d311e72),
	.w5(32'h3a94ab10),
	.w6(32'hbc5c524e),
	.w7(32'hba94d4c6),
	.w8(32'h3b8072b5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827da0),
	.w1(32'hbacebc2a),
	.w2(32'h3b47ade9),
	.w3(32'hbb567cbc),
	.w4(32'h3c28aaaf),
	.w5(32'h3b972e21),
	.w6(32'h3adda33e),
	.w7(32'hbb41b695),
	.w8(32'h3b5ab40e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c8a51),
	.w1(32'h3b9418a3),
	.w2(32'hba9a60dd),
	.w3(32'h3bf34e4a),
	.w4(32'h3cac1d6f),
	.w5(32'hb8e51897),
	.w6(32'hbb37d74b),
	.w7(32'hbbb598c5),
	.w8(32'h3cca57c2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5846fb),
	.w1(32'hbc55d366),
	.w2(32'h3aa8e11b),
	.w3(32'hbb0daa0c),
	.w4(32'hbd673a14),
	.w5(32'hbc523b28),
	.w6(32'hbbd96c8a),
	.w7(32'h3bb62c0b),
	.w8(32'hbb450726),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0dfbd6),
	.w1(32'hbadc295c),
	.w2(32'h3d80a725),
	.w3(32'h3cf3d502),
	.w4(32'h3b8804d2),
	.w5(32'h3bc960bf),
	.w6(32'hbb1b387f),
	.w7(32'hbc11a4c0),
	.w8(32'hbb8bfd10),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9084a),
	.w1(32'hba4ea2f0),
	.w2(32'hbc6d6f8b),
	.w3(32'h3b1532da),
	.w4(32'h3beee48f),
	.w5(32'h3cb3e81c),
	.w6(32'h3c00e5d8),
	.w7(32'h3bc5ab96),
	.w8(32'h3aa3480e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df2583),
	.w1(32'h39cd6e81),
	.w2(32'hbc315214),
	.w3(32'h3ca75a6b),
	.w4(32'hbc5d0c30),
	.w5(32'h3b04a544),
	.w6(32'h3912e3f4),
	.w7(32'hbc7bdb46),
	.w8(32'hbbccda3c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be745e7),
	.w1(32'hbc00c3ba),
	.w2(32'hba531493),
	.w3(32'h3c7b6152),
	.w4(32'h3b39aadc),
	.w5(32'hbbe3b63d),
	.w6(32'h3b8d0798),
	.w7(32'hbb144db8),
	.w8(32'hbbdf5605),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41cb83),
	.w1(32'hbc8e3cdb),
	.w2(32'hb9f58619),
	.w3(32'hbad6f88d),
	.w4(32'hbbc80c93),
	.w5(32'hbaff3c2e),
	.w6(32'h3ace62ec),
	.w7(32'h3aef8b69),
	.w8(32'hbc3d82c7),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cd270),
	.w1(32'hbb328c29),
	.w2(32'h3b136de6),
	.w3(32'hbb91cc15),
	.w4(32'hbb8b64ad),
	.w5(32'h3b47907f),
	.w6(32'hbbe78eef),
	.w7(32'hbb940b5c),
	.w8(32'h3ccfca5e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5ade7),
	.w1(32'hbb5305c7),
	.w2(32'hbbabca0f),
	.w3(32'h3bc395d6),
	.w4(32'hbc4fc8fe),
	.w5(32'h3c26147d),
	.w6(32'hba015cb0),
	.w7(32'hbc15962d),
	.w8(32'h3bc19415),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84ea1e),
	.w1(32'h3a9575b1),
	.w2(32'hba958801),
	.w3(32'h3b6d25f5),
	.w4(32'hbc829b91),
	.w5(32'h3bf920a7),
	.w6(32'hbc9ce96f),
	.w7(32'hb9d65a3e),
	.w8(32'h3c05e8f5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc787033),
	.w1(32'h3c24c04a),
	.w2(32'hba413920),
	.w3(32'h39c47c1b),
	.w4(32'hbbafae94),
	.w5(32'hbc0770a5),
	.w6(32'hbb46d3b3),
	.w7(32'h3b3b2fbf),
	.w8(32'hbbe4f59a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbf8ba),
	.w1(32'h3c3d1ca5),
	.w2(32'hbc03195f),
	.w3(32'hbac1f5c8),
	.w4(32'hba79da3d),
	.w5(32'h3bdb2638),
	.w6(32'hbc4efdd4),
	.w7(32'hbc35d8f3),
	.w8(32'h3ba53c38),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399be1f2),
	.w1(32'hba6db3c3),
	.w2(32'hbc246c32),
	.w3(32'hbc902615),
	.w4(32'hbc8ce78d),
	.w5(32'hbac8fa06),
	.w6(32'hba8111b0),
	.w7(32'h3c89f324),
	.w8(32'hbae01d99),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6d134),
	.w1(32'h3a98d04d),
	.w2(32'h3b2afc42),
	.w3(32'h3b28a7ee),
	.w4(32'hbc886b40),
	.w5(32'hbb9e9fa3),
	.w6(32'hbc3be6bf),
	.w7(32'hbc4d9988),
	.w8(32'hbbd62ab9),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56b718),
	.w1(32'hbbb1f442),
	.w2(32'h3bbda237),
	.w3(32'hb9c9a360),
	.w4(32'h3c518ec5),
	.w5(32'h3c20ec6a),
	.w6(32'h3c2c6eec),
	.w7(32'hbcca6a8b),
	.w8(32'hbbb72eb6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80e1bd),
	.w1(32'hbc8d9ced),
	.w2(32'h3c1b2333),
	.w3(32'hbc692d71),
	.w4(32'hbbada365),
	.w5(32'hba01d803),
	.w6(32'h3aa7e521),
	.w7(32'hbc364efe),
	.w8(32'hbcaebc4f),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba281d67),
	.w1(32'h3baeead2),
	.w2(32'h3c3c73a3),
	.w3(32'h3b820e2e),
	.w4(32'h3b8053d3),
	.w5(32'hb8f61fc3),
	.w6(32'hbc57abdf),
	.w7(32'hbb03e42c),
	.w8(32'h3b4e9bc2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc4968),
	.w1(32'h3c437aac),
	.w2(32'h3a0a7685),
	.w3(32'hba863f4b),
	.w4(32'h3b967602),
	.w5(32'hbc19805b),
	.w6(32'h3a9a84ad),
	.w7(32'h3b9985b2),
	.w8(32'h3bd1b4d3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb431d1e),
	.w1(32'hbc4fb8c1),
	.w2(32'hba6c253c),
	.w3(32'h3ae5faf6),
	.w4(32'hba77cee9),
	.w5(32'hbbb7c8e9),
	.w6(32'h3a9b3e53),
	.w7(32'hbb8e1223),
	.w8(32'hbb02bade),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b6f432),
	.w1(32'h3b9c7cba),
	.w2(32'h39807bc4),
	.w3(32'hbc2562a1),
	.w4(32'hbb20e82d),
	.w5(32'hba9aa076),
	.w6(32'h3a5e9c2a),
	.w7(32'hbb66a03f),
	.w8(32'hbc1fe713),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4509bd),
	.w1(32'hbbdcb7ca),
	.w2(32'h3b1186c3),
	.w3(32'hbba3498f),
	.w4(32'hbd1170bd),
	.w5(32'h3b9c35bc),
	.w6(32'hbc1ab597),
	.w7(32'hba72e3fe),
	.w8(32'h3c2f57d9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdda7f3),
	.w1(32'h3bc58dc5),
	.w2(32'h3ba0c372),
	.w3(32'h3be0cb10),
	.w4(32'hbb0e82ab),
	.w5(32'h3ab9380b),
	.w6(32'h3d022016),
	.w7(32'h3c46f1e8),
	.w8(32'hbcdc27e1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ff342),
	.w1(32'hbb19b8b6),
	.w2(32'hbab5f485),
	.w3(32'h3be79b6a),
	.w4(32'hbcd9327d),
	.w5(32'h3c3663c1),
	.w6(32'hbaf73d3f),
	.w7(32'hbb9081e5),
	.w8(32'h3bb509ea),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a6a58),
	.w1(32'hbb700d0c),
	.w2(32'h3ca8dbfc),
	.w3(32'hbc089c45),
	.w4(32'hbb6d9e4d),
	.w5(32'h39c6443e),
	.w6(32'h3b7191b4),
	.w7(32'h3b60666f),
	.w8(32'h3b4b483a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5a755),
	.w1(32'hbb8e1224),
	.w2(32'h3b8c6bdb),
	.w3(32'hbbdcaa42),
	.w4(32'h3ba53bbd),
	.w5(32'h3bf3dea0),
	.w6(32'hbb05cf01),
	.w7(32'hbbb70cc8),
	.w8(32'hba5ee5f4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9a33),
	.w1(32'hbb037c4f),
	.w2(32'hbba909f2),
	.w3(32'h3cc0c2de),
	.w4(32'hbbe094e5),
	.w5(32'h3b8d709e),
	.w6(32'h3b9b9b1c),
	.w7(32'hbc80e8e6),
	.w8(32'h3bc53ab4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb64b86),
	.w1(32'h3b162930),
	.w2(32'hbba64620),
	.w3(32'h3acf4af7),
	.w4(32'h3ae8882d),
	.w5(32'hbbcec075),
	.w6(32'hbc32c6b6),
	.w7(32'h3a4f673f),
	.w8(32'h3abf7cf6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46c94d),
	.w1(32'h3b58b8bd),
	.w2(32'hbae54502),
	.w3(32'h3bbe4c8a),
	.w4(32'hbbeb8fc6),
	.w5(32'h3af35f1b),
	.w6(32'hbbb08098),
	.w7(32'hbb525f0a),
	.w8(32'hbb644028),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a885870),
	.w1(32'h3ba7a69a),
	.w2(32'hbbec4065),
	.w3(32'h3a94a1c0),
	.w4(32'h3b76ad34),
	.w5(32'h3b821a8a),
	.w6(32'h3cd465dd),
	.w7(32'hbcf2b18f),
	.w8(32'hb9bd609e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a3af),
	.w1(32'h3a336055),
	.w2(32'h3b8deb11),
	.w3(32'hbafa406e),
	.w4(32'h3c6d4bfe),
	.w5(32'h3c80ce82),
	.w6(32'h3cc3b6fd),
	.w7(32'hbb032090),
	.w8(32'hbbdb8f6a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77c6aa),
	.w1(32'hb9404f9c),
	.w2(32'hbc90aec0),
	.w3(32'h3b330ed7),
	.w4(32'h39aebfca),
	.w5(32'hbb5ce059),
	.w6(32'h3bd2258b),
	.w7(32'h3bdf0fdc),
	.w8(32'h3a87a193),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6835b8),
	.w1(32'hbaea0528),
	.w2(32'h3c3a2a49),
	.w3(32'hbadf5615),
	.w4(32'h3a05b62c),
	.w5(32'hb96cdbbd),
	.w6(32'hbb3d0791),
	.w7(32'h3b4bd827),
	.w8(32'h3c8ca198),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a4260),
	.w1(32'hbb6ae184),
	.w2(32'hbabca1a7),
	.w3(32'hbb82097d),
	.w4(32'h3a9afb6e),
	.w5(32'h3934afff),
	.w6(32'hbac4f16e),
	.w7(32'hbac12bec),
	.w8(32'hbb439097),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e61298),
	.w1(32'hbc2e9942),
	.w2(32'hbc35a04b),
	.w3(32'hbb505e97),
	.w4(32'hbc3cd0c8),
	.w5(32'hbba5499e),
	.w6(32'hbdc44410),
	.w7(32'h3c361585),
	.w8(32'hbae1da14),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccdcee7),
	.w1(32'h3bbafbdb),
	.w2(32'hbb20ae3e),
	.w3(32'hbb850716),
	.w4(32'h39b40a0a),
	.w5(32'hba9f366e),
	.w6(32'hbbc84dae),
	.w7(32'h3c13f8de),
	.w8(32'h3a4f7847),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c4f1b),
	.w1(32'h3c036a43),
	.w2(32'hba1998d1),
	.w3(32'hb9bbb912),
	.w4(32'h3adf5297),
	.w5(32'h3ac2d008),
	.w6(32'h3b153806),
	.w7(32'hbc2448ac),
	.w8(32'h3b833638),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cd957),
	.w1(32'hbb9d0aa7),
	.w2(32'h3a37a880),
	.w3(32'hbd28e7cf),
	.w4(32'h3b7f71bd),
	.w5(32'h3b26a06b),
	.w6(32'h3bad23d4),
	.w7(32'h3b9fcf26),
	.w8(32'h3b26d429),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5751e5),
	.w1(32'hbadf60a5),
	.w2(32'hbb8261a9),
	.w3(32'hbadf9def),
	.w4(32'h3bd1bc59),
	.w5(32'h3c493c0a),
	.w6(32'h3b55048d),
	.w7(32'h3c4e6263),
	.w8(32'hbbade275),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10ea6c),
	.w1(32'hbc0574b1),
	.w2(32'hbbc35d6a),
	.w3(32'h3b15a5f4),
	.w4(32'hba19775d),
	.w5(32'hbb2989ed),
	.w6(32'h3b667530),
	.w7(32'hbad74c61),
	.w8(32'h3b9aa166),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e5042),
	.w1(32'hbabc752f),
	.w2(32'hbb568abd),
	.w3(32'h39425286),
	.w4(32'hbab4d241),
	.w5(32'h3bafe534),
	.w6(32'hbcb04b44),
	.w7(32'hbb43ba25),
	.w8(32'h3b480662),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda960d),
	.w1(32'hbb81452a),
	.w2(32'hbb983fc8),
	.w3(32'hbc250201),
	.w4(32'h3ba45925),
	.w5(32'hbba8c213),
	.w6(32'hba77492c),
	.w7(32'h3a7970b0),
	.w8(32'hbc34feca),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1e69e),
	.w1(32'h3a1bfb2d),
	.w2(32'h3a9c276f),
	.w3(32'hbc2f671b),
	.w4(32'hbbdcbdd4),
	.w5(32'h3b0e165c),
	.w6(32'h3c28c3f0),
	.w7(32'h3bb52d2e),
	.w8(32'hba997c1a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d8217),
	.w1(32'h3b215277),
	.w2(32'h3b4c38a0),
	.w3(32'h3b862c28),
	.w4(32'h3b4bbada),
	.w5(32'h3b9c7599),
	.w6(32'hbb218023),
	.w7(32'h390de65f),
	.w8(32'h3c8067cf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2794f6),
	.w1(32'hbbbb2d60),
	.w2(32'h3baf4456),
	.w3(32'hbd13de8b),
	.w4(32'h3a5adbf1),
	.w5(32'h3ca14ec0),
	.w6(32'h3c8684ad),
	.w7(32'hbb56bbdd),
	.w8(32'h39fc353e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01c089),
	.w1(32'hbbf55c0f),
	.w2(32'hbd4557bf),
	.w3(32'hbb90086a),
	.w4(32'h3b958193),
	.w5(32'hbb81b21f),
	.w6(32'hb74a9660),
	.w7(32'hbc600b60),
	.w8(32'h3c033047),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c598d13),
	.w1(32'hba4ff11d),
	.w2(32'h3b4326ef),
	.w3(32'h3b1dc1e2),
	.w4(32'hba7af422),
	.w5(32'h3bd00dbe),
	.w6(32'h3c085e6a),
	.w7(32'hbc1f5726),
	.w8(32'h3bad079e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b974),
	.w1(32'h3a871f15),
	.w2(32'hbae0707c),
	.w3(32'h3aed2569),
	.w4(32'h3b88f6f7),
	.w5(32'hbb729f8f),
	.w6(32'hbb2cf472),
	.w7(32'hbb982372),
	.w8(32'hbc6b286b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcaec4),
	.w1(32'hbb90793d),
	.w2(32'h3c417393),
	.w3(32'hbb00cb7a),
	.w4(32'h3b8017c1),
	.w5(32'h3bc12768),
	.w6(32'hbbb967b6),
	.w7(32'h3c299d32),
	.w8(32'h3baf1530),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b599bb0),
	.w1(32'h3d16974f),
	.w2(32'hbba9a782),
	.w3(32'hbc4fc9e2),
	.w4(32'h3ae5d311),
	.w5(32'h3ad5fb73),
	.w6(32'hbbaa6caa),
	.w7(32'h3b70e5a6),
	.w8(32'hbba5d450),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cbff1),
	.w1(32'h3be4cd41),
	.w2(32'h3c88cac4),
	.w3(32'hbbc46501),
	.w4(32'h3cfb13fc),
	.w5(32'hbc8b0eff),
	.w6(32'h3ba568d5),
	.w7(32'h3c05acf1),
	.w8(32'hbc162184),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2fa56),
	.w1(32'h3d7d4a3b),
	.w2(32'hbc75775d),
	.w3(32'h3c7adc91),
	.w4(32'h3b4da7ed),
	.w5(32'h3d1f2b49),
	.w6(32'hbc30e282),
	.w7(32'hbb578380),
	.w8(32'h3bb2f975),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bbe03),
	.w1(32'h3c1f55f1),
	.w2(32'hbc0b7835),
	.w3(32'hbc8af08a),
	.w4(32'hbb81225e),
	.w5(32'h3d15e55d),
	.w6(32'hbc31f444),
	.w7(32'hbb8b0eef),
	.w8(32'hbb95a53d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41276b),
	.w1(32'hbbf78c33),
	.w2(32'hbaa6e12f),
	.w3(32'hbc1e5b5d),
	.w4(32'hbc2c5f02),
	.w5(32'hbb8cc56c),
	.w6(32'h3be5f26e),
	.w7(32'h3bcd6f88),
	.w8(32'h3c0f3b24),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf83086),
	.w1(32'hbb76257e),
	.w2(32'hbc0d413a),
	.w3(32'h3d589f9f),
	.w4(32'h3b1008e5),
	.w5(32'hbbfc7f49),
	.w6(32'h3b518e67),
	.w7(32'h3bf6e426),
	.w8(32'h3c1e0caa),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce999e3),
	.w1(32'h3b3dabad),
	.w2(32'h3d36a20b),
	.w3(32'hbb716657),
	.w4(32'hbc09583e),
	.w5(32'hbc5a8010),
	.w6(32'h3b6e88b9),
	.w7(32'hb84c3339),
	.w8(32'hbb56cc2b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cfd64),
	.w1(32'h3b9287ff),
	.w2(32'hbc73f2b9),
	.w3(32'h3bb4e2f4),
	.w4(32'h3c2e6af9),
	.w5(32'hbc0d97fa),
	.w6(32'h3adbac4b),
	.w7(32'h3cc9119b),
	.w8(32'hbb9b998a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fe127),
	.w1(32'h3b89931b),
	.w2(32'hbaa71b85),
	.w3(32'h3a8d82cf),
	.w4(32'h3af0d0ab),
	.w5(32'h3afe2fc6),
	.w6(32'hbc94132f),
	.w7(32'h3c77accc),
	.w8(32'hbc8e1bdd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44f496),
	.w1(32'h3ba3f65f),
	.w2(32'hbaf2f82e),
	.w3(32'h3b9e483a),
	.w4(32'hbbb66743),
	.w5(32'h3c82ba4e),
	.w6(32'h3bd883c1),
	.w7(32'hbb7a117a),
	.w8(32'h3ba2f53d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e82dbc),
	.w1(32'hbb4e4a52),
	.w2(32'hbc19b87d),
	.w3(32'h381c2f7e),
	.w4(32'hbb929021),
	.w5(32'h3c97a798),
	.w6(32'hbc01f4b1),
	.w7(32'hbc40526f),
	.w8(32'h3b27248d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296174),
	.w1(32'hbb1b734c),
	.w2(32'hbc87758a),
	.w3(32'h3c3f0752),
	.w4(32'h3c546cfe),
	.w5(32'h3c86c5e2),
	.w6(32'h3b89edce),
	.w7(32'h3a35175b),
	.w8(32'h3b8469da),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843f89),
	.w1(32'h3c9716d1),
	.w2(32'h3c8a9802),
	.w3(32'h3c1e26ee),
	.w4(32'h3bad3bb2),
	.w5(32'h3b6493db),
	.w6(32'h3a9320f0),
	.w7(32'hbc7cbbf2),
	.w8(32'h3cf531f0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797dee),
	.w1(32'hbc9f6cc5),
	.w2(32'h3c4900b7),
	.w3(32'h3b95e3b0),
	.w4(32'h3ae785cb),
	.w5(32'hbb589c14),
	.w6(32'hbbe1d2e8),
	.w7(32'hbc0d23d6),
	.w8(32'h3aa9e128),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2a64),
	.w1(32'hbbc7e86a),
	.w2(32'h3dc7fa9b),
	.w3(32'h3c8f71e1),
	.w4(32'hbbc4b574),
	.w5(32'hbc0d006e),
	.w6(32'hbc655f86),
	.w7(32'h3cca7a4e),
	.w8(32'hbc5702fc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5953e7),
	.w1(32'hb8482a01),
	.w2(32'hbbc6b742),
	.w3(32'h3bf63b17),
	.w4(32'h3a52bfdf),
	.w5(32'hbc7fdece),
	.w6(32'h3965513c),
	.w7(32'h3a219641),
	.w8(32'hbc1b7778),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0034ac),
	.w1(32'hbc41fa51),
	.w2(32'hbbc2713c),
	.w3(32'h3c23a95e),
	.w4(32'hb99e1f12),
	.w5(32'hbb8125c2),
	.w6(32'hbbd38430),
	.w7(32'hbc534500),
	.w8(32'h3acc05a7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6905e),
	.w1(32'h3a85c191),
	.w2(32'h3c62a455),
	.w3(32'h3b15c193),
	.w4(32'h3ae493d2),
	.w5(32'hbb04ed70),
	.w6(32'hbc622b63),
	.w7(32'hbc1f6be6),
	.w8(32'hbbc0e845),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1143e6),
	.w1(32'h3baa6385),
	.w2(32'hbc526f37),
	.w3(32'hbcc9a7d8),
	.w4(32'h3c7f6b02),
	.w5(32'hbc1b7546),
	.w6(32'hbba61be6),
	.w7(32'hbb0b9d79),
	.w8(32'h3baef219),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca076d5),
	.w1(32'hbbcfcbda),
	.w2(32'h3c90dc54),
	.w3(32'hbac9a803),
	.w4(32'h3d2390bb),
	.w5(32'hbb0a6ab2),
	.w6(32'hbbc9feae),
	.w7(32'h3c0af422),
	.w8(32'h37bbf4e9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb80724),
	.w1(32'hbbcb96bb),
	.w2(32'h39f07920),
	.w3(32'h3c7f193a),
	.w4(32'h3c4f46bc),
	.w5(32'hbc72bf0e),
	.w6(32'h3bb8de82),
	.w7(32'h3ba75475),
	.w8(32'hbc522735),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4279fa),
	.w1(32'hbc07e67e),
	.w2(32'hbb95b605),
	.w3(32'h3c28badf),
	.w4(32'hbcb91886),
	.w5(32'h3bda8df3),
	.w6(32'h3c51bffc),
	.w7(32'h3bdf02cc),
	.w8(32'hbcc018f6),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a960f61),
	.w1(32'h3ab0c252),
	.w2(32'h3b49cc2e),
	.w3(32'h3aa664ec),
	.w4(32'h3b2adf02),
	.w5(32'hbbc718d9),
	.w6(32'h3b9f750e),
	.w7(32'hba2d1cb5),
	.w8(32'h3bf8c899),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1b8f7),
	.w1(32'h3c3c9f2c),
	.w2(32'h3c879e64),
	.w3(32'h3b7bf18b),
	.w4(32'hbbe0104b),
	.w5(32'hbbbe4369),
	.w6(32'hbbdaf83d),
	.w7(32'hbbab70fe),
	.w8(32'h3c712910),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c3a89),
	.w1(32'hbbf11647),
	.w2(32'hbafe7df6),
	.w3(32'h3b7d3096),
	.w4(32'hbbedc803),
	.w5(32'h3acf3985),
	.w6(32'h3d83a5a5),
	.w7(32'h3bb80511),
	.w8(32'hbc53ab2a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd7f93),
	.w1(32'hbbe0592a),
	.w2(32'hbc777b5c),
	.w3(32'h3c3ca68f),
	.w4(32'h3ad4f03a),
	.w5(32'h3b627da9),
	.w6(32'hbc717a05),
	.w7(32'h3c31528c),
	.w8(32'h3bbb2585),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb9617),
	.w1(32'hbc18b837),
	.w2(32'h3c800c1f),
	.w3(32'h3c7c4a37),
	.w4(32'h3a934996),
	.w5(32'h3bb3d89d),
	.w6(32'h3c23571c),
	.w7(32'h3bc9ecd6),
	.w8(32'h3c7c57bd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d318c65),
	.w1(32'hbb8268b6),
	.w2(32'hbbd626c3),
	.w3(32'hbc3f5397),
	.w4(32'hbb663bb2),
	.w5(32'h3a8041d2),
	.w6(32'hbb590c94),
	.w7(32'hbc1b7e62),
	.w8(32'h3aa528dc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8aa79),
	.w1(32'hbad08ec9),
	.w2(32'hbc06015f),
	.w3(32'hbb6fef7c),
	.w4(32'hbc601e9d),
	.w5(32'h3c0aeabb),
	.w6(32'h3c8e6b89),
	.w7(32'h3b2dd6d7),
	.w8(32'hbb8ba591),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306916),
	.w1(32'h3b9fa421),
	.w2(32'h3b23c1f7),
	.w3(32'hbb0a7d45),
	.w4(32'hbb42c7f7),
	.w5(32'h3b93bbab),
	.w6(32'h3ae5f7a6),
	.w7(32'hbb8413e7),
	.w8(32'hbba5f128),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0e6a),
	.w1(32'hbafd713f),
	.w2(32'hbc222aba),
	.w3(32'h3d9645d3),
	.w4(32'hbb6b9ca4),
	.w5(32'h3b803628),
	.w6(32'h3be632ac),
	.w7(32'h3aa845a6),
	.w8(32'h398f571d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd7e3f),
	.w1(32'hbbc1d832),
	.w2(32'h3ba61e61),
	.w3(32'hbb982b83),
	.w4(32'hbb56adb2),
	.w5(32'h3bf85e5b),
	.w6(32'h3be3342a),
	.w7(32'hbbc13c8b),
	.w8(32'hbb9eb9db),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad24249),
	.w1(32'h3bf99fc3),
	.w2(32'h3ba3d4b8),
	.w3(32'h3b30e2c3),
	.w4(32'hbc0589ef),
	.w5(32'h3c7424d9),
	.w6(32'hbc9b4ba8),
	.w7(32'h3c389146),
	.w8(32'h38eb2975),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e34f9),
	.w1(32'hb99059e4),
	.w2(32'h3a312706),
	.w3(32'h3b98c7ea),
	.w4(32'h3bf386a9),
	.w5(32'h3b0edaa8),
	.w6(32'h3b245488),
	.w7(32'h3ca9d018),
	.w8(32'h3a5d1674),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc264479),
	.w1(32'hbc211e93),
	.w2(32'hbaa2ac3d),
	.w3(32'h3b129f7d),
	.w4(32'hbc0f40e7),
	.w5(32'h3b6b17d6),
	.w6(32'h3b1215bf),
	.w7(32'h3baf6ba9),
	.w8(32'hbc04df6c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4851fe),
	.w1(32'hbb858afd),
	.w2(32'hbbfc2965),
	.w3(32'hb9eb3e20),
	.w4(32'h3b9c71e1),
	.w5(32'h3b151e9c),
	.w6(32'h3b53e7d4),
	.w7(32'h3bd7236f),
	.w8(32'hbaba2521),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978fb4f),
	.w1(32'hbae329bb),
	.w2(32'hbb92851c),
	.w3(32'hbc17b384),
	.w4(32'hbb779d43),
	.w5(32'hbbe68460),
	.w6(32'h3b971fa2),
	.w7(32'hbb8637f7),
	.w8(32'h39d6845e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82deab),
	.w1(32'h3b9dd013),
	.w2(32'h3bc318c9),
	.w3(32'h3b476af7),
	.w4(32'hbd021ac7),
	.w5(32'hbbed5d4f),
	.w6(32'hbb557738),
	.w7(32'hbbd9804d),
	.w8(32'hb9f0dda0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9086fd),
	.w1(32'h3b1c030f),
	.w2(32'hb5860e06),
	.w3(32'hbc2a6428),
	.w4(32'hb9b4eebd),
	.w5(32'hbb7d1a36),
	.w6(32'hbaa44a6d),
	.w7(32'h3b93786c),
	.w8(32'h3c19e055),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45f82),
	.w1(32'hbb74d91e),
	.w2(32'hbac678cc),
	.w3(32'h3b27c745),
	.w4(32'hbb1b3798),
	.w5(32'h3b2249d0),
	.w6(32'hbc4bb5ce),
	.w7(32'h3b7b06f5),
	.w8(32'hbcc28ddf),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56a2dc),
	.w1(32'hbb0df604),
	.w2(32'hb90b58cf),
	.w3(32'h3b8ac42e),
	.w4(32'hba8cbea7),
	.w5(32'h3b15c248),
	.w6(32'hbc231223),
	.w7(32'hbc5ff188),
	.w8(32'h3b0fb389),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a5b60),
	.w1(32'h3b2f5efa),
	.w2(32'hbc0b9a01),
	.w3(32'h3bc71017),
	.w4(32'h3bd850b3),
	.w5(32'hba3c8222),
	.w6(32'h3b0c376d),
	.w7(32'h3b7d3770),
	.w8(32'h3b90eeb7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5089c),
	.w1(32'h3b2dfaa3),
	.w2(32'h3cbeb685),
	.w3(32'hbd2fae96),
	.w4(32'h3c8b4173),
	.w5(32'hbc0ba556),
	.w6(32'h3a116488),
	.w7(32'h3c8ce0d6),
	.w8(32'h3b801f52),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb2245),
	.w1(32'h3b2e09ae),
	.w2(32'hbaaf5272),
	.w3(32'hbcc86b11),
	.w4(32'h3c151509),
	.w5(32'hbbd86558),
	.w6(32'h3c0dc1f2),
	.w7(32'hbc225063),
	.w8(32'hbc1827fc),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd0ea),
	.w1(32'h3af15fbd),
	.w2(32'hbb8a1231),
	.w3(32'hbbd644ab),
	.w4(32'h3ba20010),
	.w5(32'h391a2d42),
	.w6(32'h3bfe602a),
	.w7(32'hbadfa446),
	.w8(32'hbc06e9d8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac29ee),
	.w1(32'h3b09a726),
	.w2(32'h393ac737),
	.w3(32'hba13f5e2),
	.w4(32'h3bad457a),
	.w5(32'hbba96084),
	.w6(32'hbb4c775d),
	.w7(32'h38c62f97),
	.w8(32'hbc69cdca),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2dbf),
	.w1(32'hbb8845d0),
	.w2(32'hbc469290),
	.w3(32'h3bb0dab9),
	.w4(32'h3c18410a),
	.w5(32'hbb9475f3),
	.w6(32'hbb80cdbb),
	.w7(32'hbbd8fab5),
	.w8(32'hbb464a60),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ade9ad),
	.w1(32'hbb12c634),
	.w2(32'hba1f1331),
	.w3(32'h3a93e97e),
	.w4(32'hbb48e6df),
	.w5(32'h3ab0f565),
	.w6(32'hbbba733a),
	.w7(32'hbc1d41a2),
	.w8(32'hbcdb382c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21d2b1),
	.w1(32'h3c041f35),
	.w2(32'h3aa17a82),
	.w3(32'hbd07d8bd),
	.w4(32'h3c8783fd),
	.w5(32'hba54131d),
	.w6(32'hba5e2fd0),
	.w7(32'hbb20f1bc),
	.w8(32'hbaf59054),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bb99f),
	.w1(32'h3c9fdb27),
	.w2(32'hbc23249d),
	.w3(32'hbb38f713),
	.w4(32'h3c00f716),
	.w5(32'h3ade1db3),
	.w6(32'h3bc79627),
	.w7(32'h3c4ac3ef),
	.w8(32'h3c5c0c6a),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45962e),
	.w1(32'h3c0b3ec7),
	.w2(32'h3aaa04d4),
	.w3(32'hbc3949b6),
	.w4(32'h3b922a7c),
	.w5(32'hbae9489d),
	.w6(32'h3a5df945),
	.w7(32'hb8c7137b),
	.w8(32'hbc3f8d44),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4694d3),
	.w1(32'h3b8aab8a),
	.w2(32'hbb2d9b56),
	.w3(32'h3ba434b0),
	.w4(32'hb91d7d70),
	.w5(32'h3d183ab3),
	.w6(32'hbae5a49a),
	.w7(32'h3aba3c37),
	.w8(32'h3cf05b33),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3daf39),
	.w1(32'h3b3a8a05),
	.w2(32'hbbe961b4),
	.w3(32'hbaf3525b),
	.w4(32'hbb4e7915),
	.w5(32'hba83a958),
	.w6(32'h3b3213a4),
	.w7(32'hbba9f83c),
	.w8(32'hb9d2ea11),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96255b),
	.w1(32'h3bcd9910),
	.w2(32'hba4ea0fd),
	.w3(32'h3a01a146),
	.w4(32'h3b5a8863),
	.w5(32'h3a8ea6b6),
	.w6(32'hbb28407f),
	.w7(32'hbca0ac5b),
	.w8(32'h3b900a8c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eeed0),
	.w1(32'h3bdac547),
	.w2(32'h3af75586),
	.w3(32'hbcb6b7cb),
	.w4(32'hbb471508),
	.w5(32'hbb8674c9),
	.w6(32'h3bf148c9),
	.w7(32'hbc916376),
	.w8(32'h3adc6ef5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af471e4),
	.w1(32'h3b338466),
	.w2(32'hbc0c8631),
	.w3(32'h39872ada),
	.w4(32'h3b5f8a7b),
	.w5(32'hbb421947),
	.w6(32'h3ba4d5f8),
	.w7(32'hbb95b6e4),
	.w8(32'hb944faf0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c139aee),
	.w1(32'h3b359320),
	.w2(32'hbbbd4a90),
	.w3(32'hbc5684cc),
	.w4(32'h3b1a069a),
	.w5(32'hbc0be133),
	.w6(32'hbc23ef9c),
	.w7(32'hbb4c4f50),
	.w8(32'hba13aa4f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8338b0),
	.w1(32'h3c9dedd3),
	.w2(32'h3c3c53eb),
	.w3(32'hbb7ee4d4),
	.w4(32'h3c19dd62),
	.w5(32'hb99af266),
	.w6(32'hbbaec28f),
	.w7(32'hbb902938),
	.w8(32'hbbcd49ee),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58790c),
	.w1(32'h3cc6d0ed),
	.w2(32'h3c545745),
	.w3(32'h3c8cfd94),
	.w4(32'hbb194edf),
	.w5(32'hbc61d2de),
	.w6(32'hbbfae8c9),
	.w7(32'h3c167b82),
	.w8(32'hbc9cd640),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc329d5d),
	.w1(32'h3b9044d0),
	.w2(32'hbc8118b8),
	.w3(32'h3c5a3ee7),
	.w4(32'h3b3eebb9),
	.w5(32'hbc483990),
	.w6(32'hbb978a1f),
	.w7(32'hbba59588),
	.w8(32'h3a95b231),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15ee44),
	.w1(32'hb8a0ac74),
	.w2(32'hbaf83fcb),
	.w3(32'hbbad02ac),
	.w4(32'hbbd2e959),
	.w5(32'hbc712bbc),
	.w6(32'hbb7e43dc),
	.w7(32'hbc9f4ec4),
	.w8(32'h3c14d5bd),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5b51e),
	.w1(32'hbb06c91d),
	.w2(32'hbb73655a),
	.w3(32'hbc2abdf3),
	.w4(32'hbcc68182),
	.w5(32'hb99fe78b),
	.w6(32'hbc7bb947),
	.w7(32'h3bce3c2f),
	.w8(32'h3c33f5fe),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7af0a1),
	.w1(32'h3a78dc45),
	.w2(32'hbac60db1),
	.w3(32'h3c935241),
	.w4(32'h3bbcf0ee),
	.w5(32'h3b262981),
	.w6(32'h3a8af252),
	.w7(32'h3c879bf7),
	.w8(32'h3babe583),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1ebe2),
	.w1(32'h3d2ea13f),
	.w2(32'hbd6f480a),
	.w3(32'hba80d36d),
	.w4(32'hbb9e73a3),
	.w5(32'hbc90df56),
	.w6(32'hbae77d1a),
	.w7(32'hbbe9ab87),
	.w8(32'hbc970772),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4db9b),
	.w1(32'h3c3d0eb5),
	.w2(32'h3c65b23a),
	.w3(32'hbc020ede),
	.w4(32'h3b88b84e),
	.w5(32'hbc0be6f9),
	.w6(32'h3bdfe192),
	.w7(32'hbc6c197a),
	.w8(32'h3bbcac65),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16865),
	.w1(32'hbba19a24),
	.w2(32'hbc325b10),
	.w3(32'hbc0be808),
	.w4(32'hbbfadaf9),
	.w5(32'hbc2926ed),
	.w6(32'h3ba879c0),
	.w7(32'h3be07148),
	.w8(32'hbc4b249d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc620a6b),
	.w1(32'h3c1b12b0),
	.w2(32'hbbc065c7),
	.w3(32'h3bc5a61f),
	.w4(32'h3b944fdb),
	.w5(32'hbbb60b1e),
	.w6(32'h3c0d4275),
	.w7(32'hbbbb4a12),
	.w8(32'hba2c9f37),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c207666),
	.w1(32'hbc69b1cc),
	.w2(32'hbb065461),
	.w3(32'h3affa17c),
	.w4(32'h3c2a9945),
	.w5(32'hbc95480d),
	.w6(32'hbc7a3ba7),
	.w7(32'h3a17e3fa),
	.w8(32'hbbee197b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b329e97),
	.w1(32'h3b8474da),
	.w2(32'hbb872bfa),
	.w3(32'hbbae578e),
	.w4(32'hbbbc720f),
	.w5(32'h3c34b1b2),
	.w6(32'hbb589c25),
	.w7(32'h3c559d05),
	.w8(32'h39be2f02),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9122),
	.w1(32'h3b27ae0e),
	.w2(32'h3c67403d),
	.w3(32'h38dfed3a),
	.w4(32'hbbfdd309),
	.w5(32'h3c1dabea),
	.w6(32'hbbe080fd),
	.w7(32'hbc2ac4ad),
	.w8(32'h3c2f10c2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb414006),
	.w1(32'hbd5e96e9),
	.w2(32'hbc0f9b36),
	.w3(32'hbc456f9a),
	.w4(32'hbb06cfd1),
	.w5(32'hbca58c94),
	.w6(32'hbb6aec9c),
	.w7(32'hbb849c97),
	.w8(32'h3cab9e60),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc94bfb0),
	.w1(32'h3a877204),
	.w2(32'hbc893166),
	.w3(32'h3c7e0074),
	.w4(32'hb9c232af),
	.w5(32'h3b673e83),
	.w6(32'hbc4a0d41),
	.w7(32'hbc65cdb9),
	.w8(32'h3be4e04e),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaa948),
	.w1(32'h3b666fff),
	.w2(32'h3a9f49a6),
	.w3(32'hbc224fa4),
	.w4(32'h3b756633),
	.w5(32'hbc042f91),
	.w6(32'h3b988fe7),
	.w7(32'hbc100ad3),
	.w8(32'h3b538f4a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1fc3),
	.w1(32'hb93976a7),
	.w2(32'hbc184d9e),
	.w3(32'hbb4d409d),
	.w4(32'h3c0da20e),
	.w5(32'h3b5dd858),
	.w6(32'h3c197727),
	.w7(32'hbc530945),
	.w8(32'h3c2d7045),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8fc82),
	.w1(32'hbc2303da),
	.w2(32'h3c5b1c5e),
	.w3(32'h3b971ef8),
	.w4(32'hbb919c99),
	.w5(32'h3cca5419),
	.w6(32'h392ba4dd),
	.w7(32'h3bd8b514),
	.w8(32'h3be62d96),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f3d0a),
	.w1(32'h3bc27f02),
	.w2(32'h3d28ccfe),
	.w3(32'h3c3e56bc),
	.w4(32'hbb96ac7f),
	.w5(32'hbc7d8fb7),
	.w6(32'h3ba624cc),
	.w7(32'h3c73e840),
	.w8(32'hbc6d4d62),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe39d8),
	.w1(32'hbab692d4),
	.w2(32'h3c9274ae),
	.w3(32'hbc8c00b6),
	.w4(32'h3ba79295),
	.w5(32'hbc35a817),
	.w6(32'hbc7fc3c2),
	.w7(32'h3c766ef9),
	.w8(32'hbc7d25ac),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd834b),
	.w1(32'hbb7d7796),
	.w2(32'hbc214e28),
	.w3(32'hbc0dc794),
	.w4(32'hbca68adf),
	.w5(32'h3c7a828f),
	.w6(32'hbc03dbfa),
	.w7(32'h3b38ac10),
	.w8(32'h3b7f5ccc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc882251),
	.w1(32'hbbb11259),
	.w2(32'h3ab93858),
	.w3(32'hbc15a993),
	.w4(32'hbcae9357),
	.w5(32'hbb588754),
	.w6(32'hbc850340),
	.w7(32'h3a6bd0ec),
	.w8(32'hbccb00ed),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98b235),
	.w1(32'hbc85c90f),
	.w2(32'h3ba4d334),
	.w3(32'hba78e20d),
	.w4(32'hbc2420c8),
	.w5(32'h3b3f9a98),
	.w6(32'h3c343bac),
	.w7(32'h3c8bdcb9),
	.w8(32'h3aa2d621),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb730ba),
	.w1(32'h3c85c488),
	.w2(32'hbc67ae54),
	.w3(32'hbc0be300),
	.w4(32'hbc0602e3),
	.w5(32'hbb82f592),
	.w6(32'h3a933f27),
	.w7(32'hbb8ece56),
	.w8(32'h3b630277),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e02c7),
	.w1(32'hbc1f1476),
	.w2(32'hba4b43a7),
	.w3(32'hbbd8883c),
	.w4(32'h3c511208),
	.w5(32'h3c0166e7),
	.w6(32'h3c81069c),
	.w7(32'hbc5a33e7),
	.w8(32'h3bb9a809),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15d992),
	.w1(32'h38d68d28),
	.w2(32'h3bb8b13f),
	.w3(32'hbc7408cb),
	.w4(32'hbc97d9a1),
	.w5(32'hbb21c883),
	.w6(32'h3b98196b),
	.w7(32'h3c44f245),
	.w8(32'hbc1a04d4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dec72),
	.w1(32'h39a8e9b7),
	.w2(32'h3b757c2f),
	.w3(32'h3a8a25a2),
	.w4(32'h3ab1c5c0),
	.w5(32'h3b8d771a),
	.w6(32'h3cbd0bd4),
	.w7(32'h3b2cd7b3),
	.w8(32'hbb9ebb92),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f15f),
	.w1(32'hbbdfeda4),
	.w2(32'h3bcdb0ba),
	.w3(32'h3b9827be),
	.w4(32'h3c0f4826),
	.w5(32'hbad85360),
	.w6(32'hbcdb2602),
	.w7(32'h3b3a1303),
	.w8(32'hbbb145a5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba900d64),
	.w1(32'hbb1f976a),
	.w2(32'h3b0c4de5),
	.w3(32'h3ba78017),
	.w4(32'h3bdf2dbf),
	.w5(32'h3b2ce89f),
	.w6(32'h3cbc6991),
	.w7(32'h399d4505),
	.w8(32'h3b17f298),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule