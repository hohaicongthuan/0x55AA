module layer_8_featuremap_62(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b3a1b),
	.w1(32'hb72e5e96),
	.w2(32'h38f5107b),
	.w3(32'hb93f2aa3),
	.w4(32'hb79ae9f5),
	.w5(32'h36fd07f5),
	.w6(32'hb942bdaf),
	.w7(32'hb8afb93d),
	.w8(32'h35b63c08),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941a314),
	.w1(32'h39810886),
	.w2(32'h39b99d24),
	.w3(32'h39a36ffe),
	.w4(32'h39ae16e2),
	.w5(32'h39b843cf),
	.w6(32'h39a5211f),
	.w7(32'h39caa2b5),
	.w8(32'h39a7e602),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2ec56),
	.w1(32'h39288959),
	.w2(32'h38d125ec),
	.w3(32'h39fb0e2a),
	.w4(32'h391ad6b5),
	.w5(32'h38bddc7a),
	.w6(32'h39a29a76),
	.w7(32'h390e5e50),
	.w8(32'h38d59fad),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377dda5e),
	.w1(32'hb76103f3),
	.w2(32'h36b0c5e5),
	.w3(32'hb7ad521e),
	.w4(32'hb7f74d34),
	.w5(32'hb5e88255),
	.w6(32'hb6c882a6),
	.w7(32'hb7e2ec1d),
	.w8(32'hb64b899b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901a285),
	.w1(32'h39c31442),
	.w2(32'h3a04952c),
	.w3(32'h39247111),
	.w4(32'h39c2f1eb),
	.w5(32'h39caac87),
	.w6(32'h39be4ac3),
	.w7(32'h39cf460b),
	.w8(32'h39a44c62),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f1884),
	.w1(32'h38d9b3a6),
	.w2(32'h3712a535),
	.w3(32'h3934de0c),
	.w4(32'h3892db0b),
	.w5(32'h36071847),
	.w6(32'h398a4fdc),
	.w7(32'h395090e6),
	.w8(32'h38d0cbd5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75b0fc7),
	.w1(32'hb6d5644f),
	.w2(32'hb6b8675d),
	.w3(32'hb49a3911),
	.w4(32'hb5e5a90c),
	.w5(32'hb7b8e7fd),
	.w6(32'h35313eb0),
	.w7(32'h36695ee8),
	.w8(32'hb6b43e5b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a156478),
	.w1(32'h3a434039),
	.w2(32'h3a41db3f),
	.w3(32'h39f752ee),
	.w4(32'h3a07425d),
	.w5(32'h3a20e658),
	.w6(32'h3a4310d4),
	.w7(32'h3a425ee1),
	.w8(32'h3a11a759),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06d52f),
	.w1(32'h3a290235),
	.w2(32'h39f5c4e7),
	.w3(32'h398e021d),
	.w4(32'h398e7403),
	.w5(32'h38ec31d7),
	.w6(32'h3a17658f),
	.w7(32'h3a0d0e85),
	.w8(32'h39dfe2a6),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39951f8a),
	.w1(32'h395d295c),
	.w2(32'h391e65d7),
	.w3(32'h39d8ad53),
	.w4(32'h39c55307),
	.w5(32'h399d3174),
	.w6(32'h39aff21a),
	.w7(32'h398fd35d),
	.w8(32'h3953f129),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f61576),
	.w1(32'hb9568430),
	.w2(32'h37d02b86),
	.w3(32'hba0766a8),
	.w4(32'hb9b14d4c),
	.w5(32'hb9099446),
	.w6(32'hb9b50bb8),
	.w7(32'hb99c4bf5),
	.w8(32'hb9251902),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861cb1f),
	.w1(32'h38cf5fd9),
	.w2(32'h38cc266e),
	.w3(32'h385b9cf0),
	.w4(32'h380a1b42),
	.w5(32'h36ff70fa),
	.w6(32'hb913b29f),
	.w7(32'hb904121d),
	.w8(32'hb8869de9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b812d9),
	.w1(32'h398e2154),
	.w2(32'h399c1c28),
	.w3(32'h39c2353b),
	.w4(32'h398f2747),
	.w5(32'h39b37cf3),
	.w6(32'h39e12513),
	.w7(32'h39c00632),
	.w8(32'h39ac26c8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7751381),
	.w1(32'h364e8735),
	.w2(32'hb594d6f8),
	.w3(32'h3804b4b8),
	.w4(32'hb6893048),
	.w5(32'hb70c40c4),
	.w6(32'h37a5daae),
	.w7(32'hb7de6a90),
	.w8(32'hb76288f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61f2d6b),
	.w1(32'h36addb44),
	.w2(32'h37010ba8),
	.w3(32'h37316e99),
	.w4(32'h37894b75),
	.w5(32'h36598502),
	.w6(32'h372a7ad6),
	.w7(32'h370243ae),
	.w8(32'h3648c59e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76dfff3),
	.w1(32'hb7c790e9),
	.w2(32'h3698cb6c),
	.w3(32'hb81b2d09),
	.w4(32'h354fa3e2),
	.w5(32'h37a66cf9),
	.w6(32'h38bb32c4),
	.w7(32'h391c6b5b),
	.w8(32'h38938062),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9348701),
	.w1(32'hb8f3c9c7),
	.w2(32'h35f0286a),
	.w3(32'hb90f5a22),
	.w4(32'hb89b6327),
	.w5(32'hb91e60e6),
	.w6(32'hb97c1280),
	.w7(32'hb88d75f2),
	.w8(32'hb8b26ee4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f052c9),
	.w1(32'h399d11ea),
	.w2(32'h39af25b4),
	.w3(32'h3a4538bf),
	.w4(32'h3a020015),
	.w5(32'h39bcd797),
	.w6(32'h3a2d3b5f),
	.w7(32'h3a32de56),
	.w8(32'h39e7f8e6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86bb87),
	.w1(32'hb8cf80c5),
	.w2(32'h3a1d4822),
	.w3(32'hba918cd1),
	.w4(32'hba24194c),
	.w5(32'h38daf9cc),
	.w6(32'hb9a4d07b),
	.w7(32'hb6540ed7),
	.w8(32'h396ffbdb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d0cff),
	.w1(32'h398a6387),
	.w2(32'h38c18104),
	.w3(32'h3a2e43a1),
	.w4(32'h3a1a10f0),
	.w5(32'h39a7c0d3),
	.w6(32'h3a2ed78b),
	.w7(32'h39f7ade5),
	.w8(32'hb86baf3d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba177874),
	.w1(32'hb9f246d8),
	.w2(32'hba241320),
	.w3(32'hb989849f),
	.w4(32'hb95f4dc1),
	.w5(32'hb9fb213e),
	.w6(32'hb9f921cf),
	.w7(32'hb9b6de58),
	.w8(32'hb844160d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712bc3c),
	.w1(32'h383588b7),
	.w2(32'hb989f9e3),
	.w3(32'h39a816c4),
	.w4(32'h38f8eb5c),
	.w5(32'hb84f0240),
	.w6(32'h39eb153b),
	.w7(32'h393b5b94),
	.w8(32'hb70e33f3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8785c),
	.w1(32'h3aca74b8),
	.w2(32'h3b263d2e),
	.w3(32'hb972cb12),
	.w4(32'h3aa84990),
	.w5(32'h3af4996d),
	.w6(32'h3a4a037a),
	.w7(32'h3aea7eb9),
	.w8(32'h3ae9f89d),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9133c),
	.w1(32'h39da2997),
	.w2(32'h39cb6e20),
	.w3(32'h3a2ad322),
	.w4(32'h3a13d4b0),
	.w5(32'h397eec73),
	.w6(32'h3975194c),
	.w7(32'h38de26c1),
	.w8(32'h384cfcd6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a67197),
	.w1(32'h37809d8c),
	.w2(32'h39440bd2),
	.w3(32'hb91b117a),
	.w4(32'hb9af0fab),
	.w5(32'hb8bb2a76),
	.w6(32'hb8f55e2b),
	.w7(32'hb9357c90),
	.w8(32'hb5bf31e1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf0bbb),
	.w1(32'h39f9f788),
	.w2(32'h3a89be91),
	.w3(32'hb97f2f00),
	.w4(32'h39a3e1b4),
	.w5(32'h3a237d9c),
	.w6(32'h38aa3a52),
	.w7(32'h3a0f225f),
	.w8(32'h3a00d030),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386a311e),
	.w1(32'h38301fb5),
	.w2(32'h3710fb22),
	.w3(32'h37f046c8),
	.w4(32'h380ebe2a),
	.w5(32'h3798b770),
	.w6(32'h388cddbb),
	.w7(32'h38869339),
	.w8(32'h37c5e6aa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1e4c7),
	.w1(32'hbb842d21),
	.w2(32'h3a81d803),
	.w3(32'hbb98142f),
	.w4(32'hbbd4497e),
	.w5(32'hbbacdbc5),
	.w6(32'hbb6247d7),
	.w7(32'hbb61849f),
	.w8(32'hbbdb8949),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2fcec),
	.w1(32'h385750c9),
	.w2(32'h39b759a2),
	.w3(32'hb98e05fc),
	.w4(32'h382eeba1),
	.w5(32'h396bd27a),
	.w6(32'hb91d14d5),
	.w7(32'h3911c802),
	.w8(32'h3980cf56),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2a8cf),
	.w1(32'h38d4acbc),
	.w2(32'h390c25e1),
	.w3(32'h395fa6c8),
	.w4(32'h3947e1ae),
	.w5(32'h38c4c40b),
	.w6(32'h396c5015),
	.w7(32'h394a1218),
	.w8(32'h39456b91),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38468cb5),
	.w1(32'hb7c2d920),
	.w2(32'h3879094c),
	.w3(32'h3919d8b5),
	.w4(32'h38622108),
	.w5(32'h38abcd14),
	.w6(32'h390574c0),
	.w7(32'h38144fb9),
	.w8(32'h384a9d0f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388fa002),
	.w1(32'hb7de8ba2),
	.w2(32'hb8cfd85c),
	.w3(32'h38999221),
	.w4(32'hb8c3b5fe),
	.w5(32'hb90880ca),
	.w6(32'h3893f3bf),
	.w7(32'hb8bd9865),
	.w8(32'hb8fa7a81),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f1658),
	.w1(32'hb73b3d23),
	.w2(32'hb72b9493),
	.w3(32'h3632120f),
	.w4(32'h3525797d),
	.w5(32'hb6e90d01),
	.w6(32'h36545bef),
	.w7(32'h36b649b2),
	.w8(32'h36964fa3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63a6428),
	.w1(32'hb610a96b),
	.w2(32'hb62c5a6a),
	.w3(32'hb564040d),
	.w4(32'hb65d1c9d),
	.w5(32'hb68cf148),
	.w6(32'hb62cb689),
	.w7(32'hb6a61494),
	.w8(32'hb6838285),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c77126),
	.w1(32'h385fb512),
	.w2(32'hb8d0ae7a),
	.w3(32'h3a0db400),
	.w4(32'h399afc8b),
	.w5(32'h38056941),
	.w6(32'h39ec44a1),
	.w7(32'h39818ea9),
	.w8(32'h390205de),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce26b9),
	.w1(32'h39cf6932),
	.w2(32'h3a0f9b0e),
	.w3(32'h397951a0),
	.w4(32'h39e11a37),
	.w5(32'h3a1205fa),
	.w6(32'h39e00cfe),
	.w7(32'h3a17e113),
	.w8(32'h3a04e0fc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3747d92c),
	.w1(32'hb6698ce1),
	.w2(32'hb711cf67),
	.w3(32'h3678a593),
	.w4(32'h379e0fae),
	.w5(32'h3707bb48),
	.w6(32'hb4471cfd),
	.w7(32'h381e4bc6),
	.w8(32'h370faccc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac6e51),
	.w1(32'h3a1e189c),
	.w2(32'h3a5a7b33),
	.w3(32'h39cfa4aa),
	.w4(32'h3a21022b),
	.w5(32'h3a271e54),
	.w6(32'h39e80514),
	.w7(32'h3a2fbf9f),
	.w8(32'h3a189a5c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370f4ae0),
	.w1(32'hb6c77477),
	.w2(32'hb762e804),
	.w3(32'h36392173),
	.w4(32'hb70c7d6e),
	.w5(32'hb7243a2e),
	.w6(32'h361a174c),
	.w7(32'hb6d0537f),
	.w8(32'h35ce1623),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d198a),
	.w1(32'hb821eeac),
	.w2(32'hb7f59df4),
	.w3(32'hb83f6fc8),
	.w4(32'hb8331426),
	.w5(32'hb7fc1269),
	.w6(32'hb858fe03),
	.w7(32'hb85262c1),
	.w8(32'hb807108b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1205b),
	.w1(32'h39c23307),
	.w2(32'h3a1eb959),
	.w3(32'h3a70acd1),
	.w4(32'h3a37dcec),
	.w5(32'h3a19e685),
	.w6(32'h3a83b436),
	.w7(32'h3a6e20f3),
	.w8(32'h39a34908),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e658ac),
	.w1(32'h39a18bf1),
	.w2(32'h39931a2d),
	.w3(32'hba6adf1a),
	.w4(32'hba2995d5),
	.w5(32'hba1dd187),
	.w6(32'hba03e7aa),
	.w7(32'h38e85078),
	.w8(32'hbaf26c06),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb870d65),
	.w1(32'hbb4c0ca7),
	.w2(32'hb90803e6),
	.w3(32'hbb684c19),
	.w4(32'h3755975b),
	.w5(32'hbb654a4d),
	.w6(32'h3b56799e),
	.w7(32'hb88f257c),
	.w8(32'h396265cf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f09ec),
	.w1(32'h3a2a1f61),
	.w2(32'h39f74444),
	.w3(32'hb98b019d),
	.w4(32'hb7fcf242),
	.w5(32'h39765c2d),
	.w6(32'hb9c17745),
	.w7(32'h39ea4af5),
	.w8(32'h3a684b6f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f1d07),
	.w1(32'h3a93cad3),
	.w2(32'h3afc97a7),
	.w3(32'hb9c540b7),
	.w4(32'hb7e3e3c7),
	.w5(32'h3a51b796),
	.w6(32'hb9518323),
	.w7(32'h3a79c949),
	.w8(32'hba95f248),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2da714),
	.w1(32'h38f9c145),
	.w2(32'h3a34f353),
	.w3(32'h39566a5c),
	.w4(32'h3aad57b9),
	.w5(32'h3afd4d4c),
	.w6(32'hbacd6240),
	.w7(32'hb9cbbdd9),
	.w8(32'hbb7877dd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e68bb),
	.w1(32'hbaab5a24),
	.w2(32'hbbeecd11),
	.w3(32'hba835a1e),
	.w4(32'hba82b1b1),
	.w5(32'h3b363930),
	.w6(32'hbb3fe136),
	.w7(32'hba7d139c),
	.w8(32'hbaa3ae63),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a17d7),
	.w1(32'h393f008f),
	.w2(32'h3b065fe5),
	.w3(32'hba2b3e4f),
	.w4(32'hbae337e0),
	.w5(32'hba686ac4),
	.w6(32'hba4e9a48),
	.w7(32'h386afbab),
	.w8(32'h3ac08ed7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd4593),
	.w1(32'h39b70199),
	.w2(32'h3af46238),
	.w3(32'h3b472fe4),
	.w4(32'h3b325fe2),
	.w5(32'h3b81ae14),
	.w6(32'h3b101cc4),
	.w7(32'h3aecd3bd),
	.w8(32'h3a0a7005),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac13099),
	.w1(32'h3aa4fec8),
	.w2(32'h3ad31bcc),
	.w3(32'h3a2bb5da),
	.w4(32'h3a9417fc),
	.w5(32'h3abe29bb),
	.w6(32'hba00d3e7),
	.w7(32'h3a2fbc48),
	.w8(32'h39a95461),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cd2d8),
	.w1(32'h3a4f1f31),
	.w2(32'h3aa35a8c),
	.w3(32'h395c2c22),
	.w4(32'h39eba3d5),
	.w5(32'h3a39c450),
	.w6(32'h392d85b5),
	.w7(32'h3a8be63f),
	.w8(32'h3916053c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384a439c),
	.w1(32'h3b07ba3f),
	.w2(32'h3b4b9060),
	.w3(32'hbab50923),
	.w4(32'hb94211e2),
	.w5(32'h3a8b9cb2),
	.w6(32'hb7b8d415),
	.w7(32'h3afcec84),
	.w8(32'hbad7a531),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64e48f),
	.w1(32'hba12874d),
	.w2(32'hbc0d08a0),
	.w3(32'hbb84e7c4),
	.w4(32'h3a6dba28),
	.w5(32'hbb9b041e),
	.w6(32'h3b7de4cf),
	.w7(32'hbb1db448),
	.w8(32'h3ac4e64b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac982a6),
	.w1(32'hba71395d),
	.w2(32'h3a8e38ec),
	.w3(32'hb9bbeb8e),
	.w4(32'hbafdffb7),
	.w5(32'hb8dcb9bc),
	.w6(32'h394cb4e4),
	.w7(32'hb94acb52),
	.w8(32'h3b69d000),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcecdfb),
	.w1(32'hbb57ff32),
	.w2(32'hbb5d9a1f),
	.w3(32'h3b0e539a),
	.w4(32'h39ac178e),
	.w5(32'hba8ba297),
	.w6(32'h3a06df06),
	.w7(32'hbab04acd),
	.w8(32'hbb23a73a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba731b9),
	.w1(32'hbb297958),
	.w2(32'hbbbf142e),
	.w3(32'hbb9882f1),
	.w4(32'hbbb9acfb),
	.w5(32'hbbbf597f),
	.w6(32'hbbd337a6),
	.w7(32'hbbaee42e),
	.w8(32'h39e29cb5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac14c1c),
	.w1(32'hba7d1a95),
	.w2(32'h3a2a8908),
	.w3(32'h398189b3),
	.w4(32'h39be29b3),
	.w5(32'hb99467dd),
	.w6(32'hbb1de843),
	.w7(32'hbac88e93),
	.w8(32'hb9c73a6a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf263e6),
	.w1(32'hbb787f1c),
	.w2(32'h39ee9131),
	.w3(32'hbaf89213),
	.w4(32'h38915521),
	.w5(32'hb8a7a6be),
	.w6(32'h3b59d24b),
	.w7(32'h3b1a54bc),
	.w8(32'h3b19d8d3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba164732),
	.w1(32'hb9b1ef9d),
	.w2(32'h3a06e77e),
	.w3(32'hb9dd7590),
	.w4(32'h38be217c),
	.w5(32'h3a7dcd6d),
	.w6(32'h3993c3bd),
	.w7(32'h3a64413e),
	.w8(32'hbb5a44f6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2da77f),
	.w1(32'hbab14313),
	.w2(32'hbad43e40),
	.w3(32'hbb1facb3),
	.w4(32'hbb77d623),
	.w5(32'hbb14bd75),
	.w6(32'hbaca7123),
	.w7(32'hbb5222a8),
	.w8(32'hbb008a69),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb687f3c),
	.w1(32'h3a247d09),
	.w2(32'hbb6bc82a),
	.w3(32'h3b14efa7),
	.w4(32'h3b3aaed9),
	.w5(32'hbaaec6b0),
	.w6(32'hbafcd07a),
	.w7(32'hbb9699a2),
	.w8(32'hba873e21),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf9f35),
	.w1(32'hbaceb6c8),
	.w2(32'hbad0fc48),
	.w3(32'hbaf110d5),
	.w4(32'hba915843),
	.w5(32'hbae0ffb2),
	.w6(32'hbb259eaa),
	.w7(32'hbb0b1d45),
	.w8(32'h3aa534d0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02043b),
	.w1(32'h3a27da22),
	.w2(32'h3aad6edd),
	.w3(32'h3a572908),
	.w4(32'h3a0f94d2),
	.w5(32'h3a946d89),
	.w6(32'hb9b90ec1),
	.w7(32'h3a7076c8),
	.w8(32'hb905e264),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a53aa),
	.w1(32'h39d78dd4),
	.w2(32'hba210240),
	.w3(32'hba7cd035),
	.w4(32'hb9f456e5),
	.w5(32'hba23242c),
	.w6(32'hb9f10b2a),
	.w7(32'h3b1088cd),
	.w8(32'h39baab9b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5db599),
	.w1(32'h3a54e000),
	.w2(32'h3aaf38bd),
	.w3(32'h3974036a),
	.w4(32'h3a217b3b),
	.w5(32'h3a9939a8),
	.w6(32'h37e74024),
	.w7(32'h3a9eacbc),
	.w8(32'hb8db0f51),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d3ff2),
	.w1(32'h3a305705),
	.w2(32'h3a1c7ff6),
	.w3(32'h39a45fa6),
	.w4(32'h39632af0),
	.w5(32'h395801df),
	.w6(32'h39a2c1ca),
	.w7(32'h3a2d9501),
	.w8(32'h39be3258),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921d3ed),
	.w1(32'h39cc515c),
	.w2(32'h3a13ae82),
	.w3(32'hb7a2f4a6),
	.w4(32'hb8de780b),
	.w5(32'h3951fd66),
	.w6(32'hb8da3428),
	.w7(32'h39c8fa23),
	.w8(32'hbb37c569),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2784d4),
	.w1(32'h379f6ef5),
	.w2(32'hbac49b42),
	.w3(32'hb9b2dd20),
	.w4(32'h3b0cf61d),
	.w5(32'h37851edc),
	.w6(32'hba4da39e),
	.w7(32'hbb046519),
	.w8(32'h3a1a1234),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f0b44),
	.w1(32'h3a46f445),
	.w2(32'h3a8687f6),
	.w3(32'hb794a2de),
	.w4(32'h39a6ced3),
	.w5(32'h3a2014ef),
	.w6(32'hb981f1f2),
	.w7(32'h3a284829),
	.w8(32'h38978be9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d712c),
	.w1(32'hba3cf191),
	.w2(32'hbaa9456a),
	.w3(32'hbb5d8aee),
	.w4(32'hbb119d51),
	.w5(32'hbb18d783),
	.w6(32'hbaf06bda),
	.w7(32'hb9d9950e),
	.w8(32'hba5fe75d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39887382),
	.w1(32'h39e2f9c8),
	.w2(32'h3a0138a3),
	.w3(32'hba1cf4c6),
	.w4(32'hb947e6e9),
	.w5(32'h392e57c4),
	.w6(32'hb99d48cd),
	.w7(32'h3a0b7ff9),
	.w8(32'h391d3e34),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab757a7),
	.w1(32'h3a948d8d),
	.w2(32'h3aa4a8d1),
	.w3(32'h3a69c2c6),
	.w4(32'h3a914ed5),
	.w5(32'h3a6240c8),
	.w6(32'hba1dde39),
	.w7(32'h390bf319),
	.w8(32'hb7f83275),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13d023),
	.w1(32'h3a0e407e),
	.w2(32'h3a412167),
	.w3(32'hb9ed8ebe),
	.w4(32'hb946f40a),
	.w5(32'h39edb902),
	.w6(32'hb98eac39),
	.w7(32'h3a35ea91),
	.w8(32'h3a5e9391),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb5e7),
	.w1(32'h3b6f3b9c),
	.w2(32'h3a2ba0d5),
	.w3(32'h3b939817),
	.w4(32'h3bc4f270),
	.w5(32'h3b8ff413),
	.w6(32'h39bdf486),
	.w7(32'hbb425759),
	.w8(32'hba98349b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d485e),
	.w1(32'hb9f3254d),
	.w2(32'hb96cf607),
	.w3(32'hba9d0299),
	.w4(32'hbac12a8a),
	.w5(32'hba99acf8),
	.w6(32'hbac25585),
	.w7(32'hba14600a),
	.w8(32'h38b8bc88),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d91172),
	.w1(32'h3a2b422a),
	.w2(32'h3a9d1d78),
	.w3(32'hb9da9d19),
	.w4(32'h39f0d905),
	.w5(32'h3a50796c),
	.w6(32'hb80d0cbb),
	.w7(32'h3a8f1d67),
	.w8(32'h39a8106e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42913a),
	.w1(32'hb818e581),
	.w2(32'h3855fcf6),
	.w3(32'hbab6047b),
	.w4(32'hba640f6f),
	.w5(32'hba53d1d1),
	.w6(32'hb9d2e123),
	.w7(32'h39299e73),
	.w8(32'h399d79ce),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa7662),
	.w1(32'hb9baf780),
	.w2(32'hba1f9a79),
	.w3(32'hbb14f9ab),
	.w4(32'hbab61720),
	.w5(32'hbacf4a4b),
	.w6(32'hb9e95ad7),
	.w7(32'h3a71f34b),
	.w8(32'hb8faa909),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d64105),
	.w1(32'h39180ea5),
	.w2(32'hb843b914),
	.w3(32'hba9843f8),
	.w4(32'hb9f5989c),
	.w5(32'hba7c6e93),
	.w6(32'hb9c26ab0),
	.w7(32'h398d1341),
	.w8(32'h39f9a186),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39692a1c),
	.w1(32'h3a6df140),
	.w2(32'h39943c46),
	.w3(32'hba3f3dd4),
	.w4(32'hba869361),
	.w5(32'hba67e65b),
	.w6(32'h398ac4f9),
	.w7(32'hb9f72e4f),
	.w8(32'hbb1e91b4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c72a8a),
	.w1(32'h3bc194b7),
	.w2(32'h3b2c18c3),
	.w3(32'hbb0467f8),
	.w4(32'hbaae0bf7),
	.w5(32'hbbab44f9),
	.w6(32'hb9a76b59),
	.w7(32'hba285a9e),
	.w8(32'hba866ba2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba662136),
	.w1(32'hb9cd3198),
	.w2(32'h37776b92),
	.w3(32'hbb0e064f),
	.w4(32'hbaebe274),
	.w5(32'hba8e0514),
	.w6(32'hbacc9d41),
	.w7(32'hb9c3267a),
	.w8(32'hb8c46a34),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f3c8),
	.w1(32'h3aa4a614),
	.w2(32'h3adbf545),
	.w3(32'h38108073),
	.w4(32'hb9730356),
	.w5(32'hb8b934d3),
	.w6(32'hbae67119),
	.w7(32'hba319e09),
	.w8(32'hbbb39812),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0d0a3),
	.w1(32'hbb59b239),
	.w2(32'hbb8fb292),
	.w3(32'hbbdfcb9e),
	.w4(32'hbb937496),
	.w5(32'hbbb9df04),
	.w6(32'hbb9d701c),
	.w7(32'hbb08426a),
	.w8(32'hba141107),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4616dc),
	.w1(32'hb92af798),
	.w2(32'h3ace4ca3),
	.w3(32'hbb256755),
	.w4(32'hbb0de561),
	.w5(32'hba837716),
	.w6(32'hba90e0b3),
	.w7(32'hba7e2c52),
	.w8(32'h3a5199db),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a461d61),
	.w1(32'h3a85bc48),
	.w2(32'h3abec6b0),
	.w3(32'hba1982e9),
	.w4(32'h39820c8a),
	.w5(32'h3a3235c6),
	.w6(32'hba147e8e),
	.w7(32'h3a223af9),
	.w8(32'h3b18e03b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8cc8c),
	.w1(32'h39a332ab),
	.w2(32'h3b17481d),
	.w3(32'h3b7e10a8),
	.w4(32'h3b63bab8),
	.w5(32'h3ba988b9),
	.w6(32'h3b378112),
	.w7(32'h3b1251eb),
	.w8(32'h39999ed0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1104f),
	.w1(32'h39ca5068),
	.w2(32'h3b195f06),
	.w3(32'h3a1e9e11),
	.w4(32'h3a5c86ab),
	.w5(32'h3b0ee54c),
	.w6(32'hba89e663),
	.w7(32'h3addcf64),
	.w8(32'hbb3734c8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf539a3),
	.w1(32'hb85e8883),
	.w2(32'hbaf4d8c3),
	.w3(32'hbb741cd2),
	.w4(32'hbbb5cee9),
	.w5(32'hbbba0848),
	.w6(32'hbb49c21f),
	.w7(32'hbb80fac8),
	.w8(32'h3b0baa23),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac82fcf),
	.w1(32'h391f79de),
	.w2(32'h3afc0409),
	.w3(32'h3b5c7699),
	.w4(32'h3b45fd16),
	.w5(32'h3b905d50),
	.w6(32'h3b166ff7),
	.w7(32'h3ad9bc1b),
	.w8(32'h3ab8047b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9194e),
	.w1(32'h38e9b94c),
	.w2(32'h3ae84f13),
	.w3(32'h3b3160b6),
	.w4(32'h3b21e012),
	.w5(32'h3b80895b),
	.w6(32'h3aeede65),
	.w7(32'h3ac2e285),
	.w8(32'hb990272c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd073),
	.w1(32'hba7bd523),
	.w2(32'h3905134d),
	.w3(32'hbaa7cb90),
	.w4(32'hbb284a89),
	.w5(32'hbaa2645d),
	.w6(32'hba81cb19),
	.w7(32'hbafe8a79),
	.w8(32'hbb2a99f8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7c29),
	.w1(32'hba0f2789),
	.w2(32'h3a7f83d8),
	.w3(32'hba9c03b5),
	.w4(32'hbaaaf040),
	.w5(32'hbaf392d8),
	.w6(32'h3b33dda8),
	.w7(32'hb85e6cb9),
	.w8(32'hb9722e49),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ded0d),
	.w1(32'h3a3e045a),
	.w2(32'h3a2151a7),
	.w3(32'h39e4be38),
	.w4(32'h39d7c2c3),
	.w5(32'h397e035e),
	.w6(32'h39920ea3),
	.w7(32'h3a0aac58),
	.w8(32'hba356dc4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec5526),
	.w1(32'hba7caa72),
	.w2(32'hbbaf39d7),
	.w3(32'h3b11c81d),
	.w4(32'h3ba69e09),
	.w5(32'hbb273aa1),
	.w6(32'hbac39c74),
	.w7(32'hba9826ea),
	.w8(32'hbadccfc3),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b377ef3),
	.w1(32'h3aa607fa),
	.w2(32'h3ba6641c),
	.w3(32'hbb9fa700),
	.w4(32'hbbc4d691),
	.w5(32'hbb73d90e),
	.w6(32'hbaab3191),
	.w7(32'hbb11711d),
	.w8(32'h3b670238),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3e0e0),
	.w1(32'h3a2f597f),
	.w2(32'h3989ea9c),
	.w3(32'h3ba7a1f9),
	.w4(32'h3bf5c4da),
	.w5(32'h3b69ba78),
	.w6(32'h3b9cf52d),
	.w7(32'h3b6052e6),
	.w8(32'hbb5cf69a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d2c7),
	.w1(32'h3bb49cb3),
	.w2(32'hbad0f301),
	.w3(32'hbbc7fdfb),
	.w4(32'hbbccd58c),
	.w5(32'hbb4f8842),
	.w6(32'hbb6c359d),
	.w7(32'hbb5acc06),
	.w8(32'h397df5d8),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa31d07),
	.w1(32'hb94727af),
	.w2(32'hba2985fc),
	.w3(32'hbadcb09b),
	.w4(32'hba8e3054),
	.w5(32'hbababf87),
	.w6(32'hb9711cd4),
	.w7(32'h3a6a9596),
	.w8(32'h3a828098),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeecc8f),
	.w1(32'h3aa05122),
	.w2(32'h3af47f7a),
	.w3(32'hb86bcf44),
	.w4(32'h3a0e54bf),
	.w5(32'h3abb4e2f),
	.w6(32'hb59d394d),
	.w7(32'h3acf094c),
	.w8(32'hbacace2e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d007),
	.w1(32'hb90a05ff),
	.w2(32'hba32d5e6),
	.w3(32'hbaf0946a),
	.w4(32'hbb561b6a),
	.w5(32'hbae9f3fc),
	.w6(32'hbab267d9),
	.w7(32'hbb221877),
	.w8(32'hb92174bc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaafb0),
	.w1(32'h3a2eab51),
	.w2(32'h3a8c43d9),
	.w3(32'h399703a6),
	.w4(32'h3930d6f3),
	.w5(32'h3a01896c),
	.w6(32'hb7ebae89),
	.w7(32'h3a196f6b),
	.w8(32'h38373576),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d9590f),
	.w1(32'h39ad869c),
	.w2(32'h3a2809f1),
	.w3(32'hbb1264c7),
	.w4(32'hba0918f8),
	.w5(32'hbab8424c),
	.w6(32'hbaadea2d),
	.w7(32'h3923cc99),
	.w8(32'hba8bda1d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a977baa),
	.w1(32'h392aa8a0),
	.w2(32'h3900760f),
	.w3(32'hbb0474af),
	.w4(32'hbb552bcb),
	.w5(32'hbb2c4933),
	.w6(32'hbaccd57a),
	.w7(32'hbb40978f),
	.w8(32'h3a6011c6),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ddb85),
	.w1(32'h391dbcb2),
	.w2(32'h3a572ce9),
	.w3(32'h3ac68a72),
	.w4(32'h3aadff28),
	.w5(32'h3af9bb04),
	.w6(32'h3a8d7b60),
	.w7(32'h3a54c4da),
	.w8(32'h3a52d094),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fce88c),
	.w1(32'h3a58be88),
	.w2(32'h3a9012c5),
	.w3(32'hba29479f),
	.w4(32'h39b1aaf4),
	.w5(32'h3a0781c0),
	.w6(32'h398ed231),
	.w7(32'h39ead927),
	.w8(32'hbab699d5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd14e),
	.w1(32'hbaf0412c),
	.w2(32'hbaa1967e),
	.w3(32'hbaa92e59),
	.w4(32'hbaa8f78e),
	.w5(32'hbb4a98b5),
	.w6(32'hba86be22),
	.w7(32'hb9024976),
	.w8(32'h39deb7cc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e3eb8),
	.w1(32'hb9739d18),
	.w2(32'hb911eb1e),
	.w3(32'h386a7771),
	.w4(32'hb8678e9a),
	.w5(32'hb7447f60),
	.w6(32'h39e2dd1d),
	.w7(32'hb83f1924),
	.w8(32'h3a4545ac),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58dcd7),
	.w1(32'h3a2ee65f),
	.w2(32'h3a0e46dd),
	.w3(32'h39df4604),
	.w4(32'h3a1f55b6),
	.w5(32'h39f26e43),
	.w6(32'h39ce006a),
	.w7(32'h39af4966),
	.w8(32'hba26ec2c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab76b41),
	.w1(32'hbac04166),
	.w2(32'hba74fb88),
	.w3(32'hba823f77),
	.w4(32'hba6f50c0),
	.w5(32'hba3b7452),
	.w6(32'hba425c43),
	.w7(32'hb9d54e61),
	.w8(32'h3aa8bfc4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f2fbfa),
	.w1(32'hbb64d440),
	.w2(32'hbb1c7c7f),
	.w3(32'hba919b90),
	.w4(32'hbb656ccd),
	.w5(32'hbadffe50),
	.w6(32'h3a803368),
	.w7(32'h3a4aa795),
	.w8(32'h3a36b443),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79f713),
	.w1(32'hb9336683),
	.w2(32'h3a6ddf4b),
	.w3(32'h3a800fdc),
	.w4(32'h39a07976),
	.w5(32'h39b9ac08),
	.w6(32'h3a307fb7),
	.w7(32'h3aa39180),
	.w8(32'hb9acb8ea),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c8c8e),
	.w1(32'hba2cbae3),
	.w2(32'hb9e23463),
	.w3(32'hb9cf5579),
	.w4(32'hba142eb3),
	.w5(32'hb986d747),
	.w6(32'hb92effbf),
	.w7(32'hb99777b4),
	.w8(32'h3a4b846c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df546c),
	.w1(32'h39159d46),
	.w2(32'h39ae2bed),
	.w3(32'h3994615b),
	.w4(32'h396a12ff),
	.w5(32'h3982b82f),
	.w6(32'h39c1ee08),
	.w7(32'h39e3af78),
	.w8(32'h394943ab),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862c1dc),
	.w1(32'hb9016b39),
	.w2(32'hb74607d5),
	.w3(32'hb9651ac7),
	.w4(32'hb9890892),
	.w5(32'hb8b4b60e),
	.w6(32'h3555863a),
	.w7(32'hb8052fea),
	.w8(32'h3a11647e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959c99f),
	.w1(32'hb9d997fb),
	.w2(32'hb9636535),
	.w3(32'hba35bbe1),
	.w4(32'hba353bf1),
	.w5(32'hb9b086e1),
	.w6(32'hb94cd9fb),
	.w7(32'hb9726114),
	.w8(32'h3b0056ce),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af11b9a),
	.w1(32'h3ae2471a),
	.w2(32'h3ab7f888),
	.w3(32'h3ae4ee8e),
	.w4(32'h3a29d87c),
	.w5(32'h3abe7b37),
	.w6(32'h3aecb348),
	.w7(32'h3b2c9ee0),
	.w8(32'hba1ce57b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2956b),
	.w1(32'hbaed0a1e),
	.w2(32'hba8f198d),
	.w3(32'hbae3f1ca),
	.w4(32'hbaea678f),
	.w5(32'hba6fd92e),
	.w6(32'hbb08a425),
	.w7(32'hbb002761),
	.w8(32'h3a518c34),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae8d9d),
	.w1(32'hbb5e2ccc),
	.w2(32'hbae45a3f),
	.w3(32'h39fed1b6),
	.w4(32'hbb15b100),
	.w5(32'hbadad759),
	.w6(32'hba52be76),
	.w7(32'h39b08f51),
	.w8(32'hb940db4a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb087480),
	.w1(32'hbb10c6fd),
	.w2(32'hbad25bdd),
	.w3(32'hbac1eec9),
	.w4(32'hbb37e83c),
	.w5(32'hbadaccc3),
	.w6(32'h3907e7ba),
	.w7(32'hb9943cf2),
	.w8(32'h3a3a0055),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cc7c72),
	.w1(32'hb88a4d75),
	.w2(32'h3b0c4e30),
	.w3(32'h39c4ad82),
	.w4(32'h3a9cbb2f),
	.w5(32'h3ab99fd5),
	.w6(32'h3a4b27df),
	.w7(32'h3a89ff88),
	.w8(32'hbaff9c5a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2dc51),
	.w1(32'hba71ecb7),
	.w2(32'h395a82a6),
	.w3(32'h3a8a31f5),
	.w4(32'h39c5fc1a),
	.w5(32'hbaebc151),
	.w6(32'h3a8ac7f1),
	.w7(32'h3b26dec4),
	.w8(32'h3a92641c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39202701),
	.w1(32'h38913426),
	.w2(32'h39b78b71),
	.w3(32'hb794e919),
	.w4(32'h384535a4),
	.w5(32'h37ddefe4),
	.w6(32'h387f5d85),
	.w7(32'h381dcf5d),
	.w8(32'hba82aeff),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d81d6),
	.w1(32'hba2d30ff),
	.w2(32'hba9d293c),
	.w3(32'hba25a243),
	.w4(32'hbac8e807),
	.w5(32'hba6bd1c0),
	.w6(32'hba15f1e3),
	.w7(32'hba4be1f4),
	.w8(32'h390d799a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51d9cf),
	.w1(32'hbaf1bb4d),
	.w2(32'h3a4c1cd2),
	.w3(32'h3a690fca),
	.w4(32'h3a999aae),
	.w5(32'hb6a63827),
	.w6(32'hba3c162a),
	.w7(32'hbaefb0fc),
	.w8(32'h38d50f52),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06b5f0),
	.w1(32'hbb20618d),
	.w2(32'hbb13c5dc),
	.w3(32'hba4ce778),
	.w4(32'hbaba7479),
	.w5(32'hbb0f453b),
	.w6(32'hb9b87d50),
	.w7(32'hba82afeb),
	.w8(32'h3a30f5b8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fd1af),
	.w1(32'h39f02465),
	.w2(32'h39852c86),
	.w3(32'h3a61665a),
	.w4(32'h3a38cc70),
	.w5(32'h39d430c7),
	.w6(32'h3a029933),
	.w7(32'h39831e95),
	.w8(32'hbab9f9da),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7a73a),
	.w1(32'h3a18f29d),
	.w2(32'hbab786cc),
	.w3(32'h3a923eab),
	.w4(32'h3a265f93),
	.w5(32'h3a52d1f5),
	.w6(32'hba1f5ad9),
	.w7(32'h3a2aa62d),
	.w8(32'h39ca0211),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule