module layer_10_featuremap_434(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fd48b),
	.w1(32'hbbc65903),
	.w2(32'hbac7f0d9),
	.w3(32'hbb31ab62),
	.w4(32'hbc1ee755),
	.w5(32'hbb9bdd08),
	.w6(32'hbb2fa146),
	.w7(32'hbc00844e),
	.w8(32'hbb9ac9c7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b010232),
	.w1(32'h3894a2be),
	.w2(32'hbc0434b8),
	.w3(32'h3959a277),
	.w4(32'h3bccc643),
	.w5(32'hbaede1cb),
	.w6(32'h3a2b8748),
	.w7(32'h3b93241a),
	.w8(32'hbb902597),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc555f9c),
	.w1(32'hbb661554),
	.w2(32'hbad1ea8f),
	.w3(32'hbc24f08f),
	.w4(32'hbbbc4b61),
	.w5(32'hba9ee2ed),
	.w6(32'hbc34beac),
	.w7(32'hb93be4a8),
	.w8(32'hbb9ed16c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911cc02),
	.w1(32'hbadb790a),
	.w2(32'h3a9c887d),
	.w3(32'h39c549c9),
	.w4(32'h3a902e7c),
	.w5(32'h3c2106b8),
	.w6(32'h3b07f2a0),
	.w7(32'h3b13d5ab),
	.w8(32'h3bbacc6e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6fb30),
	.w1(32'hbb3e9533),
	.w2(32'hbadb9358),
	.w3(32'h3c3fec89),
	.w4(32'hbb3e10a1),
	.w5(32'hb89e7914),
	.w6(32'h3c10c311),
	.w7(32'hbb7adf7e),
	.w8(32'hba1b643c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892232),
	.w1(32'h3ae9d8c4),
	.w2(32'hbadfc3ac),
	.w3(32'hbb9e096e),
	.w4(32'h3aba1b84),
	.w5(32'hba626d1b),
	.w6(32'hbb6cfefc),
	.w7(32'h3ba81855),
	.w8(32'h3b96c477),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3169a9),
	.w1(32'hbc2b0023),
	.w2(32'hbc4495ef),
	.w3(32'hbb40a626),
	.w4(32'hbc051d07),
	.w5(32'hbc2a6a9c),
	.w6(32'h3a8cf6b9),
	.w7(32'hba0dc26b),
	.w8(32'hba0281be),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292cea),
	.w1(32'hbb569c5c),
	.w2(32'hb9d473da),
	.w3(32'hbbadd3da),
	.w4(32'hbacfadf6),
	.w5(32'hba97e508),
	.w6(32'hbbd39ca8),
	.w7(32'h3b101db0),
	.w8(32'h3b4feb7b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbe54b),
	.w1(32'hba5aaf0f),
	.w2(32'h3bb24613),
	.w3(32'h3b9af726),
	.w4(32'hbb601c28),
	.w5(32'h3b5087fe),
	.w6(32'h3bcadd07),
	.w7(32'hbbace2e6),
	.w8(32'hba83f242),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc787db),
	.w1(32'h3bd16b93),
	.w2(32'h3a99d502),
	.w3(32'hb9653c8e),
	.w4(32'hbb671f86),
	.w5(32'hbbacf51a),
	.w6(32'hbaf395e0),
	.w7(32'hbbe0d281),
	.w8(32'hbbc2f9e0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33153a),
	.w1(32'h3b9706e7),
	.w2(32'h3c1cae44),
	.w3(32'h39c08092),
	.w4(32'hbbc5ef34),
	.w5(32'h3b3b6906),
	.w6(32'hba60dc6b),
	.w7(32'hbbdb36a9),
	.w8(32'hbbaee3cd),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf8eea),
	.w1(32'h3b8a1ca2),
	.w2(32'h3b27f11a),
	.w3(32'h39f45a4a),
	.w4(32'h3c037e97),
	.w5(32'h3c0d5ba8),
	.w6(32'hbb6e2943),
	.w7(32'h3b08647e),
	.w8(32'h3b58d4c2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba492b1),
	.w1(32'hbae4e2db),
	.w2(32'hbc5f4348),
	.w3(32'hbb26e143),
	.w4(32'h3b537932),
	.w5(32'hbc97b435),
	.w6(32'hbb98ffa9),
	.w7(32'hbc220ff6),
	.w8(32'hbcc47c81),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b47d9),
	.w1(32'h3b13aa6d),
	.w2(32'hbb94441e),
	.w3(32'hbcc2af74),
	.w4(32'hbba9077a),
	.w5(32'hbb609241),
	.w6(32'hbcd49722),
	.w7(32'hbc2e9fea),
	.w8(32'hbc4ed7d1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9faa19),
	.w1(32'hbb127993),
	.w2(32'hb90b17f4),
	.w3(32'hbb60e716),
	.w4(32'h3af14133),
	.w5(32'h3b5b2e7f),
	.w6(32'hbc081535),
	.w7(32'h3afd09e8),
	.w8(32'h3a662717),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92962a),
	.w1(32'h3a9b8591),
	.w2(32'h3bb6c042),
	.w3(32'h3b99dbdd),
	.w4(32'h3b8243b0),
	.w5(32'h3b0ff459),
	.w6(32'h3a577d22),
	.w7(32'hba09320a),
	.w8(32'h3a5e8723),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8baef6),
	.w1(32'h3acc5ec5),
	.w2(32'h3a055ae7),
	.w3(32'h3b6e48e4),
	.w4(32'h3bc53ff2),
	.w5(32'h3c040a3f),
	.w6(32'hbb27fc61),
	.w7(32'h3c9ae335),
	.w8(32'h3ca6ab69),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24d7ea),
	.w1(32'hbc2f4bba),
	.w2(32'hbb8487f4),
	.w3(32'h3b46d818),
	.w4(32'hbc1d9203),
	.w5(32'hbb6adb61),
	.w6(32'h3c29b91c),
	.w7(32'hbbc77d9c),
	.w8(32'hbb210fd5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6834be),
	.w1(32'h3aa0482b),
	.w2(32'h3bb3f491),
	.w3(32'h3b65571c),
	.w4(32'h3b583aa2),
	.w5(32'h3c17dd7c),
	.w6(32'h3bc86711),
	.w7(32'h3b3967a2),
	.w8(32'h3c0446bb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde23fb),
	.w1(32'h3a8ef269),
	.w2(32'hba9cd870),
	.w3(32'h3bcb09b4),
	.w4(32'h3bcbbc9c),
	.w5(32'h3534be5c),
	.w6(32'h3bb3ba58),
	.w7(32'h3b9f3114),
	.w8(32'h3b373a52),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f33c3),
	.w1(32'hbaf79d6c),
	.w2(32'hbbdabed8),
	.w3(32'hbb5a29cd),
	.w4(32'hbb8a6970),
	.w5(32'hbbcfafb5),
	.w6(32'hbbe54c78),
	.w7(32'hbb3ab5a8),
	.w8(32'hbbce1dcb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65c427),
	.w1(32'h3b063c2f),
	.w2(32'hbbc70d43),
	.w3(32'h3b1becdc),
	.w4(32'h3c179ea2),
	.w5(32'hba9d8de9),
	.w6(32'h3b1be911),
	.w7(32'h3b803893),
	.w8(32'hbb2f3f79),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f18d8),
	.w1(32'hb9a56e0e),
	.w2(32'hbb2d7fe4),
	.w3(32'hbb4b5a2b),
	.w4(32'h3ae6e67f),
	.w5(32'h3b7e31e0),
	.w6(32'h3a0bb4fb),
	.w7(32'hba8bf09d),
	.w8(32'h3b000884),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24466f),
	.w1(32'h3aa5a706),
	.w2(32'h3b00ea62),
	.w3(32'hb9482cec),
	.w4(32'h3c88fcd6),
	.w5(32'h3c8c0df8),
	.w6(32'h3ac22206),
	.w7(32'h3ae970d2),
	.w8(32'h3b39d991),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43be5e),
	.w1(32'hbb446fdd),
	.w2(32'hbbd876fc),
	.w3(32'h3abaa928),
	.w4(32'h3b37ab50),
	.w5(32'h3b831629),
	.w6(32'hbc2a970b),
	.w7(32'hbae2c215),
	.w8(32'hbb630fc7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ec310),
	.w1(32'hbbe03bc1),
	.w2(32'hbbe70c15),
	.w3(32'h3a3e36bb),
	.w4(32'hbba27dec),
	.w5(32'hbc305d31),
	.w6(32'hbb3ab10b),
	.w7(32'h3a007303),
	.w8(32'hbb0584d9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d0135),
	.w1(32'hbba55f40),
	.w2(32'hbbdfc3e1),
	.w3(32'h3af9ac33),
	.w4(32'hbc268a9d),
	.w5(32'hbc4fb391),
	.w6(32'h3bd4cc15),
	.w7(32'hbb54e0d5),
	.w8(32'hbbabca9b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacb1ad),
	.w1(32'hbc2455c4),
	.w2(32'hbb11d552),
	.w3(32'hbc20fde5),
	.w4(32'hbbd496da),
	.w5(32'h3b062dc3),
	.w6(32'hbb4dec3a),
	.w7(32'hbba1e8d7),
	.w8(32'h3bc6c1a9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc7ae),
	.w1(32'hba6a6979),
	.w2(32'hbb96fc42),
	.w3(32'h3847651b),
	.w4(32'hbb9c3397),
	.w5(32'hbaca3cea),
	.w6(32'hb8f7823a),
	.w7(32'hbb4cf5f2),
	.w8(32'h3bc011e5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b6384),
	.w1(32'hbaecf756),
	.w2(32'hba389fd2),
	.w3(32'hbb2eadab),
	.w4(32'hbb48266e),
	.w5(32'hbae39b8d),
	.w6(32'h3c0ae602),
	.w7(32'hbb6cfefc),
	.w8(32'hbb28f07a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa61eba),
	.w1(32'h398ff890),
	.w2(32'hbba2595e),
	.w3(32'hb9c1a077),
	.w4(32'hbac6f51b),
	.w5(32'hbb8e67e0),
	.w6(32'hbaf1f77b),
	.w7(32'h391c2ceb),
	.w8(32'h36309725),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb105ebc),
	.w1(32'h39f15591),
	.w2(32'hbb89b7a2),
	.w3(32'hbadd2eb0),
	.w4(32'hbbd5d447),
	.w5(32'hbbc95677),
	.w6(32'hbb4bc9dc),
	.w7(32'h3b142505),
	.w8(32'hbb4dea5d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dda3f),
	.w1(32'hba5da69c),
	.w2(32'hbbb16fdc),
	.w3(32'hbc2aa6a2),
	.w4(32'h39a93391),
	.w5(32'hbb325f5a),
	.w6(32'hbb874429),
	.w7(32'h3b10ce85),
	.w8(32'h3b19115c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbf24e),
	.w1(32'hbbd4bdd4),
	.w2(32'hbbe472ad),
	.w3(32'hbacd04ee),
	.w4(32'hbbc68ef7),
	.w5(32'hbbf5519e),
	.w6(32'h3b510453),
	.w7(32'hbb96844f),
	.w8(32'h3a48ac7c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d187b),
	.w1(32'hbb73d34c),
	.w2(32'hbb2bdbdb),
	.w3(32'h37ac68c9),
	.w4(32'hbb0daf6a),
	.w5(32'h3acd9103),
	.w6(32'hbae0d9da),
	.w7(32'hbbbd218d),
	.w8(32'h3b835737),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b370f),
	.w1(32'h3aa90909),
	.w2(32'h38bacddb),
	.w3(32'h3affdc6a),
	.w4(32'h3a0b41d0),
	.w5(32'hba7817be),
	.w6(32'hb9550689),
	.w7(32'hbb47bacf),
	.w8(32'hbbf6b80c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabca42a),
	.w1(32'hbbe00b7f),
	.w2(32'hbbef6529),
	.w3(32'hbb1cf54d),
	.w4(32'hbc161ba5),
	.w5(32'hbbbddd89),
	.w6(32'hbb2e6e5a),
	.w7(32'hbbbc1667),
	.w8(32'hbbf32612),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f383),
	.w1(32'h3b618ec5),
	.w2(32'hbc6167f4),
	.w3(32'h3b403387),
	.w4(32'hbb850727),
	.w5(32'hbc83758a),
	.w6(32'h3b331835),
	.w7(32'hbaeb2524),
	.w8(32'hbc62771e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc799995),
	.w1(32'hbc01f2ee),
	.w2(32'hbad1f1f1),
	.w3(32'hbc928cd3),
	.w4(32'hbc4f1af1),
	.w5(32'hbbd3f634),
	.w6(32'hbc5472ba),
	.w7(32'hbc84b46f),
	.w8(32'hbc4dccac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cf9f8),
	.w1(32'h3b93d3ca),
	.w2(32'h3b3918b2),
	.w3(32'h3b252023),
	.w4(32'h3b3762d0),
	.w5(32'h3aef77c4),
	.w6(32'hbbcc5c64),
	.w7(32'h3bb9b10c),
	.w8(32'h3b9485a5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e85a2),
	.w1(32'hba383f22),
	.w2(32'hb8906875),
	.w3(32'h3aead481),
	.w4(32'h39082c7b),
	.w5(32'h39d8b868),
	.w6(32'h3be55072),
	.w7(32'hb95d65f1),
	.w8(32'h3bf4715a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf86cd),
	.w1(32'h3b93c4e0),
	.w2(32'h3b4d2bf5),
	.w3(32'hbbbb0923),
	.w4(32'h3b611931),
	.w5(32'h3c000a1b),
	.w6(32'hbb399098),
	.w7(32'h3a5b4cec),
	.w8(32'hb8e0567c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad63124),
	.w1(32'h39c4220b),
	.w2(32'h3aa3d8c0),
	.w3(32'h3b88c0e1),
	.w4(32'h3b792e1c),
	.w5(32'h3ba51ab5),
	.w6(32'hbaa1a8ab),
	.w7(32'h39c45fe7),
	.w8(32'hba5e729d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4529),
	.w1(32'hbb949ece),
	.w2(32'hbafc9646),
	.w3(32'h3aad6add),
	.w4(32'hbb27d781),
	.w5(32'h3816bfaf),
	.w6(32'h3aa37b35),
	.w7(32'h3a074b1a),
	.w8(32'h3ba5b574),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8805f),
	.w1(32'hb8dd56f9),
	.w2(32'h3b32921a),
	.w3(32'h3c45b1db),
	.w4(32'h3b58e25a),
	.w5(32'h3b9fe41c),
	.w6(32'h3c74fa49),
	.w7(32'h3b1cd83d),
	.w8(32'h3b84d5cd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2027fd),
	.w1(32'h3bd63d26),
	.w2(32'h3c2ce55f),
	.w3(32'h3abdf3c1),
	.w4(32'h3bb0dd28),
	.w5(32'h3bbceb7b),
	.w6(32'h39b8c971),
	.w7(32'h3ab7e3a2),
	.w8(32'h3b725833),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe8d69),
	.w1(32'hbb77dcce),
	.w2(32'hbb4b45c6),
	.w3(32'h3baa7f4f),
	.w4(32'hbc119827),
	.w5(32'hbc3babe0),
	.w6(32'h38856516),
	.w7(32'hbc9cc968),
	.w8(32'hbcb85c2b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0b99),
	.w1(32'hba85fa2a),
	.w2(32'h3b2fd02b),
	.w3(32'hbbfa81c3),
	.w4(32'hbbe24a66),
	.w5(32'hba40ecf7),
	.w6(32'hbc8d68eb),
	.w7(32'hbae87db9),
	.w8(32'h3a90e119),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f0fc7),
	.w1(32'hbb888cb8),
	.w2(32'h3aa1f0ff),
	.w3(32'h3b8cddca),
	.w4(32'hbb408a46),
	.w5(32'h3b744f63),
	.w6(32'h3b27f644),
	.w7(32'hbc062978),
	.w8(32'h39c54878),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53bffd),
	.w1(32'hbae067ba),
	.w2(32'h3b913aa6),
	.w3(32'h3a35f5f8),
	.w4(32'hbbd631f1),
	.w5(32'h3aa1d6e5),
	.w6(32'h3b5cce76),
	.w7(32'h3ae64025),
	.w8(32'h3b80cf95),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b096127),
	.w1(32'hbad048f5),
	.w2(32'h3a8e45f2),
	.w3(32'h3bae2575),
	.w4(32'hbb21c9d5),
	.w5(32'h3bfb1e2f),
	.w6(32'h3abb0588),
	.w7(32'hbb4547d1),
	.w8(32'h3ba193c1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75b312),
	.w1(32'hbb63fcf3),
	.w2(32'h3b7f654a),
	.w3(32'h3b2cc6fe),
	.w4(32'hba5dc3f0),
	.w5(32'h3bb2c70a),
	.w6(32'h3ae53aa8),
	.w7(32'hbb6d2b68),
	.w8(32'hba77c7aa),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2249c5),
	.w1(32'hba765ad0),
	.w2(32'hb917a48e),
	.w3(32'h3bcd30d2),
	.w4(32'hbb9f5693),
	.w5(32'hbae6f50b),
	.w6(32'hba422c7b),
	.w7(32'hbbdb5092),
	.w8(32'hbb0c4203),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc86022),
	.w1(32'h3ba7117e),
	.w2(32'hbb259861),
	.w3(32'h3b6fb099),
	.w4(32'h3bde11dd),
	.w5(32'h3b3b10e1),
	.w6(32'hbb3e9fed),
	.w7(32'h3b7e0391),
	.w8(32'h3b2df529),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba54e56),
	.w1(32'h3b8ee51f),
	.w2(32'hbb99a1cc),
	.w3(32'h3b376f44),
	.w4(32'hb9dbea90),
	.w5(32'hbb93f870),
	.w6(32'h3b724a7f),
	.w7(32'h3b80702c),
	.w8(32'hbb9393d0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b6ec),
	.w1(32'h3bcff339),
	.w2(32'h3c0a1da8),
	.w3(32'hbbb31be5),
	.w4(32'h3bf80a4b),
	.w5(32'h3c587edd),
	.w6(32'h3a4eedc1),
	.w7(32'h39334de6),
	.w8(32'h3ad93436),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2038d6),
	.w1(32'h3b875581),
	.w2(32'h3a230511),
	.w3(32'h3c610e8f),
	.w4(32'h3b45cc42),
	.w5(32'hbb09991d),
	.w6(32'h3c0c6e16),
	.w7(32'h3aab34ef),
	.w8(32'hbac8cbe4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15952),
	.w1(32'hbb322fbb),
	.w2(32'hbbce97bf),
	.w3(32'hbbc67f20),
	.w4(32'h3b2ba5b2),
	.w5(32'hbc08246a),
	.w6(32'hbbf1f60b),
	.w7(32'h38c261a7),
	.w8(32'hbb8a9e22),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2e0d3),
	.w1(32'h3b9a8c7b),
	.w2(32'hba927e73),
	.w3(32'hbbbac130),
	.w4(32'h3c741446),
	.w5(32'h3c0fb345),
	.w6(32'hbb95dcc2),
	.w7(32'h3c40e8eb),
	.w8(32'h3c0c4b18),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab98cdf),
	.w1(32'hbac6d4e0),
	.w2(32'hbb918bbf),
	.w3(32'h3c003a16),
	.w4(32'hba9cad24),
	.w5(32'hbb85c7b4),
	.w6(32'h3c32474f),
	.w7(32'hbb8c4674),
	.w8(32'hbbf3391a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd482d),
	.w1(32'hbb1a48fe),
	.w2(32'hbb36c012),
	.w3(32'h3ac13e2e),
	.w4(32'hbbd2623e),
	.w5(32'hbc3cca57),
	.w6(32'hbb1c50c7),
	.w7(32'hbafc224a),
	.w8(32'hbb904080),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf6711),
	.w1(32'h39008ddb),
	.w2(32'h3a9c1e41),
	.w3(32'h3a93a68a),
	.w4(32'h3b4ebcc6),
	.w5(32'h3bc09bb8),
	.w6(32'h3b9d92d6),
	.w7(32'h3c047bcb),
	.w8(32'h3bba847b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49734b),
	.w1(32'h3bd400e4),
	.w2(32'h3c30a553),
	.w3(32'h3af8b8b5),
	.w4(32'h3c565680),
	.w5(32'h3c9dbcf5),
	.w6(32'h3a8ccdd8),
	.w7(32'h3c09aaf5),
	.w8(32'h3c386d69),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a925c83),
	.w1(32'h3c01e19f),
	.w2(32'h3c177d31),
	.w3(32'h3a8e6503),
	.w4(32'h3c22a955),
	.w5(32'h3c423f37),
	.w6(32'h3b771cca),
	.w7(32'h3aebc34b),
	.w8(32'h3b63a327),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35963f),
	.w1(32'hbbc76fb5),
	.w2(32'hb9555472),
	.w3(32'hbb0e7058),
	.w4(32'hbb21a583),
	.w5(32'h3aa5366d),
	.w6(32'hbb5b47d9),
	.w7(32'hbc1a00b2),
	.w8(32'hbb4f295e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad88fe8),
	.w1(32'hbc07392d),
	.w2(32'hbc1080eb),
	.w3(32'h3ba70a82),
	.w4(32'hbbbba387),
	.w5(32'hbb24c3f5),
	.w6(32'h3ab52959),
	.w7(32'hbbc3783e),
	.w8(32'hbbe87eb0),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a82ac),
	.w1(32'h3c68178b),
	.w2(32'h3c0ca650),
	.w3(32'h3b1bc872),
	.w4(32'h3b88c207),
	.w5(32'h3a25d21f),
	.w6(32'hbb97efcf),
	.w7(32'h3b545f13),
	.w8(32'h3983fe15),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9cb47),
	.w1(32'h3a930035),
	.w2(32'h3bfaf6db),
	.w3(32'hbb411f1b),
	.w4(32'h3bc6235f),
	.w5(32'h3bc6f090),
	.w6(32'hbb909655),
	.w7(32'h3bbe1f1f),
	.w8(32'h3beb9ab1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befa204),
	.w1(32'hbbae199d),
	.w2(32'hbb7570fc),
	.w3(32'h3c335949),
	.w4(32'hbbedfecb),
	.w5(32'hbbaf7fe9),
	.w6(32'h3bd957ad),
	.w7(32'hbb869470),
	.w8(32'hbb97b27e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1560fb),
	.w1(32'hbafc18c0),
	.w2(32'hba92d305),
	.w3(32'h3b9a5d52),
	.w4(32'h3ad51b83),
	.w5(32'h3b30e114),
	.w6(32'h3bbd05b4),
	.w7(32'h3b0ee18b),
	.w8(32'h3ad5a3f2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa12a9c),
	.w1(32'hbb0cfb8a),
	.w2(32'hbb0493e0),
	.w3(32'h3b8803d2),
	.w4(32'hbb550132),
	.w5(32'hbb7cb2f3),
	.w6(32'h3ae9fdff),
	.w7(32'hbb1f68e6),
	.w8(32'hb9968118),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3da5b),
	.w1(32'h3b6878a7),
	.w2(32'h3a63ec4d),
	.w3(32'hbb3e353b),
	.w4(32'h3aa9c847),
	.w5(32'h3a17b7af),
	.w6(32'hb803406d),
	.w7(32'hbba627b4),
	.w8(32'hbb9b3020),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e38f3),
	.w1(32'hba151eeb),
	.w2(32'hba7ed404),
	.w3(32'hbb3f2ca7),
	.w4(32'h3b1507fc),
	.w5(32'h3b305bd8),
	.w6(32'hbad5ffd7),
	.w7(32'h3b10472e),
	.w8(32'hbb11ae1d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a828282),
	.w1(32'hbb83a578),
	.w2(32'hbb74fa18),
	.w3(32'h3b1afcc1),
	.w4(32'hbb2f7131),
	.w5(32'hbad6e1f9),
	.w6(32'h3b3eaa6e),
	.w7(32'hbb2d062c),
	.w8(32'hbac84b4f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab87520),
	.w1(32'hbb273c86),
	.w2(32'hbae90d02),
	.w3(32'hbaabec6d),
	.w4(32'hbb03b5a6),
	.w5(32'hbb0dfe1a),
	.w6(32'hba52fb0a),
	.w7(32'hbaae630f),
	.w8(32'hbac3c54d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280d48),
	.w1(32'h3affcf13),
	.w2(32'h3a278b37),
	.w3(32'hbb914491),
	.w4(32'h3b02da5e),
	.w5(32'h39dd409e),
	.w6(32'hbb9e2dac),
	.w7(32'h3a7c211a),
	.w8(32'h3b0c21af),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74adc6),
	.w1(32'hba901b28),
	.w2(32'hbb215e7e),
	.w3(32'h3a7a5cef),
	.w4(32'hb952aa34),
	.w5(32'h3ad3ad96),
	.w6(32'h3add8a2c),
	.w7(32'h391ad49b),
	.w8(32'h3a0426b9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9744),
	.w1(32'hbb5d9009),
	.w2(32'hbb86d21f),
	.w3(32'hbaafc593),
	.w4(32'hbb0e192b),
	.w5(32'hbac8f473),
	.w6(32'hbb7ed2b9),
	.w7(32'hb6ea448f),
	.w8(32'hbb4ee467),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939de24),
	.w1(32'h3a9a7027),
	.w2(32'h38012cb3),
	.w3(32'hbb5b259c),
	.w4(32'h3ba8ebcd),
	.w5(32'hb9aae933),
	.w6(32'hbba5f86d),
	.w7(32'h3b5c4aaf),
	.w8(32'hba347b27),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0925dd),
	.w1(32'hba21b1c6),
	.w2(32'h39417c69),
	.w3(32'h3b47b345),
	.w4(32'hbb0d2ed2),
	.w5(32'hba3db43c),
	.w6(32'hbab7cb04),
	.w7(32'hbb386410),
	.w8(32'hbb6e62c4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07b5b2),
	.w1(32'h3b8074ca),
	.w2(32'hb9b0bdef),
	.w3(32'hbaa1d904),
	.w4(32'h3b5a582a),
	.w5(32'h3adb9241),
	.w6(32'hbb2f1b58),
	.w7(32'h3b75ab75),
	.w8(32'h3a336ac5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cd88b),
	.w1(32'h378b812e),
	.w2(32'hbaab2b1e),
	.w3(32'h3b96e9e2),
	.w4(32'h3a847a68),
	.w5(32'hb8a0b8c4),
	.w6(32'h3a39e2f3),
	.w7(32'h3af4419a),
	.w8(32'h38d49b4b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd019),
	.w1(32'h378bd2d2),
	.w2(32'hb8826ab1),
	.w3(32'hba8ef250),
	.w4(32'hb9ba96e5),
	.w5(32'hbb4f49df),
	.w6(32'hba6cf0cd),
	.w7(32'hbb7816f7),
	.w8(32'hbb731540),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4e5b),
	.w1(32'hbaa9fbe2),
	.w2(32'hbb0998f5),
	.w3(32'hbb90f244),
	.w4(32'h3b4c5c96),
	.w5(32'h3b9e68d7),
	.w6(32'hbb65215c),
	.w7(32'h3b3f697d),
	.w8(32'h3a3c6c22),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f199d6),
	.w1(32'hb987a6af),
	.w2(32'hbb30c387),
	.w3(32'h3b8d5f4e),
	.w4(32'h3aa2ffbf),
	.w5(32'h3a302857),
	.w6(32'h3a2a1ca9),
	.w7(32'h3990844c),
	.w8(32'hba1da340),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c1d9e),
	.w1(32'hbb86ed2b),
	.w2(32'hbb424766),
	.w3(32'hbaebb925),
	.w4(32'hbb24fc1f),
	.w5(32'h3a1e7161),
	.w6(32'hb892db33),
	.w7(32'hb98027db),
	.w8(32'hba8d58eb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb167301),
	.w1(32'h3ad0682d),
	.w2(32'h391b0cde),
	.w3(32'hb9ee6da7),
	.w4(32'h3911231b),
	.w5(32'hbaccb384),
	.w6(32'h394e1d8f),
	.w7(32'h3b1f8abb),
	.w8(32'hbb07d84d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9038f2),
	.w1(32'h3b06798c),
	.w2(32'h3af6e5d3),
	.w3(32'h3927792d),
	.w4(32'h3a7607ad),
	.w5(32'h3b10d04e),
	.w6(32'hbaeff00f),
	.w7(32'hba9d8860),
	.w8(32'hbb862c02),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7fc0e),
	.w1(32'hbab3995d),
	.w2(32'hbb742f5f),
	.w3(32'hb9d5fdd3),
	.w4(32'h39a6259c),
	.w5(32'hbafc8431),
	.w6(32'h38e7db1b),
	.w7(32'hba71fd92),
	.w8(32'hba84c518),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb151737),
	.w1(32'hbb4c0831),
	.w2(32'hbb25d827),
	.w3(32'hbaa2dd62),
	.w4(32'hbb162a98),
	.w5(32'hbb4a8eb5),
	.w6(32'hbb253e68),
	.w7(32'h3a11304a),
	.w8(32'hba97ec88),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56ac3c),
	.w1(32'hbadaee36),
	.w2(32'hbb91609d),
	.w3(32'hb9ae247a),
	.w4(32'hbb345286),
	.w5(32'hbb18a861),
	.w6(32'hbb290377),
	.w7(32'hbb53b7d6),
	.w8(32'hbb808dd9),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843e54),
	.w1(32'hbb327bfb),
	.w2(32'hbb3c21a7),
	.w3(32'hbba7c3e3),
	.w4(32'hbb11ded3),
	.w5(32'hba049339),
	.w6(32'hbbc040ef),
	.w7(32'hba965fcf),
	.w8(32'hb9a08674),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09ccdd),
	.w1(32'h3b105ed6),
	.w2(32'h3babae82),
	.w3(32'hbb70c233),
	.w4(32'h3bad2aae),
	.w5(32'h3b8dd917),
	.w6(32'hbac42a76),
	.w7(32'h3a1679c4),
	.w8(32'h3b1daab3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d9f03),
	.w1(32'h39d5b57c),
	.w2(32'h3b30d774),
	.w3(32'h3b1578c2),
	.w4(32'h3abd1bdd),
	.w5(32'h3b0da11a),
	.w6(32'h3a9058d2),
	.w7(32'h3abe2c1e),
	.w8(32'h3a8cfc3e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4817f9),
	.w1(32'hb9ed98c8),
	.w2(32'hbaa66937),
	.w3(32'h3b2137a9),
	.w4(32'hba3750a9),
	.w5(32'h39ba0dac),
	.w6(32'h3b12e611),
	.w7(32'hba03b73d),
	.w8(32'hba691115),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff32df),
	.w1(32'hba8069d8),
	.w2(32'h3aa4e912),
	.w3(32'hbbb2e6bb),
	.w4(32'hbb844db3),
	.w5(32'hbb135f28),
	.w6(32'hbb365f9b),
	.w7(32'hbbfc544e),
	.w8(32'hbb5fcd4c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285b85),
	.w1(32'h3ab8b9a1),
	.w2(32'hb9da35a7),
	.w3(32'hb9b33351),
	.w4(32'h3aab52a8),
	.w5(32'h3a436b55),
	.w6(32'hbad24509),
	.w7(32'h3a2f5c20),
	.w8(32'hbb4d6e96),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9152f2),
	.w1(32'h3809903f),
	.w2(32'hba6ad19f),
	.w3(32'hbae96115),
	.w4(32'hbb0bb141),
	.w5(32'h3b2c885b),
	.w6(32'h3a5cf9bb),
	.w7(32'hbb596d91),
	.w8(32'h3b3efd6c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb567781),
	.w1(32'hba549156),
	.w2(32'hbb2429ea),
	.w3(32'h3b5ec640),
	.w4(32'h389fb344),
	.w5(32'h387f2266),
	.w6(32'h3b07a6e2),
	.w7(32'hbae0fdfa),
	.w8(32'hba98cfa3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a794f),
	.w1(32'hbbe310b3),
	.w2(32'hbbb3874c),
	.w3(32'hba21f434),
	.w4(32'hbba1a713),
	.w5(32'hbb3cc11c),
	.w6(32'hbb0ea2a2),
	.w7(32'h3b50ae42),
	.w8(32'h3b047fbd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb711083),
	.w1(32'h3b4e72f1),
	.w2(32'h39b33b87),
	.w3(32'hbb63aa47),
	.w4(32'h3af114e9),
	.w5(32'hba3d9ef8),
	.w6(32'hbabe4703),
	.w7(32'hba5242d8),
	.w8(32'hbb85f8b6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39946af6),
	.w1(32'hbb3b47b7),
	.w2(32'hbaf1df43),
	.w3(32'hbab76d1b),
	.w4(32'hbab3789b),
	.w5(32'hbb23dea1),
	.w6(32'h3926a5ad),
	.w7(32'h3a91e55c),
	.w8(32'hb90abf8c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ece214),
	.w1(32'h3b0f75b8),
	.w2(32'h3b2bb9a4),
	.w3(32'hba22fb13),
	.w4(32'hbacff214),
	.w5(32'h39aae388),
	.w6(32'hbad2af5f),
	.w7(32'hbb0875b9),
	.w8(32'hbaa29c23),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1323a),
	.w1(32'h39bd35c8),
	.w2(32'hbb2a33eb),
	.w3(32'h3a33b792),
	.w4(32'h3b4747ee),
	.w5(32'hbabb927e),
	.w6(32'h3a8e7957),
	.w7(32'h3b83df4c),
	.w8(32'hba5159f3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fda39),
	.w1(32'hb9ae3603),
	.w2(32'h3b2c0e44),
	.w3(32'hbad033f7),
	.w4(32'h3b21e4f9),
	.w5(32'h3ac73eba),
	.w6(32'h3a087983),
	.w7(32'hb9d61efb),
	.w8(32'h3855b8ae),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb130757),
	.w1(32'h3af580b4),
	.w2(32'hb9ac1e5b),
	.w3(32'hbb1edd77),
	.w4(32'h3b1e5d35),
	.w5(32'h3a1b401b),
	.w6(32'hba12f990),
	.w7(32'h3ad2bed9),
	.w8(32'h3a82ba97),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fc01f),
	.w1(32'hb8e81f98),
	.w2(32'h3a01c2ea),
	.w3(32'hb94eac85),
	.w4(32'h3a73793a),
	.w5(32'hba744ec6),
	.w6(32'h39c258cc),
	.w7(32'h3a4360f8),
	.w8(32'hba137d17),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bb062),
	.w1(32'hbb6dc9e7),
	.w2(32'hbb721ca2),
	.w3(32'hbad17e72),
	.w4(32'hbb3bec8a),
	.w5(32'h3ac1a0ce),
	.w6(32'hbb0d995d),
	.w7(32'hbb6b11a9),
	.w8(32'hb9f6fe93),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35428a),
	.w1(32'hb823f868),
	.w2(32'h3ac07c04),
	.w3(32'hbb4ca217),
	.w4(32'h3a6225b1),
	.w5(32'hbaabb93e),
	.w6(32'hbadc81d9),
	.w7(32'h39994988),
	.w8(32'hbb13a9dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba655163),
	.w1(32'hbaac6f40),
	.w2(32'h3b3bf5b9),
	.w3(32'hbb3b5c97),
	.w4(32'hbad8e9a9),
	.w5(32'hba0bfccc),
	.w6(32'hba2a660d),
	.w7(32'hbb25e836),
	.w8(32'hba563d36),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba711a1c),
	.w1(32'h3a7ba0aa),
	.w2(32'hbafa54c5),
	.w3(32'hbbcc882a),
	.w4(32'hb9245e0b),
	.w5(32'hb8ba4aee),
	.w6(32'hbba05b17),
	.w7(32'hbb1eba9d),
	.w8(32'hbaed1ca5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28493f),
	.w1(32'hbb47ccbc),
	.w2(32'hbb9e85e4),
	.w3(32'h3a52f152),
	.w4(32'hbb5f48d1),
	.w5(32'hbb84aa29),
	.w6(32'hba653dbf),
	.w7(32'hba8aa186),
	.w8(32'hbaf19ab1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaccc33),
	.w1(32'h389674fd),
	.w2(32'h3a01802d),
	.w3(32'hba96658b),
	.w4(32'hbaf8a2c5),
	.w5(32'h3b778bae),
	.w6(32'hbaf257c9),
	.w7(32'hb93b14c9),
	.w8(32'hb9cb3d56),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a6dd9),
	.w1(32'h3a372ee8),
	.w2(32'h393fc178),
	.w3(32'h3a31f0eb),
	.w4(32'h3b817276),
	.w5(32'hba9f246a),
	.w6(32'hba338edb),
	.w7(32'h3b6ca93e),
	.w8(32'h3944c0f0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b53ef),
	.w1(32'h3afbe2fe),
	.w2(32'h3ad9bbfc),
	.w3(32'h3995cbfe),
	.w4(32'h39cbb295),
	.w5(32'hb7ed1ebc),
	.w6(32'hbadb93b2),
	.w7(32'hba950ae4),
	.w8(32'hbafa9c9f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba463942),
	.w1(32'hbaa607cf),
	.w2(32'hbb52e2e8),
	.w3(32'hb9ea86e0),
	.w4(32'hb99acc58),
	.w5(32'hbb77d0ba),
	.w6(32'hba0330e3),
	.w7(32'hba64425e),
	.w8(32'hbacb156f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0b653),
	.w1(32'h3b7ceb53),
	.w2(32'h3b6de8fa),
	.w3(32'hba8134a5),
	.w4(32'h3b5523ba),
	.w5(32'h3bb8c096),
	.w6(32'h3a584263),
	.w7(32'hbb09ad51),
	.w8(32'h37e998bd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd4221),
	.w1(32'h3a47939d),
	.w2(32'h3bb3caab),
	.w3(32'hbad53779),
	.w4(32'h3b0b954b),
	.w5(32'h3b8b685c),
	.w6(32'hbb570bb1),
	.w7(32'h3ab4710d),
	.w8(32'h3b961fd0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b2c4c),
	.w1(32'h393e82fb),
	.w2(32'hbac5b4dd),
	.w3(32'h3ab67586),
	.w4(32'hba663342),
	.w5(32'hba92eff7),
	.w6(32'h3acf20f3),
	.w7(32'hba016f93),
	.w8(32'hbb0ee0e0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1858ba),
	.w1(32'h3c26ee40),
	.w2(32'h3bd9e94f),
	.w3(32'hbad3c57b),
	.w4(32'h3ba2883b),
	.w5(32'h3bdf9ca7),
	.w6(32'hbb160a9f),
	.w7(32'h3aff90bb),
	.w8(32'h3b56da2f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8cfb2),
	.w1(32'h37865244),
	.w2(32'hbaf16f76),
	.w3(32'hbad7cafa),
	.w4(32'h3b783ac5),
	.w5(32'h3b19a5ce),
	.w6(32'h3a2a6ca7),
	.w7(32'h3b4cc1ed),
	.w8(32'h3ab4395b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85022e7),
	.w1(32'hbb93061b),
	.w2(32'hbb35f937),
	.w3(32'h3ab41c7d),
	.w4(32'hbb073695),
	.w5(32'hbb12f2e7),
	.w6(32'hba8cad3a),
	.w7(32'hbb935f9f),
	.w8(32'hb9063112),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392defa0),
	.w1(32'h3a4ed681),
	.w2(32'h391261ed),
	.w3(32'hba5aab35),
	.w4(32'hbb48dc41),
	.w5(32'hbb2e8467),
	.w6(32'h3ac11354),
	.w7(32'hbb3789a1),
	.w8(32'hbb86da60),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f808f),
	.w1(32'hbb305869),
	.w2(32'hbb9e3c4a),
	.w3(32'hbb803b88),
	.w4(32'hbafffc6b),
	.w5(32'hbb1f04af),
	.w6(32'hbae17ffe),
	.w7(32'hbaa63bad),
	.w8(32'hbb700572),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7be400),
	.w1(32'hbb171029),
	.w2(32'hba20d6ff),
	.w3(32'hbb2c0e49),
	.w4(32'hbaed7605),
	.w5(32'hbac73314),
	.w6(32'hbaff4637),
	.w7(32'hbb921feb),
	.w8(32'hbb920ce0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e37d6),
	.w1(32'h3a15c75d),
	.w2(32'h3ae2dc78),
	.w3(32'hbba34d63),
	.w4(32'h3b1c190b),
	.w5(32'h3b25bb94),
	.w6(32'hbb9e20d2),
	.w7(32'h3a61a9d6),
	.w8(32'h39eb1f42),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf55cc),
	.w1(32'hbc155b25),
	.w2(32'hbbe2c3f5),
	.w3(32'h3adbd4c4),
	.w4(32'hbbb74ccb),
	.w5(32'hbba73145),
	.w6(32'h3a52bf08),
	.w7(32'hbb07d3a0),
	.w8(32'h3a7fc870),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3027fb),
	.w1(32'h38208c65),
	.w2(32'hbaadfd47),
	.w3(32'hbaab50ee),
	.w4(32'hbadeea3c),
	.w5(32'hb99566ed),
	.w6(32'h3969b5e0),
	.w7(32'hbaf6e0d5),
	.w8(32'hba7579fa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0062b1),
	.w1(32'h391ed607),
	.w2(32'hba24fc74),
	.w3(32'hba6eafbb),
	.w4(32'hbb12182c),
	.w5(32'hba448fb8),
	.w6(32'h397d475b),
	.w7(32'hba54eae2),
	.w8(32'hba87bc28),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad68800),
	.w1(32'hbb65c28f),
	.w2(32'hbaf33b06),
	.w3(32'hbb00c504),
	.w4(32'hbb8e3ebc),
	.w5(32'hbabd7ff5),
	.w6(32'hbb183e24),
	.w7(32'hbbab5d3d),
	.w8(32'hbb445134),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e80d4),
	.w1(32'h399e1733),
	.w2(32'hbb4baa3f),
	.w3(32'hbabe6010),
	.w4(32'h3b007204),
	.w5(32'hb9dd80cb),
	.w6(32'hbb35fd9d),
	.w7(32'hb9a39fbf),
	.w8(32'hbad7f2b7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab423ad),
	.w1(32'h3aada0e6),
	.w2(32'h3abe9486),
	.w3(32'hbb0a6e47),
	.w4(32'h3b3f4a1e),
	.w5(32'hbb1806e5),
	.w6(32'hba81f45a),
	.w7(32'h3abaac5c),
	.w8(32'hbb0a6ed0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16fda5),
	.w1(32'hbae9c2f7),
	.w2(32'hbb2c3732),
	.w3(32'h3ad1a22d),
	.w4(32'hbad656d1),
	.w5(32'hbb2389f1),
	.w6(32'h3a583153),
	.w7(32'hbaae3661),
	.w8(32'hbb0a414d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e3756),
	.w1(32'hbb27b708),
	.w2(32'hba077495),
	.w3(32'hbad12f87),
	.w4(32'hbb038b75),
	.w5(32'h3846108f),
	.w6(32'hbad1b36b),
	.w7(32'h3a2d5a94),
	.w8(32'hba9330fd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f8ca),
	.w1(32'hbaab19d1),
	.w2(32'hbb8ee096),
	.w3(32'hbaebd8ea),
	.w4(32'hbb2c9c88),
	.w5(32'hbb6ecb2f),
	.w6(32'hbaf00034),
	.w7(32'hbb5dffc5),
	.w8(32'hbb92e61f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4488a8),
	.w1(32'hbab25fdc),
	.w2(32'hbaee6ed7),
	.w3(32'hbb3f2375),
	.w4(32'hbb12a92e),
	.w5(32'hbb163fe6),
	.w6(32'hbb3d94f1),
	.w7(32'h39d1c100),
	.w8(32'hb7f10477),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39324229),
	.w1(32'hbade0c58),
	.w2(32'hbaa64f03),
	.w3(32'h3ae56ea2),
	.w4(32'h3b1f0ed0),
	.w5(32'h3933be84),
	.w6(32'h3ae273ee),
	.w7(32'h3b19603b),
	.w8(32'hba37baa0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8352cb),
	.w1(32'hba8ef5d0),
	.w2(32'h3afcbf66),
	.w3(32'h3b215a55),
	.w4(32'h3b751a94),
	.w5(32'h3ac59441),
	.w6(32'h3b4f98ba),
	.w7(32'h3ae4e981),
	.w8(32'hba82726c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab073c4),
	.w1(32'hba8f98d7),
	.w2(32'hba9bf990),
	.w3(32'hbb1e8c8c),
	.w4(32'hbad8b40c),
	.w5(32'hbaf9ab73),
	.w6(32'h39b5ee4e),
	.w7(32'hbaac141a),
	.w8(32'hba80b156),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb499296),
	.w1(32'hb974d552),
	.w2(32'hbb0bb96e),
	.w3(32'hbbc2fcaa),
	.w4(32'h3ad8ea74),
	.w5(32'hb8c35508),
	.w6(32'hbb202de3),
	.w7(32'h3b3e9174),
	.w8(32'h3a39f2df),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84849a),
	.w1(32'h3a800010),
	.w2(32'h3a355736),
	.w3(32'h3a476b29),
	.w4(32'h3b8b603e),
	.w5(32'h3ae217ac),
	.w6(32'hba78e56f),
	.w7(32'h3b2a35d9),
	.w8(32'h3a96de88),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bc30d),
	.w1(32'hb5f42f6b),
	.w2(32'h3a2a3f2b),
	.w3(32'h3944db1c),
	.w4(32'h3ab04bf7),
	.w5(32'hba902d94),
	.w6(32'hb9d2680e),
	.w7(32'hba2441dc),
	.w8(32'hbabd0e18),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a906c41),
	.w1(32'hbb1b5a57),
	.w2(32'hbb5035a9),
	.w3(32'hbb10be17),
	.w4(32'hbb1e178f),
	.w5(32'h390c29b0),
	.w6(32'hba2cb016),
	.w7(32'hbb1eb185),
	.w8(32'hba3051d7),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf62220),
	.w1(32'hba888cb2),
	.w2(32'hbadefaff),
	.w3(32'hbb049ee4),
	.w4(32'hbaa1b153),
	.w5(32'h3961a028),
	.w6(32'hbb2bc560),
	.w7(32'hb9a5eb62),
	.w8(32'h396eb6dd),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9538a6d),
	.w1(32'h3864c6d6),
	.w2(32'hba0fda80),
	.w3(32'h38969bde),
	.w4(32'hba14dccd),
	.w5(32'h3a8f5cf0),
	.w6(32'hb91a6974),
	.w7(32'hbae23427),
	.w8(32'hba64042e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df313b),
	.w1(32'h3aa2a1f4),
	.w2(32'h3b7ae359),
	.w3(32'hb938dd20),
	.w4(32'h3aab409a),
	.w5(32'h39e62919),
	.w6(32'hbb38c690),
	.w7(32'h3ad33c7d),
	.w8(32'hba6c70c6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20efac),
	.w1(32'h38310346),
	.w2(32'hbb5889ab),
	.w3(32'h3933aecf),
	.w4(32'h3b27bb89),
	.w5(32'hb6d86080),
	.w6(32'hbb38e559),
	.w7(32'h3b415f77),
	.w8(32'hba5c91c4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb736c0f),
	.w1(32'hb782d2cd),
	.w2(32'hbabfbce3),
	.w3(32'hbb3c6ec3),
	.w4(32'hbae678fd),
	.w5(32'h3a55c232),
	.w6(32'hbab56ced),
	.w7(32'hbaae9101),
	.w8(32'hbb3c55ca),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004bf2),
	.w1(32'h39ab1f0b),
	.w2(32'h380990f2),
	.w3(32'hbab962bc),
	.w4(32'h3b269ef9),
	.w5(32'h3a83c85a),
	.w6(32'hbb377876),
	.w7(32'hb96beb24),
	.w8(32'hba9fcec8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0735ef),
	.w1(32'hbb6b42bc),
	.w2(32'h39846c24),
	.w3(32'hbac2d1bb),
	.w4(32'hba5a03c4),
	.w5(32'h3b62f913),
	.w6(32'hbb73719b),
	.w7(32'h3a95c730),
	.w8(32'h3bb0c003),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c2b4a),
	.w1(32'hbb42abd7),
	.w2(32'h39515900),
	.w3(32'h3b6e52de),
	.w4(32'hbae07602),
	.w5(32'h3b2efda6),
	.w6(32'h3b31eb21),
	.w7(32'hba53d4ff),
	.w8(32'hb8ed8dd2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad726bb),
	.w1(32'hbb46de57),
	.w2(32'hbb6d8fbb),
	.w3(32'h3776e2f9),
	.w4(32'hb9b3ce3b),
	.w5(32'hbb2e9a8f),
	.w6(32'h3b643b1a),
	.w7(32'h3af1d82b),
	.w8(32'hb9f7cd0d),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6af1d),
	.w1(32'hba0869bc),
	.w2(32'hba33eba9),
	.w3(32'h3af5bd23),
	.w4(32'hb9b9feb1),
	.w5(32'hbaabcf13),
	.w6(32'h3b86a82d),
	.w7(32'hba2327ed),
	.w8(32'hbb4046c0),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaef286),
	.w1(32'hbb9aee8d),
	.w2(32'hbbbcea2a),
	.w3(32'hba2a9dd8),
	.w4(32'hbb69e432),
	.w5(32'hbac1f5f5),
	.w6(32'hb8a511e5),
	.w7(32'hba06eee2),
	.w8(32'h3b1c1c24),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39958214),
	.w1(32'h3872ecf1),
	.w2(32'hbb01a73e),
	.w3(32'h3b6df65d),
	.w4(32'hbb2a941b),
	.w5(32'hb9a91385),
	.w6(32'h3bd3c93b),
	.w7(32'hbb69184b),
	.w8(32'hba482307),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae958d0),
	.w1(32'hbb3689e8),
	.w2(32'hbad0e8a1),
	.w3(32'h3a85503a),
	.w4(32'hbb1f55a6),
	.w5(32'hba9f1a67),
	.w6(32'h3a1f7cd3),
	.w7(32'hbb3c4e17),
	.w8(32'hbb815b72),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a26f7),
	.w1(32'hbb1066d8),
	.w2(32'hbb9492e7),
	.w3(32'hbb37570f),
	.w4(32'hbb18f7a8),
	.w5(32'hba06c6e7),
	.w6(32'hbb2e6ff3),
	.w7(32'hbb96009a),
	.w8(32'hbb507a90),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfff59a),
	.w1(32'hba3bbda4),
	.w2(32'hb9a2d1af),
	.w3(32'hbae61785),
	.w4(32'h3a54ee1e),
	.w5(32'hba3383a8),
	.w6(32'hbb63b8c5),
	.w7(32'h3adc27fc),
	.w8(32'hba223ec3),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab09094),
	.w1(32'hbb014d7b),
	.w2(32'hbbc76f03),
	.w3(32'hb92e00ca),
	.w4(32'hbb408659),
	.w5(32'hba78323a),
	.w6(32'hbb4df11f),
	.w7(32'hba2b8656),
	.w8(32'hba912040),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fde0d),
	.w1(32'h3b25da24),
	.w2(32'hbaf9e278),
	.w3(32'h3996375d),
	.w4(32'h3b165203),
	.w5(32'hb9c3cb7a),
	.w6(32'hbb91f1d3),
	.w7(32'h3a8d0fbe),
	.w8(32'hba95aa37),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f8f41),
	.w1(32'hba2fa563),
	.w2(32'hbb4f9408),
	.w3(32'hbb3bb67a),
	.w4(32'hba068cc0),
	.w5(32'hbace0111),
	.w6(32'hbafa6b0a),
	.w7(32'h3b1d3d5c),
	.w8(32'hbb164802),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5bcd),
	.w1(32'hba95531a),
	.w2(32'hbb0d587a),
	.w3(32'h3a313814),
	.w4(32'hbafdbe0f),
	.w5(32'h3a847db5),
	.w6(32'h3ab728a1),
	.w7(32'hba9bf934),
	.w8(32'hbb900e1d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f84bf4),
	.w1(32'h3a6f3b71),
	.w2(32'h3a8caa64),
	.w3(32'hbad88ff3),
	.w4(32'h3b2168b3),
	.w5(32'hbafb66fa),
	.w6(32'hb990b1fb),
	.w7(32'hba2095aa),
	.w8(32'hba9738dd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31ebe5),
	.w1(32'hb9f9f687),
	.w2(32'h3a869677),
	.w3(32'hbabaef61),
	.w4(32'h3b090857),
	.w5(32'hba7b9e72),
	.w6(32'hba2751a7),
	.w7(32'h3a9fabe7),
	.w8(32'hbaae6dfd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa8264),
	.w1(32'h3afffaf8),
	.w2(32'h3b4be210),
	.w3(32'h3ae77216),
	.w4(32'h3b095683),
	.w5(32'h3b365caa),
	.w6(32'hbabb760d),
	.w7(32'h3a2073a0),
	.w8(32'hb997e626),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43e39c),
	.w1(32'h3b0b3cc3),
	.w2(32'hbae2635a),
	.w3(32'h3b360536),
	.w4(32'h3a3359a7),
	.w5(32'hbb3c9aa4),
	.w6(32'h3a96140a),
	.w7(32'h3b1f0799),
	.w8(32'hbb2f2695),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e4141),
	.w1(32'hb9f80fb2),
	.w2(32'h3b72c8c5),
	.w3(32'hbb5ddb79),
	.w4(32'hbb27238f),
	.w5(32'h3a535b7d),
	.w6(32'hbb4f1b85),
	.w7(32'hbb3d970a),
	.w8(32'h38e4f332),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977f48e),
	.w1(32'hbb4488ef),
	.w2(32'hbb6cc75f),
	.w3(32'hbaed5765),
	.w4(32'hbac3aaaa),
	.w5(32'hbaae12eb),
	.w6(32'hbaabc0ed),
	.w7(32'hbb084e77),
	.w8(32'hbb37b19a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee0270),
	.w1(32'hb93218e9),
	.w2(32'h3b89e454),
	.w3(32'hbb168446),
	.w4(32'h3a43e48a),
	.w5(32'h3b2a7635),
	.w6(32'hba1540de),
	.w7(32'h3b84c4d7),
	.w8(32'h3b07f693),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a78fa),
	.w1(32'h3af271ac),
	.w2(32'h3b041d51),
	.w3(32'h3b083afe),
	.w4(32'h3992e0a3),
	.w5(32'h38148e4f),
	.w6(32'h3b68a7fc),
	.w7(32'hb9feae12),
	.w8(32'hba36d2f1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7c50),
	.w1(32'h3909d858),
	.w2(32'hbb046367),
	.w3(32'hba1f316b),
	.w4(32'h3b107017),
	.w5(32'hbb405ad2),
	.w6(32'hbaa16d1d),
	.w7(32'h3883d1b2),
	.w8(32'hbb19fcf0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abdba0a),
	.w1(32'h3b4b8cab),
	.w2(32'h3af6de0b),
	.w3(32'h3b214d71),
	.w4(32'h3b31558b),
	.w5(32'h3b3f7a15),
	.w6(32'h3ab287aa),
	.w7(32'h3b8ac70f),
	.w8(32'h3b09676d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0eb78),
	.w1(32'hbb5ad792),
	.w2(32'hbb4b8526),
	.w3(32'h39f271f1),
	.w4(32'hbb1048f5),
	.w5(32'hbac01f07),
	.w6(32'h3a7d5781),
	.w7(32'hba632d66),
	.w8(32'hbabc1518),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75a9f0),
	.w1(32'hbb05629c),
	.w2(32'hbad31ce0),
	.w3(32'hbb12f550),
	.w4(32'hbb08b753),
	.w5(32'hba87045c),
	.w6(32'h399f8b08),
	.w7(32'hba2b71f6),
	.w8(32'hb8f0d70f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae60ca4),
	.w1(32'hb999f912),
	.w2(32'hba9c2510),
	.w3(32'hba6e3244),
	.w4(32'hbb0a23dc),
	.w5(32'h38f3ef8f),
	.w6(32'hb9b1f279),
	.w7(32'hbb558bb9),
	.w8(32'hba304dca),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b890b),
	.w1(32'h3aea7800),
	.w2(32'h3b78536b),
	.w3(32'hbb9beda0),
	.w4(32'h39ee9373),
	.w5(32'h3b3ae668),
	.w6(32'hbab2f181),
	.w7(32'h3a644f07),
	.w8(32'h3aaa7d08),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d95fad),
	.w1(32'hba1d2dcf),
	.w2(32'hba36f7c8),
	.w3(32'h3a392bb4),
	.w4(32'h3a82b9a5),
	.w5(32'h3a8d6298),
	.w6(32'h3b424a64),
	.w7(32'hbb15abb9),
	.w8(32'h3990a1e5),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23dc02),
	.w1(32'h3b924ccd),
	.w2(32'h3b84eace),
	.w3(32'h3af0ab42),
	.w4(32'h3b7a15f5),
	.w5(32'h3b9f715f),
	.w6(32'hb9cf67b7),
	.w7(32'hbab227c3),
	.w8(32'h3af31b43),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e288),
	.w1(32'hbb015d07),
	.w2(32'hbb1ca474),
	.w3(32'h3b42d2e1),
	.w4(32'hbb141e9e),
	.w5(32'h3ac88ea1),
	.w6(32'hbb4b977f),
	.w7(32'h38231dec),
	.w8(32'h3b399f5f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb2e31),
	.w1(32'h39578c22),
	.w2(32'h3b8826b4),
	.w3(32'hbaa186da),
	.w4(32'hb9e7ce9c),
	.w5(32'h3af22d3e),
	.w6(32'hb94ea1d0),
	.w7(32'hbafbe877),
	.w8(32'hba6e0731),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38dbe4),
	.w1(32'h3ad4e2b9),
	.w2(32'h3adb03c4),
	.w3(32'hba431b1b),
	.w4(32'h3adc54d7),
	.w5(32'h3a4851c7),
	.w6(32'h3ae30980),
	.w7(32'h3a5e086a),
	.w8(32'hba807430),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85cd36),
	.w1(32'h3b38c100),
	.w2(32'h3a77c6e9),
	.w3(32'h3bae433b),
	.w4(32'h3b71f961),
	.w5(32'hba4c0d07),
	.w6(32'h3b203426),
	.w7(32'hb9494b60),
	.w8(32'hbb8c937e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5be8b),
	.w1(32'hbad1e90d),
	.w2(32'hbb95a8a5),
	.w3(32'h3b85bb4b),
	.w4(32'h3a22627b),
	.w5(32'hbb019d2a),
	.w6(32'h3b1ed4be),
	.w7(32'h39e355d0),
	.w8(32'hbb3b955c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f7b3),
	.w1(32'h39ead513),
	.w2(32'hbb2560db),
	.w3(32'hbb16b6d1),
	.w4(32'h3b2b1ca6),
	.w5(32'hbb3a5316),
	.w6(32'hbb2c0f77),
	.w7(32'h3ab6ddf6),
	.w8(32'hbb6b9cad),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f60da0),
	.w1(32'hbafa84b3),
	.w2(32'hbb3ad8da),
	.w3(32'h3a324abd),
	.w4(32'hba721e3f),
	.w5(32'hbac63ba7),
	.w6(32'hba9d69ae),
	.w7(32'h3aacf408),
	.w8(32'hba7e1246),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d5997),
	.w1(32'hbb7d0c08),
	.w2(32'hbb2c6a94),
	.w3(32'hbb4cb6ac),
	.w4(32'hbb5dc4ae),
	.w5(32'hba5965e7),
	.w6(32'hbb1269fe),
	.w7(32'hbacea3e9),
	.w8(32'h3b2e482d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af176),
	.w1(32'hbb08fb4e),
	.w2(32'hbb11f9e2),
	.w3(32'h39a517b3),
	.w4(32'hbaa36e93),
	.w5(32'hba80efd2),
	.w6(32'h3a3beb96),
	.w7(32'h37330b04),
	.w8(32'h3a5b8e80),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb278ac2),
	.w1(32'hbb524533),
	.w2(32'hbb79271b),
	.w3(32'h3acadb66),
	.w4(32'hbb177d0d),
	.w5(32'hbb423ed2),
	.w6(32'h3b485f6f),
	.w7(32'hbb919f56),
	.w8(32'h3909957e),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac88c93),
	.w1(32'hbb622734),
	.w2(32'hbb631e73),
	.w3(32'hbb80f6d3),
	.w4(32'hbb5270ba),
	.w5(32'hba8a4534),
	.w6(32'hbaf0dd30),
	.w7(32'hbb7e1a43),
	.w8(32'hbb3f913f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fd289),
	.w1(32'h3a6c51cc),
	.w2(32'hba9f333f),
	.w3(32'hbb1f3a21),
	.w4(32'hba1f8112),
	.w5(32'h3a8e7f6d),
	.w6(32'hbb6b0218),
	.w7(32'hbab3ab2a),
	.w8(32'hbae5d39f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba918ad2),
	.w1(32'h3b2f4f5d),
	.w2(32'h3a8c2e2b),
	.w3(32'hbb2c9028),
	.w4(32'h3b03ce41),
	.w5(32'hbb13bb0a),
	.w6(32'hbb456ad7),
	.w7(32'hba788884),
	.w8(32'hbac029c1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb411533),
	.w1(32'hba9f79a1),
	.w2(32'hbb6d2df6),
	.w3(32'hba5def65),
	.w4(32'h3b00112d),
	.w5(32'hbad2812b),
	.w6(32'hb9811227),
	.w7(32'h3b811814),
	.w8(32'hb9a4f842),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93f760),
	.w1(32'h3b077e32),
	.w2(32'h3a2155fe),
	.w3(32'hbb3755c8),
	.w4(32'h3b118ee0),
	.w5(32'h3a8cd87a),
	.w6(32'hb9ecb1c5),
	.w7(32'h3b4fdbf5),
	.w8(32'h3a5d504f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8f60),
	.w1(32'hb9413384),
	.w2(32'h3b32db1a),
	.w3(32'h3a91b8a3),
	.w4(32'h3a5d7039),
	.w5(32'h3a352148),
	.w6(32'h3a39a9c7),
	.w7(32'hb9c66208),
	.w8(32'hb9759868),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b2bf8),
	.w1(32'hbb106adc),
	.w2(32'hbb1f7bb9),
	.w3(32'h3b3e75ac),
	.w4(32'hba7acc31),
	.w5(32'hb9b09bdd),
	.w6(32'h3ab06a1f),
	.w7(32'hbaf690b1),
	.w8(32'hbafa21fa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63793a),
	.w1(32'h3ab47c42),
	.w2(32'hba583faa),
	.w3(32'hbacbe4a9),
	.w4(32'hbadd520f),
	.w5(32'h3ab28989),
	.w6(32'hba6fbb39),
	.w7(32'hbb100a8b),
	.w8(32'hbb80a9ae),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a6bf8),
	.w1(32'h3b773310),
	.w2(32'h3a65448a),
	.w3(32'hbb0c6de9),
	.w4(32'h3aebc14e),
	.w5(32'h3ad89f68),
	.w6(32'hbb64302e),
	.w7(32'h3a2aeb89),
	.w8(32'h3ae97cfd),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4b1a2),
	.w1(32'hbac5b8ee),
	.w2(32'hbb14af9b),
	.w3(32'h3b154ec9),
	.w4(32'hb994b08e),
	.w5(32'hba11350e),
	.w6(32'h3ba36740),
	.w7(32'hbb3ffbd1),
	.w8(32'hbb5d2945),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f4aaf),
	.w1(32'hbafc944d),
	.w2(32'hbaffa54b),
	.w3(32'hbad5f00d),
	.w4(32'hbaf9ad60),
	.w5(32'hba73e2cf),
	.w6(32'hba6e993a),
	.w7(32'hbb232c5e),
	.w8(32'hbb09b504),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0647a4),
	.w1(32'hb964fc5d),
	.w2(32'hbac7ab6e),
	.w3(32'hbaf3b2ea),
	.w4(32'hbb0bd4a5),
	.w5(32'hb9f39b39),
	.w6(32'hbaa2d24c),
	.w7(32'hba8f0a8c),
	.w8(32'hba8c8dd7),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1763ab),
	.w1(32'hb9c2cdda),
	.w2(32'hb9b34827),
	.w3(32'h3929aae5),
	.w4(32'hba023c34),
	.w5(32'hbb0a9541),
	.w6(32'hb91278ff),
	.w7(32'hbb29051f),
	.w8(32'hbb35a637),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94966b0),
	.w1(32'hb8e78b14),
	.w2(32'h3a4d9889),
	.w3(32'hbb31a701),
	.w4(32'h3962ffe1),
	.w5(32'hba7ed79f),
	.w6(32'hbb0fbe9b),
	.w7(32'hba9fe49b),
	.w8(32'hbaaaeb98),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d27a5),
	.w1(32'hba23644d),
	.w2(32'h3af24b74),
	.w3(32'hbad643f1),
	.w4(32'hb9d07ec4),
	.w5(32'h3993eb2d),
	.w6(32'hba8d27e5),
	.w7(32'h39ccb0da),
	.w8(32'hb9c1b326),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84ca91),
	.w1(32'hb8bc3754),
	.w2(32'h39695e89),
	.w3(32'h39c2974d),
	.w4(32'h3ace86ca),
	.w5(32'h3ae00500),
	.w6(32'hbb342576),
	.w7(32'h39d022d7),
	.w8(32'h3a27b91b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38013118),
	.w1(32'h398947b8),
	.w2(32'hbb243b3e),
	.w3(32'h3a8ef901),
	.w4(32'hbaa87fdf),
	.w5(32'hbb9fb691),
	.w6(32'hb99acbb6),
	.w7(32'hbaa47e85),
	.w8(32'hbb32de06),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29af66),
	.w1(32'hbb70e6ab),
	.w2(32'hbb58fd40),
	.w3(32'hbb85d985),
	.w4(32'hbb12dd1a),
	.w5(32'hb92cafca),
	.w6(32'hbb7cc7ab),
	.w7(32'hbb0f1edf),
	.w8(32'hbb457bb4),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba853405),
	.w1(32'h3a185f33),
	.w2(32'h3aa7d3bc),
	.w3(32'hbb3c5ebd),
	.w4(32'hb8a256e7),
	.w5(32'h3a3c5b1f),
	.w6(32'hbada5b5b),
	.w7(32'h396a7825),
	.w8(32'h39292bb9),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f887a),
	.w1(32'hbaaef061),
	.w2(32'hba86f333),
	.w3(32'h3a6e3b81),
	.w4(32'hba8c9f05),
	.w5(32'hbadc01a4),
	.w6(32'h3934a5d2),
	.w7(32'h39f623ca),
	.w8(32'hbb270a05),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59cba7),
	.w1(32'h3b9cff5b),
	.w2(32'h3b8bb6e3),
	.w3(32'hbad168b0),
	.w4(32'h3b8a5405),
	.w5(32'h3ade491e),
	.w6(32'hbaa5e5e6),
	.w7(32'h3b82e1c2),
	.w8(32'h3b831dfa),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb3986),
	.w1(32'h394ccb46),
	.w2(32'hb904d653),
	.w3(32'h3ad1c52a),
	.w4(32'h398c3eea),
	.w5(32'hba5de804),
	.w6(32'h3b3af06d),
	.w7(32'hb8074581),
	.w8(32'hb9a471d6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab61c44),
	.w1(32'hbaa02db8),
	.w2(32'hba80e1b1),
	.w3(32'hb9a34cb4),
	.w4(32'hbab271c4),
	.w5(32'hba30e221),
	.w6(32'h3a8a946c),
	.w7(32'hbae49b43),
	.w8(32'hb9a8f96a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba275f3d),
	.w1(32'hba94ef15),
	.w2(32'hbac7a663),
	.w3(32'hb78bf1ea),
	.w4(32'hb99d596c),
	.w5(32'hbb19d437),
	.w6(32'h38d034ae),
	.w7(32'hbaed050a),
	.w8(32'hbb9af27c),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fa6b),
	.w1(32'hba94e930),
	.w2(32'hb9fd0876),
	.w3(32'hbb6ed587),
	.w4(32'hbb09cc36),
	.w5(32'h39ea6bc8),
	.w6(32'h39a2c058),
	.w7(32'hbaf8a863),
	.w8(32'hba384a93),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934b253),
	.w1(32'hb9dd49e4),
	.w2(32'hbbc3a3bb),
	.w3(32'hbac43946),
	.w4(32'hb94642bc),
	.w5(32'hbb97a94d),
	.w6(32'hba43f38f),
	.w7(32'hbba02a98),
	.w8(32'hbbca2432),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb560a8a),
	.w1(32'hbad2f3a1),
	.w2(32'h3afb947d),
	.w3(32'hbb884d12),
	.w4(32'hb9b47d6e),
	.w5(32'h3b472703),
	.w6(32'hbb2fe2bd),
	.w7(32'h3a8ead67),
	.w8(32'h3b412669),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2917b3),
	.w1(32'hbac0b28d),
	.w2(32'hbac30c1c),
	.w3(32'h3a62e999),
	.w4(32'hbae1dc30),
	.w5(32'hba91012c),
	.w6(32'h395eb660),
	.w7(32'hba15883d),
	.w8(32'hbafa213d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63d35b),
	.w1(32'hb9c7504c),
	.w2(32'hb97e153e),
	.w3(32'hba47114f),
	.w4(32'hbacd1401),
	.w5(32'hb95a0855),
	.w6(32'hbac4d30d),
	.w7(32'hba529e9f),
	.w8(32'hbb432a7a),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9a924),
	.w1(32'hbab30ccb),
	.w2(32'hb85a71dc),
	.w3(32'hbb348f76),
	.w4(32'hba0bc491),
	.w5(32'h3989019e),
	.w6(32'hbba4f9c1),
	.w7(32'h3a027dad),
	.w8(32'h378982ff),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a612d08),
	.w1(32'hbac27e4d),
	.w2(32'hba628351),
	.w3(32'h3a4929c2),
	.w4(32'hba9c3b53),
	.w5(32'h3a9e2d04),
	.w6(32'h38a22d6a),
	.w7(32'hbaaf315f),
	.w8(32'h3925961d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a255),
	.w1(32'hba7a4467),
	.w2(32'h387dc87e),
	.w3(32'hbb251d6d),
	.w4(32'hb91f81bf),
	.w5(32'h3ae05cbb),
	.w6(32'hbb0cfcb4),
	.w7(32'hbaed83bf),
	.w8(32'hbac1f0fe),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9661209),
	.w1(32'h3ab85671),
	.w2(32'h3a843ce9),
	.w3(32'hbaa2ac75),
	.w4(32'h3a994d1c),
	.w5(32'h3a8b8ae7),
	.w6(32'hba826df1),
	.w7(32'hba15092c),
	.w8(32'hba32e96a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4768be),
	.w1(32'h3b08fdeb),
	.w2(32'h3a5f08de),
	.w3(32'h3a97fdaa),
	.w4(32'h3acd5412),
	.w5(32'h3951597d),
	.w6(32'hba144a11),
	.w7(32'hba6b478c),
	.w8(32'hba65215f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab56f03),
	.w1(32'h3ac0137c),
	.w2(32'h3a400245),
	.w3(32'hbaba8ef9),
	.w4(32'hb9fc15a1),
	.w5(32'h3b009606),
	.w6(32'hba991b28),
	.w7(32'hb90f0520),
	.w8(32'hbac0465a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a061aea),
	.w1(32'hba8e15b3),
	.w2(32'hba85660a),
	.w3(32'h3a6d789b),
	.w4(32'hbb127707),
	.w5(32'hbb625b2e),
	.w6(32'h394e6814),
	.w7(32'hbac479e0),
	.w8(32'hbae7787b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6b491),
	.w1(32'hbb0a2d7b),
	.w2(32'hbb4f49e6),
	.w3(32'hbb252935),
	.w4(32'hbb924feb),
	.w5(32'hbb2cd1e8),
	.w6(32'hba90ae08),
	.w7(32'hbb7b683c),
	.w8(32'hbb852f68),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade0a9d),
	.w1(32'h3a49b504),
	.w2(32'hbad53d70),
	.w3(32'hbb104079),
	.w4(32'h38b40536),
	.w5(32'hbb16175b),
	.w6(32'hbab2ae01),
	.w7(32'h3abcc563),
	.w8(32'hbb1253d2),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa37665),
	.w1(32'hbab53fe4),
	.w2(32'hb92dace3),
	.w3(32'hbb12f786),
	.w4(32'hbafb8b76),
	.w5(32'h390c4785),
	.w6(32'hbb3966ac),
	.w7(32'hbb342d94),
	.w8(32'hbaa49e57),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba232d16),
	.w1(32'h3950f519),
	.w2(32'h39fc77a9),
	.w3(32'hbb2d5898),
	.w4(32'hba7fe596),
	.w5(32'h3b289d15),
	.w6(32'hbb18f6fc),
	.w7(32'hbab7e2d6),
	.w8(32'hbaba7a56),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397dd5c1),
	.w1(32'hba2045b1),
	.w2(32'h37c42234),
	.w3(32'h3a50ef8f),
	.w4(32'hba413166),
	.w5(32'h3a2596ad),
	.w6(32'hbb1e503c),
	.w7(32'h38ed3cfc),
	.w8(32'h3a00db3d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d32cb),
	.w1(32'hb914f777),
	.w2(32'hba08ff90),
	.w3(32'hb98aef95),
	.w4(32'hba963cd8),
	.w5(32'hba04b07d),
	.w6(32'h3948b71a),
	.w7(32'hbaf452ca),
	.w8(32'hba65eb53),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e33bcd),
	.w1(32'h3726b974),
	.w2(32'hbaf3858e),
	.w3(32'h39594db4),
	.w4(32'hbafa23be),
	.w5(32'hbb3d7cc4),
	.w6(32'h37b656c3),
	.w7(32'h39e228be),
	.w8(32'hbab998fb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26884d),
	.w1(32'hbaa5407b),
	.w2(32'hba2464b1),
	.w3(32'hbb2650e1),
	.w4(32'hba7abaca),
	.w5(32'hb9c2c7c8),
	.w6(32'hbaf9a0e5),
	.w7(32'hba606936),
	.w8(32'h3ab71688),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77b598),
	.w1(32'h3a171db3),
	.w2(32'h3a4e0eb7),
	.w3(32'hbadc7d4c),
	.w4(32'h3a0e3838),
	.w5(32'h386fb8b2),
	.w6(32'h378ad7f7),
	.w7(32'hbaa359a2),
	.w8(32'hba9b6438),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a8c654),
	.w1(32'h3a8663d4),
	.w2(32'hb9269eb3),
	.w3(32'h3a35f2a1),
	.w4(32'h380d4732),
	.w5(32'hb9d59fa2),
	.w6(32'h389f216d),
	.w7(32'hba5cccb6),
	.w8(32'hbac9062d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d207),
	.w1(32'h39a53394),
	.w2(32'h39f76a58),
	.w3(32'hba90f076),
	.w4(32'h38bcd378),
	.w5(32'hbabecd6c),
	.w6(32'hbaad0c0f),
	.w7(32'h39c18210),
	.w8(32'h3aac66f7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08fe0d),
	.w1(32'hb9e96583),
	.w2(32'hb9ac15b4),
	.w3(32'h3ac83607),
	.w4(32'hba91f209),
	.w5(32'h39cec6ec),
	.w6(32'h3b56282f),
	.w7(32'hbafdd90b),
	.w8(32'hbaa0d3ca),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95bd94),
	.w1(32'h39cab30f),
	.w2(32'h3a2082df),
	.w3(32'hba49776c),
	.w4(32'h3a25d181),
	.w5(32'h3afb9096),
	.w6(32'hbb2c629a),
	.w7(32'h3a7c33ab),
	.w8(32'h3ab9c38a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a3cfe),
	.w1(32'hba429a4c),
	.w2(32'hbb5fabab),
	.w3(32'h3b5f95b8),
	.w4(32'h39b1376f),
	.w5(32'h3a861a56),
	.w6(32'h3a99f47a),
	.w7(32'h379c4b08),
	.w8(32'hbaa71330),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a0fca),
	.w1(32'hbb894334),
	.w2(32'hbb0b5711),
	.w3(32'hbabe2e3d),
	.w4(32'hbb7cdd64),
	.w5(32'hbaeb8690),
	.w6(32'hbb32e72d),
	.w7(32'hbb490b08),
	.w8(32'hbb12e463),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f80e4d),
	.w1(32'hbac346c9),
	.w2(32'hbaf6e96d),
	.w3(32'hbb06a2b3),
	.w4(32'hbaaefcca),
	.w5(32'hba9fdec4),
	.w6(32'hbb2a5178),
	.w7(32'hbb155507),
	.w8(32'hbb4ea7ec),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440565),
	.w1(32'h39c3c22c),
	.w2(32'hba355a90),
	.w3(32'hbb210e0e),
	.w4(32'hb9feb048),
	.w5(32'hbb5d2476),
	.w6(32'hbad559d4),
	.w7(32'h394cf3ae),
	.w8(32'hbadf8202),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae893e9),
	.w1(32'h3931e661),
	.w2(32'hb87d158e),
	.w3(32'hbad7b8dd),
	.w4(32'hbad876a9),
	.w5(32'hb958a0a4),
	.w6(32'hba82e8d2),
	.w7(32'hbae5d134),
	.w8(32'hbb0f558b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f5ea6),
	.w1(32'h379914ed),
	.w2(32'h3ad844c3),
	.w3(32'hb7bde9af),
	.w4(32'h39b27d5d),
	.w5(32'h3b086036),
	.w6(32'hb9677a6e),
	.w7(32'h387a31ff),
	.w8(32'h37c8e1f2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb798029e),
	.w1(32'hba888c4c),
	.w2(32'h3a26cecc),
	.w3(32'h3a84c089),
	.w4(32'hbb1d4dee),
	.w5(32'h3a12dffe),
	.w6(32'hb9ee5e24),
	.w7(32'hbb54801a),
	.w8(32'hba179436),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55e534),
	.w1(32'hb90af8e6),
	.w2(32'hba8d96ae),
	.w3(32'hba925cdd),
	.w4(32'h38cabfb2),
	.w5(32'h3acb0993),
	.w6(32'hbaea56d7),
	.w7(32'h394a536f),
	.w8(32'h3a6fa687),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ae72a),
	.w1(32'hb9e21813),
	.w2(32'hba8c2e49),
	.w3(32'h3a979144),
	.w4(32'hb9b13552),
	.w5(32'hbacab2c1),
	.w6(32'hba47ab10),
	.w7(32'hb9a48174),
	.w8(32'hba21fde1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba035df3),
	.w1(32'hbacb99ab),
	.w2(32'hba310a64),
	.w3(32'hba93511b),
	.w4(32'hbab0af4e),
	.w5(32'hb870242e),
	.w6(32'h3a15f951),
	.w7(32'h3a2ad4db),
	.w8(32'h398b4cc9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c8127),
	.w1(32'hba9a9a91),
	.w2(32'hbac60d5e),
	.w3(32'hbab029d1),
	.w4(32'hbb188247),
	.w5(32'hbb05147a),
	.w6(32'hba237142),
	.w7(32'hba5b6ab7),
	.w8(32'hba05ecff),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a951196),
	.w1(32'hb96e4902),
	.w2(32'hbab0e94f),
	.w3(32'h39f2ccb9),
	.w4(32'hba720dae),
	.w5(32'hba981000),
	.w6(32'hb7d5ad8a),
	.w7(32'hba9bf66e),
	.w8(32'hba8d9b0b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025283),
	.w1(32'hbaac5b27),
	.w2(32'hba8cc961),
	.w3(32'hbb1877ba),
	.w4(32'hba06f3f7),
	.w5(32'h3abd88a6),
	.w6(32'hbb3cc209),
	.w7(32'hbabdaa87),
	.w8(32'h3a16468b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf60ce5),
	.w1(32'hb9a031e2),
	.w2(32'hba519726),
	.w3(32'h3a4cd948),
	.w4(32'hbb3c4724),
	.w5(32'hbae4f90c),
	.w6(32'hbaf96c80),
	.w7(32'hbb17c146),
	.w8(32'hbb03176a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7c87f),
	.w1(32'h3b38f28d),
	.w2(32'h3a98061e),
	.w3(32'hbab9842c),
	.w4(32'h39612d4c),
	.w5(32'hb95b87ba),
	.w6(32'hba3e5002),
	.w7(32'hb6c1cbd6),
	.w8(32'hba812cb2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f7292),
	.w1(32'hb9a41caa),
	.w2(32'h36696e77),
	.w3(32'h3ae6e470),
	.w4(32'hba348e7e),
	.w5(32'h3b3a8e49),
	.w6(32'h3a89ebf9),
	.w7(32'h3a7f387b),
	.w8(32'h3aa6e7cb),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a665bf7),
	.w1(32'hbae29ec9),
	.w2(32'hbadb8ab7),
	.w3(32'h3afc0618),
	.w4(32'hbb27f65c),
	.w5(32'hbb1116cd),
	.w6(32'h3b1e6555),
	.w7(32'hbb310ae5),
	.w8(32'hbb167944),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f1375),
	.w1(32'hbb1f6461),
	.w2(32'hbb7c7dcc),
	.w3(32'hb9647429),
	.w4(32'hbaa86b3c),
	.w5(32'hbacd3317),
	.w6(32'hba6818ca),
	.w7(32'hbaed0b8a),
	.w8(32'hbb68bec5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61929),
	.w1(32'h3b1998ff),
	.w2(32'h3a78fca2),
	.w3(32'hbbe58b1c),
	.w4(32'h3b04cd09),
	.w5(32'hb899bcdf),
	.w6(32'hbbc68fac),
	.w7(32'hbac38ac5),
	.w8(32'hbb1a88e1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule