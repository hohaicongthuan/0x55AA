module layer_6_featuremap_64(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b282998),
	.w1(32'h3a52c434),
	.w2(32'hba7534b5),
	.w3(32'h390ed790),
	.w4(32'hba4f01c4),
	.w5(32'hbaf693bb),
	.w6(32'h3b0a4bdc),
	.w7(32'h3c0d4d5f),
	.w8(32'hbadb746b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389146b2),
	.w1(32'h3b5e21b4),
	.w2(32'hbb0429c6),
	.w3(32'hbc2001e9),
	.w4(32'hbbd0da78),
	.w5(32'hbbd73fc3),
	.w6(32'h3aa0d6f9),
	.w7(32'hbbb9a281),
	.w8(32'hbb84ccac),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ea6b4),
	.w1(32'h3adcf9ef),
	.w2(32'hbb844cf3),
	.w3(32'hbbdc0155),
	.w4(32'hba2eb514),
	.w5(32'h3b6ccefb),
	.w6(32'h3bc10f23),
	.w7(32'hbb3a7be1),
	.w8(32'h3c551aba),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba789141),
	.w1(32'h3b662572),
	.w2(32'hbb29c59f),
	.w3(32'h39c254ea),
	.w4(32'hbb075138),
	.w5(32'hbac53a29),
	.w6(32'hbb178fcb),
	.w7(32'hb9b40a8b),
	.w8(32'hbb8706ff),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86ff65),
	.w1(32'hbc783566),
	.w2(32'h3d2af237),
	.w3(32'hbcb18b14),
	.w4(32'h3d02a21f),
	.w5(32'h3b58b6c4),
	.w6(32'h3d104edd),
	.w7(32'hbd8acd16),
	.w8(32'h3d1bda84),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccba2af),
	.w1(32'hbb26ceab),
	.w2(32'h3b2d30af),
	.w3(32'hbbbe91c8),
	.w4(32'hbb2bdfd2),
	.w5(32'h3a91c10d),
	.w6(32'hbae87c1c),
	.w7(32'h3b3520a3),
	.w8(32'hbab66206),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357691c5),
	.w1(32'h3bb4c92b),
	.w2(32'h3b95cb07),
	.w3(32'hbbbab279),
	.w4(32'h3a8c2fd5),
	.w5(32'h3b1c0d89),
	.w6(32'hbb142f4f),
	.w7(32'h3a708110),
	.w8(32'h3c3986e0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3463a6),
	.w1(32'hba9a6fad),
	.w2(32'h3c5030b0),
	.w3(32'hbc512bf6),
	.w4(32'h3b5c0fd8),
	.w5(32'hbb8ad2ad),
	.w6(32'h3c2b13dd),
	.w7(32'hbbb74563),
	.w8(32'h3cc71296),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28091c),
	.w1(32'hbd03ffef),
	.w2(32'h3db1441d),
	.w3(32'hbc6ebd83),
	.w4(32'h3cf4af34),
	.w5(32'hbc370ef1),
	.w6(32'h3d5fb7d6),
	.w7(32'hbde9ef19),
	.w8(32'h3d89fa2e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ec6ff),
	.w1(32'h3ac33694),
	.w2(32'h3b85cdf6),
	.w3(32'hb96600c9),
	.w4(32'h39b0c401),
	.w5(32'h3a800faf),
	.w6(32'h3aa92ab3),
	.w7(32'h3be8f957),
	.w8(32'h3b3f13f0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc5494),
	.w1(32'h3ba1d2c0),
	.w2(32'hbb0fa20e),
	.w3(32'h3b04918b),
	.w4(32'h3bd95a5d),
	.w5(32'h3b9db823),
	.w6(32'h3bd7c5d8),
	.w7(32'h3bb83ea0),
	.w8(32'h3b035d53),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22ad53),
	.w1(32'hba5bcf64),
	.w2(32'h3a548800),
	.w3(32'h3a9498ce),
	.w4(32'hbbada7f2),
	.w5(32'h3b4a6399),
	.w6(32'hbb9e5265),
	.w7(32'hbba8485a),
	.w8(32'hb9e45356),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be902cf),
	.w1(32'h3b82cfe7),
	.w2(32'hbb7cb5d8),
	.w3(32'hba8d7ee3),
	.w4(32'hba981581),
	.w5(32'h3b8a4eaa),
	.w6(32'h3b512043),
	.w7(32'hbbbec679),
	.w8(32'h3b20d9fc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b205555),
	.w1(32'hbca21ed0),
	.w2(32'h3c9f23db),
	.w3(32'hbc0373ca),
	.w4(32'hbd0f8f8a),
	.w5(32'h3cfa26b4),
	.w6(32'h3bf3dbb0),
	.w7(32'h3bf84e33),
	.w8(32'hbc032c33),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc413128),
	.w1(32'hbb84e06a),
	.w2(32'hbbda10f3),
	.w3(32'hbbb7c25d),
	.w4(32'hbb94fe9a),
	.w5(32'h3b9c03cc),
	.w6(32'h399b7e71),
	.w7(32'hbb5107be),
	.w8(32'hba97f449),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a0e0e),
	.w1(32'h3ac546a6),
	.w2(32'hbb73869a),
	.w3(32'h3a92c457),
	.w4(32'hba1fc693),
	.w5(32'h3acf73a5),
	.w6(32'hba9474d0),
	.w7(32'h3b6164e5),
	.w8(32'hbb394931),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfeda8a),
	.w1(32'hbc4e5550),
	.w2(32'hbc5eb63e),
	.w3(32'hbb9865c1),
	.w4(32'hbc84b0ee),
	.w5(32'hbad80407),
	.w6(32'hbb47ce70),
	.w7(32'hbc942eba),
	.w8(32'hbce99b0b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b166),
	.w1(32'h3ab4c7d3),
	.w2(32'hba9c099e),
	.w3(32'hbb010e32),
	.w4(32'h3a0afeea),
	.w5(32'hbb47ce91),
	.w6(32'hbb827421),
	.w7(32'h3bd28f9d),
	.w8(32'hba24a6bf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6531bb),
	.w1(32'hb8bdfee7),
	.w2(32'h3b0a20f3),
	.w3(32'h39e7e62c),
	.w4(32'h3a526f40),
	.w5(32'hba3e650c),
	.w6(32'h3a377a6a),
	.w7(32'h3a53b032),
	.w8(32'hb950e78f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5f42),
	.w1(32'hbca0c637),
	.w2(32'h3c60d4bc),
	.w3(32'h3bbcd5d4),
	.w4(32'h3c093dce),
	.w5(32'hbc2b6d1d),
	.w6(32'h3c3e9021),
	.w7(32'h3bc5a38b),
	.w8(32'h3b494017),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f971b),
	.w1(32'h3a8e6566),
	.w2(32'hbb2b5bf6),
	.w3(32'hba1e2241),
	.w4(32'hb905e731),
	.w5(32'hb8f4eba7),
	.w6(32'h3a54066f),
	.w7(32'hbb161949),
	.w8(32'hbb48f240),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add9495),
	.w1(32'h3ac98aa8),
	.w2(32'hbb180ca5),
	.w3(32'h3b9eff14),
	.w4(32'hbbd23a2e),
	.w5(32'h3b8ef589),
	.w6(32'h38d6e6a6),
	.w7(32'h3aefebbb),
	.w8(32'hbc09ff1d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07e006),
	.w1(32'h3b33724c),
	.w2(32'hbc019cc0),
	.w3(32'hbb8621e6),
	.w4(32'hbc81db26),
	.w5(32'h3bdde2f2),
	.w6(32'h3b5da0c5),
	.w7(32'h3b116f63),
	.w8(32'hbc814993),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2632c6),
	.w1(32'hbc094744),
	.w2(32'h3b9f70c4),
	.w3(32'hba5a21dc),
	.w4(32'hbbdaf396),
	.w5(32'h3a704593),
	.w6(32'h3ba10575),
	.w7(32'h3c2d7510),
	.w8(32'hbbfe1561),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c414237),
	.w1(32'h3b0f50d8),
	.w2(32'hb8344c66),
	.w3(32'hbb2b9a45),
	.w4(32'hbbc6b719),
	.w5(32'h3b23f3f5),
	.w6(32'hbb5a2e52),
	.w7(32'hbc84917a),
	.w8(32'hbc425ed6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01cb8c),
	.w1(32'h3c269c14),
	.w2(32'h3c5f83bf),
	.w3(32'h3c0e3295),
	.w4(32'h3bc9e96d),
	.w5(32'h3c5a87d4),
	.w6(32'h3c0ebedc),
	.w7(32'h3c4c8646),
	.w8(32'hbb7c455c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dae7a),
	.w1(32'hbb859bcf),
	.w2(32'hbbc6838d),
	.w3(32'hbb3aee2d),
	.w4(32'hbc476341),
	.w5(32'h3a375224),
	.w6(32'hbc3dfd27),
	.w7(32'hbbbec786),
	.w8(32'hbbd1c721),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f84f5),
	.w1(32'h39c5a26d),
	.w2(32'h3a09b788),
	.w3(32'hbb90d840),
	.w4(32'hbaa964bb),
	.w5(32'hba5aca1d),
	.w6(32'hbb139891),
	.w7(32'hbb2021c5),
	.w8(32'h3b8c56ea),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b048e60),
	.w1(32'hbb3bccc3),
	.w2(32'hbb4339fe),
	.w3(32'h3955572e),
	.w4(32'hba0e8ea5),
	.w5(32'hbaeae88f),
	.w6(32'hbaec7910),
	.w7(32'hbb163a75),
	.w8(32'h389082e8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becea23),
	.w1(32'h3d975da9),
	.w2(32'hbbad87c5),
	.w3(32'h3cbe6eb7),
	.w4(32'h3d2c72e8),
	.w5(32'hbd394696),
	.w6(32'hbccf9419),
	.w7(32'h3d3c5778),
	.w8(32'h3da31d4d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0e28b),
	.w1(32'hbc080f1f),
	.w2(32'h3d096226),
	.w3(32'hbceb103b),
	.w4(32'h3ca32381),
	.w5(32'hbbdc0c41),
	.w6(32'h3cebceb3),
	.w7(32'hbd473f24),
	.w8(32'h3ca1d746),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73f61d),
	.w1(32'h3b9e4864),
	.w2(32'h3c15962d),
	.w3(32'h3b79ad50),
	.w4(32'h3c20aa0a),
	.w5(32'h3c8bf8f5),
	.w6(32'h3b8a8182),
	.w7(32'h3c9295ec),
	.w8(32'h3c94d3cb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1932b),
	.w1(32'h3bec8274),
	.w2(32'hbca1d4a7),
	.w3(32'h3b9d87d2),
	.w4(32'hbc16ee08),
	.w5(32'h3be31e60),
	.w6(32'hbc680927),
	.w7(32'h3c53ba86),
	.w8(32'hbc2dcb01),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cdd0a),
	.w1(32'hbc744533),
	.w2(32'h3dc25c0e),
	.w3(32'h3cabdef6),
	.w4(32'h3ce68cd5),
	.w5(32'h3d5408cd),
	.w6(32'h3dad04e7),
	.w7(32'h3dc9349b),
	.w8(32'h3c6b3713),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d891496),
	.w1(32'h3ab880a8),
	.w2(32'h3a875814),
	.w3(32'h3af20b7f),
	.w4(32'hbb2d52e8),
	.w5(32'h3aa14461),
	.w6(32'h3b44a37a),
	.w7(32'h3b369f7f),
	.w8(32'hba9175d1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10bbf7),
	.w1(32'h3bd038d3),
	.w2(32'h39a2b8a3),
	.w3(32'h3b1ef1b6),
	.w4(32'h3afebb68),
	.w5(32'h3c02cb93),
	.w6(32'h3aaabc2b),
	.w7(32'hba80d4f5),
	.w8(32'hbabeb806),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb170d6),
	.w1(32'hbbba08f1),
	.w2(32'hb84e863f),
	.w3(32'hbbadc21e),
	.w4(32'hbb560a51),
	.w5(32'h39044057),
	.w6(32'h3b61469e),
	.w7(32'h3b8a3bc7),
	.w8(32'hbb59da63),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed28b5),
	.w1(32'h3ad23937),
	.w2(32'h3b52dec0),
	.w3(32'h3aaa08fc),
	.w4(32'h3aba4a14),
	.w5(32'h3a755cf3),
	.w6(32'h3abda08a),
	.w7(32'h3b226d1d),
	.w8(32'h3a55505a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636f29),
	.w1(32'hbc9679d6),
	.w2(32'hbb21ed3c),
	.w3(32'hbc4de97c),
	.w4(32'hbb261e4a),
	.w5(32'hbc125181),
	.w6(32'hbbb2f970),
	.w7(32'hbca722b5),
	.w8(32'hbc8fb12b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10cd9d),
	.w1(32'hbc842697),
	.w2(32'h3d403a01),
	.w3(32'hbc5fe903),
	.w4(32'h3d21e4f0),
	.w5(32'hbcff5763),
	.w6(32'h3d124b6e),
	.w7(32'hbd959be7),
	.w8(32'h3daa7139),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1528ab),
	.w1(32'h3b7f91af),
	.w2(32'h3a12de03),
	.w3(32'hbbfa7843),
	.w4(32'h3bd512b8),
	.w5(32'h3b8eac38),
	.w6(32'h3c3be7b8),
	.w7(32'hbb0b3055),
	.w8(32'hbb8c9e32),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a511),
	.w1(32'hba8ce4d2),
	.w2(32'hbb4dfbe3),
	.w3(32'h395765e8),
	.w4(32'hba7a2160),
	.w5(32'hbae96335),
	.w6(32'hbab697c0),
	.w7(32'h3a66b2a7),
	.w8(32'hbac9fef5),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6839c7),
	.w1(32'hbba5a089),
	.w2(32'hbb7b3904),
	.w3(32'hb9179ad4),
	.w4(32'hbaf8f7a7),
	.w5(32'h3b67ef60),
	.w6(32'h39cd3396),
	.w7(32'h3b873d60),
	.w8(32'h3b43d83f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17d2c7),
	.w1(32'h3b83d53f),
	.w2(32'h3c0aef20),
	.w3(32'h3beee0d4),
	.w4(32'h3b80dced),
	.w5(32'h3bdbc84b),
	.w6(32'hba30e76b),
	.w7(32'hbbb3c3a0),
	.w8(32'h3b0109d8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9afd74),
	.w1(32'h3a76be5c),
	.w2(32'hbbd6ba74),
	.w3(32'h383b2d05),
	.w4(32'hbac90e69),
	.w5(32'hbb72492e),
	.w6(32'hba567356),
	.w7(32'hbb956746),
	.w8(32'hbb45c9c4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94a07f),
	.w1(32'hbc922164),
	.w2(32'hbd23d3f6),
	.w3(32'hbbed6e68),
	.w4(32'hbca98443),
	.w5(32'hbce319b5),
	.w6(32'hbcfc9bd0),
	.w7(32'hbc1c6679),
	.w8(32'hbc326e1e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21dd5a),
	.w1(32'h3be8a189),
	.w2(32'h3ba63ef6),
	.w3(32'hbc3f9216),
	.w4(32'hbad03c3c),
	.w5(32'hbac6dd1a),
	.w6(32'h3aee11fb),
	.w7(32'hbc2155d2),
	.w8(32'h3b8df3c8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bc5ba),
	.w1(32'hbcbe3538),
	.w2(32'hbc5a5bdc),
	.w3(32'h3a1b0889),
	.w4(32'hbba8414a),
	.w5(32'h3c018d3d),
	.w6(32'hbb212424),
	.w7(32'hbc23641f),
	.w8(32'h3ba0f472),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62764f),
	.w1(32'h3b8026e3),
	.w2(32'hb9abe956),
	.w3(32'h3ac99d3b),
	.w4(32'h3b442c50),
	.w5(32'h3b8ab16c),
	.w6(32'h3b24b2f0),
	.w7(32'h38cab69d),
	.w8(32'h3b70fb0b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b364d60),
	.w1(32'h3d02e230),
	.w2(32'hbd410478),
	.w3(32'h3c46f6de),
	.w4(32'hbced34a2),
	.w5(32'h3c953bd3),
	.w6(32'hbd5a0c7f),
	.w7(32'h3d81deba),
	.w8(32'hbd4acbe1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4a6395),
	.w1(32'h3b77f2f6),
	.w2(32'hba2bed5a),
	.w3(32'hbab7132c),
	.w4(32'h3adee30b),
	.w5(32'h3a95d9f7),
	.w6(32'h395ea3dc),
	.w7(32'h3b8ebed5),
	.w8(32'hbb9115ee),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1c3bb),
	.w1(32'h3a7bb1f2),
	.w2(32'h3a28d921),
	.w3(32'hb9bdd3b6),
	.w4(32'hba71fa55),
	.w5(32'hbac9e0ef),
	.w6(32'h3971448c),
	.w7(32'hb901446d),
	.w8(32'h3b13ead6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8a0bc),
	.w1(32'h3b7ba564),
	.w2(32'h3b0b4c6b),
	.w3(32'h3b7e78aa),
	.w4(32'hba9c7ce5),
	.w5(32'h3b4c562b),
	.w6(32'h3bbeee69),
	.w7(32'hba48e7d5),
	.w8(32'h38f9bb05),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405867),
	.w1(32'h3b8f0fc8),
	.w2(32'h3b5a0014),
	.w3(32'h3b5f2b9f),
	.w4(32'h3b509e9b),
	.w5(32'h3bb710a3),
	.w6(32'h3c33f14e),
	.w7(32'h3bde9f4e),
	.w8(32'h3c23a761),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2bc61),
	.w1(32'h3b9289ff),
	.w2(32'h3b197651),
	.w3(32'h39b9a046),
	.w4(32'hbacad788),
	.w5(32'hbb109fd0),
	.w6(32'h3afc6bf5),
	.w7(32'h3b534b4b),
	.w8(32'hba6ea298),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94c39e),
	.w1(32'h3b09bc09),
	.w2(32'h3b561350),
	.w3(32'h3a69984d),
	.w4(32'h3ab170bd),
	.w5(32'h3a400785),
	.w6(32'hbcdeff0b),
	.w7(32'hbce962d2),
	.w8(32'hbd0231d3),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1433be),
	.w1(32'hbb96c4e6),
	.w2(32'hbaef1d42),
	.w3(32'hbb81fc3f),
	.w4(32'hbb637a9b),
	.w5(32'hbb1119ad),
	.w6(32'hbb80dfa2),
	.w7(32'hbaff4e5b),
	.w8(32'hbae031bf),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a39980),
	.w1(32'hbbb7a46d),
	.w2(32'h39b12cb6),
	.w3(32'hbb381de6),
	.w4(32'h3b91bcf0),
	.w5(32'hba9abc7c),
	.w6(32'h3c99cdf9),
	.w7(32'h3cd7ba75),
	.w8(32'h3ccd4361),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c0fcc),
	.w1(32'h3ace347a),
	.w2(32'h3b133be0),
	.w3(32'hba633607),
	.w4(32'hba09f111),
	.w5(32'h3a3a90c0),
	.w6(32'h3acdbd1d),
	.w7(32'h3b0d83b7),
	.w8(32'h3b65a73a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4f5b),
	.w1(32'h3b98b598),
	.w2(32'h3bc070ee),
	.w3(32'hbc2a72d2),
	.w4(32'hbc1dac76),
	.w5(32'h39ba3cfd),
	.w6(32'h3c27ea42),
	.w7(32'h3c4299c9),
	.w8(32'h3c66b51c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b8ed),
	.w1(32'h3b6b86d3),
	.w2(32'h3b1c857f),
	.w3(32'hba33fa4b),
	.w4(32'hbab5b111),
	.w5(32'hba84f55c),
	.w6(32'h3b6b91c2),
	.w7(32'h3bb157c1),
	.w8(32'h3bdd819f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9b772),
	.w1(32'h3b6d0e08),
	.w2(32'hbb5cac23),
	.w3(32'hbb0d9327),
	.w4(32'hbafa302e),
	.w5(32'h3a85b4da),
	.w6(32'hb97151c5),
	.w7(32'hbba7e2f7),
	.w8(32'hbab4e598),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd87a),
	.w1(32'hbc555047),
	.w2(32'hbc863e2a),
	.w3(32'hbbda8135),
	.w4(32'hbbc4cd45),
	.w5(32'hbc0bea3f),
	.w6(32'hbce20b2d),
	.w7(32'hbca55cc1),
	.w8(32'hbcbb21e5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978f7bc),
	.w1(32'h3b5b1116),
	.w2(32'h3c1af69b),
	.w3(32'hbbe2d172),
	.w4(32'hbb8d346a),
	.w5(32'hbba53afa),
	.w6(32'hb92b694a),
	.w7(32'h3b8e5fe2),
	.w8(32'h3bb1d938),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule