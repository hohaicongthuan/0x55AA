module layer_10_featuremap_262(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2562f),
	.w1(32'h3c0b0396),
	.w2(32'h3b43c3fc),
	.w3(32'hbb8a2607),
	.w4(32'h3aff453b),
	.w5(32'hba851b85),
	.w6(32'hbb50b915),
	.w7(32'hbb5529e6),
	.w8(32'hbbcd8f25),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d06b5),
	.w1(32'hbbc453f3),
	.w2(32'hbb5c4477),
	.w3(32'hbb7a38bb),
	.w4(32'hbb456981),
	.w5(32'hbadaa19e),
	.w6(32'hbbc36de6),
	.w7(32'hbbe9ce15),
	.w8(32'h3af97ffd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41d94f),
	.w1(32'h3b2401a9),
	.w2(32'h3bfadba3),
	.w3(32'h3aa43a38),
	.w4(32'h38c2bc23),
	.w5(32'hbae8e739),
	.w6(32'h3aa84d6e),
	.w7(32'h3bcf1fde),
	.w8(32'hbb8ebc6e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872e91),
	.w1(32'hbb6759d8),
	.w2(32'hbb83d5b6),
	.w3(32'h3a7c649f),
	.w4(32'hb92d426f),
	.w5(32'h3b088c60),
	.w6(32'hba9aa1e3),
	.w7(32'hbad1d4e0),
	.w8(32'hbb3d46ba),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29ef8b),
	.w1(32'hbb83840d),
	.w2(32'h3b12e5c0),
	.w3(32'hbb02f145),
	.w4(32'hbb37ea13),
	.w5(32'hbae8bf14),
	.w6(32'h39dbc51c),
	.w7(32'hb9326a54),
	.w8(32'hbaa5c1c4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33fb13),
	.w1(32'h3b020f84),
	.w2(32'h3b1440ba),
	.w3(32'hba8e9da8),
	.w4(32'h3aac7bed),
	.w5(32'hba48700e),
	.w6(32'h3a678b85),
	.w7(32'hba66e56b),
	.w8(32'hbba03dda),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a55f),
	.w1(32'hbb3481f9),
	.w2(32'hb98871c8),
	.w3(32'hbba28459),
	.w4(32'hbb43621b),
	.w5(32'hb9947a45),
	.w6(32'hbb7718ce),
	.w7(32'hbb22b3dd),
	.w8(32'hbbe82fd7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092dd9),
	.w1(32'hbb02871f),
	.w2(32'hbb6ae9f1),
	.w3(32'hba09d0bc),
	.w4(32'h3c1117de),
	.w5(32'hb937d567),
	.w6(32'hbbb81a5b),
	.w7(32'hba08f882),
	.w8(32'hbb29089e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a918e6d),
	.w1(32'h3b3bd536),
	.w2(32'h3b38dea4),
	.w3(32'hba8b20b2),
	.w4(32'hbb247f36),
	.w5(32'hb7f83f7e),
	.w6(32'hbb549ae3),
	.w7(32'hbb23b97e),
	.w8(32'h3ae26f3a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900765e),
	.w1(32'h3ae65e88),
	.w2(32'h3b0cbfc9),
	.w3(32'hbb370fa0),
	.w4(32'hbafd09cf),
	.w5(32'hb943ce43),
	.w6(32'h3b673f94),
	.w7(32'hb948f7ec),
	.w8(32'h3ab9bf8f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510cb8),
	.w1(32'h3acf50fa),
	.w2(32'h39dbc1c5),
	.w3(32'hba21f260),
	.w4(32'h3adf65d6),
	.w5(32'hbabe974b),
	.w6(32'h3ab47d80),
	.w7(32'hba9f79a0),
	.w8(32'hbb363fed),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad64083),
	.w1(32'h3bcc77c0),
	.w2(32'h3bc87cbb),
	.w3(32'h3a0dac82),
	.w4(32'h3b908b3f),
	.w5(32'hbb5d0fa4),
	.w6(32'hbadbb293),
	.w7(32'h3b5dfcf9),
	.w8(32'h38eb2e66),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79c35fb),
	.w1(32'h3b6829c7),
	.w2(32'hbb5882f1),
	.w3(32'hba4d37ed),
	.w4(32'h3b876247),
	.w5(32'hb92a4abe),
	.w6(32'hbb8d797f),
	.w7(32'hbb1522d7),
	.w8(32'h3abb18ce),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54a8d5),
	.w1(32'h3c0fed3f),
	.w2(32'h3bf0ae07),
	.w3(32'hbb9c63cd),
	.w4(32'hbaeae232),
	.w5(32'hba799bab),
	.w6(32'h3b81dad2),
	.w7(32'h3b5f6604),
	.w8(32'hbb6f2ecf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe061),
	.w1(32'h3b45b436),
	.w2(32'h3a33ee8a),
	.w3(32'h3acaee49),
	.w4(32'h3ad1542c),
	.w5(32'hbafeca7e),
	.w6(32'h3ba01645),
	.w7(32'h3b8cdfc5),
	.w8(32'hbb2f0d26),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5505b),
	.w1(32'hba9690b2),
	.w2(32'hba977497),
	.w3(32'hbb4647d2),
	.w4(32'hbaeb595a),
	.w5(32'hbba134b4),
	.w6(32'hbbc3d43d),
	.w7(32'h391affb0),
	.w8(32'hbb982101),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46c060),
	.w1(32'hb908f165),
	.w2(32'hbbc2e8bb),
	.w3(32'h397a634c),
	.w4(32'hba1492a8),
	.w5(32'hba886346),
	.w6(32'hbbbfa29a),
	.w7(32'hbbbab629),
	.w8(32'h3a19fc1a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b4760),
	.w1(32'h3afae521),
	.w2(32'h3ac06ee9),
	.w3(32'h379c39ff),
	.w4(32'h3adfca51),
	.w5(32'hbacb5760),
	.w6(32'h3ad62e0d),
	.w7(32'h3a0fbf91),
	.w8(32'h3b2b55ff),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ebacb),
	.w1(32'h3b2ec521),
	.w2(32'h3aa76802),
	.w3(32'hba3fd9d3),
	.w4(32'h3b3d44ee),
	.w5(32'h3b29c2ad),
	.w6(32'h3b1b5ea8),
	.w7(32'hb94779d9),
	.w8(32'h3b3b32da),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b71a),
	.w1(32'h3a90f73c),
	.w2(32'h3bd03446),
	.w3(32'hbaaa48b6),
	.w4(32'hba81a1c1),
	.w5(32'hbb4d61cb),
	.w6(32'h3bdc8c2a),
	.w7(32'h3ba943ce),
	.w8(32'hbb94981e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba096c32),
	.w1(32'h3b1828e7),
	.w2(32'hbad9c53a),
	.w3(32'hbb220b44),
	.w4(32'hbb15138d),
	.w5(32'h3bbc54ff),
	.w6(32'hbb39c7a6),
	.w7(32'hbb137658),
	.w8(32'hb9ebfe15),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25dbfb),
	.w1(32'hbb5e8243),
	.w2(32'hbb07a418),
	.w3(32'h3b6c5c63),
	.w4(32'h393ef3ec),
	.w5(32'hbb804681),
	.w6(32'h39fdeac7),
	.w7(32'h3a527bb3),
	.w8(32'hba80008d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8dd18),
	.w1(32'h3b281c55),
	.w2(32'hba4afd16),
	.w3(32'hba643ee8),
	.w4(32'hbb352c98),
	.w5(32'hbb5fc524),
	.w6(32'hbb1d044b),
	.w7(32'hbb9f01e8),
	.w8(32'hbb4a39fa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09b0d4),
	.w1(32'hba8c7dc8),
	.w2(32'h3ac261ae),
	.w3(32'hbb8156e0),
	.w4(32'hbbe4f507),
	.w5(32'h3b68eb77),
	.w6(32'hbba407ee),
	.w7(32'hbbf0fcb0),
	.w8(32'h3c8f106c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f9802),
	.w1(32'h3af93b16),
	.w2(32'h3c30d9a6),
	.w3(32'hbab261de),
	.w4(32'hbba1c518),
	.w5(32'hbb4b5a0e),
	.w6(32'h3c45f7b7),
	.w7(32'h3b2a1601),
	.w8(32'hba463cff),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cf8ee),
	.w1(32'h398bedb9),
	.w2(32'hbabe139a),
	.w3(32'h3b0747e0),
	.w4(32'h3b067336),
	.w5(32'h3b80baa8),
	.w6(32'h3aee7b34),
	.w7(32'hba48c9cf),
	.w8(32'hb91bb47a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf785f),
	.w1(32'hbb361a1d),
	.w2(32'h3a50455e),
	.w3(32'h3b8444a4),
	.w4(32'h3b7eabe3),
	.w5(32'h3ae44c67),
	.w6(32'hbb1ee327),
	.w7(32'h3b3e4e99),
	.w8(32'h3c0ac61d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b8b5),
	.w1(32'h3c34a7b3),
	.w2(32'h3bf2b910),
	.w3(32'hbbc6bc1e),
	.w4(32'hbafdbd6c),
	.w5(32'hbafdc3a4),
	.w6(32'hbb8a6aa0),
	.w7(32'hbaf83e6f),
	.w8(32'h3be27bdc),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76cb22),
	.w1(32'h3a5b4806),
	.w2(32'h3b13f943),
	.w3(32'hbbf6419a),
	.w4(32'hbbf51523),
	.w5(32'hbc051507),
	.w6(32'h3c6f0771),
	.w7(32'h3b68b8e0),
	.w8(32'h3b11c5ce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e815f),
	.w1(32'h3bfc1cfc),
	.w2(32'h3b966f39),
	.w3(32'hbbda8af6),
	.w4(32'hbb9ac80b),
	.w5(32'h3b96a768),
	.w6(32'h3b849bed),
	.w7(32'hba99c686),
	.w8(32'h3c3c9504),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d3d9f),
	.w1(32'h3b9133f4),
	.w2(32'h3c4c51c9),
	.w3(32'hbaa84bb7),
	.w4(32'hbb2e4af9),
	.w5(32'h3baf5cdf),
	.w6(32'h3bf897b8),
	.w7(32'hbb5477ff),
	.w8(32'h3b255427),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b768af5),
	.w1(32'h3b67e1e6),
	.w2(32'h39665334),
	.w3(32'h3b57ff4f),
	.w4(32'h3b268f4a),
	.w5(32'hb79751e0),
	.w6(32'h3c2e2ba7),
	.w7(32'h3bb4edb6),
	.w8(32'h3ada97dd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a03c0c),
	.w1(32'hbb2b9596),
	.w2(32'h3ba4836c),
	.w3(32'h3a9645a2),
	.w4(32'h3b63490d),
	.w5(32'hbb1898dc),
	.w6(32'h39671a4e),
	.w7(32'h3b5b086d),
	.w8(32'hbb002953),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a305f7f),
	.w1(32'hb94ac554),
	.w2(32'hbad22c34),
	.w3(32'hba4e7822),
	.w4(32'h3a8a4e47),
	.w5(32'h3bf4f444),
	.w6(32'h3a0e6fd9),
	.w7(32'hbb912ad1),
	.w8(32'h3bc71927),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8b655),
	.w1(32'h3aedaee5),
	.w2(32'h3b9f3397),
	.w3(32'hbab3d9ee),
	.w4(32'h3ae1f8a9),
	.w5(32'hbb473178),
	.w6(32'h3c090d6d),
	.w7(32'h3bacc4b9),
	.w8(32'hbb5f0622),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a486326),
	.w1(32'h3b1b546b),
	.w2(32'h3b9907c7),
	.w3(32'hba9ea596),
	.w4(32'h3a25d0d7),
	.w5(32'h3b66eb65),
	.w6(32'hbbb648e1),
	.w7(32'hbc19fa8d),
	.w8(32'h3c4161c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4bfb),
	.w1(32'hbad5efea),
	.w2(32'h3b8adf11),
	.w3(32'hbb9ec385),
	.w4(32'hb95cc703),
	.w5(32'h3b5cc363),
	.w6(32'h3c1079d9),
	.w7(32'h3a118242),
	.w8(32'h3b02f179),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce04b5),
	.w1(32'hbb64d02a),
	.w2(32'h38f01828),
	.w3(32'h3aa531d5),
	.w4(32'hbacb6f44),
	.w5(32'h3a561463),
	.w6(32'hbb0f56f7),
	.w7(32'hbae528d9),
	.w8(32'h3c21c124),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1569),
	.w1(32'hbbdde5f2),
	.w2(32'h3af01ad3),
	.w3(32'hbb431dc1),
	.w4(32'hbb77ec90),
	.w5(32'hbba97904),
	.w6(32'h3cacb75a),
	.w7(32'h3aed4e74),
	.w8(32'hbbeb3749),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb930cd1),
	.w1(32'hbb0ce230),
	.w2(32'hbb971dde),
	.w3(32'hbb8595af),
	.w4(32'hbb93c49a),
	.w5(32'hb9c4de68),
	.w6(32'hb9dcaac8),
	.w7(32'hbab7f3d3),
	.w8(32'hba505303),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ba3d),
	.w1(32'h3b789aae),
	.w2(32'hbad45670),
	.w3(32'hbbbfdbec),
	.w4(32'h3883ab2c),
	.w5(32'hba3fda8a),
	.w6(32'hba5e56bf),
	.w7(32'hba6b5d68),
	.w8(32'hbb08257d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f0444),
	.w1(32'hbb5077f0),
	.w2(32'hbb5d6ad1),
	.w3(32'h39811db8),
	.w4(32'h3a0aac30),
	.w5(32'hbb35ae0a),
	.w6(32'hba371cb1),
	.w7(32'hb8781d23),
	.w8(32'h34188e72),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3960ecdc),
	.w1(32'hbb102046),
	.w2(32'h3b91342a),
	.w3(32'hbaab8f6f),
	.w4(32'hbb63ef8c),
	.w5(32'h39847b66),
	.w6(32'hba16e76b),
	.w7(32'h3b11c53e),
	.w8(32'hbc09a9c4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf9a5a),
	.w1(32'hb9f92a7a),
	.w2(32'h3b5f627c),
	.w3(32'hba964c3e),
	.w4(32'h3b89d9c2),
	.w5(32'hbba19e51),
	.w6(32'hbb4580c9),
	.w7(32'hb81a7286),
	.w8(32'hbc054ac1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8f93),
	.w1(32'hbb248319),
	.w2(32'hba001309),
	.w3(32'hbb0d9226),
	.w4(32'hba2c811e),
	.w5(32'h3b5fcbe3),
	.w6(32'hbb56a136),
	.w7(32'hbb74a14b),
	.w8(32'h3ba12f77),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beffe76),
	.w1(32'h3b8026ef),
	.w2(32'h38dfce7d),
	.w3(32'h3b7d0027),
	.w4(32'h3ae785d1),
	.w5(32'h3ad43c82),
	.w6(32'h3bc58e8f),
	.w7(32'h3aa52fb8),
	.w8(32'hbaaa5f19),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e50f25),
	.w1(32'h397c1aed),
	.w2(32'h39fd0d93),
	.w3(32'h3ae423f6),
	.w4(32'h3b60f09b),
	.w5(32'h3b8c7760),
	.w6(32'hbb0363fa),
	.w7(32'h3a788e5f),
	.w8(32'h3b5346d6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0e1a),
	.w1(32'hba6b6a80),
	.w2(32'h3b146962),
	.w3(32'hbb007df3),
	.w4(32'hbb6909c0),
	.w5(32'h3ab0216f),
	.w6(32'h3b09210f),
	.w7(32'h3aa86c36),
	.w8(32'h3c07d127),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d4495),
	.w1(32'h3b342e24),
	.w2(32'h3aba0c59),
	.w3(32'h3aed5831),
	.w4(32'h3b4badb5),
	.w5(32'h3bede4f3),
	.w6(32'h3b13a1d6),
	.w7(32'hbb502af3),
	.w8(32'h3b2b4a85),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9abc82),
	.w1(32'hba0ceb5a),
	.w2(32'h3a96bc0d),
	.w3(32'h3b618323),
	.w4(32'h3b4fc517),
	.w5(32'hba5c8568),
	.w6(32'h3b2b597b),
	.w7(32'h3bd2dbac),
	.w8(32'hbbf74246),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4758c),
	.w1(32'hb8117146),
	.w2(32'hbb846b9a),
	.w3(32'hbb91220a),
	.w4(32'hbb8bc195),
	.w5(32'hbb37279b),
	.w6(32'hb9014b1c),
	.w7(32'hbb936043),
	.w8(32'hbbb56a95),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac22ee7),
	.w1(32'hbb3e83e3),
	.w2(32'hbb2000a5),
	.w3(32'h3b3a2e2c),
	.w4(32'hb9e79008),
	.w5(32'hba8ae92b),
	.w6(32'hbb955ce9),
	.w7(32'hbb7c8760),
	.w8(32'hbb1f3977),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba227ab),
	.w1(32'h3bfc5d7d),
	.w2(32'hb8ef27b0),
	.w3(32'hbb4544c3),
	.w4(32'hbb1b868e),
	.w5(32'hba339b09),
	.w6(32'hbb0dee67),
	.w7(32'hbb2108cb),
	.w8(32'h3a934da2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39f56a),
	.w1(32'hbb2d1470),
	.w2(32'hb824e01c),
	.w3(32'hbc20c2df),
	.w4(32'h3b386da4),
	.w5(32'h398bc1e4),
	.w6(32'hbb77c525),
	.w7(32'h3af691c7),
	.w8(32'h3a812801),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad08c2d),
	.w1(32'hba39c969),
	.w2(32'hba9b77c4),
	.w3(32'hbae7e7b0),
	.w4(32'hbb3d343d),
	.w5(32'h3b6316f2),
	.w6(32'h3af2b05e),
	.w7(32'hba110e63),
	.w8(32'h3beed314),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eedd6),
	.w1(32'hbb97c4a8),
	.w2(32'h3b08c85c),
	.w3(32'hba4da6ef),
	.w4(32'hbb68bfd1),
	.w5(32'h39e14014),
	.w6(32'h3c6942fe),
	.w7(32'h3be05d0c),
	.w8(32'h3bc61dcc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cbe41),
	.w1(32'h3abff675),
	.w2(32'h3b0bac53),
	.w3(32'hbb1b872f),
	.w4(32'hbae712f7),
	.w5(32'hbb04cc22),
	.w6(32'h3bd03e2a),
	.w7(32'h3a9b1dcd),
	.w8(32'h39d046fb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a09c0),
	.w1(32'h3b311ef8),
	.w2(32'hbbbbe9dd),
	.w3(32'hbc0488f7),
	.w4(32'hba9558d1),
	.w5(32'h3bb128e7),
	.w6(32'hbb061b94),
	.w7(32'hbaeecee8),
	.w8(32'h3a8055b3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb7e11),
	.w1(32'hbaaa260a),
	.w2(32'hbae6d751),
	.w3(32'h3b3e88ca),
	.w4(32'h3af3280e),
	.w5(32'h3bce3b3c),
	.w6(32'h39eff960),
	.w7(32'h3ba2e2d8),
	.w8(32'hbaad7810),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1c08f),
	.w1(32'hbc4852b6),
	.w2(32'hbbefe157),
	.w3(32'h3be0a93d),
	.w4(32'h3b39dc61),
	.w5(32'h3c0ca5da),
	.w6(32'hbade71bf),
	.w7(32'h3b8975af),
	.w8(32'h3c370e7c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b79d),
	.w1(32'hbb77d483),
	.w2(32'hba80ad5e),
	.w3(32'h3bb49628),
	.w4(32'h3b254ce8),
	.w5(32'hbb612668),
	.w6(32'h3ce58d20),
	.w7(32'h3c6f5ca7),
	.w8(32'h3a86f7f9),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac60ea9),
	.w1(32'h3a4344c3),
	.w2(32'hbb4e1133),
	.w3(32'h38810ca3),
	.w4(32'h3b4cb2b5),
	.w5(32'h3b7490d0),
	.w6(32'h3aafff9f),
	.w7(32'h3aa57f7d),
	.w8(32'h3a3963e5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c417),
	.w1(32'hba8a6604),
	.w2(32'h3b293388),
	.w3(32'hb792c364),
	.w4(32'h3b016fd4),
	.w5(32'h3b460a37),
	.w6(32'h39c463f0),
	.w7(32'h3b543743),
	.w8(32'h3bad6a2a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac97b02),
	.w1(32'h3b8fc485),
	.w2(32'h3b71cacb),
	.w3(32'hbbc5215c),
	.w4(32'hb9f4c244),
	.w5(32'h3a149164),
	.w6(32'h3bcc75d3),
	.w7(32'h3aed57be),
	.w8(32'h3b8744b5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d88df),
	.w1(32'hbb6a18ea),
	.w2(32'h3ae867bd),
	.w3(32'hbb6ee690),
	.w4(32'hbbb942c7),
	.w5(32'hb9fa591b),
	.w6(32'h3bc67541),
	.w7(32'h3b8c4189),
	.w8(32'hb979b949),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd495b9),
	.w1(32'hba04ce33),
	.w2(32'h3ac7c97c),
	.w3(32'hbb3392ff),
	.w4(32'hbae93c4a),
	.w5(32'h37a8998b),
	.w6(32'h3aa1accd),
	.w7(32'hb9a06bcd),
	.w8(32'hbaa71c96),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398458b2),
	.w1(32'h3be3090a),
	.w2(32'h3a6f2a76),
	.w3(32'h39cb4ba2),
	.w4(32'h3c08ccb6),
	.w5(32'hbaffa71b),
	.w6(32'h3acfcd05),
	.w7(32'h3b4d4e4a),
	.w8(32'hb9a1ad3c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8449bc),
	.w1(32'hbb677afc),
	.w2(32'hbc07853b),
	.w3(32'hbb8cc2eb),
	.w4(32'hbc0b5abc),
	.w5(32'h3aaa88fd),
	.w6(32'hba0201b1),
	.w7(32'hbc264edb),
	.w8(32'h3b156bdf),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b199862),
	.w1(32'h3875c5f8),
	.w2(32'h3b076395),
	.w3(32'h39b894a6),
	.w4(32'hbb0bdcd9),
	.w5(32'h3b16b8a7),
	.w6(32'h395cef41),
	.w7(32'h3ad37d62),
	.w8(32'h3a9e8582),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1003d8),
	.w1(32'h3b5c4346),
	.w2(32'hb9aef110),
	.w3(32'h3bd79d6c),
	.w4(32'h3b5e2a7e),
	.w5(32'h3977f3af),
	.w6(32'h3b9ac758),
	.w7(32'hbb8f869e),
	.w8(32'hbb4ee179),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb523ada),
	.w1(32'hbb7702ef),
	.w2(32'h3a21d4d1),
	.w3(32'hb9839b46),
	.w4(32'h3aa74094),
	.w5(32'h3af85bf6),
	.w6(32'hbb061659),
	.w7(32'h39ccd5b5),
	.w8(32'h3bc74f17),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ce4a),
	.w1(32'h3a866a51),
	.w2(32'hbb4a6d5e),
	.w3(32'h3a9e47ed),
	.w4(32'h39ba14ca),
	.w5(32'hbb54637b),
	.w6(32'h38a4fe78),
	.w7(32'hbc075fb0),
	.w8(32'h3a1a7cdf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb626b8f),
	.w1(32'hbb834d43),
	.w2(32'h3b52c011),
	.w3(32'hbac0a41e),
	.w4(32'hbad9c788),
	.w5(32'hbb9c0442),
	.w6(32'hbbc05877),
	.w7(32'hbc0fbbbf),
	.w8(32'h3a04d0b7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f83672),
	.w1(32'h37978387),
	.w2(32'h3b9b4f47),
	.w3(32'hbbcd05c7),
	.w4(32'h3b03bef3),
	.w5(32'hbac1802c),
	.w6(32'h3ba23577),
	.w7(32'hbb434cec),
	.w8(32'hbb3b2c88),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a791270),
	.w1(32'h3b807e2b),
	.w2(32'h3ad0fb30),
	.w3(32'hbb1fbe4c),
	.w4(32'h3acd61c5),
	.w5(32'hbb983122),
	.w6(32'h3965f2d4),
	.w7(32'hbae3f6fd),
	.w8(32'h3b1cd133),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba547328),
	.w1(32'h3b78a010),
	.w2(32'h3b4d5b3a),
	.w3(32'hbb0452e3),
	.w4(32'hbb313826),
	.w5(32'hbaed3bc4),
	.w6(32'h39df3a90),
	.w7(32'hbbc5af10),
	.w8(32'hb8a37969),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae35bda),
	.w1(32'h3b1bc2bb),
	.w2(32'h3a01b357),
	.w3(32'hbb2bd812),
	.w4(32'hb934b566),
	.w5(32'h3a1345f3),
	.w6(32'hba52983f),
	.w7(32'hbb146ec0),
	.w8(32'hb918bc9d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80c961),
	.w1(32'h3a6736c1),
	.w2(32'hb8a0df1e),
	.w3(32'h3b860074),
	.w4(32'h3b01ff67),
	.w5(32'h3b6e0ee4),
	.w6(32'h3b2364af),
	.w7(32'hbb098c9d),
	.w8(32'h3b18630d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ccc6),
	.w1(32'h3b6d58c4),
	.w2(32'hb9d7bd1b),
	.w3(32'h3bbaa540),
	.w4(32'h3bc08740),
	.w5(32'hbad41f7f),
	.w6(32'h3b0a96b4),
	.w7(32'h3b32d5a1),
	.w8(32'hbb090178),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b191ccf),
	.w1(32'h3af26643),
	.w2(32'hbac5911a),
	.w3(32'hbb3828c9),
	.w4(32'h3a32ea23),
	.w5(32'h3b6ce512),
	.w6(32'hba94adec),
	.w7(32'hbc0cc70f),
	.w8(32'hbac73613),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b44b5),
	.w1(32'h38fa31fc),
	.w2(32'h3952e371),
	.w3(32'h3b78f492),
	.w4(32'h3b083443),
	.w5(32'hbada2a72),
	.w6(32'hbb1b3357),
	.w7(32'h3a89ef9e),
	.w8(32'h3b8b2c80),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b184127),
	.w1(32'h3b547797),
	.w2(32'h3bc20ffe),
	.w3(32'h3940be2f),
	.w4(32'h3af4a444),
	.w5(32'hbba00d55),
	.w6(32'h3b8dc7ba),
	.w7(32'hbb036812),
	.w8(32'h3a1f6e66),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae82418),
	.w1(32'hb9fbee8c),
	.w2(32'h3a440155),
	.w3(32'hba5ceb32),
	.w4(32'hba9d83bc),
	.w5(32'hbafecf38),
	.w6(32'hbb570cc3),
	.w7(32'hbafbb14a),
	.w8(32'h3b08e824),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09f3a0),
	.w1(32'h3b62e562),
	.w2(32'hba8dde58),
	.w3(32'h3c01cad4),
	.w4(32'h38e8966b),
	.w5(32'hbb08f2a9),
	.w6(32'h3b6ee4a3),
	.w7(32'hbb14d7e3),
	.w8(32'h3b5c81fa),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92535d),
	.w1(32'h3ab254c9),
	.w2(32'h39c784e9),
	.w3(32'hbb1ba702),
	.w4(32'hba04d729),
	.w5(32'h3b317b33),
	.w6(32'hbb57b625),
	.w7(32'hbb25d8a0),
	.w8(32'h3b884aca),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed779),
	.w1(32'hbabc4e0f),
	.w2(32'hbb023e16),
	.w3(32'hbb232d88),
	.w4(32'hba98104e),
	.w5(32'h3a5edac6),
	.w6(32'h3b8503c0),
	.w7(32'hbad8c744),
	.w8(32'hbaf5d74e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cfbff),
	.w1(32'hbaacadd9),
	.w2(32'h3bb71d6d),
	.w3(32'hb901e7f3),
	.w4(32'h3b5f52bd),
	.w5(32'h3b9a8d63),
	.w6(32'hbb26c9ad),
	.w7(32'h3ba23378),
	.w8(32'h3bf91ea9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f3f9c),
	.w1(32'hb8966fa8),
	.w2(32'h3b29bf0b),
	.w3(32'h3aae8212),
	.w4(32'hbb18ee53),
	.w5(32'h3a3fbd02),
	.w6(32'h3c09f665),
	.w7(32'h3b616a25),
	.w8(32'hbba6b4ff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aeb3f),
	.w1(32'hbae94220),
	.w2(32'hbb0e0948),
	.w3(32'h399c7277),
	.w4(32'hba74fe92),
	.w5(32'hbb1b44b5),
	.w6(32'hbb2b98f1),
	.w7(32'hb67a2869),
	.w8(32'hb922a988),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5999dd),
	.w1(32'h3c370139),
	.w2(32'hbb2f3421),
	.w3(32'hbb7d160e),
	.w4(32'h3a797a0b),
	.w5(32'h3b8c5974),
	.w6(32'hbab44328),
	.w7(32'hbbf98318),
	.w8(32'hbb84529d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b582010),
	.w1(32'h3b351918),
	.w2(32'h3b1e25b4),
	.w3(32'hbb1c9797),
	.w4(32'hbb6db20a),
	.w5(32'hbbc65e6a),
	.w6(32'h3a5700bb),
	.w7(32'hbbe11675),
	.w8(32'hbb5fbb5e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d389f),
	.w1(32'h3bade6da),
	.w2(32'h3b0edb60),
	.w3(32'hbad70a3d),
	.w4(32'hb96319a9),
	.w5(32'hbb82b587),
	.w6(32'h3a113298),
	.w7(32'h3a38b7e8),
	.w8(32'hb9e24f1e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48b642),
	.w1(32'hbb0dd16f),
	.w2(32'h38b781df),
	.w3(32'hb98a9c81),
	.w4(32'h3aa324d3),
	.w5(32'h3b34ecaa),
	.w6(32'h3ac8e848),
	.w7(32'h3b2d1041),
	.w8(32'h39be3471),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5402a4),
	.w1(32'h3b8e1f42),
	.w2(32'h3ae72203),
	.w3(32'h3abd84e8),
	.w4(32'hb992bbb1),
	.w5(32'h3b5a69c9),
	.w6(32'h3b502d08),
	.w7(32'h3aad1490),
	.w8(32'h3bf67e73),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170ac3),
	.w1(32'h3b68bfde),
	.w2(32'h3b43b652),
	.w3(32'h3a94ec74),
	.w4(32'h3a941802),
	.w5(32'hb8bc74c4),
	.w6(32'h3a09a8e4),
	.w7(32'hb9f08b57),
	.w8(32'hbaf2349f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becece5),
	.w1(32'h3b3ec77a),
	.w2(32'hb9b41251),
	.w3(32'h3b24e5c9),
	.w4(32'h39bd6ce9),
	.w5(32'hbaf5b371),
	.w6(32'hbb15cbd3),
	.w7(32'h3b5b9413),
	.w8(32'hba962e64),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf43872),
	.w1(32'hba0c8423),
	.w2(32'hbab2c1d7),
	.w3(32'hba51d0b2),
	.w4(32'hba942836),
	.w5(32'hba81e76c),
	.w6(32'h3aa7c429),
	.w7(32'hbb295d89),
	.w8(32'h3b0bae5a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb4b2),
	.w1(32'h39998bc6),
	.w2(32'h3966a2b7),
	.w3(32'hbb063274),
	.w4(32'hbaca79e3),
	.w5(32'hba7cc41a),
	.w6(32'hbbd5f251),
	.w7(32'hbbd6b1be),
	.w8(32'hbb1cf3a3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a95a0),
	.w1(32'h3aa7c08c),
	.w2(32'h3b3e039f),
	.w3(32'hba44a0cc),
	.w4(32'h3ae7d52b),
	.w5(32'h3b916d7f),
	.w6(32'hbb699ef1),
	.w7(32'h39d0d13a),
	.w8(32'h3b342f3b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ea37),
	.w1(32'hbbf43416),
	.w2(32'hbab537ae),
	.w3(32'hbb8dbcb3),
	.w4(32'hbb836a7a),
	.w5(32'h3a8e25ce),
	.w6(32'h3a4d1fc9),
	.w7(32'h37ef6c83),
	.w8(32'h3ab58c7c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb540f65),
	.w1(32'hbb2fd41e),
	.w2(32'h3bdd2f25),
	.w3(32'hbb06ecf9),
	.w4(32'hb9f9f78d),
	.w5(32'hbbb8d203),
	.w6(32'hbb40ca4e),
	.w7(32'h3c0c5ccd),
	.w8(32'hbb0b836c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a028780),
	.w1(32'hbb80c773),
	.w2(32'hbb90227f),
	.w3(32'hbc442ac3),
	.w4(32'hbb571acb),
	.w5(32'hbb30fa2c),
	.w6(32'hb946366b),
	.w7(32'hbb71a6ae),
	.w8(32'hbbfdf3c1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906a89),
	.w1(32'hbaf6568d),
	.w2(32'h3bfd10ec),
	.w3(32'hbbafc097),
	.w4(32'hbb5efa36),
	.w5(32'h3a14ff8d),
	.w6(32'hbaa585f4),
	.w7(32'h398d5268),
	.w8(32'h3b532050),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ac35e),
	.w1(32'hbbe8db00),
	.w2(32'hbbb244ae),
	.w3(32'hbb3f9ec7),
	.w4(32'hbbe11424),
	.w5(32'hb8c99d87),
	.w6(32'h392e1794),
	.w7(32'h3a1e4015),
	.w8(32'h3b0fd308),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2c898),
	.w1(32'hbba96108),
	.w2(32'h3bcc07c8),
	.w3(32'h3b30f8eb),
	.w4(32'hbb90f4a1),
	.w5(32'h39beb847),
	.w6(32'hba3033c9),
	.w7(32'hbb1a3d79),
	.w8(32'h3af781a4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5109a7),
	.w1(32'hba8919ef),
	.w2(32'h3b767818),
	.w3(32'h3a87ba19),
	.w4(32'h386ba258),
	.w5(32'hbaf2413e),
	.w6(32'h39f00e56),
	.w7(32'h3aa69823),
	.w8(32'h3b06e638),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbcf81),
	.w1(32'h3a7c714f),
	.w2(32'hbbf34d5c),
	.w3(32'h3bc2c874),
	.w4(32'hb9cdd092),
	.w5(32'hb9ee8565),
	.w6(32'h3c8fd146),
	.w7(32'hbbe82284),
	.w8(32'hba4f8471),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b525d17),
	.w1(32'hbc04bd63),
	.w2(32'h3b5f4972),
	.w3(32'hbbed462b),
	.w4(32'h3ad5bf0c),
	.w5(32'hbb13f27f),
	.w6(32'hbc2a1396),
	.w7(32'h394008ce),
	.w8(32'hbb8e69d0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff60a),
	.w1(32'hbb8104dc),
	.w2(32'h3b7b613e),
	.w3(32'hbb490f92),
	.w4(32'h3a5453e9),
	.w5(32'h3a6392b1),
	.w6(32'hbbf140a6),
	.w7(32'h3b596ad1),
	.w8(32'hbb98f9d1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72d51a),
	.w1(32'h397edd8e),
	.w2(32'h3b761e89),
	.w3(32'hbb7468cb),
	.w4(32'h3a912e85),
	.w5(32'h3c088770),
	.w6(32'hbb884958),
	.w7(32'hbaa1af4a),
	.w8(32'h3b5282e0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813cb88),
	.w1(32'hbab3d166),
	.w2(32'hbb058065),
	.w3(32'h3acca643),
	.w4(32'h3bb836c3),
	.w5(32'hbc472c16),
	.w6(32'h39a95ad9),
	.w7(32'h3ad6bf56),
	.w8(32'hbc7a9f43),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80b7c5c),
	.w1(32'h3c90d27e),
	.w2(32'h3b839b5d),
	.w3(32'h3b53f918),
	.w4(32'h3bff49a3),
	.w5(32'h3ae4059f),
	.w6(32'h3d0bd506),
	.w7(32'h3ba4a1c7),
	.w8(32'hbb6bc2e7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959293),
	.w1(32'h3b76a231),
	.w2(32'h3ba38e49),
	.w3(32'h3b86aa51),
	.w4(32'h3ac60f09),
	.w5(32'h3c28db42),
	.w6(32'h3b2bf37a),
	.w7(32'h38156c7d),
	.w8(32'h3c3701e4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0339f),
	.w1(32'h3b87721c),
	.w2(32'h3c151fa1),
	.w3(32'h3b8c9e16),
	.w4(32'hbbc0db91),
	.w5(32'h3b1d4014),
	.w6(32'h382ded26),
	.w7(32'hba83d59c),
	.w8(32'hbadf858e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2f594),
	.w1(32'h3bfb3380),
	.w2(32'h39f76994),
	.w3(32'hba7b13e9),
	.w4(32'hbb3ec9e0),
	.w5(32'hbc001bae),
	.w6(32'h3b88dd2e),
	.w7(32'hb6361852),
	.w8(32'hbc354d61),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba99395),
	.w1(32'h3bb0d992),
	.w2(32'hbb8d8abb),
	.w3(32'hbc1b0d87),
	.w4(32'h3c2bd9a6),
	.w5(32'hbb0ed553),
	.w6(32'h3ca48717),
	.w7(32'h3c56394f),
	.w8(32'hb8ae2fc2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a180b0c),
	.w1(32'hbab65608),
	.w2(32'hbb3dfd7c),
	.w3(32'h3a280bf5),
	.w4(32'hba76113c),
	.w5(32'hbada2073),
	.w6(32'hba3434f1),
	.w7(32'hbb0317b3),
	.w8(32'h3b32b9d7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2377bd),
	.w1(32'h3b05708a),
	.w2(32'h3b80bb04),
	.w3(32'hbb9a92b9),
	.w4(32'hbc307779),
	.w5(32'hb78ec2d9),
	.w6(32'hbb53e592),
	.w7(32'h39472b60),
	.w8(32'hbb778588),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc1ad5),
	.w1(32'hbb5469b6),
	.w2(32'h3bb78da1),
	.w3(32'hbb36a0a5),
	.w4(32'h3ac8a9ba),
	.w5(32'h3bcf1382),
	.w6(32'hbbce62ef),
	.w7(32'h3b1a18ad),
	.w8(32'h3ab25290),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02eca5),
	.w1(32'hbb97b3e7),
	.w2(32'hbaa23cea),
	.w3(32'hbb26405e),
	.w4(32'hbbb24931),
	.w5(32'hbc0fdc9a),
	.w6(32'hbb6c306c),
	.w7(32'h3a931589),
	.w8(32'hbc83af86),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53d267),
	.w1(32'h3c59b10e),
	.w2(32'h3bc5beda),
	.w3(32'h3a8a75c3),
	.w4(32'h3c4ae5a4),
	.w5(32'hbaeda6cb),
	.w6(32'h3ca0bae6),
	.w7(32'h3cc98555),
	.w8(32'hbaff9d95),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fade3),
	.w1(32'h3c06634f),
	.w2(32'hbb15ee23),
	.w3(32'h3bd82e47),
	.w4(32'h3a8edd29),
	.w5(32'h3b87c464),
	.w6(32'h3c86e2e8),
	.w7(32'h3a38d8dc),
	.w8(32'h3b6c4a86),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c67e16),
	.w1(32'hbb4dc619),
	.w2(32'h3906fdc5),
	.w3(32'h3b2aad2c),
	.w4(32'h3b9611e7),
	.w5(32'hbbad0728),
	.w6(32'hbb9c2765),
	.w7(32'hba7a2760),
	.w8(32'hbc0ed274),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab49da4),
	.w1(32'h3b534179),
	.w2(32'hb886782b),
	.w3(32'hbb0cd55f),
	.w4(32'hba65e678),
	.w5(32'h3aee93e1),
	.w6(32'h3a141f6e),
	.w7(32'hbb04cd35),
	.w8(32'h3a6d9acf),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfd858),
	.w1(32'h38dbbf60),
	.w2(32'hba9bfccb),
	.w3(32'h3acf4840),
	.w4(32'h3c1c674b),
	.w5(32'h3bf1195b),
	.w6(32'hbae2f731),
	.w7(32'h3b93c815),
	.w8(32'hbb014ef0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc347e0c),
	.w1(32'h3bfdfb3e),
	.w2(32'h3bc309e2),
	.w3(32'h3b619f56),
	.w4(32'hbc077aa5),
	.w5(32'hba761a11),
	.w6(32'h3b8ab31c),
	.w7(32'hbad411a4),
	.w8(32'hbb40dbb1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8479b3),
	.w1(32'hbb180a93),
	.w2(32'hb9a6c29c),
	.w3(32'hbafdf8ec),
	.w4(32'h3b95fd72),
	.w5(32'hbb03bb1d),
	.w6(32'hbbed162d),
	.w7(32'h3b058b6f),
	.w8(32'hbbd77913),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f686a),
	.w1(32'h3ba45251),
	.w2(32'hbbd64f15),
	.w3(32'h3b4d0ae2),
	.w4(32'hbbdc987f),
	.w5(32'h3c2d0ecb),
	.w6(32'h3bd3656b),
	.w7(32'hbb8f7dd5),
	.w8(32'h3bf52c82),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa88335),
	.w1(32'h3ae55c90),
	.w2(32'h3ac3cc08),
	.w3(32'h3b9674e5),
	.w4(32'h3ad4eab6),
	.w5(32'hbbd2de19),
	.w6(32'hb8696fb3),
	.w7(32'hbae4276f),
	.w8(32'hbad57e22),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d147e),
	.w1(32'h3a227260),
	.w2(32'h3bdfd082),
	.w3(32'hba3432b8),
	.w4(32'h398f2de4),
	.w5(32'hbb2c5412),
	.w6(32'h3ae3d6c2),
	.w7(32'h3b08e591),
	.w8(32'hbab5f1ba),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff07d0),
	.w1(32'h3c1d2ccc),
	.w2(32'hbaf1cdf7),
	.w3(32'hba3350a8),
	.w4(32'h3bcb6800),
	.w5(32'hb77d8013),
	.w6(32'h3c9fdcb2),
	.w7(32'h3c593569),
	.w8(32'hb9527a57),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96ad54),
	.w1(32'hbb20c5a0),
	.w2(32'hbb6e0632),
	.w3(32'hbb1c3ce2),
	.w4(32'hbadf6d43),
	.w5(32'h3b9b6dc5),
	.w6(32'hb9207d7e),
	.w7(32'h3a2db096),
	.w8(32'hbb7d9f28),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06c9cf),
	.w1(32'hbb082d6e),
	.w2(32'hbba9eb77),
	.w3(32'hbbd477ac),
	.w4(32'hbbc102b4),
	.w5(32'hbb0abd75),
	.w6(32'hbbe18230),
	.w7(32'hbb9cab8a),
	.w8(32'hbb977f34),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb242823),
	.w1(32'hbbe0ac3d),
	.w2(32'hba33ba92),
	.w3(32'hbbafdd81),
	.w4(32'hbaa23225),
	.w5(32'hb915d75a),
	.w6(32'hbbeaf56a),
	.w7(32'h38d02161),
	.w8(32'hbab6ebc3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb486ec5),
	.w1(32'h3b851291),
	.w2(32'h3b2e516d),
	.w3(32'h3adca398),
	.w4(32'h3b7d895c),
	.w5(32'hba7720b2),
	.w6(32'h3bc68cbf),
	.w7(32'h3b4c9cb0),
	.w8(32'h394f5952),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3865c),
	.w1(32'h3a8285a9),
	.w2(32'hba5d5652),
	.w3(32'hbab0ac73),
	.w4(32'hbb67e796),
	.w5(32'hbaab7c27),
	.w6(32'hba801252),
	.w7(32'hbb2dfc5b),
	.w8(32'hbbade538),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03a0a9),
	.w1(32'h3b8a887c),
	.w2(32'h3bbb1665),
	.w3(32'h3b487918),
	.w4(32'h3aff745e),
	.w5(32'hbb6313dc),
	.w6(32'h3a73e9fc),
	.w7(32'h3a59368e),
	.w8(32'hbba49f1c),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41fe44),
	.w1(32'hbba245b4),
	.w2(32'hba5cf9ac),
	.w3(32'hbbd9d915),
	.w4(32'hbaeebc91),
	.w5(32'h39743dd8),
	.w6(32'hbbc20f96),
	.w7(32'hb9a26fc6),
	.w8(32'hbaaa78ee),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8952a),
	.w1(32'hbbe2ebb5),
	.w2(32'hbb046db3),
	.w3(32'hbbbc4af3),
	.w4(32'hbb81f1bc),
	.w5(32'h3ad80017),
	.w6(32'hbb61aa04),
	.w7(32'hba97a8cb),
	.w8(32'h3bdc10cb),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1797b3),
	.w1(32'hb93c8ffc),
	.w2(32'hbb02b72c),
	.w3(32'hbb9fa0bd),
	.w4(32'hbbceac1c),
	.w5(32'h3b2f2a34),
	.w6(32'hbb28a6b3),
	.w7(32'hba476ce8),
	.w8(32'h3b2a32ac),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054f01),
	.w1(32'h3b533504),
	.w2(32'h3b37b1a2),
	.w3(32'h39816b86),
	.w4(32'h3a9c4e1b),
	.w5(32'hbaeab1f8),
	.w6(32'hbab31467),
	.w7(32'hbb1d5b1a),
	.w8(32'h3aeb5f98),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06ee86),
	.w1(32'h3bb49704),
	.w2(32'hbbb82f31),
	.w3(32'h3c179a25),
	.w4(32'hbc37c34d),
	.w5(32'h3b07af6e),
	.w6(32'h3cd47fd6),
	.w7(32'hbc4503cb),
	.w8(32'h38d611e4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3647fc6c),
	.w1(32'hb8f59393),
	.w2(32'hbb603ce5),
	.w3(32'hbac9c7df),
	.w4(32'h3acf81ec),
	.w5(32'h3bbc483b),
	.w6(32'hb97f892f),
	.w7(32'h3a2bdc8f),
	.w8(32'h3bf02d3d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f4ef),
	.w1(32'hbaf410cf),
	.w2(32'h3b20d974),
	.w3(32'hb4799422),
	.w4(32'h3b6c40c7),
	.w5(32'h3b799b42),
	.w6(32'hbaa92a30),
	.w7(32'h3b00ef69),
	.w8(32'hbadb3844),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94dde8),
	.w1(32'hb994cadf),
	.w2(32'h3bb55f48),
	.w3(32'h3b19bec2),
	.w4(32'h3b43c700),
	.w5(32'h3a9bc4fa),
	.w6(32'hbb9ef19c),
	.w7(32'h3a06ffcd),
	.w8(32'hb96296bb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28bef3),
	.w1(32'hbb0a4399),
	.w2(32'hbb015511),
	.w3(32'hba0cbd33),
	.w4(32'hbb84d9ca),
	.w5(32'h3ba86724),
	.w6(32'h3a3528fc),
	.w7(32'hbb22d6ec),
	.w8(32'h3b88b5f5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a0da0),
	.w1(32'hbc07dad2),
	.w2(32'hba779472),
	.w3(32'h3a746cd7),
	.w4(32'h3a12faf5),
	.w5(32'h3b0f3f45),
	.w6(32'hbb761aed),
	.w7(32'hbae98914),
	.w8(32'hbc059162),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63324f),
	.w1(32'h3c63f0c3),
	.w2(32'h3c907634),
	.w3(32'h3c5bc782),
	.w4(32'h3adc2ab5),
	.w5(32'hbbbc917f),
	.w6(32'h3c1b2e8b),
	.w7(32'h3c043f43),
	.w8(32'hbbc8dfc6),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6be77),
	.w1(32'h3af7525a),
	.w2(32'h3ba69be4),
	.w3(32'hba9adb54),
	.w4(32'h3ae96aa8),
	.w5(32'hb961946b),
	.w6(32'h3c0598e9),
	.w7(32'h3ad8d5b9),
	.w8(32'h38b57a99),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93744c1),
	.w1(32'hbae951e3),
	.w2(32'h39990f92),
	.w3(32'hba86aa2f),
	.w4(32'h3a9729f8),
	.w5(32'h3bf45669),
	.w6(32'hbb9ede15),
	.w7(32'h39e2fdb3),
	.w8(32'h3bcfac40),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97753c),
	.w1(32'hbba44b45),
	.w2(32'h3be929fc),
	.w3(32'hbbe0df52),
	.w4(32'hbb8f017d),
	.w5(32'hba097c78),
	.w6(32'hbb19736f),
	.w7(32'hbb7389cf),
	.w8(32'h3b0bd6f9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3015d2),
	.w1(32'h3b87e716),
	.w2(32'h3c1dc739),
	.w3(32'h3911ad1b),
	.w4(32'h3bf4039d),
	.w5(32'h3b9c4ac9),
	.w6(32'h3c0f83ec),
	.w7(32'h3c0a0750),
	.w8(32'h3b50d33b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b720083),
	.w1(32'hbb24b6fd),
	.w2(32'hbae17823),
	.w3(32'hbbed07bc),
	.w4(32'h3a9f9361),
	.w5(32'h3aa5184a),
	.w6(32'h3ba7a4ab),
	.w7(32'h3cbf17e5),
	.w8(32'hbbc90425),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb640414),
	.w1(32'hbbeb9800),
	.w2(32'hba3b1742),
	.w3(32'hbb0579cc),
	.w4(32'h3a6b87cb),
	.w5(32'h3b0cfec9),
	.w6(32'hbb7b38d7),
	.w7(32'h3ac13195),
	.w8(32'h3abfba30),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa3a0e),
	.w1(32'h3b79ec6b),
	.w2(32'h3c177fb2),
	.w3(32'h3b027546),
	.w4(32'h3c094043),
	.w5(32'h3b495c8a),
	.w6(32'h3b25ea7d),
	.w7(32'h3c4aba3f),
	.w8(32'hbb5205c5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7dc38),
	.w1(32'h3beebfa0),
	.w2(32'h3c06bfe8),
	.w3(32'h3b8c7651),
	.w4(32'h3bcbb949),
	.w5(32'hbb131841),
	.w6(32'h3af492ba),
	.w7(32'h3b13efd4),
	.w8(32'hbc0dd256),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19b799),
	.w1(32'hbb81f769),
	.w2(32'hbc47b7c2),
	.w3(32'hbbc4682d),
	.w4(32'hbc78c749),
	.w5(32'hbb304064),
	.w6(32'h38f70e8b),
	.w7(32'hbc5068df),
	.w8(32'hbba33ec0),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb76b524),
	.w1(32'h3c1d0105),
	.w2(32'h3890682a),
	.w3(32'h3c225d32),
	.w4(32'h3b0fc5b9),
	.w5(32'h3b0a1582),
	.w6(32'h3c8250c1),
	.w7(32'h3b982eb1),
	.w8(32'hba613565),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fb256),
	.w1(32'h3baaeab9),
	.w2(32'hbb048d3f),
	.w3(32'hbaae3c9b),
	.w4(32'hbb116039),
	.w5(32'h3a337c32),
	.w6(32'hbbb4c299),
	.w7(32'hbb189642),
	.w8(32'hbb36ba04),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c0aa8),
	.w1(32'hbbbac079),
	.w2(32'hbb7e1cb3),
	.w3(32'hbc0ddafd),
	.w4(32'hbbb384ca),
	.w5(32'hbc4b438b),
	.w6(32'hbb8f5afb),
	.w7(32'h3bcbf74a),
	.w8(32'hbc5237ff),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84e88a),
	.w1(32'hbb05521e),
	.w2(32'hbc0110c1),
	.w3(32'hbb37e0ab),
	.w4(32'hbb09afae),
	.w5(32'h3a131416),
	.w6(32'h3b8c66b4),
	.w7(32'hbb5ea7c4),
	.w8(32'h3b650b76),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8959b7),
	.w1(32'hbabe25d1),
	.w2(32'hbb114763),
	.w3(32'hbb5e0926),
	.w4(32'hbb8651ad),
	.w5(32'h3bb86037),
	.w6(32'hba5e9304),
	.w7(32'hbaa7b3ca),
	.w8(32'h3bf4447d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aff15),
	.w1(32'hbc1a250c),
	.w2(32'h3aa4ae88),
	.w3(32'hbc192ad0),
	.w4(32'hbaaa9990),
	.w5(32'hba923e11),
	.w6(32'hbc263d1f),
	.w7(32'h3c6e5ede),
	.w8(32'hbb982ee2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954c9f),
	.w1(32'hbb267164),
	.w2(32'hbacee977),
	.w3(32'hbba5514b),
	.w4(32'hba32a1d5),
	.w5(32'hbb84707e),
	.w6(32'h3b28a621),
	.w7(32'hbb08dcd9),
	.w8(32'h3b9254aa),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50ec2b),
	.w1(32'hbb79a605),
	.w2(32'h3b305eae),
	.w3(32'hbbccc2d2),
	.w4(32'hbbc72dca),
	.w5(32'hb9711c0d),
	.w6(32'hbbd10422),
	.w7(32'h3bbcd5ae),
	.w8(32'hbb33433a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eba37),
	.w1(32'hbae1ad83),
	.w2(32'h3bcb8758),
	.w3(32'h3aaacc30),
	.w4(32'h3b18ca3f),
	.w5(32'hbb279e04),
	.w6(32'hb9cf03d5),
	.w7(32'h3b9c7d4e),
	.w8(32'hbb49411c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5f8f2),
	.w1(32'h3b3c687a),
	.w2(32'h3ba36f36),
	.w3(32'hbb3ab50c),
	.w4(32'hb9e91cbb),
	.w5(32'hbb9a285c),
	.w6(32'hbc07754b),
	.w7(32'hbbb2d267),
	.w8(32'hbb06d7a9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf399e),
	.w1(32'hbaee3e77),
	.w2(32'hbb280215),
	.w3(32'h3b1a3c0e),
	.w4(32'hbb14dce6),
	.w5(32'hba73a64f),
	.w6(32'h3a5a0cb5),
	.w7(32'hba8d7e8b),
	.w8(32'h3bb0f14a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88717e),
	.w1(32'h3be41d0d),
	.w2(32'h3b53ad8f),
	.w3(32'hba845a25),
	.w4(32'hbacf6a6e),
	.w5(32'hbaa2947d),
	.w6(32'h3c691a90),
	.w7(32'h3bc629d1),
	.w8(32'hbb844c13),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00bb6),
	.w1(32'hbbdd22b6),
	.w2(32'hba5e203e),
	.w3(32'hbb47c429),
	.w4(32'h3af5da7a),
	.w5(32'h3bc1bf9a),
	.w6(32'hbbb0048d),
	.w7(32'h3b41c875),
	.w8(32'h3b55314e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866672),
	.w1(32'hbab8d14f),
	.w2(32'h3acc2af1),
	.w3(32'h3ba4f61a),
	.w4(32'h3bbba3d7),
	.w5(32'hb9bf810c),
	.w6(32'h3a376076),
	.w7(32'h3b9ad123),
	.w8(32'hbb1b804b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07d100),
	.w1(32'hbb93a8ed),
	.w2(32'h3b0fac55),
	.w3(32'hbb80adf8),
	.w4(32'h3bb3fbb4),
	.w5(32'hb894cc9e),
	.w6(32'hbbf09f7d),
	.w7(32'h3ab67037),
	.w8(32'hbad7972e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba403c38),
	.w1(32'hbb1f2005),
	.w2(32'hba1d1c4b),
	.w3(32'hbad6005b),
	.w4(32'h3a06ff4f),
	.w5(32'h3adc0d09),
	.w6(32'hbafc274c),
	.w7(32'h3bfedc67),
	.w8(32'h3b15922d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0b1ab),
	.w1(32'h3b72d7aa),
	.w2(32'h38e0cf5d),
	.w3(32'h3b217000),
	.w4(32'h3b9bda36),
	.w5(32'h3ace7065),
	.w6(32'hbb4e0086),
	.w7(32'h3a5858fd),
	.w8(32'h3b8549b1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25b6a5),
	.w1(32'hbafa5f58),
	.w2(32'h3976008d),
	.w3(32'hbb873909),
	.w4(32'h3a9a9eb8),
	.w5(32'hbbb2166d),
	.w6(32'hba8648c0),
	.w7(32'h3b976af7),
	.w8(32'hbbc27329),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e94fe),
	.w1(32'h3ac9bcb6),
	.w2(32'h3bc7ef4a),
	.w3(32'h3ae51aa9),
	.w4(32'h3b7cb540),
	.w5(32'hba2f4ff8),
	.w6(32'hb9b24370),
	.w7(32'h3a5848ab),
	.w8(32'hbb2eeef0),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd065f2),
	.w1(32'h3b7cf5a4),
	.w2(32'h3b605ace),
	.w3(32'hbb602e67),
	.w4(32'h3b2ba112),
	.w5(32'hbac2fecf),
	.w6(32'hbb2681f5),
	.w7(32'hba58687e),
	.w8(32'hbaddae58),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb894755),
	.w1(32'hbb81adc4),
	.w2(32'hba815881),
	.w3(32'h3aa7ee00),
	.w4(32'h3b02944d),
	.w5(32'h3a8d45a3),
	.w6(32'hbb40fe41),
	.w7(32'h3a2fcf1e),
	.w8(32'hbc5ac1c0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f897),
	.w1(32'h3c96ada9),
	.w2(32'h3b1d44f4),
	.w3(32'h3ba435a1),
	.w4(32'h3c29d2e7),
	.w5(32'h3b299080),
	.w6(32'h3ce1803c),
	.w7(32'h3c4f90fe),
	.w8(32'h3abb6faf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99729a1),
	.w1(32'h3b609168),
	.w2(32'h3be8feb5),
	.w3(32'h39a9dfc3),
	.w4(32'hbac85a33),
	.w5(32'hbc02fbbe),
	.w6(32'h3a1d9ca1),
	.w7(32'h3afb2f7f),
	.w8(32'hbc1e5627),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f7eb7),
	.w1(32'hbb1dc8a0),
	.w2(32'hbc6acd78),
	.w3(32'hbb45a842),
	.w4(32'hbc25552d),
	.w5(32'hb9584608),
	.w6(32'h3c5d7740),
	.w7(32'hbbdf5fa7),
	.w8(32'hb94930b9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28a462),
	.w1(32'h3b9fc9ab),
	.w2(32'hbaec1291),
	.w3(32'h3b89fa48),
	.w4(32'hb993cf44),
	.w5(32'h3a9976ec),
	.w6(32'h3bc69a85),
	.w7(32'hbb49d53e),
	.w8(32'hbbc124e7),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44814),
	.w1(32'h3a7d57ed),
	.w2(32'h3b930e5a),
	.w3(32'hb8b0d8d9),
	.w4(32'h3a632484),
	.w5(32'hbb16e83c),
	.w6(32'hbb6cb3bd),
	.w7(32'hba986cf9),
	.w8(32'hbb037a9c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ca4d0),
	.w1(32'hbbd20f0f),
	.w2(32'h3ab0ec14),
	.w3(32'hbbdf4fbf),
	.w4(32'h3aa4880d),
	.w5(32'h3c24bd66),
	.w6(32'hbc25ab4e),
	.w7(32'h3c106214),
	.w8(32'h3c8c3681),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c720b89),
	.w1(32'hb8c99b2a),
	.w2(32'h3c25bf81),
	.w3(32'h3b08f4a8),
	.w4(32'h3c3daa59),
	.w5(32'h3aec637a),
	.w6(32'h3986a661),
	.w7(32'h3c84a548),
	.w8(32'hbb1bebf9),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231a4e),
	.w1(32'h3c22f313),
	.w2(32'h3b25fc83),
	.w3(32'h3c325414),
	.w4(32'hbb66755e),
	.w5(32'hba1eff5d),
	.w6(32'h3ca78c3b),
	.w7(32'hbbe0463d),
	.w8(32'hbadac01f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa649),
	.w1(32'hbac3eb6b),
	.w2(32'h3908bd62),
	.w3(32'h3a98a132),
	.w4(32'h38b267c1),
	.w5(32'hbb8fb3b0),
	.w6(32'hb93f22f4),
	.w7(32'hb9f6c8a7),
	.w8(32'hbb3ad80c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93dbd3),
	.w1(32'hbc11cc0b),
	.w2(32'hb9199bb4),
	.w3(32'hbbb770d9),
	.w4(32'hbb2a44c0),
	.w5(32'hba921bf2),
	.w6(32'hbc900e59),
	.w7(32'h3b093350),
	.w8(32'hba24e601),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84942c),
	.w1(32'h3b310cb2),
	.w2(32'h3b067e3f),
	.w3(32'h3a9db3a1),
	.w4(32'h3b96c5d6),
	.w5(32'h3b8f3268),
	.w6(32'hba132ba9),
	.w7(32'h3a2612c4),
	.w8(32'hb992b705),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994ad54),
	.w1(32'hbb3f08ca),
	.w2(32'h3b0b62cb),
	.w3(32'hb98d4788),
	.w4(32'h3baa115e),
	.w5(32'hbb493d2c),
	.w6(32'hbbf03ded),
	.w7(32'h3aab8cc5),
	.w8(32'hbb8062b1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9f91),
	.w1(32'hbb96fd2b),
	.w2(32'hbafc6ae5),
	.w3(32'hbc3b193f),
	.w4(32'hbb337161),
	.w5(32'h3aa3c475),
	.w6(32'hbc0795e8),
	.w7(32'h3b653bac),
	.w8(32'h3afe5148),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b962336),
	.w1(32'hbbb3e3cc),
	.w2(32'hba5a6c75),
	.w3(32'hbbfca9c5),
	.w4(32'h3a0dcd53),
	.w5(32'h3b25c584),
	.w6(32'hbb152813),
	.w7(32'h3a0b23f9),
	.w8(32'h3b03906e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83acb1),
	.w1(32'h3bb8912d),
	.w2(32'h3af3f417),
	.w3(32'h3a6beb31),
	.w4(32'h3bbb0f87),
	.w5(32'hbbd40903),
	.w6(32'h3b8bce76),
	.w7(32'h3b95a6d4),
	.w8(32'hbb90cf99),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0247),
	.w1(32'hbb753888),
	.w2(32'hbb8d5930),
	.w3(32'hbb216bd5),
	.w4(32'h3b3972e8),
	.w5(32'hba9276d8),
	.w6(32'hbbd66e1d),
	.w7(32'hbb61e7bd),
	.w8(32'hbb2e0c9b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f0706),
	.w1(32'h3b188da4),
	.w2(32'hbb0d071e),
	.w3(32'hb9ae4a2b),
	.w4(32'h3b14be21),
	.w5(32'hbc5a0f01),
	.w6(32'h3b0fc892),
	.w7(32'h3a9c879d),
	.w8(32'hbc996393),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0baeb),
	.w1(32'hbb3ca811),
	.w2(32'h3b867c01),
	.w3(32'hbbe85106),
	.w4(32'hbab68c36),
	.w5(32'hba5ee88a),
	.w6(32'hbaf4649e),
	.w7(32'hbbbc4152),
	.w8(32'hbc218989),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4a161),
	.w1(32'h3a9aa0f9),
	.w2(32'hba8cd15d),
	.w3(32'h3b76cd6f),
	.w4(32'h3b3aa6b2),
	.w5(32'h3bcafa5f),
	.w6(32'h3c496ce4),
	.w7(32'h3b1b3134),
	.w8(32'h3bd57227),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fdbfe),
	.w1(32'hbae15621),
	.w2(32'hb9a3c2cf),
	.w3(32'h3b44c526),
	.w4(32'h3bb493cb),
	.w5(32'h3b02c37e),
	.w6(32'hbc12d6e7),
	.w7(32'hba717911),
	.w8(32'h3b357658),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba727261),
	.w1(32'hbb2cc985),
	.w2(32'h3b2e8662),
	.w3(32'h39dfe1ee),
	.w4(32'h3aa445fb),
	.w5(32'h3b3147fa),
	.w6(32'hbb80ec8c),
	.w7(32'h3b828281),
	.w8(32'hbaa1e6f9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b2e3),
	.w1(32'h3c03cb70),
	.w2(32'hb9d06942),
	.w3(32'hb8834bd0),
	.w4(32'hbb1c3d33),
	.w5(32'h3b00dd50),
	.w6(32'h3b6f55c9),
	.w7(32'hbbbe21e9),
	.w8(32'h3ae9e754),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33edbe),
	.w1(32'hbb47de2d),
	.w2(32'h3a469779),
	.w3(32'hbb83375b),
	.w4(32'hbb762ded),
	.w5(32'hbaf4bb37),
	.w6(32'hbb8a7f04),
	.w7(32'hbb6f9948),
	.w8(32'hbae0439e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9796e),
	.w1(32'hbb3751d2),
	.w2(32'h3a907703),
	.w3(32'hbafbd040),
	.w4(32'hbb9a2ffe),
	.w5(32'h3b7f7443),
	.w6(32'hbb5ecc82),
	.w7(32'h3b595477),
	.w8(32'h3ad0e886),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80a4dd),
	.w1(32'hbb7cab44),
	.w2(32'hbb840221),
	.w3(32'hbabcfd5e),
	.w4(32'hbbbaddf7),
	.w5(32'hbaa157e9),
	.w6(32'hbb0e8bd7),
	.w7(32'hbbcef219),
	.w8(32'hba1a294b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb918c),
	.w1(32'h3a95af49),
	.w2(32'h3b17956e),
	.w3(32'hbb1ed2ec),
	.w4(32'hbb439a99),
	.w5(32'hbb4ab798),
	.w6(32'h3a329004),
	.w7(32'hbac7358c),
	.w8(32'hbab6b692),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01e5ee),
	.w1(32'hbb0adc14),
	.w2(32'h3c1e365b),
	.w3(32'hbbbb2806),
	.w4(32'hbb8f3fd5),
	.w5(32'h3c01a7ea),
	.w6(32'hbbaee2d4),
	.w7(32'h3aec606c),
	.w8(32'h3bec6eb6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a895785),
	.w1(32'hbab2969f),
	.w2(32'h3a9db728),
	.w3(32'h3b358500),
	.w4(32'hbb1560ef),
	.w5(32'h3b6680af),
	.w6(32'hba6e6531),
	.w7(32'hbb1197d1),
	.w8(32'h3b1f1548),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e3a95),
	.w1(32'hbb406531),
	.w2(32'hbb121568),
	.w3(32'hbb3dae20),
	.w4(32'h3a1e3cfb),
	.w5(32'h3b8f7306),
	.w6(32'hbb0a2a8b),
	.w7(32'h3a6224c2),
	.w8(32'hbad0fefc),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81cd1f),
	.w1(32'h3b9638df),
	.w2(32'h3bb472ce),
	.w3(32'h3aba3bd4),
	.w4(32'h3ba5a6f9),
	.w5(32'hbbd43918),
	.w6(32'hbb191034),
	.w7(32'h3872e7f6),
	.w8(32'hbb8d19ee),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7bce3),
	.w1(32'hbb88ffc6),
	.w2(32'h3b00618a),
	.w3(32'h39cc77fd),
	.w4(32'h3b5ff1e5),
	.w5(32'h3baf2200),
	.w6(32'h3b83de3a),
	.w7(32'h3c0bc280),
	.w8(32'h3b89a8ea),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abeff96),
	.w1(32'hbb465f37),
	.w2(32'hba8a7333),
	.w3(32'h3b2a784b),
	.w4(32'h3a1b23ec),
	.w5(32'h3afc49a6),
	.w6(32'hba92acb9),
	.w7(32'h3a7a7db6),
	.w8(32'h3ad3933d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6d259),
	.w1(32'h3b2f5eaa),
	.w2(32'h3b9d0a49),
	.w3(32'h3b8ff655),
	.w4(32'h3ab29a88),
	.w5(32'hbc10f2ba),
	.w6(32'h3c7a3ed8),
	.w7(32'h3b85e6d6),
	.w8(32'hbbbea46e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc35280),
	.w1(32'h3b9fb326),
	.w2(32'h3bdb4bd0),
	.w3(32'h3a91f6c2),
	.w4(32'h3bbc69df),
	.w5(32'h3ba2f8b8),
	.w6(32'h3c5029d8),
	.w7(32'h3c7116b5),
	.w8(32'h3b8d15bb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1bae6),
	.w1(32'hbb59cf4d),
	.w2(32'h3a342279),
	.w3(32'hba78cda6),
	.w4(32'h3774dbb2),
	.w5(32'h3a7fde07),
	.w6(32'h3b9289b2),
	.w7(32'h3adc381a),
	.w8(32'hbadb443d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db6f4),
	.w1(32'hbae63f5b),
	.w2(32'h3b79af34),
	.w3(32'hbb34e6b4),
	.w4(32'h3b6b0810),
	.w5(32'h3a909198),
	.w6(32'hbb1fbf2d),
	.w7(32'h3b7655ac),
	.w8(32'h3a861aa0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3e219),
	.w1(32'h3c13dda9),
	.w2(32'h3b1592ee),
	.w3(32'h3b0f7800),
	.w4(32'h3c5a57f8),
	.w5(32'hbbae8b9d),
	.w6(32'h3c48362e),
	.w7(32'h3be5a2fa),
	.w8(32'hbb8d8191),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc136e67),
	.w1(32'hbb4c9fc2),
	.w2(32'h3b506aff),
	.w3(32'hbbc5c40a),
	.w4(32'hbbbaf128),
	.w5(32'h3af5c167),
	.w6(32'hbba63fb9),
	.w7(32'h39a4db30),
	.w8(32'hb9828767),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15328d),
	.w1(32'h3a95ae45),
	.w2(32'h3b1dad54),
	.w3(32'h3ba05779),
	.w4(32'h3ba58e01),
	.w5(32'h38d251e2),
	.w6(32'h3a864a94),
	.w7(32'h3af4eeef),
	.w8(32'hbb6e3b55),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd9fff),
	.w1(32'h3b49efc7),
	.w2(32'h3a0c5cc0),
	.w3(32'hba391092),
	.w4(32'hbad97ba5),
	.w5(32'hbbdc46bc),
	.w6(32'h3c9bfae0),
	.w7(32'h39793d6e),
	.w8(32'hbb571ed9),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb756171),
	.w1(32'h3ae8d871),
	.w2(32'h3b516a67),
	.w3(32'hbb6572dd),
	.w4(32'h3ba4b312),
	.w5(32'hbac6b147),
	.w6(32'h3a9d0450),
	.w7(32'h3b62122f),
	.w8(32'hbb9703bb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7893),
	.w1(32'hbb0aa636),
	.w2(32'hbb112323),
	.w3(32'h3a4868b8),
	.w4(32'h3af2690f),
	.w5(32'h3bbb7f73),
	.w6(32'h3c3a59d1),
	.w7(32'h3b487047),
	.w8(32'h3a051371),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac638b),
	.w1(32'hbbcf67a8),
	.w2(32'hbb9f6360),
	.w3(32'hbb520d78),
	.w4(32'hb9a10257),
	.w5(32'hbb6e1767),
	.w6(32'hbb8a2ce3),
	.w7(32'hba788cf5),
	.w8(32'hbc04c909),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69ca69),
	.w1(32'h3a8acad1),
	.w2(32'hbb22fdb3),
	.w3(32'h3ba7fcfe),
	.w4(32'hbab4d5eb),
	.w5(32'hbb438489),
	.w6(32'h3c0ab603),
	.w7(32'hbabc96f4),
	.w8(32'hbbb34aa0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb631589),
	.w1(32'hba80273c),
	.w2(32'h3b0ea86d),
	.w3(32'hbab12088),
	.w4(32'h3a3dc451),
	.w5(32'h3b81ff7a),
	.w6(32'h3ab68725),
	.w7(32'h3b059883),
	.w8(32'h3acfbd61),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91675d),
	.w1(32'hbc092b93),
	.w2(32'hbb5c3add),
	.w3(32'hbb2c1559),
	.w4(32'h3b7f77f4),
	.w5(32'hbb93d965),
	.w6(32'hbb85ecb0),
	.w7(32'h399119cd),
	.w8(32'h3891ecd9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47397f),
	.w1(32'hbb940c34),
	.w2(32'hbaf94740),
	.w3(32'hbbce41bc),
	.w4(32'hbb168b57),
	.w5(32'hb930c054),
	.w6(32'hbbe47edd),
	.w7(32'h3b700fa6),
	.w8(32'hbb810586),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc08d54),
	.w1(32'hba3c20f2),
	.w2(32'hb8c78571),
	.w3(32'hba812cd6),
	.w4(32'hbaef14fc),
	.w5(32'hbaa4caa2),
	.w6(32'h3b813fe3),
	.w7(32'h3bb339f4),
	.w8(32'hba9ef36d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6dd6c),
	.w1(32'hbb15a81f),
	.w2(32'hb9da7285),
	.w3(32'hbb23784a),
	.w4(32'h3b199333),
	.w5(32'hbb03a1c1),
	.w6(32'hbb659b76),
	.w7(32'h3b112935),
	.w8(32'h3ad2f28e),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9925705),
	.w1(32'h3c4ca7c5),
	.w2(32'h3bfacd59),
	.w3(32'hbbe54c3d),
	.w4(32'hb871b1e1),
	.w5(32'h3a9be36b),
	.w6(32'h3c08c634),
	.w7(32'h3c0717b1),
	.w8(32'h3a049540),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6e62e),
	.w1(32'hba2d49b1),
	.w2(32'hb80d69af),
	.w3(32'hba6bf101),
	.w4(32'h3b15ac02),
	.w5(32'hbb937ef5),
	.w6(32'hbb66e290),
	.w7(32'hba83b152),
	.w8(32'hbb9cd35f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa65e26),
	.w1(32'hbaa1af88),
	.w2(32'h3b8a998f),
	.w3(32'hbb982496),
	.w4(32'hbba0db58),
	.w5(32'h3947274b),
	.w6(32'hbb99c998),
	.w7(32'hbbba1110),
	.w8(32'hbb14bced),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9c2f7),
	.w1(32'h3bc67f00),
	.w2(32'h3ac439bb),
	.w3(32'hbb420296),
	.w4(32'h398e1acd),
	.w5(32'h3b81e5ef),
	.w6(32'h3bc0234e),
	.w7(32'h3be110bb),
	.w8(32'h3c0690e6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7a88f),
	.w1(32'h3bc3b34e),
	.w2(32'h3c1f4be6),
	.w3(32'hbad24be3),
	.w4(32'h3c45542a),
	.w5(32'hbbf5e9b5),
	.w6(32'h3b628335),
	.w7(32'h3c04d81b),
	.w8(32'hbbbf96a7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb531e36),
	.w1(32'hbc068941),
	.w2(32'hbbd2b4d9),
	.w3(32'hbbafda45),
	.w4(32'hbbccbdcd),
	.w5(32'h39ab0ed3),
	.w6(32'hbba7b1a3),
	.w7(32'hbc019cfd),
	.w8(32'h3bb12df5),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3166bd),
	.w1(32'h3bafef73),
	.w2(32'h39cb54d2),
	.w3(32'hbb302fa9),
	.w4(32'h3ac62bb2),
	.w5(32'hbacb416e),
	.w6(32'h3b1398fb),
	.w7(32'h3b003bc9),
	.w8(32'hbb072096),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6be5c4),
	.w1(32'h3c8a92d6),
	.w2(32'h3bcf8c00),
	.w3(32'hbbc113ea),
	.w4(32'h3a84ad21),
	.w5(32'h3b6a29ae),
	.w6(32'h3bc41dd3),
	.w7(32'h38908f7f),
	.w8(32'hba38082a),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9b4dd),
	.w1(32'h3aaf24f0),
	.w2(32'h3a709c43),
	.w3(32'hbafad8ff),
	.w4(32'hba842c7b),
	.w5(32'hbbd75936),
	.w6(32'hba8b58c4),
	.w7(32'h3ba0b860),
	.w8(32'hbbfa1913),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cac13),
	.w1(32'hbbc8f599),
	.w2(32'hbbde0329),
	.w3(32'hbbf14ecf),
	.w4(32'hbae81674),
	.w5(32'hbab4f5a7),
	.w6(32'hbc28136a),
	.w7(32'hbbc8352e),
	.w8(32'hbabf6324),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df65c),
	.w1(32'hbb2b184d),
	.w2(32'hbbd47835),
	.w3(32'h39f112fb),
	.w4(32'hbbab1b9d),
	.w5(32'h386f7db8),
	.w6(32'h3b0615a0),
	.w7(32'hbb4719b6),
	.w8(32'hbbe72dac),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db3323),
	.w1(32'hba60f630),
	.w2(32'h3bad5f44),
	.w3(32'hbbb7ccc8),
	.w4(32'h3950b18e),
	.w5(32'hba08676c),
	.w6(32'hbb763ab9),
	.w7(32'hb9f101c4),
	.w8(32'hbb16974f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab86b24),
	.w1(32'h3bb1a16f),
	.w2(32'h3ba6cdb2),
	.w3(32'hbb0f5232),
	.w4(32'hb8dfdd9e),
	.w5(32'hbbe233c5),
	.w6(32'h3b9c649c),
	.w7(32'h3bdb2c52),
	.w8(32'hbbeb9b0a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cb60),
	.w1(32'hb9d2e702),
	.w2(32'hbbd02cb2),
	.w3(32'hbaa22082),
	.w4(32'hbb18eeec),
	.w5(32'hb9c5ba5e),
	.w6(32'h3afc0302),
	.w7(32'hbb5fae65),
	.w8(32'h3b1862b1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdf1c2),
	.w1(32'h3babe800),
	.w2(32'h3a6e5486),
	.w3(32'hbb34b409),
	.w4(32'hbba1f5c6),
	.w5(32'h3a13559c),
	.w6(32'hbb2dc206),
	.w7(32'hbaabaf8b),
	.w8(32'h3bbdca97),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4d040),
	.w1(32'h3b4ca517),
	.w2(32'hb7ad22cb),
	.w3(32'h3b5e3784),
	.w4(32'h3b11e2df),
	.w5(32'hbbb1a3bc),
	.w6(32'h3b88731a),
	.w7(32'h3b98e477),
	.w8(32'hbc02a04c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba85333),
	.w1(32'h3a96fb53),
	.w2(32'h3bd9bd61),
	.w3(32'hbbd8e966),
	.w4(32'hbb44c206),
	.w5(32'hbb01093a),
	.w6(32'h39c9ff14),
	.w7(32'hb800246c),
	.w8(32'hbb00b7a6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e3e45),
	.w1(32'hbade5ece),
	.w2(32'h3a2463f8),
	.w3(32'hbb21ae10),
	.w4(32'h386cea99),
	.w5(32'h3806753c),
	.w6(32'hbb9a9df0),
	.w7(32'h3a58b876),
	.w8(32'h3b4e7716),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94bc73),
	.w1(32'h38ffc302),
	.w2(32'h3b6c02fc),
	.w3(32'h3bed76f9),
	.w4(32'hbac116fb),
	.w5(32'h3bbb5c2a),
	.w6(32'hbbf9910c),
	.w7(32'h3b0268fb),
	.w8(32'h3bac7813),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee1e39),
	.w1(32'h3bbb1339),
	.w2(32'hba33ad9b),
	.w3(32'h3b2e4157),
	.w4(32'hbaa4bad2),
	.w5(32'hbc3f2d41),
	.w6(32'hbb279552),
	.w7(32'h3b7418e9),
	.w8(32'hbc19f517),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f91ff),
	.w1(32'hbba5040f),
	.w2(32'hbb8f9f8f),
	.w3(32'hbc89b986),
	.w4(32'hba3f02e4),
	.w5(32'hb90ae78a),
	.w6(32'hbc2c284a),
	.w7(32'hbbd710ca),
	.w8(32'h3a9fc1f1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454f72),
	.w1(32'hbb794918),
	.w2(32'h3b5a1971),
	.w3(32'hbbc46398),
	.w4(32'hbc0d46d9),
	.w5(32'hbaec5b25),
	.w6(32'hbbc51926),
	.w7(32'hba5f738c),
	.w8(32'hbb88d0a5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836599),
	.w1(32'hbb3411dc),
	.w2(32'h3a9a84f0),
	.w3(32'h3be340ca),
	.w4(32'h3bf16174),
	.w5(32'hbc5c0ba2),
	.w6(32'h3b927b8b),
	.w7(32'h3be4899a),
	.w8(32'hbb23032a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba16a63),
	.w1(32'h3a8e6829),
	.w2(32'hbb821a6e),
	.w3(32'h3a8758fa),
	.w4(32'h3c29e7a7),
	.w5(32'h3c2fd78b),
	.w6(32'h3b72258e),
	.w7(32'h3b3a42eb),
	.w8(32'hba5f3995),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0383a7),
	.w1(32'h3bad3c26),
	.w2(32'h3b2d114a),
	.w3(32'h3c05ef73),
	.w4(32'hbb9a6a81),
	.w5(32'hbb56664b),
	.w6(32'h3c9e8bb0),
	.w7(32'hbc2130ed),
	.w8(32'hbc606e9d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9dd22),
	.w1(32'hbaca16ec),
	.w2(32'hbbc58f74),
	.w3(32'hbad9b892),
	.w4(32'hbb26b17c),
	.w5(32'hbb13bdfd),
	.w6(32'hbafa2b71),
	.w7(32'h3a724e8f),
	.w8(32'hbaa683a9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd18469),
	.w1(32'hbba625fb),
	.w2(32'hbb993cd5),
	.w3(32'hbb2823f5),
	.w4(32'h3b177eba),
	.w5(32'h3bac32e2),
	.w6(32'hba464429),
	.w7(32'h3a48e86a),
	.w8(32'h3aceae7e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01a14d),
	.w1(32'h3abb0f93),
	.w2(32'h3b29995c),
	.w3(32'h3a9d13f2),
	.w4(32'h39c78f4d),
	.w5(32'h3b0d2947),
	.w6(32'h3a10a873),
	.w7(32'h3a99903e),
	.w8(32'h3b821eea),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be314bf),
	.w1(32'h3b095498),
	.w2(32'h3b1078ec),
	.w3(32'h3b20f080),
	.w4(32'h38cff445),
	.w5(32'hbc169428),
	.w6(32'hba93d004),
	.w7(32'h3aff8937),
	.w8(32'hbbe31828),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule