module layer_8_featuremap_130(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc188717),
	.w1(32'hbc5c2e76),
	.w2(32'hbbd0e544),
	.w3(32'hbc174d45),
	.w4(32'hbc18e7a4),
	.w5(32'h3b8b3c75),
	.w6(32'h3c55c453),
	.w7(32'hbc128769),
	.w8(32'h3c933099),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69adfb),
	.w1(32'hbc1c9e17),
	.w2(32'h3b45801c),
	.w3(32'hb8bb08b2),
	.w4(32'h3c8348f3),
	.w5(32'h3c053ba9),
	.w6(32'h3b5b2c1f),
	.w7(32'hbbd26af4),
	.w8(32'hbb09e329),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983c14b),
	.w1(32'h3c3d1f4e),
	.w2(32'hbb1e31a8),
	.w3(32'h3c15631a),
	.w4(32'hbb1f38d6),
	.w5(32'hbbc2df4b),
	.w6(32'h3b86083f),
	.w7(32'hbc057759),
	.w8(32'hbbc28686),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bebb8),
	.w1(32'hbbc6f2be),
	.w2(32'hbcd79af6),
	.w3(32'hbbaa6edd),
	.w4(32'h3a992d17),
	.w5(32'h3a50a395),
	.w6(32'h3c209d2b),
	.w7(32'h3d086bd4),
	.w8(32'h3d126d18),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd089096),
	.w1(32'hbcbc6f3f),
	.w2(32'hbbf45e63),
	.w3(32'hbbb8f5a5),
	.w4(32'h3b6d1d63),
	.w5(32'h3b801d4c),
	.w6(32'h3c3558e4),
	.w7(32'hbbf15b3f),
	.w8(32'hbc728d6e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd2615),
	.w1(32'hbc9b8fbf),
	.w2(32'h3a89d89a),
	.w3(32'hbbcd58fe),
	.w4(32'h3bf7c1a8),
	.w5(32'h3c49ee0b),
	.w6(32'hbbeaeda6),
	.w7(32'hbc9ca838),
	.w8(32'hbc331375),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc764ed4),
	.w1(32'hbc051c8e),
	.w2(32'h3ab6ccd5),
	.w3(32'h3bb6bd11),
	.w4(32'h3c903bfd),
	.w5(32'h3b0dd058),
	.w6(32'h3c265b9f),
	.w7(32'h3a185b7c),
	.w8(32'hbc48bde2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fdd59),
	.w1(32'hbac6dd1b),
	.w2(32'hbbaf09f6),
	.w3(32'h390acec2),
	.w4(32'hbba261b5),
	.w5(32'hbb2e2ebc),
	.w6(32'h3ba786bd),
	.w7(32'hbb463ae1),
	.w8(32'h3ae2ea83),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33d647),
	.w1(32'hbbd48cbf),
	.w2(32'hbc134357),
	.w3(32'hbc737ac9),
	.w4(32'hbc1b58c2),
	.w5(32'hbc029bfa),
	.w6(32'h3ae117d0),
	.w7(32'h3b325bdb),
	.w8(32'h3ccde8ee),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0452e7),
	.w1(32'hbc08f63a),
	.w2(32'h3bb197a0),
	.w3(32'hbc8b2f83),
	.w4(32'hba4b5c1c),
	.w5(32'hba92967a),
	.w6(32'h3b2f90d3),
	.w7(32'hbba88a8c),
	.w8(32'h3c9866ce),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f5ff7),
	.w1(32'hbcc38d4e),
	.w2(32'hbc529795),
	.w3(32'hbc367d2f),
	.w4(32'hbc455f7c),
	.w5(32'h3ac0e90b),
	.w6(32'h3c133634),
	.w7(32'hbc17391f),
	.w8(32'hbc8a0c9d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3347a),
	.w1(32'h3ca1e5b4),
	.w2(32'hbc47e12d),
	.w3(32'hbb923bec),
	.w4(32'hbc076db8),
	.w5(32'hbc0e3920),
	.w6(32'hb968526a),
	.w7(32'hbc00663b),
	.w8(32'hbb9a0e39),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4d846),
	.w1(32'hbbf9fdfc),
	.w2(32'hb98de643),
	.w3(32'hbbc6319f),
	.w4(32'hbb4a149f),
	.w5(32'h3bd744ef),
	.w6(32'h3c6769a1),
	.w7(32'hb7d6cd5c),
	.w8(32'h3b30b640),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a3801),
	.w1(32'h3a82e38e),
	.w2(32'h3a22d7f6),
	.w3(32'h3be5a487),
	.w4(32'hbb7185fe),
	.w5(32'h3ac6d642),
	.w6(32'h3b3c0922),
	.w7(32'h3a345448),
	.w8(32'h3b98eaf2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817dc96),
	.w1(32'hbaf9a158),
	.w2(32'hba09d7ae),
	.w3(32'h3b7e73f2),
	.w4(32'hbb3086a9),
	.w5(32'h3b1edeec),
	.w6(32'h3b94dd4a),
	.w7(32'hbb0f7025),
	.w8(32'h3b94cb10),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74f5f2),
	.w1(32'hbb83dce4),
	.w2(32'h3a94d4cc),
	.w3(32'h3b1ca2b9),
	.w4(32'h3a897fa0),
	.w5(32'hb9e53f75),
	.w6(32'h3b0a0050),
	.w7(32'h3bf80a76),
	.w8(32'h3cc3beea),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eec9f),
	.w1(32'hbcbe47c6),
	.w2(32'hbc040236),
	.w3(32'hbc748640),
	.w4(32'hbb484e1b),
	.w5(32'hbc34a5ca),
	.w6(32'h3c4d18f6),
	.w7(32'hbc4bbe8b),
	.w8(32'hbc9d6cc3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb206c4),
	.w1(32'h3a92baa6),
	.w2(32'h3aedccae),
	.w3(32'hbc2080a5),
	.w4(32'h3b1b3d48),
	.w5(32'h3b2ddd2a),
	.w6(32'hbc185623),
	.w7(32'hbb29cd25),
	.w8(32'hbc3301f3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e810),
	.w1(32'hbb4deef4),
	.w2(32'hbc0ab933),
	.w3(32'h3b9f3c7c),
	.w4(32'hbba023a8),
	.w5(32'h3b3f7748),
	.w6(32'hbc8206de),
	.w7(32'h3c05db07),
	.w8(32'hbb27bfca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd51a9),
	.w1(32'hbc09b5f1),
	.w2(32'hbcac484b),
	.w3(32'hbbbf715f),
	.w4(32'hbc418948),
	.w5(32'hbcb2909c),
	.w6(32'hbbcc32ac),
	.w7(32'hbbf54d5f),
	.w8(32'hbca44ce5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bd3dc),
	.w1(32'hbc97b859),
	.w2(32'hbaa0d6d3),
	.w3(32'hbb79cc29),
	.w4(32'h3a251252),
	.w5(32'hbb8ce719),
	.w6(32'hbcb35841),
	.w7(32'hbc8cb014),
	.w8(32'hbc2301a1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01dc47),
	.w1(32'h3c5ba4ee),
	.w2(32'hbc8ff67e),
	.w3(32'hbb1de6ee),
	.w4(32'h3a612d65),
	.w5(32'h3b7c2808),
	.w6(32'hbc369db4),
	.w7(32'h3bb39884),
	.w8(32'hbbcf1168),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfae083),
	.w1(32'hbb8a49b8),
	.w2(32'hbac33801),
	.w3(32'hba22377e),
	.w4(32'hbcabce8b),
	.w5(32'hbbc47492),
	.w6(32'h3a8aee70),
	.w7(32'hbc0a2d68),
	.w8(32'h3cb23c9b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d3f73),
	.w1(32'hbc0567f5),
	.w2(32'h3b80b79f),
	.w3(32'hbc7a748d),
	.w4(32'hb9319c9b),
	.w5(32'hbaf979d6),
	.w6(32'h3be2fb2a),
	.w7(32'hbbbe3104),
	.w8(32'hbbdb3fdc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bcdf3),
	.w1(32'hbae0e2a4),
	.w2(32'h3b82323e),
	.w3(32'h3b832f97),
	.w4(32'hbaab4cbf),
	.w5(32'hba4f1ee8),
	.w6(32'h3bb65278),
	.w7(32'hba9549cf),
	.w8(32'h3b650a2f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69bf4d),
	.w1(32'h3a88ff26),
	.w2(32'hbcba47d9),
	.w3(32'hba43f3a9),
	.w4(32'h3c36b635),
	.w5(32'h3ca96d57),
	.w6(32'h3b245b47),
	.w7(32'h3c85d2fa),
	.w8(32'h3d35208f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf8ee21),
	.w1(32'hbcb7f60d),
	.w2(32'hbc5f34ef),
	.w3(32'h3b160fef),
	.w4(32'h3c2b2e3e),
	.w5(32'hbc25fc8c),
	.w6(32'h3ce176f8),
	.w7(32'h3b0cfe65),
	.w8(32'h3ab376a5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c012cf3),
	.w1(32'h3b28cf9e),
	.w2(32'hbcb5f52e),
	.w3(32'h3d210192),
	.w4(32'hbd2af8a6),
	.w5(32'hbd14a4a4),
	.w6(32'hbcc4ad61),
	.w7(32'h3c95fabe),
	.w8(32'h3d9021f8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bb7e3),
	.w1(32'hbc30593d),
	.w2(32'h3c3efbec),
	.w3(32'hbccecc3e),
	.w4(32'h3bd183c4),
	.w5(32'hbc46c883),
	.w6(32'h3cdca160),
	.w7(32'hbc1fec39),
	.w8(32'hbc9f8db6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68e213),
	.w1(32'h3c1c266d),
	.w2(32'h3cd0e332),
	.w3(32'hbaf2607c),
	.w4(32'h3c333efa),
	.w5(32'h3d0f52b2),
	.w6(32'h3c1eccdf),
	.w7(32'hbd6ad694),
	.w8(32'hbdb3039f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3108aa),
	.w1(32'h3c9630cf),
	.w2(32'h3a49828b),
	.w3(32'h3d095bcf),
	.w4(32'h3805ae43),
	.w5(32'h3bdf4443),
	.w6(32'hbd29c1e8),
	.w7(32'hbad7c6fd),
	.w8(32'h3bb31d00),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f86b0),
	.w1(32'h3b0e8623),
	.w2(32'hbc800370),
	.w3(32'h3bb6ab5f),
	.w4(32'hbcca35c2),
	.w5(32'hbcce48de),
	.w6(32'h3b1f2689),
	.w7(32'h3bb02da6),
	.w8(32'h3bb104a1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0689),
	.w1(32'hbc993e01),
	.w2(32'h3c9135ff),
	.w3(32'hbcb301ad),
	.w4(32'h3c543f71),
	.w5(32'h3cc8382d),
	.w6(32'hbc69ff8f),
	.w7(32'hbcc32ff4),
	.w8(32'hbd395422),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81973a),
	.w1(32'h3c9c1b8b),
	.w2(32'hbc028495),
	.w3(32'h3c895545),
	.w4(32'h3b5d2479),
	.w5(32'h3bd1d1ec),
	.w6(32'hbd003d73),
	.w7(32'h3a803dcb),
	.w8(32'h3c4c4d25),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27cfd2),
	.w1(32'h3c4922c2),
	.w2(32'h3bc6035b),
	.w3(32'h3b4710d8),
	.w4(32'hb95eb56d),
	.w5(32'h3b2194e0),
	.w6(32'h3a8676ef),
	.w7(32'h39a6e35b),
	.w8(32'hbb021960),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa59ec),
	.w1(32'hbbc9c514),
	.w2(32'h3c42fcac),
	.w3(32'hba8f3c6f),
	.w4(32'h3b4d4c5a),
	.w5(32'h3bd5211c),
	.w6(32'hbc258ce9),
	.w7(32'hbc9344a3),
	.w8(32'hbbd23dd1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc105d7f),
	.w1(32'hbc184795),
	.w2(32'hbc252173),
	.w3(32'h3c92d20e),
	.w4(32'hbc8b69fd),
	.w5(32'hbc1a1bfa),
	.w6(32'h3c2cd3a0),
	.w7(32'h3c6764f6),
	.w8(32'h3ce57488),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11efba),
	.w1(32'hbc5a0c4e),
	.w2(32'hbc61a215),
	.w3(32'hbc237ec2),
	.w4(32'hbc00aebe),
	.w5(32'h3a3199f6),
	.w6(32'hb90020e0),
	.w7(32'hbac4bf8e),
	.w8(32'hbb01f174),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb2d37),
	.w1(32'hbbb8c9cb),
	.w2(32'hbba5af39),
	.w3(32'hbc0af15b),
	.w4(32'hbbb2f1de),
	.w5(32'hbc902882),
	.w6(32'hbacad1fa),
	.w7(32'h3bf717cf),
	.w8(32'hbc29812f),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f4e66),
	.w1(32'hbb671efd),
	.w2(32'h3b23734c),
	.w3(32'hbc91007f),
	.w4(32'h3b541ff8),
	.w5(32'hbb31889d),
	.w6(32'hbab93757),
	.w7(32'hba3c365e),
	.w8(32'h3a9da1b6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71939a),
	.w1(32'h3b6ac872),
	.w2(32'hbc2bfecb),
	.w3(32'h3b91ac35),
	.w4(32'hbbd5ef96),
	.w5(32'hbc942bb5),
	.w6(32'h3bcb6203),
	.w7(32'h3c633a9d),
	.w8(32'hbb893e92),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa08ce6),
	.w1(32'hbc2bd2d4),
	.w2(32'hbcdc642d),
	.w3(32'hbc069ec4),
	.w4(32'h3bb06f6c),
	.w5(32'h3c541d3d),
	.w6(32'hbba72f1b),
	.w7(32'hbc039733),
	.w8(32'h3d79884e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97e123),
	.w1(32'hbc723f9a),
	.w2(32'h3d0da11c),
	.w3(32'hbc8af308),
	.w4(32'h3bc2d570),
	.w5(32'hbb9a3c38),
	.w6(32'h3ca6eea8),
	.w7(32'hbcd5c9b9),
	.w8(32'hbd5daae4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e08af),
	.w1(32'h3c99377e),
	.w2(32'hbb4a767a),
	.w3(32'hbc02e6ae),
	.w4(32'hbba77707),
	.w5(32'h3bd8f2dd),
	.w6(32'hbccc69c5),
	.w7(32'hbb03152f),
	.w8(32'h3b8e9b1f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55c1d5),
	.w1(32'hbb9b0f57),
	.w2(32'h3c862dab),
	.w3(32'h3bd81ca8),
	.w4(32'h3acfa458),
	.w5(32'hbc3b06d6),
	.w6(32'h3ac56f99),
	.w7(32'hbbef5d01),
	.w8(32'hbc821785),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27b364),
	.w1(32'h3c6ad0dd),
	.w2(32'h3c0ed492),
	.w3(32'hbbef95ce),
	.w4(32'hbb2e65a9),
	.w5(32'h3c3745e4),
	.w6(32'h3bdfb4ba),
	.w7(32'hbcaad731),
	.w8(32'h3bb1d725),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9940bf),
	.w1(32'hbbb18eac),
	.w2(32'hba90a4ca),
	.w3(32'h3bb5b511),
	.w4(32'h3cadcad6),
	.w5(32'h3c598f1d),
	.w6(32'h3bfd3c01),
	.w7(32'hbbd4d87f),
	.w8(32'hbcf9e5d2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc340312),
	.w1(32'hb9c68236),
	.w2(32'hbbb31f6b),
	.w3(32'h3b0184db),
	.w4(32'h3c27f1a6),
	.w5(32'h3bfacf51),
	.w6(32'hbd095097),
	.w7(32'hba30446e),
	.w8(32'hbc8e083b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ef59c),
	.w1(32'h3bc1abf1),
	.w2(32'hbcf79a70),
	.w3(32'h3bc195e5),
	.w4(32'h3987658b),
	.w5(32'h392beed2),
	.w6(32'hbb89d280),
	.w7(32'hbba6efa5),
	.w8(32'h3c4f5f38),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd180fec),
	.w1(32'hbca4577a),
	.w2(32'hbc754d1c),
	.w3(32'h39a16373),
	.w4(32'hbc51816a),
	.w5(32'hbc690878),
	.w6(32'h3bed78d1),
	.w7(32'hbbfc4bdd),
	.w8(32'hbc154509),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f71fde),
	.w1(32'hbc0e4677),
	.w2(32'hbbd56e04),
	.w3(32'hbc3df85e),
	.w4(32'h3c24f6c0),
	.w5(32'h3c8bf5be),
	.w6(32'hbc1e8ba4),
	.w7(32'h3c492349),
	.w8(32'h3bb41439),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84e8d1),
	.w1(32'hbc9e48d9),
	.w2(32'hbba73c44),
	.w3(32'hbae2d96d),
	.w4(32'hbc220586),
	.w5(32'hba5861ee),
	.w6(32'h3c0bd731),
	.w7(32'h3c5c7de7),
	.w8(32'h3bbd6e3d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fbb9e),
	.w1(32'h3c557492),
	.w2(32'hbbac39b8),
	.w3(32'hbc38f275),
	.w4(32'hbc462f74),
	.w5(32'hbca7005a),
	.w6(32'hbc020f07),
	.w7(32'h3c40495b),
	.w8(32'hbc573381),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6ffd7),
	.w1(32'h3bcd442f),
	.w2(32'h3b34c18c),
	.w3(32'hb9ab36d9),
	.w4(32'hba9c5916),
	.w5(32'h3c16cd8e),
	.w6(32'hbc1724ce),
	.w7(32'hbb651a7b),
	.w8(32'h3b0e89db),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20b582),
	.w1(32'hb9a6fbe6),
	.w2(32'h3ca58ad5),
	.w3(32'h3bdb5053),
	.w4(32'hbb4b1adb),
	.w5(32'h3bf50d5a),
	.w6(32'h3b64c342),
	.w7(32'h3af6e593),
	.w8(32'h3cd1c360),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c803bcb),
	.w1(32'h3c4913f2),
	.w2(32'hbb3d43e3),
	.w3(32'h3c382d3d),
	.w4(32'hbb312865),
	.w5(32'hbae3d827),
	.w6(32'hbb9d0153),
	.w7(32'hbadbfa20),
	.w8(32'hbaa09fe8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aabc3),
	.w1(32'hbb447d84),
	.w2(32'hbc007e66),
	.w3(32'h3b77bc62),
	.w4(32'h3b25af51),
	.w5(32'h3b3e68f4),
	.w6(32'h3c0054b3),
	.w7(32'h3a08564d),
	.w8(32'h3c287d24),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4bed3),
	.w1(32'hbb624db1),
	.w2(32'h3c8a2ce0),
	.w3(32'h3c078aa5),
	.w4(32'h3b9631d2),
	.w5(32'hb9ab9e73),
	.w6(32'h3c03d8ce),
	.w7(32'hbc105c5a),
	.w8(32'hbce77cf4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d7d97),
	.w1(32'hbbf05fa4),
	.w2(32'h3a1e2026),
	.w3(32'hbbf2bfde),
	.w4(32'hbad648bf),
	.w5(32'h3c05af8d),
	.w6(32'hbc4715b9),
	.w7(32'hbab54dde),
	.w8(32'h3c0136e6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07f4ba),
	.w1(32'h3a7942cf),
	.w2(32'hbc297445),
	.w3(32'h3c0b8a32),
	.w4(32'hbc90df31),
	.w5(32'hbc982372),
	.w6(32'h3bdc0b26),
	.w7(32'h3ced0cf4),
	.w8(32'h3d83aeda),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbd428),
	.w1(32'hbbdb1750),
	.w2(32'h3c7c1ff9),
	.w3(32'hbca7260c),
	.w4(32'hbc16b72f),
	.w5(32'hbcb9d6db),
	.w6(32'h3c841789),
	.w7(32'hba8df6d5),
	.w8(32'h3c5f03fa),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac0aa8),
	.w1(32'h3c810285),
	.w2(32'hb9caf94e),
	.w3(32'hbc016c45),
	.w4(32'hbc061890),
	.w5(32'hbc100581),
	.w6(32'h3c37d131),
	.w7(32'hbb33bb75),
	.w8(32'hbb294245),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9faa29),
	.w1(32'h3a048ed6),
	.w2(32'h3bcc831c),
	.w3(32'hbae25c31),
	.w4(32'h3c403c9c),
	.w5(32'h3c50b1a4),
	.w6(32'h3b0e053d),
	.w7(32'h3c446cda),
	.w8(32'hbc636fad),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b735153),
	.w1(32'hbb452ac2),
	.w2(32'hbb9b9116),
	.w3(32'h3b723683),
	.w4(32'h3a1d6630),
	.w5(32'h3b307014),
	.w6(32'hbc3d5819),
	.w7(32'h3a7dfc9f),
	.w8(32'hbc56d7bf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ac2c4),
	.w1(32'hbb35a9d8),
	.w2(32'h3bb3276e),
	.w3(32'h3babd913),
	.w4(32'h3b265d11),
	.w5(32'h3bb2547b),
	.w6(32'hbbd918a5),
	.w7(32'hbc9284fb),
	.w8(32'h3c0976de),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26cc18),
	.w1(32'h3bf56355),
	.w2(32'h3c570287),
	.w3(32'hbba1709e),
	.w4(32'h3ba60050),
	.w5(32'h3c43768f),
	.w6(32'hbc0e8277),
	.w7(32'hbc471aa9),
	.w8(32'hbc50a726),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ca693),
	.w1(32'h3c465a03),
	.w2(32'hbbe531c4),
	.w3(32'h3c9b1426),
	.w4(32'h38349bb8),
	.w5(32'h3a308bbb),
	.w6(32'h3b4e5e24),
	.w7(32'hbc11c135),
	.w8(32'hbbf60216),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8890d2),
	.w1(32'h3b0b45a2),
	.w2(32'hbacf73a1),
	.w3(32'hbb764215),
	.w4(32'h3bbed045),
	.w5(32'h3c23ca79),
	.w6(32'h3bd352a1),
	.w7(32'hb99d3ba6),
	.w8(32'h3cb0fd3a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd14b5a),
	.w1(32'h3bb0d742),
	.w2(32'h3bbde0b2),
	.w3(32'h3c463a90),
	.w4(32'hba1f2491),
	.w5(32'h3a628d29),
	.w6(32'h3a0b0281),
	.w7(32'h3c71fe6b),
	.w8(32'h3d2509b0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1b8ca4),
	.w1(32'h3c139333),
	.w2(32'h3c0df086),
	.w3(32'hba33ae7f),
	.w4(32'h3c91fad3),
	.w5(32'h3c8115f5),
	.w6(32'h3b1761f2),
	.w7(32'hbc1d0f3c),
	.w8(32'hbcc07690),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8618a),
	.w1(32'h3c7780b3),
	.w2(32'hb9414566),
	.w3(32'h3ca05776),
	.w4(32'h3b9785b3),
	.w5(32'h3b87c36a),
	.w6(32'hbcd8b913),
	.w7(32'hbbef0db5),
	.w8(32'hbb960c46),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8e722),
	.w1(32'h3c740e42),
	.w2(32'hbbf0cc50),
	.w3(32'h3c6a2f04),
	.w4(32'hba4795a7),
	.w5(32'hbbb96137),
	.w6(32'hbc715231),
	.w7(32'hbb3d1e3e),
	.w8(32'hbb7123ec),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae9d5b),
	.w1(32'hbc0d2918),
	.w2(32'hbc1c5448),
	.w3(32'hbac8cb49),
	.w4(32'hbc253f0b),
	.w5(32'h3b7dfee7),
	.w6(32'hbabaeea5),
	.w7(32'hbbd8dc90),
	.w8(32'hbb7eb9b9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40695),
	.w1(32'hbc05dc56),
	.w2(32'hbb805aa0),
	.w3(32'h3be355db),
	.w4(32'hbc0909c2),
	.w5(32'h3b9facec),
	.w6(32'hbc5753c0),
	.w7(32'h3c824c5c),
	.w8(32'h3c3dc2ed),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c153e),
	.w1(32'hbb2e5e83),
	.w2(32'hbc925cc1),
	.w3(32'h3c320bc5),
	.w4(32'hba7eaef2),
	.w5(32'h3a1385ce),
	.w6(32'hbbfbede6),
	.w7(32'hbc1dd5d3),
	.w8(32'hbc9679bd),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce747b0),
	.w1(32'hbcde11c6),
	.w2(32'hba2f09a4),
	.w3(32'h398ac08f),
	.w4(32'hba19dbaf),
	.w5(32'h3bc31402),
	.w6(32'hbc47d7c9),
	.w7(32'hbbb664bc),
	.w8(32'hbb5dfe93),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a958b),
	.w1(32'h3bb9d7fb),
	.w2(32'h38e3b10e),
	.w3(32'h3c8fbe6f),
	.w4(32'h3a0e2d41),
	.w5(32'hbafa21d6),
	.w6(32'hbbc697d2),
	.w7(32'hba41f681),
	.w8(32'h3a6a0be9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b640b2a),
	.w1(32'hbad34007),
	.w2(32'hbb40c0a9),
	.w3(32'h39a01f83),
	.w4(32'hbbf5fa66),
	.w5(32'h3985ee8c),
	.w6(32'hba5a11f6),
	.w7(32'hbad07e33),
	.w8(32'h3b6aef5a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ccf0c),
	.w1(32'h3afa4466),
	.w2(32'h3b4fa4f8),
	.w3(32'h396871fe),
	.w4(32'hbae41bb7),
	.w5(32'h3bae1ba2),
	.w6(32'hbb568c4a),
	.w7(32'hbb2d59de),
	.w8(32'h3afbaa2d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab41bf1),
	.w1(32'hbae0667e),
	.w2(32'h3b43a3f4),
	.w3(32'hba5d3bf2),
	.w4(32'hbb8d25fd),
	.w5(32'h393572ee),
	.w6(32'hba6d356c),
	.w7(32'h3ac5d7cd),
	.w8(32'h3babcaab),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6116c1),
	.w1(32'h3b336f1f),
	.w2(32'h3b0b3ca0),
	.w3(32'h3b6e74ba),
	.w4(32'h3ac83127),
	.w5(32'h3c82a80e),
	.w6(32'h3be7e4b0),
	.w7(32'h3b69129d),
	.w8(32'h3c4965e6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4abfcf),
	.w1(32'h3b0cd8be),
	.w2(32'hbb841fc5),
	.w3(32'h3b83a847),
	.w4(32'hba2b7eec),
	.w5(32'hbba6ca32),
	.w6(32'h3a1a66d0),
	.w7(32'hbc061286),
	.w8(32'hbbacbb64),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe49ba4),
	.w1(32'hbb524ae5),
	.w2(32'hbb7b3326),
	.w3(32'hbb875fb6),
	.w4(32'hbafef9b9),
	.w5(32'hbb0a6758),
	.w6(32'hbba33a77),
	.w7(32'h3908c321),
	.w8(32'hbb6f4301),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba09768),
	.w1(32'h3b3810b5),
	.w2(32'h3b86bef8),
	.w3(32'h3bff4f31),
	.w4(32'h3c3f9d37),
	.w5(32'h3ca3e959),
	.w6(32'h3c8e63e2),
	.w7(32'h3c1be1cc),
	.w8(32'h3bc1f391),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba020285),
	.w1(32'hbc07b601),
	.w2(32'h3b89de9c),
	.w3(32'h3bc60bdd),
	.w4(32'hba02179f),
	.w5(32'h3be00dcd),
	.w6(32'hbb037790),
	.w7(32'h3c072ea1),
	.w8(32'h3c055baf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6903c),
	.w1(32'hbb2af007),
	.w2(32'h3b74a0b2),
	.w3(32'h3a264595),
	.w4(32'h3a6d3441),
	.w5(32'h3ab3cc65),
	.w6(32'h3b7520ce),
	.w7(32'h3b40aafb),
	.w8(32'hba14e58f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce72cf),
	.w1(32'hbbab64e2),
	.w2(32'h3b5a5808),
	.w3(32'hbbd0d4a6),
	.w4(32'hba3d27a7),
	.w5(32'hbb844b88),
	.w6(32'hbb843c88),
	.w7(32'h3bae0cab),
	.w8(32'h3be5fc7c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5a971),
	.w1(32'h3bb1fae0),
	.w2(32'hbbbac6ad),
	.w3(32'hbb0790fb),
	.w4(32'hbba9a74c),
	.w5(32'h3a63e82d),
	.w6(32'h3bbb6fd7),
	.w7(32'hbbb346bb),
	.w8(32'h3af376a5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27b79a),
	.w1(32'h3b4bd41d),
	.w2(32'hbac38010),
	.w3(32'h3b059ad1),
	.w4(32'h3b79c4be),
	.w5(32'hbc07454c),
	.w6(32'h3b515f1f),
	.w7(32'hbb4638eb),
	.w8(32'hbc246897),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5faf7),
	.w1(32'hba92248c),
	.w2(32'h3bc35349),
	.w3(32'hbb70d394),
	.w4(32'h3bdb62f8),
	.w5(32'h3bbbfa19),
	.w6(32'hbbbdfda4),
	.w7(32'h3c1b9b5c),
	.w8(32'hbab849b6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0af2),
	.w1(32'hbc40057c),
	.w2(32'h3be372bb),
	.w3(32'hbbd54b77),
	.w4(32'h3a7234ee),
	.w5(32'h3b45de42),
	.w6(32'hbc05e1d5),
	.w7(32'h3c34dce8),
	.w8(32'h3b52b124),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e19ca),
	.w1(32'h3a8e1975),
	.w2(32'h3ba8ff1c),
	.w3(32'h3b87b6c1),
	.w4(32'hbb26ac5f),
	.w5(32'hbb6b8837),
	.w6(32'h3c182fa8),
	.w7(32'h3c40c2f8),
	.w8(32'hb8851b23),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dd6a9),
	.w1(32'hbb6ddbd1),
	.w2(32'h3b5e0a7a),
	.w3(32'hbb0ea840),
	.w4(32'h3c0e1770),
	.w5(32'h3c171ff8),
	.w6(32'h3b572c08),
	.w7(32'h3bca3e4d),
	.w8(32'h3bb8fb6a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dea18),
	.w1(32'h3ab4cda5),
	.w2(32'h3c0e27d3),
	.w3(32'h3ba626cd),
	.w4(32'h3aeeac28),
	.w5(32'h3b6b4c04),
	.w6(32'h3b778774),
	.w7(32'h3bae52b1),
	.w8(32'h3c680125),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2873e7),
	.w1(32'h3c7f3148),
	.w2(32'h3b2b9846),
	.w3(32'h3bd729e6),
	.w4(32'h3b8a41b0),
	.w5(32'h3beb2e5b),
	.w6(32'h3c176fea),
	.w7(32'h3b8a3ec6),
	.w8(32'h3be872a1),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2a1a),
	.w1(32'h3abdaf51),
	.w2(32'h3b67a112),
	.w3(32'h3b386eef),
	.w4(32'hbc08985f),
	.w5(32'hbb4804f7),
	.w6(32'h3b1ab1d3),
	.w7(32'hbbf1094d),
	.w8(32'h3b0c2211),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd13715),
	.w1(32'hbaa5e4a1),
	.w2(32'h398cbeb9),
	.w3(32'hbba1cf7f),
	.w4(32'h3ae68de5),
	.w5(32'h3c0f0291),
	.w6(32'h3a835e4c),
	.w7(32'hbb452240),
	.w8(32'h3bc8d6ee),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc043e),
	.w1(32'hbbbd9c46),
	.w2(32'h3aedbd4e),
	.w3(32'h3bcc86d5),
	.w4(32'h3b9b8df7),
	.w5(32'h3c4be847),
	.w6(32'hba86bdb6),
	.w7(32'hb90189b9),
	.w8(32'h3beed2d5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c124c1e),
	.w1(32'h3b914b62),
	.w2(32'h3b8a7841),
	.w3(32'h3bcd1470),
	.w4(32'h3bc3cab8),
	.w5(32'hbabb913e),
	.w6(32'h3b0d7f1f),
	.w7(32'h3b59b371),
	.w8(32'hbb54b6ad),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c9c39c),
	.w1(32'h3b65f73a),
	.w2(32'h3be6d36d),
	.w3(32'hba73444a),
	.w4(32'h3bfdc695),
	.w5(32'h3b4b0c5f),
	.w6(32'h395ddc65),
	.w7(32'h3af07158),
	.w8(32'h3b90aca0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5439a3),
	.w1(32'h3a62c0a8),
	.w2(32'hbbda915c),
	.w3(32'hbb22d0be),
	.w4(32'hbaaabbd4),
	.w5(32'h3afe4704),
	.w6(32'hbbbd32ff),
	.w7(32'hbc0c8b0c),
	.w8(32'hbb3331ca),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e897e),
	.w1(32'hbbd1d4ca),
	.w2(32'h3b01bbbe),
	.w3(32'h3ace0fc4),
	.w4(32'h3a9ae588),
	.w5(32'hbb934ba8),
	.w6(32'hbaf531fc),
	.w7(32'h3b34fc98),
	.w8(32'hbb29f747),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0aab1),
	.w1(32'hbb749928),
	.w2(32'hbb52f94c),
	.w3(32'h3a96ce13),
	.w4(32'h392ceb92),
	.w5(32'hbbc64f62),
	.w6(32'h3ac6a252),
	.w7(32'hbb4e11c5),
	.w8(32'hbbf77843),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5e7f),
	.w1(32'h3a47fbe9),
	.w2(32'h3be4ec25),
	.w3(32'hbb5caa02),
	.w4(32'hb8d877b1),
	.w5(32'hba96b0c0),
	.w6(32'hbbc683e2),
	.w7(32'h3c74e6cc),
	.w8(32'h3c60fb4c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef143e),
	.w1(32'h3b3bdd12),
	.w2(32'hbacd1dad),
	.w3(32'hbac0e74e),
	.w4(32'hba6b3c55),
	.w5(32'hbb3c1de4),
	.w6(32'h3c32ff0b),
	.w7(32'hbb7a10c3),
	.w8(32'h3ba90ffe),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8ec24),
	.w1(32'hbab8ebf0),
	.w2(32'h3bed8bd0),
	.w3(32'h3bf4d8a0),
	.w4(32'h3b032da9),
	.w5(32'hb9866af3),
	.w6(32'h3bf0b213),
	.w7(32'h3c8e73a0),
	.w8(32'h3b77e280),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28452c),
	.w1(32'h3acc0c95),
	.w2(32'hba331fe9),
	.w3(32'hbb58cf88),
	.w4(32'h3bceaa08),
	.w5(32'hbb82a879),
	.w6(32'h3b8fc4b7),
	.w7(32'h3c34cf3e),
	.w8(32'hbb988a9d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aac835),
	.w1(32'h3c0b8f33),
	.w2(32'h3a8e7273),
	.w3(32'h3b2f2cc8),
	.w4(32'h3a38d964),
	.w5(32'hbb34c223),
	.w6(32'h3b1195d1),
	.w7(32'h3994d6da),
	.w8(32'h3ab05ee3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d7707),
	.w1(32'h3babb2fb),
	.w2(32'h3afc7779),
	.w3(32'hb8e8198f),
	.w4(32'hbb23bcfe),
	.w5(32'h3a937c96),
	.w6(32'h3b94daed),
	.w7(32'hba86af52),
	.w8(32'hbb82087a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7453b),
	.w1(32'h3aac9bca),
	.w2(32'h3c3023a4),
	.w3(32'h3939ea8c),
	.w4(32'h3c115afb),
	.w5(32'hbbc6145a),
	.w6(32'hbb17ba3f),
	.w7(32'h3c1dc652),
	.w8(32'hbbb5f459),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf2cf7),
	.w1(32'h3c8952cc),
	.w2(32'hbb0bbcf8),
	.w3(32'hbb82ba4b),
	.w4(32'h3bdfb61e),
	.w5(32'h3bdfb0bd),
	.w6(32'h3c0ab808),
	.w7(32'h3be48dde),
	.w8(32'h3a8d369a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ceb0c),
	.w1(32'hbacb0f70),
	.w2(32'h3aa727aa),
	.w3(32'h3b81552c),
	.w4(32'h3a751fb9),
	.w5(32'h3b8e8552),
	.w6(32'h3b8b1418),
	.w7(32'h3ae1fb66),
	.w8(32'h3b952c2d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b47ad),
	.w1(32'h3a81bf26),
	.w2(32'hb977d841),
	.w3(32'hbbe9d605),
	.w4(32'h3ac0d554),
	.w5(32'hbbeccfd0),
	.w6(32'hba42b619),
	.w7(32'h3b6916ce),
	.w8(32'hbc10f44b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6c10c),
	.w1(32'h3b973982),
	.w2(32'hbbb30410),
	.w3(32'hbb37a5a6),
	.w4(32'hbb57f473),
	.w5(32'hba8ab2f7),
	.w6(32'h3ab91331),
	.w7(32'hbb30e1ab),
	.w8(32'h3a9b24e0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa818e8),
	.w1(32'h3ac39fce),
	.w2(32'h3c186209),
	.w3(32'hba9a4dde),
	.w4(32'hba87990d),
	.w5(32'hbac3578c),
	.w6(32'h3b94d933),
	.w7(32'h3b012182),
	.w8(32'h3bbb2777),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c5e6),
	.w1(32'h3bec6253),
	.w2(32'h3c1157db),
	.w3(32'h3ba627eb),
	.w4(32'h3c40d8fc),
	.w5(32'h3c754d81),
	.w6(32'h3c164c1d),
	.w7(32'h3c2ee4e7),
	.w8(32'h3bd37962),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0801b),
	.w1(32'h3b77e489),
	.w2(32'hbabce233),
	.w3(32'h3b8e9f60),
	.w4(32'hbc398e87),
	.w5(32'hba396ee4),
	.w6(32'hb9d12460),
	.w7(32'hbbfbba7f),
	.w8(32'h3b6af127),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd423),
	.w1(32'hbb850adf),
	.w2(32'h39a507f2),
	.w3(32'h3c2fafc9),
	.w4(32'hbac8cf18),
	.w5(32'hba739457),
	.w6(32'h3a13b3b7),
	.w7(32'h3aa810ee),
	.w8(32'h3b62a6b8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8efb99),
	.w1(32'h3b944ec9),
	.w2(32'h3b92ce15),
	.w3(32'h3958c467),
	.w4(32'hb9d9bcb7),
	.w5(32'hbab3c833),
	.w6(32'h3b5e9734),
	.w7(32'h3af6f8ef),
	.w8(32'hbb1a53e6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393263d6),
	.w1(32'h3b79df6d),
	.w2(32'h39b59232),
	.w3(32'h3ae5b35a),
	.w4(32'hba9abca5),
	.w5(32'hbb9b0ba0),
	.w6(32'h3baf3bb5),
	.w7(32'hbaa63bba),
	.w8(32'hbba04630),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d7931),
	.w1(32'h3b038032),
	.w2(32'h3caf6e44),
	.w3(32'hbb23a79a),
	.w4(32'h3b3018f3),
	.w5(32'h3c85bc6a),
	.w6(32'hbace9681),
	.w7(32'h3c8bdbbe),
	.w8(32'h3d05013d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c4714),
	.w1(32'h3b3a39ec),
	.w2(32'h3b8f51e6),
	.w3(32'h3c71026f),
	.w4(32'h3b5da08a),
	.w5(32'h3a84ef24),
	.w6(32'h3c96b6f7),
	.w7(32'h3bc4c838),
	.w8(32'h3a1caa0d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6857c3),
	.w1(32'h3940f0ea),
	.w2(32'h3ad129bd),
	.w3(32'h3bb4fa9a),
	.w4(32'h3a429a03),
	.w5(32'hbadaa77a),
	.w6(32'h3b6daf69),
	.w7(32'h389183b0),
	.w8(32'h3aa7e37c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f0eb3),
	.w1(32'h3b80e580),
	.w2(32'h39d6c6b2),
	.w3(32'hb94d8084),
	.w4(32'h3b537605),
	.w5(32'hba226f28),
	.w6(32'h3b6ca244),
	.w7(32'h3afe0808),
	.w8(32'hbbba8ac7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb640064),
	.w1(32'hbb03278a),
	.w2(32'h3bd44f23),
	.w3(32'hbaaa397d),
	.w4(32'h3b90e891),
	.w5(32'hba54ff2a),
	.w6(32'hbba9806c),
	.w7(32'h3c0f1652),
	.w8(32'h3962b21a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad845ba),
	.w1(32'hbac07047),
	.w2(32'hbb677030),
	.w3(32'h3b869650),
	.w4(32'hba8166dc),
	.w5(32'h3b991759),
	.w6(32'h3b6cb861),
	.w7(32'hbba340a5),
	.w8(32'hba8c7c03),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba083143),
	.w1(32'hbb8a0be5),
	.w2(32'hbb2246ec),
	.w3(32'h3a11e579),
	.w4(32'hbb6dcf9a),
	.w5(32'hbaf271bc),
	.w6(32'hbb514704),
	.w7(32'hbbc8ba7b),
	.w8(32'h3af7b7d6),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2603),
	.w1(32'hbb400d4b),
	.w2(32'hb8faefb7),
	.w3(32'h3b822c3d),
	.w4(32'hbb6a290f),
	.w5(32'hbac653c2),
	.w6(32'hbb16f635),
	.w7(32'hbb5db7e8),
	.w8(32'h3a91df79),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule