module layer_8_featuremap_24(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb21faa),
	.w1(32'h3bddc100),
	.w2(32'h3b92cb57),
	.w3(32'h3bb85cf9),
	.w4(32'h3c08f3db),
	.w5(32'h3bff5114),
	.w6(32'h3baa2045),
	.w7(32'h3bd4f58f),
	.w8(32'h3ba85e34),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955c11),
	.w1(32'hbbb71810),
	.w2(32'hbbd53e19),
	.w3(32'hbb49cf50),
	.w4(32'hbb90cf50),
	.w5(32'hbbaa440b),
	.w6(32'hba45eacf),
	.w7(32'hbb130097),
	.w8(32'hbb80608d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09bf12),
	.w1(32'hbb86cead),
	.w2(32'hbbaaeeaf),
	.w3(32'h3a3cdb7f),
	.w4(32'hbb2b0445),
	.w5(32'hbb7520c9),
	.w6(32'h3b3d5084),
	.w7(32'h3a7aa9e3),
	.w8(32'hbb0a0d52),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b797098),
	.w1(32'h3b751290),
	.w2(32'h3bb098fc),
	.w3(32'h3b6901f9),
	.w4(32'h3b9bd8ea),
	.w5(32'h3b83a030),
	.w6(32'h3c11c4eb),
	.w7(32'h3c07f883),
	.w8(32'h3bb62405),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f7aef),
	.w1(32'hb9f34754),
	.w2(32'h3a864cc5),
	.w3(32'h398872c6),
	.w4(32'h37bc2f1c),
	.w5(32'h3ad9a1ff),
	.w6(32'hb6bc5b1f),
	.w7(32'h396903a9),
	.w8(32'hb8e7b959),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09b389),
	.w1(32'hbbb4d019),
	.w2(32'hbb04e973),
	.w3(32'hbb87ce1f),
	.w4(32'hbb684ec5),
	.w5(32'hbb6bcdd9),
	.w6(32'hbb12b1bd),
	.w7(32'hba9da4bf),
	.w8(32'hbb8abbe2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c40d6f),
	.w1(32'hb9d89322),
	.w2(32'hb98f587f),
	.w3(32'hb9f1e031),
	.w4(32'hba571fbc),
	.w5(32'hba523f28),
	.w6(32'h39a50512),
	.w7(32'h39b3d9ac),
	.w8(32'h3ab4bddb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913c4db),
	.w1(32'hbb8ca90d),
	.w2(32'hbbbab2a7),
	.w3(32'h3be434e5),
	.w4(32'h3b87b3c3),
	.w5(32'h3b0afe6a),
	.w6(32'h3bc3ebf5),
	.w7(32'h3b8f2761),
	.w8(32'h3a9064b3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba388e4f),
	.w1(32'hbac0c5ea),
	.w2(32'hba39efc9),
	.w3(32'h3af69d88),
	.w4(32'h389b06d5),
	.w5(32'h3a3fd8fd),
	.w6(32'h3b84ebdc),
	.w7(32'h3b7c1f1c),
	.w8(32'h3b3c4fb0),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62f70d),
	.w1(32'hbba64c97),
	.w2(32'hbc28a72b),
	.w3(32'hba9c7c73),
	.w4(32'hbb20c6d6),
	.w5(32'hbbc6a703),
	.w6(32'h3af409c9),
	.w7(32'hbb4a41f6),
	.w8(32'hbaca1c43),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06cad6),
	.w1(32'h3c0f7fd3),
	.w2(32'h3bf24108),
	.w3(32'h3bda511d),
	.w4(32'h3c08d5fb),
	.w5(32'h3c02ffe7),
	.w6(32'h3b83b76e),
	.w7(32'h3ba558b8),
	.w8(32'h3badacf4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d3597),
	.w1(32'h3a6b6635),
	.w2(32'h3a96f91e),
	.w3(32'h3b25d623),
	.w4(32'h3b601cab),
	.w5(32'h3b2acc99),
	.w6(32'h3aa056bb),
	.w7(32'h3b205775),
	.w8(32'h3ac0ecaa),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f72205),
	.w1(32'hbbb71376),
	.w2(32'hbbd89b05),
	.w3(32'h3aca5f0b),
	.w4(32'hbb59e2c3),
	.w5(32'hbb9d5915),
	.w6(32'h3b6e9c78),
	.w7(32'h38bb87a4),
	.w8(32'hbb0ead48),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb899fc6c),
	.w1(32'h3a048406),
	.w2(32'h3a726506),
	.w3(32'hbaafcd56),
	.w4(32'h3a1d6610),
	.w5(32'h3a1fac74),
	.w6(32'h3a441427),
	.w7(32'h3b5d9543),
	.w8(32'h3b0332fe),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99788d3),
	.w1(32'h3834cec2),
	.w2(32'h397bab6f),
	.w3(32'hba1a390e),
	.w4(32'h398f9881),
	.w5(32'h394bbb17),
	.w6(32'h39dadb7f),
	.w7(32'h3abfc49e),
	.w8(32'h39679d2c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e2d75),
	.w1(32'h3a8297c8),
	.w2(32'h3a809bbc),
	.w3(32'hb9602a4c),
	.w4(32'h39abb569),
	.w5(32'hb8dd46ec),
	.w6(32'h3abd9200),
	.w7(32'h391668e3),
	.w8(32'hbb16ce73),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ff471),
	.w1(32'h3b20fda8),
	.w2(32'h39972760),
	.w3(32'h3b96f172),
	.w4(32'h3befccb7),
	.w5(32'hbb112bd9),
	.w6(32'hbb16dd7b),
	.w7(32'hb9f469cb),
	.w8(32'h3aaec665),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a0876),
	.w1(32'hbaa56c23),
	.w2(32'hbaaf4a15),
	.w3(32'h3ba40cb2),
	.w4(32'h3b133397),
	.w5(32'h3ae3b47d),
	.w6(32'h3b7a892b),
	.w7(32'h3ac26afd),
	.w8(32'h3b854233),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9868d2),
	.w1(32'h3c8eabe5),
	.w2(32'h39cf4b1c),
	.w3(32'h3c51c0ab),
	.w4(32'h3c650a13),
	.w5(32'h3b042864),
	.w6(32'h3c290475),
	.w7(32'h3c579f01),
	.w8(32'hbbe68e49),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f70ba),
	.w1(32'hba2f88be),
	.w2(32'hbb41a4d5),
	.w3(32'h3a9b16bd),
	.w4(32'hba8e79c6),
	.w5(32'h3b80264f),
	.w6(32'hbba49a99),
	.w7(32'hbc02939e),
	.w8(32'h3b1b023b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac69918),
	.w1(32'h39a5467c),
	.w2(32'h3b908f30),
	.w3(32'hbb995459),
	.w4(32'hb9fb99be),
	.w5(32'h3b540b89),
	.w6(32'hbb902b23),
	.w7(32'hbb639726),
	.w8(32'hba91f63e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8b15a),
	.w1(32'hbbcaeec1),
	.w2(32'hbb8f372b),
	.w3(32'h3b6ab34a),
	.w4(32'hba870b6d),
	.w5(32'h3a694ea7),
	.w6(32'h3bda87cf),
	.w7(32'h3bb36e5c),
	.w8(32'h3b12e875),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37efca),
	.w1(32'h3c8c137d),
	.w2(32'h3bc3b9e8),
	.w3(32'h3c4d54f0),
	.w4(32'h3c92bf67),
	.w5(32'h3c28b4a5),
	.w6(32'h3b0a535f),
	.w7(32'h3bc161a2),
	.w8(32'h3b9e30c7),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95a097),
	.w1(32'hbb4b06e1),
	.w2(32'hba8c2832),
	.w3(32'h3b33ef18),
	.w4(32'h3a0d253e),
	.w5(32'h3b894d9a),
	.w6(32'h3b716b05),
	.w7(32'h3b93c2f4),
	.w8(32'h3b8f9370),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b95c),
	.w1(32'h3b8d5dd1),
	.w2(32'h3c0e8437),
	.w3(32'h3c15af1f),
	.w4(32'h3a767d4f),
	.w5(32'h3bdd9849),
	.w6(32'h3c375d5a),
	.w7(32'h3ab093c7),
	.w8(32'h3bab0989),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83a60b),
	.w1(32'h3b949320),
	.w2(32'h3b98e396),
	.w3(32'h3b92a24e),
	.w4(32'h3bd993d3),
	.w5(32'h3c042a58),
	.w6(32'hb99ed890),
	.w7(32'h3a8e48a0),
	.w8(32'h3b285791),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb817550c),
	.w1(32'h3a311fb6),
	.w2(32'h3ac83fc4),
	.w3(32'h3985fedf),
	.w4(32'h3a75959d),
	.w5(32'h3b19bb93),
	.w6(32'hbaf84543),
	.w7(32'hbae79607),
	.w8(32'hb9a805fa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e17b25d),
	.w1(32'h3dcc6065),
	.w2(32'h3d644f8b),
	.w3(32'h3db1f05c),
	.w4(32'h3d64f3f1),
	.w5(32'h3c7a6b0c),
	.w6(32'h3d48f5aa),
	.w7(32'hbc8c41cf),
	.w8(32'hbbb71a10),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88ede6),
	.w1(32'h398bec8b),
	.w2(32'hbc08a757),
	.w3(32'hb9c021fe),
	.w4(32'h3b9a8a24),
	.w5(32'hbb94d510),
	.w6(32'hbbbbd328),
	.w7(32'hbbe5872a),
	.w8(32'hbaf365bd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a642529),
	.w1(32'h37aefb32),
	.w2(32'h3a4e75e8),
	.w3(32'h3af07965),
	.w4(32'h3a941410),
	.w5(32'h3b2dfccf),
	.w6(32'h3b4b0c54),
	.w7(32'h3b14d416),
	.w8(32'h398466e3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d150f),
	.w1(32'h3b384e14),
	.w2(32'h3a45416d),
	.w3(32'hbb869a50),
	.w4(32'h39c44aa0),
	.w5(32'hbb2b5034),
	.w6(32'hbbd454ea),
	.w7(32'hbb8507fe),
	.w8(32'hbb57cf5f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe0aac),
	.w1(32'hba1a09e7),
	.w2(32'h3ad425eb),
	.w3(32'h3a8ac0aa),
	.w4(32'hba7a0916),
	.w5(32'h3ae52571),
	.w6(32'h3a7e62cc),
	.w7(32'hbb199fa2),
	.w8(32'hbb78ff8e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f7f3),
	.w1(32'hbb875a23),
	.w2(32'hbb8e52b6),
	.w3(32'hba881f3b),
	.w4(32'h3af79229),
	.w5(32'hb9bec622),
	.w6(32'h3af8e27e),
	.w7(32'h3ac39a60),
	.w8(32'h370691a9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e831),
	.w1(32'h3c013a64),
	.w2(32'h3b908c41),
	.w3(32'h3a3ce68a),
	.w4(32'hba96dc7a),
	.w5(32'hb9a059b2),
	.w6(32'hba38ceec),
	.w7(32'h3ab9f223),
	.w8(32'hb9732a92),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56c9df),
	.w1(32'hbbde8134),
	.w2(32'hbbe0d1e7),
	.w3(32'hbb8cbfab),
	.w4(32'hbbd3ab97),
	.w5(32'hbbb3a6f1),
	.w6(32'hbb0f4f5a),
	.w7(32'hbb32cbf0),
	.w8(32'hbb92fee3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1b1d9),
	.w1(32'h3ac09342),
	.w2(32'hbb4fb0c3),
	.w3(32'h3bc028ef),
	.w4(32'h3b62965b),
	.w5(32'hb9954ac1),
	.w6(32'h3ba56998),
	.w7(32'h3b2a1b32),
	.w8(32'hbb48b881),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38385f03),
	.w1(32'h3a17774b),
	.w2(32'h3abb3bd6),
	.w3(32'h37da9a7f),
	.w4(32'hba395b6b),
	.w5(32'h39b976f9),
	.w6(32'hb9bbc1ac),
	.w7(32'hba9082e2),
	.w8(32'h3ab010d7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826eae),
	.w1(32'hbb86750b),
	.w2(32'hbaff48d6),
	.w3(32'hbb10c4d1),
	.w4(32'hbb44f526),
	.w5(32'hbadde2ef),
	.w6(32'hb9c33d74),
	.w7(32'hba832a0a),
	.w8(32'hba426353),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cc3b3),
	.w1(32'hb8231db7),
	.w2(32'h39e65d3b),
	.w3(32'hba47cb39),
	.w4(32'h39f12979),
	.w5(32'h397aff4a),
	.w6(32'h3a0527da),
	.w7(32'h3b1620e2),
	.w8(32'hba0e2377),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ff38f),
	.w1(32'h3924b7ae),
	.w2(32'h39c8eeb0),
	.w3(32'hb9902fea),
	.w4(32'hb993e737),
	.w5(32'h39f255fd),
	.w6(32'h3a0bd7c7),
	.w7(32'h39c7a699),
	.w8(32'h39e26867),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a6903),
	.w1(32'h3c353d1e),
	.w2(32'h3c696f64),
	.w3(32'h3ce5d7ae),
	.w4(32'h3cb2989a),
	.w5(32'h3cb6b2e3),
	.w6(32'h3ccd0c77),
	.w7(32'h3c8a181f),
	.w8(32'h3c8557f4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345b70),
	.w1(32'h3a689ae1),
	.w2(32'hbb2ff598),
	.w3(32'h3b46f5f6),
	.w4(32'h3a642483),
	.w5(32'hbb0604cb),
	.w6(32'h3b757d66),
	.w7(32'hb956d16e),
	.w8(32'hbb481845),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6259b6),
	.w1(32'hbac4388e),
	.w2(32'hbb815d11),
	.w3(32'hb9f46c7e),
	.w4(32'hba9f7101),
	.w5(32'hbb0d8c22),
	.w6(32'h3a465692),
	.w7(32'hbb31ac3f),
	.w8(32'hbb1218ee),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6780),
	.w1(32'h3ba1cc9a),
	.w2(32'h3b7156ce),
	.w3(32'h3bbcc984),
	.w4(32'h3b9fcc23),
	.w5(32'h3b9d89f5),
	.w6(32'h3bf5a42c),
	.w7(32'h3b8f62fe),
	.w8(32'h3b0b1c41),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcb1ef),
	.w1(32'h3b924ec7),
	.w2(32'h3b251f6b),
	.w3(32'h3b7d1ee8),
	.w4(32'h3c05213b),
	.w5(32'h3bb049a5),
	.w6(32'h3ae30c15),
	.w7(32'h3b3f66b9),
	.w8(32'h3a114877),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873895),
	.w1(32'hbb04c04c),
	.w2(32'hbb9972b8),
	.w3(32'h3bc0c1cf),
	.w4(32'hba93bcbb),
	.w5(32'hbb8c5c8d),
	.w6(32'h3bb0fa4b),
	.w7(32'h3941a6b7),
	.w8(32'hba860afe),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa56c26),
	.w1(32'hbadc1c53),
	.w2(32'hba36644f),
	.w3(32'hba5853a6),
	.w4(32'h39bc7c60),
	.w5(32'hb8824b8a),
	.w6(32'h3a40c277),
	.w7(32'hb9d7fbe7),
	.w8(32'h3a9e0eed),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b204a53),
	.w1(32'h3b79359d),
	.w2(32'h3aa135c6),
	.w3(32'h3ba00c6e),
	.w4(32'h3bdc33a5),
	.w5(32'h3bc1b14a),
	.w6(32'h3a9d70f7),
	.w7(32'h3ba28fdf),
	.w8(32'h3b879f4b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b595d76),
	.w1(32'h3b7d65d4),
	.w2(32'h3b5fa44d),
	.w3(32'h3b77730f),
	.w4(32'h3b8a9368),
	.w5(32'h3b8f675b),
	.w6(32'h3b461050),
	.w7(32'h3b63e570),
	.w8(32'hb9d74333),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295840),
	.w1(32'h3bc7b7b0),
	.w2(32'h3bcd4485),
	.w3(32'h3b279922),
	.w4(32'h3babe521),
	.w5(32'h3bd688cd),
	.w6(32'h3b862697),
	.w7(32'h3bd2e848),
	.w8(32'h3be01523),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5114f2),
	.w1(32'hbc841248),
	.w2(32'hbc8c8ce9),
	.w3(32'hbc3e28de),
	.w4(32'hbc847bc5),
	.w5(32'hbc87362a),
	.w6(32'hbc09fae4),
	.w7(32'hbc6dbe02),
	.w8(32'hbc86151b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c872ead),
	.w1(32'h3ca91719),
	.w2(32'h3bdc9081),
	.w3(32'h3c94a9cb),
	.w4(32'h3cce6858),
	.w5(32'h3c658f60),
	.w6(32'h3c37775c),
	.w7(32'h3c6139a1),
	.w8(32'h3bf3c8ec),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce7d8),
	.w1(32'h3b9e759a),
	.w2(32'h3b8b1ca3),
	.w3(32'h3baa8888),
	.w4(32'h3ba754ff),
	.w5(32'h3b83fb04),
	.w6(32'h3a0cefe4),
	.w7(32'h3b2e2f57),
	.w8(32'h3be70b9a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea1b7f),
	.w1(32'h3c05ac09),
	.w2(32'h3b7b1eaa),
	.w3(32'h3c014454),
	.w4(32'h3c034e40),
	.w5(32'h3bede1f1),
	.w6(32'h3bab8463),
	.w7(32'h3bc50e60),
	.w8(32'h3b474861),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39232ef6),
	.w1(32'hba7dd11d),
	.w2(32'hba00a2d9),
	.w3(32'h39f74834),
	.w4(32'h3a030c47),
	.w5(32'hb8132288),
	.w6(32'hb7815406),
	.w7(32'hb9da8ec7),
	.w8(32'h3aaf6a72),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62a6fb),
	.w1(32'h3c3fddd3),
	.w2(32'h3bbc6ae0),
	.w3(32'h3bf1fe53),
	.w4(32'h3c25e94e),
	.w5(32'h3ba83984),
	.w6(32'h3bb620d9),
	.w7(32'h3bb67fe5),
	.w8(32'h3a37763d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae26b83),
	.w1(32'hba3c7aac),
	.w2(32'hbb1edd8d),
	.w3(32'hba412fc5),
	.w4(32'hba3c4441),
	.w5(32'hbb36601b),
	.w6(32'hbb1955ef),
	.w7(32'hbaf270ce),
	.w8(32'hbb79ac7b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b709ca4),
	.w1(32'h3a9828b2),
	.w2(32'hbbc610e9),
	.w3(32'h3c08770d),
	.w4(32'h3be2d33c),
	.w5(32'h39af2e70),
	.w6(32'h3c12eab3),
	.w7(32'h3b4cee8d),
	.w8(32'hbb8d4267),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbf2fe),
	.w1(32'h3bd22492),
	.w2(32'h3ba1f220),
	.w3(32'hbb157247),
	.w4(32'h3b69c33e),
	.w5(32'h3b754e00),
	.w6(32'hbab43761),
	.w7(32'h3b114a36),
	.w8(32'h3b04e633),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ceb79),
	.w1(32'h3bc5358c),
	.w2(32'h3ba1d265),
	.w3(32'h3b7dde07),
	.w4(32'h3bb67cde),
	.w5(32'h3bcb9e6d),
	.w6(32'h3bc883c9),
	.w7(32'h3b87acc8),
	.w8(32'h3bc307a4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5f206),
	.w1(32'hb9b06686),
	.w2(32'h3a3ab3f3),
	.w3(32'h3b08b7ac),
	.w4(32'h3aa93e46),
	.w5(32'h3b163a17),
	.w6(32'h3b70f88f),
	.w7(32'h3b20217c),
	.w8(32'h3ad8210f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3446),
	.w1(32'hbadc8552),
	.w2(32'h3a1bc70a),
	.w3(32'h3a967794),
	.w4(32'h3ab801e4),
	.w5(32'h3b0325f7),
	.w6(32'hbb1dcee5),
	.w7(32'h3a7f9e7c),
	.w8(32'h3a264470),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3977c),
	.w1(32'h3b5c838e),
	.w2(32'h3b224196),
	.w3(32'h3c4a59b6),
	.w4(32'h3bebc045),
	.w5(32'h3c0f8d6f),
	.w6(32'h3ba13ea3),
	.w7(32'hb9017572),
	.w8(32'hb9f3b4d5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39910a36),
	.w1(32'hb9955fb3),
	.w2(32'hbada04c6),
	.w3(32'h3aa88cab),
	.w4(32'h3a006580),
	.w5(32'hba7bd799),
	.w6(32'h3b067b06),
	.w7(32'h3b71a99f),
	.w8(32'hba9e8b14),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba63df32),
	.w1(32'h39d1e3d8),
	.w2(32'h39fbee76),
	.w3(32'hba967392),
	.w4(32'hba30ea20),
	.w5(32'h3a22e5ff),
	.w6(32'hb9bada3d),
	.w7(32'hba3ee609),
	.w8(32'h39de4498),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af93dfe),
	.w1(32'h3af7c1fe),
	.w2(32'hbaa743d5),
	.w3(32'h3b9a5973),
	.w4(32'h3b126de6),
	.w5(32'h3a3f0217),
	.w6(32'h3ba6077a),
	.w7(32'h3acef1f7),
	.w8(32'hb93e8c8c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a5b82),
	.w1(32'h3a047bb1),
	.w2(32'hba998dd1),
	.w3(32'h3b062de6),
	.w4(32'h39342eea),
	.w5(32'h39a598d9),
	.w6(32'h3b819bc3),
	.w7(32'h3ac23fc3),
	.w8(32'hbaa3e1a4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847a009),
	.w1(32'hb7de7127),
	.w2(32'hb8d9c14f),
	.w3(32'h3ad67a8a),
	.w4(32'hb80ac6cb),
	.w5(32'h3ada75a0),
	.w6(32'hbaee6ee2),
	.w7(32'hbb77c3e8),
	.w8(32'hbb316036),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c240),
	.w1(32'hbb17f39f),
	.w2(32'hbaab8b22),
	.w3(32'hbb2f2466),
	.w4(32'hbb550fc6),
	.w5(32'hba9466ea),
	.w6(32'hbb5e23e4),
	.w7(32'hbb63ae26),
	.w8(32'hbbf815da),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ab83d),
	.w1(32'h3c647b7d),
	.w2(32'h3c64fcf8),
	.w3(32'h3bc949bb),
	.w4(32'h3c80309d),
	.w5(32'h3c78efaf),
	.w6(32'h3bb1d169),
	.w7(32'h3c0371b4),
	.w8(32'h3bf4533e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2895e),
	.w1(32'hb9954430),
	.w2(32'hba83f156),
	.w3(32'hbaddee5d),
	.w4(32'hba5bf55c),
	.w5(32'hba98997d),
	.w6(32'hba2a7014),
	.w7(32'hbac37cb0),
	.w8(32'hbb0d3365),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e0697),
	.w1(32'hba089f51),
	.w2(32'h3b406eaa),
	.w3(32'h3b66f54e),
	.w4(32'h3b3f213c),
	.w5(32'h3bca080a),
	.w6(32'h3b075b82),
	.w7(32'h3aac0e50),
	.w8(32'h3ba8904e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46770d),
	.w1(32'h3b6cf4a2),
	.w2(32'h3b0ce938),
	.w3(32'h39161b71),
	.w4(32'h3af37295),
	.w5(32'h3ab73a8d),
	.w6(32'h3a43eb97),
	.w7(32'h3a00c672),
	.w8(32'h3aa18366),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838f38),
	.w1(32'hb9f6eff4),
	.w2(32'hba7d4ecc),
	.w3(32'h3c010814),
	.w4(32'h3823053b),
	.w5(32'h3b0479a5),
	.w6(32'h3c02b8ec),
	.w7(32'h3a072f07),
	.w8(32'h3b16c832),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba043e36),
	.w1(32'hba633c51),
	.w2(32'hba647f78),
	.w3(32'hb94d0528),
	.w4(32'hba4bde2e),
	.w5(32'hba059ef3),
	.w6(32'hb9288ffd),
	.w7(32'hb9a33aeb),
	.w8(32'hb81e7ea1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967c21),
	.w1(32'h3bea32eb),
	.w2(32'h3b67123c),
	.w3(32'h3b322c1e),
	.w4(32'h3bb1aa41),
	.w5(32'h3b0baf32),
	.w6(32'hbb056b12),
	.w7(32'h39f61c04),
	.w8(32'h3ad89d3f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb808af8c),
	.w1(32'h3a269cb0),
	.w2(32'h39ee6e95),
	.w3(32'h3982b61f),
	.w4(32'h39ce7baa),
	.w5(32'h3a1b3c60),
	.w6(32'h3998452a),
	.w7(32'h38b0b12c),
	.w8(32'hbbf14ad6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab78fb5),
	.w1(32'h3b87f4e0),
	.w2(32'h3a23ed04),
	.w3(32'h3a18fae5),
	.w4(32'h3b72eba4),
	.w5(32'h3b13b0bb),
	.w6(32'h3a763b89),
	.w7(32'h3810cd03),
	.w8(32'hbacd5e19),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d486),
	.w1(32'hbc001bab),
	.w2(32'hbc31e617),
	.w3(32'hba8b07ac),
	.w4(32'hbbabfa55),
	.w5(32'hbbed9a63),
	.w6(32'hbb344c08),
	.w7(32'hbbeca37e),
	.w8(32'hbbeb4311),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a7a42),
	.w1(32'h3b19aec8),
	.w2(32'h3a2f0ae6),
	.w3(32'h3b2495da),
	.w4(32'h3b2e8ee7),
	.w5(32'h3a2e4b3b),
	.w6(32'h3b86cf28),
	.w7(32'h3b114b72),
	.w8(32'hb9e52c9f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c32c),
	.w1(32'hba3c38be),
	.w2(32'hbb112c1a),
	.w3(32'hba93adae),
	.w4(32'hba4f1470),
	.w5(32'hba9a1b9c),
	.w6(32'hba26533b),
	.w7(32'hbb211357),
	.w8(32'hb957bc78),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84c5a8),
	.w1(32'h3bbebc3e),
	.w2(32'h3bf6df92),
	.w3(32'h3bbb6a3a),
	.w4(32'h3c065221),
	.w5(32'h3c22322c),
	.w6(32'h3bc3630a),
	.w7(32'h3bf9d8a9),
	.w8(32'h3ba46ad6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac55cd),
	.w1(32'h3acc16d6),
	.w2(32'h3b32b7c7),
	.w3(32'h3bf64914),
	.w4(32'h3bcd99af),
	.w5(32'h3bf7f844),
	.w6(32'h3b6c3901),
	.w7(32'h3b890a55),
	.w8(32'h3baffd8b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c242177),
	.w1(32'h3c000ee2),
	.w2(32'h3c5c4642),
	.w3(32'h3cb1b9c4),
	.w4(32'h3c672392),
	.w5(32'h3cae4fd1),
	.w6(32'h3cac86fb),
	.w7(32'h3c305584),
	.w8(32'h3c8575f4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d010e),
	.w1(32'h3c16eba8),
	.w2(32'h3c241ba8),
	.w3(32'h3c85d7b0),
	.w4(32'h3c5dc541),
	.w5(32'h3c686099),
	.w6(32'h3bf5f0b8),
	.w7(32'h3b364253),
	.w8(32'h3b19feea),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5d5da),
	.w1(32'h3bd8e2e2),
	.w2(32'h3c0432bb),
	.w3(32'h3b1b3258),
	.w4(32'h3be69deb),
	.w5(32'h3c37106d),
	.w6(32'hbb0371fc),
	.w7(32'h3a0df959),
	.w8(32'h3bfdf134),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3717ff),
	.w1(32'h3b54c909),
	.w2(32'h3b679f66),
	.w3(32'h3ae67e09),
	.w4(32'h3b199de5),
	.w5(32'h3b312eaa),
	.w6(32'h3b50be05),
	.w7(32'h3b613249),
	.w8(32'hb980ef6d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba5634),
	.w1(32'hba97f4a7),
	.w2(32'hba3ff0af),
	.w3(32'hba08480d),
	.w4(32'hbab592d8),
	.w5(32'hb9cdbc9f),
	.w6(32'hb9aa7302),
	.w7(32'hb8ffcd12),
	.w8(32'h3a275a43),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39827ea5),
	.w1(32'hba857de1),
	.w2(32'hba91610b),
	.w3(32'hbabd59ec),
	.w4(32'hbadd000c),
	.w5(32'hbadf37f3),
	.w6(32'hbaeb2c1f),
	.w7(32'hbac8016d),
	.w8(32'h3b5d51a9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8483ab),
	.w1(32'h3baf29f1),
	.w2(32'h3bc30648),
	.w3(32'h3b9a527a),
	.w4(32'h3be94aaf),
	.w5(32'h3bb37955),
	.w6(32'h3b846ed1),
	.w7(32'h3b8a49cb),
	.w8(32'h3b640460),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e780),
	.w1(32'h3c1a38b2),
	.w2(32'h3c39d5a7),
	.w3(32'h3c056715),
	.w4(32'h3c2d3888),
	.w5(32'h3c3a3d78),
	.w6(32'h3ba0a661),
	.w7(32'h3bb77a7f),
	.w8(32'h3c0bad87),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39f1ab),
	.w1(32'h39a95b03),
	.w2(32'hb97bc978),
	.w3(32'hba889b8c),
	.w4(32'hbb561fd6),
	.w5(32'hbb4d571c),
	.w6(32'h39282d1c),
	.w7(32'hbb6f85d9),
	.w8(32'hbb0f3c92),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b284343),
	.w1(32'hbaa81f08),
	.w2(32'h3afcf78d),
	.w3(32'h3bb5ba72),
	.w4(32'h3ab12931),
	.w5(32'h3b865a0d),
	.w6(32'h3b8bd582),
	.w7(32'h3acaf88d),
	.w8(32'hba3ad344),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8d20),
	.w1(32'h3b8f5d3b),
	.w2(32'h3bb4c3b9),
	.w3(32'h3ba9836c),
	.w4(32'h3bf800b7),
	.w5(32'h3c0d5f70),
	.w6(32'h3ba9d36b),
	.w7(32'h3bb09294),
	.w8(32'h3bf73db3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce535e),
	.w1(32'hbbdf4280),
	.w2(32'hbb6866f3),
	.w3(32'hb9ff5b5b),
	.w4(32'h3b12bc86),
	.w5(32'h3b822848),
	.w6(32'hba4cf78c),
	.w7(32'h3b1e0393),
	.w8(32'h3bb30dd2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1e513),
	.w1(32'hbb8e8470),
	.w2(32'hbbc79c42),
	.w3(32'h3b29cbfb),
	.w4(32'hbb60afb5),
	.w5(32'hbbe6efc1),
	.w6(32'h3a8dc787),
	.w7(32'hbb1accd5),
	.w8(32'hbb752056),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b055e5c),
	.w1(32'h3b6d7b78),
	.w2(32'hbab4b7b9),
	.w3(32'h3b8c9b0d),
	.w4(32'h3bc55fce),
	.w5(32'h3b44367e),
	.w6(32'hbbaaf02b),
	.w7(32'hbadb6e9a),
	.w8(32'hbb79f29a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a191eff),
	.w1(32'h3b0fc1ef),
	.w2(32'h3b062aef),
	.w3(32'h393dcfde),
	.w4(32'h3aa87b39),
	.w5(32'h39927cd9),
	.w6(32'hba3d75d8),
	.w7(32'h3a2cb6f2),
	.w8(32'hbbdf8d0c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc40eef),
	.w1(32'hbb4fd7b1),
	.w2(32'hbb503654),
	.w3(32'hbbd0f492),
	.w4(32'hbb7c1eb5),
	.w5(32'hbb644eb0),
	.w6(32'hbb904ec1),
	.w7(32'hbb85515c),
	.w8(32'hb7635dfd),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b72828),
	.w1(32'hb92bc1f3),
	.w2(32'hb9dddb47),
	.w3(32'hba076dd8),
	.w4(32'hb99ed3ec),
	.w5(32'hb8df454c),
	.w6(32'h3a06848f),
	.w7(32'h39d6e1e3),
	.w8(32'hb987b482),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38749c26),
	.w1(32'hb911cbc5),
	.w2(32'hba35ab15),
	.w3(32'hbad4cf8f),
	.w4(32'hbaf6c8d7),
	.w5(32'hbaa1196d),
	.w6(32'hb9d30dae),
	.w7(32'hba7ff314),
	.w8(32'hb9f45cf8),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4b2c2),
	.w1(32'h3a4e7acf),
	.w2(32'h3aa694b0),
	.w3(32'h3b2a252d),
	.w4(32'h3b2e3d71),
	.w5(32'h3b433450),
	.w6(32'h3b4186ea),
	.w7(32'h3b5388b4),
	.w8(32'hbb14f783),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddbfb1),
	.w1(32'hbc0004b8),
	.w2(32'hbbb09816),
	.w3(32'hbbf0425d),
	.w4(32'hbc033537),
	.w5(32'hbb845029),
	.w6(32'hbbe6d70c),
	.w7(32'hbc076a0a),
	.w8(32'h3b05941b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc92ef),
	.w1(32'h3b8f4d24),
	.w2(32'h3abc576b),
	.w3(32'h3c03e693),
	.w4(32'h3b2fcad8),
	.w5(32'h3b12276b),
	.w6(32'h3c1b0a81),
	.w7(32'h3ba52e2c),
	.w8(32'h3b7aa698),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4fb6f),
	.w1(32'h39e954bc),
	.w2(32'h3b158116),
	.w3(32'h3aa0b525),
	.w4(32'h39e7ff82),
	.w5(32'h3b38ef15),
	.w6(32'h3b0d45e9),
	.w7(32'h3b0d29e9),
	.w8(32'h3ac23b74),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d7156),
	.w1(32'h3c77d865),
	.w2(32'h3c8e36c8),
	.w3(32'h3c4086d9),
	.w4(32'h3c70b560),
	.w5(32'h3c98d009),
	.w6(32'h3bf301b4),
	.w7(32'h3c079b94),
	.w8(32'h3c3adddc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadcfb2),
	.w1(32'h39676e9e),
	.w2(32'h3b9335bd),
	.w3(32'hba358f94),
	.w4(32'h3b38ba8b),
	.w5(32'h3baccf79),
	.w6(32'hba0c48c5),
	.w7(32'h3b8e0d47),
	.w8(32'h3ba8622c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b683f82),
	.w1(32'hbad0103b),
	.w2(32'h398d169c),
	.w3(32'h3bb55b56),
	.w4(32'h3b1fc004),
	.w5(32'h3b81c6ae),
	.w6(32'h3b451a79),
	.w7(32'h3b22c9d1),
	.w8(32'h3b68c577),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab394eb),
	.w1(32'hba28d15c),
	.w2(32'h3a5b5a2b),
	.w3(32'hba4afe06),
	.w4(32'h39284dbf),
	.w5(32'h3a35ced5),
	.w6(32'hbb097379),
	.w7(32'hb963f064),
	.w8(32'hba5dccb3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d0ab2),
	.w1(32'hb7c46cd5),
	.w2(32'hb940b0fc),
	.w3(32'h3b4c8b48),
	.w4(32'h3b987f27),
	.w5(32'h3b0a0656),
	.w6(32'h39a3d0bc),
	.w7(32'h3af0aabe),
	.w8(32'hbbccec7b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6b3a7),
	.w1(32'h3c610f3a),
	.w2(32'h3aaf29ad),
	.w3(32'hb905ffc7),
	.w4(32'hba9a4d38),
	.w5(32'h39f87e70),
	.w6(32'hba7cb053),
	.w7(32'hbb1f7734),
	.w8(32'hbbdfd008),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b73190),
	.w1(32'h3a8f85b9),
	.w2(32'h3b7ef880),
	.w3(32'hbb0743c8),
	.w4(32'hb992a5af),
	.w5(32'h384855a4),
	.w6(32'hbb47b689),
	.w7(32'hbb9a5784),
	.w8(32'h3aebfe0d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e971a),
	.w1(32'hbb4ec9f5),
	.w2(32'hbad918da),
	.w3(32'h39ca7517),
	.w4(32'hbb408c0f),
	.w5(32'hbaa8a544),
	.w6(32'hba3404a0),
	.w7(32'hbb0bf4f5),
	.w8(32'hba8b1244),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d65ac1),
	.w1(32'h3a3fc001),
	.w2(32'h3a0b61d0),
	.w3(32'h3ae4d789),
	.w4(32'h3b1002cc),
	.w5(32'h3aaab53e),
	.w6(32'h39e3a9d8),
	.w7(32'h3a441476),
	.w8(32'h38c0a5bd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3faf3c),
	.w1(32'h3a6ecbfd),
	.w2(32'h398a8fed),
	.w3(32'h3adc230b),
	.w4(32'h3b07dc44),
	.w5(32'h39a2bb99),
	.w6(32'h3a5e23d8),
	.w7(32'h3ad506f9),
	.w8(32'h39e36c8c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac19fa3),
	.w1(32'h38986309),
	.w2(32'h3abf9a82),
	.w3(32'h3b299070),
	.w4(32'h3b0dc29b),
	.w5(32'h3a422b05),
	.w6(32'hb8dca640),
	.w7(32'hb980c45e),
	.w8(32'h3a912ae5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c5d63),
	.w1(32'hbbb7b1a8),
	.w2(32'h39b1c280),
	.w3(32'hbb649cd2),
	.w4(32'hbb8e2463),
	.w5(32'hba87c062),
	.w6(32'hbb9e8da0),
	.w7(32'hbbe0bab6),
	.w8(32'h3b9a7bce),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d5a02),
	.w1(32'h3c10eb0d),
	.w2(32'h3bf7e026),
	.w3(32'h3c343fcd),
	.w4(32'h3c3563d1),
	.w5(32'h3c23f7ba),
	.w6(32'h3b9d6a68),
	.w7(32'h3b94010f),
	.w8(32'hb9ceb2e5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13ce38),
	.w1(32'h3c6cda6d),
	.w2(32'h397d3f9b),
	.w3(32'hbafc3b04),
	.w4(32'h3c01d9b9),
	.w5(32'hb9f01f6f),
	.w6(32'h3beeb417),
	.w7(32'hba2520c4),
	.w8(32'hbb8cb5f0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e638b),
	.w1(32'hbafc667c),
	.w2(32'h3a30645f),
	.w3(32'hbae7d267),
	.w4(32'h3a830ee2),
	.w5(32'h3a2d1134),
	.w6(32'hbb1613d2),
	.w7(32'h3acb3e10),
	.w8(32'hbacc010b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20d3b7),
	.w1(32'hb98be0a2),
	.w2(32'hbac9bace),
	.w3(32'h3ba73d94),
	.w4(32'h3b6277ea),
	.w5(32'h3bafa36a),
	.w6(32'hbabd3685),
	.w7(32'hbb5ae110),
	.w8(32'h39f3c158),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba63388),
	.w1(32'h3baf810c),
	.w2(32'h3b4eef2d),
	.w3(32'hbb306bf4),
	.w4(32'h3c243a2c),
	.w5(32'h3b90a79b),
	.w6(32'h3b12b03a),
	.w7(32'hba68b341),
	.w8(32'h3b505353),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb04cb),
	.w1(32'hba42c137),
	.w2(32'h3ae63422),
	.w3(32'h3a9110bd),
	.w4(32'hb929bcda),
	.w5(32'h3a3f060b),
	.w6(32'h36145d1d),
	.w7(32'h3a61e0d4),
	.w8(32'h39674105),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e295),
	.w1(32'hbab08fcd),
	.w2(32'hbbec85de),
	.w3(32'hbb02e2ea),
	.w4(32'hbbbd8447),
	.w5(32'hbc114ae5),
	.w6(32'hba7b5a87),
	.w7(32'hbbbf4b2f),
	.w8(32'hbb92aa25),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62970d),
	.w1(32'h3ab79cef),
	.w2(32'h3a41e646),
	.w3(32'hbb08986f),
	.w4(32'h3aebe5b9),
	.w5(32'hbb2a5357),
	.w6(32'hbba57eb7),
	.w7(32'hba4d1351),
	.w8(32'hbb6535fb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a71d4),
	.w1(32'h39f1a9cd),
	.w2(32'hb9af95f0),
	.w3(32'hbaa349e7),
	.w4(32'h39ed3bef),
	.w5(32'hbac08b10),
	.w6(32'hbac46c93),
	.w7(32'hbacbe484),
	.w8(32'hba2d5e96),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f74fe),
	.w1(32'hbb220239),
	.w2(32'h3a927708),
	.w3(32'h3c075bbf),
	.w4(32'h3b01d6b2),
	.w5(32'h3b246881),
	.w6(32'h3bc38de1),
	.w7(32'h3afe995b),
	.w8(32'h3b7ec5d7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985bb06),
	.w1(32'h3b7ef6cf),
	.w2(32'hba0eafdc),
	.w3(32'hba0abbe3),
	.w4(32'h3bb78513),
	.w5(32'hb992b388),
	.w6(32'h3be4b315),
	.w7(32'hb9f21fb6),
	.w8(32'hbac82437),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule