module layer_10_featuremap_303(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b1da3),
	.w1(32'hba954e50),
	.w2(32'h3960ab5a),
	.w3(32'hba5eabd6),
	.w4(32'h37fedb1f),
	.w5(32'hb9d3607a),
	.w6(32'hbac59f0d),
	.w7(32'hb98d824b),
	.w8(32'hb852d538),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add0b1c),
	.w1(32'h39ae2263),
	.w2(32'h3a97b309),
	.w3(32'h3a4613e8),
	.w4(32'hb9d2b1ee),
	.w5(32'h39cd3e42),
	.w6(32'h3ad4af9f),
	.w7(32'h395f3aa9),
	.w8(32'h3a65f1d8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df44a2),
	.w1(32'h39ba8e9a),
	.w2(32'h3995b42b),
	.w3(32'h392a8bb3),
	.w4(32'h39ee84c9),
	.w5(32'hba263683),
	.w6(32'hba08cc23),
	.w7(32'hba06cc5b),
	.w8(32'hba141ee9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c521f),
	.w1(32'hb9ba6bcb),
	.w2(32'hb9148660),
	.w3(32'hb8fb4afd),
	.w4(32'hb9156451),
	.w5(32'hbac73fc5),
	.w6(32'h39a9744f),
	.w7(32'hb8bcd1e0),
	.w8(32'hbab3962c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada4ee3),
	.w1(32'hbaf0204c),
	.w2(32'hb9dde22c),
	.w3(32'hbb2e9652),
	.w4(32'hbaf3a6f6),
	.w5(32'hba644cee),
	.w6(32'hba459046),
	.w7(32'hba89f19f),
	.w8(32'hba8933ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10fd42),
	.w1(32'hb9a4077e),
	.w2(32'h397a0c29),
	.w3(32'hba21beee),
	.w4(32'hb9432eaa),
	.w5(32'hb9dec836),
	.w6(32'hba27f3d7),
	.w7(32'hb90dab85),
	.w8(32'hb924ccac),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980f2d9),
	.w1(32'h39da33be),
	.w2(32'h3b4b335e),
	.w3(32'hb82961e2),
	.w4(32'h3b334ee1),
	.w5(32'h3b6f6514),
	.w6(32'h39c27a6e),
	.w7(32'h3b0d2bd9),
	.w8(32'h3b19c74f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c6147),
	.w1(32'h3b0e9372),
	.w2(32'h3ad0554c),
	.w3(32'h3bd329f5),
	.w4(32'h3b835977),
	.w5(32'h3a966ef6),
	.w6(32'h3bc8ff20),
	.w7(32'h3b49537b),
	.w8(32'h3b06817d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a454377),
	.w1(32'h38b2aba2),
	.w2(32'h3a4f457a),
	.w3(32'h3a32937a),
	.w4(32'h3a4a048b),
	.w5(32'h39c0e78e),
	.w6(32'h3a3da744),
	.w7(32'h3a7b9a22),
	.w8(32'h3a71b788),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b879f14),
	.w1(32'h3b19a676),
	.w2(32'h3bf6cb13),
	.w3(32'h3b891c58),
	.w4(32'h3a79de14),
	.w5(32'h3bae6bbb),
	.w6(32'h3bbcd6e4),
	.w7(32'h3b024e53),
	.w8(32'h3bc09942),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1691ee),
	.w1(32'hb9f10160),
	.w2(32'hb99d07f8),
	.w3(32'hb96dfb92),
	.w4(32'hb90d2367),
	.w5(32'h3a38d598),
	.w6(32'h39918485),
	.w7(32'hb9cdaa76),
	.w8(32'hb8e8d663),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff236c),
	.w1(32'hbaac22c8),
	.w2(32'h3b3bf992),
	.w3(32'h3ab78744),
	.w4(32'hba9193b4),
	.w5(32'h3b081afa),
	.w6(32'h39d1f99b),
	.w7(32'hbb138fea),
	.w8(32'h3a23c405),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58acdc),
	.w1(32'h3a8da030),
	.w2(32'h3b313cfb),
	.w3(32'h3b096383),
	.w4(32'hba35480d),
	.w5(32'h3b2bcc28),
	.w6(32'h3ad7434c),
	.w7(32'hb798124f),
	.w8(32'h3b6aab11),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969af81),
	.w1(32'h3a076425),
	.w2(32'h3a1cf40c),
	.w3(32'h39f0e397),
	.w4(32'h3a951fe7),
	.w5(32'h3a1b9db5),
	.w6(32'hba3e8ea9),
	.w7(32'hb7dfa336),
	.w8(32'h39c0da02),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa780bb),
	.w1(32'hba0f5f38),
	.w2(32'h3b3cecb7),
	.w3(32'h39ada729),
	.w4(32'hba93fc12),
	.w5(32'h3a1295e1),
	.w6(32'h3b0aa782),
	.w7(32'h38a60f04),
	.w8(32'h3ae15074),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56ff5c),
	.w1(32'h3b05636c),
	.w2(32'h3b888ba7),
	.w3(32'h3b297c2a),
	.w4(32'h39d18fbf),
	.w5(32'h3b05cf8f),
	.w6(32'h3b5a786d),
	.w7(32'h3b25c2d1),
	.w8(32'h3b77fe32),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c779ca),
	.w1(32'hba742767),
	.w2(32'hb9a0b06f),
	.w3(32'h3989dd44),
	.w4(32'hba3ea357),
	.w5(32'hb8a674ce),
	.w6(32'h3978acaf),
	.w7(32'hba5442bf),
	.w8(32'hb9d4087b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e9143),
	.w1(32'h3b26d7e6),
	.w2(32'h3b303c2b),
	.w3(32'h3bc3cca1),
	.w4(32'h3b59a3c2),
	.w5(32'h3baeef6d),
	.w6(32'h3b95992a),
	.w7(32'h3b245a68),
	.w8(32'h3b916c91),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c544a),
	.w1(32'h3ac78d38),
	.w2(32'h3aa350d8),
	.w3(32'h3b59d891),
	.w4(32'h3b41b48f),
	.w5(32'h3b516c3b),
	.w6(32'h3b1b76bd),
	.w7(32'h3af60727),
	.w8(32'h3b367f0e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab29241),
	.w1(32'hb98ca401),
	.w2(32'h3a12e72f),
	.w3(32'h37ca1e81),
	.w4(32'hba34f4fa),
	.w5(32'hba0b155d),
	.w6(32'hb92aca93),
	.w7(32'hb900e86f),
	.w8(32'hba839ff9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed50d0),
	.w1(32'hba484906),
	.w2(32'h37baa287),
	.w3(32'hba489992),
	.w4(32'h38306f2a),
	.w5(32'hb9824fa4),
	.w6(32'hbab0656f),
	.w7(32'hba114341),
	.w8(32'hb8120c1f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57c8d7),
	.w1(32'hbaca9019),
	.w2(32'hb8f7725f),
	.w3(32'hba240e41),
	.w4(32'hbaacf82d),
	.w5(32'h3a0a9e06),
	.w6(32'hb958353f),
	.w7(32'hbae29418),
	.w8(32'hb97ad6fc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c509),
	.w1(32'h38611ae0),
	.w2(32'h3ba5a0f0),
	.w3(32'h3ba81eef),
	.w4(32'h3afc54b6),
	.w5(32'h3c057daa),
	.w6(32'h3bf3bbd5),
	.w7(32'h3bc1b79b),
	.w8(32'h3c559804),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b856989),
	.w1(32'h3a859b98),
	.w2(32'h3bc984e0),
	.w3(32'h3ae7300a),
	.w4(32'hba624c2a),
	.w5(32'h3bbb2468),
	.w6(32'h3b7232f3),
	.w7(32'hb9a6058d),
	.w8(32'h3bb5a044),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b453a07),
	.w1(32'hbb453ad7),
	.w2(32'h3b3fb00e),
	.w3(32'h3b0b7679),
	.w4(32'hbb59fbe7),
	.w5(32'h3aad2cf5),
	.w6(32'h3b92553d),
	.w7(32'hbab507db),
	.w8(32'h3b66ba2c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba7aa1),
	.w1(32'hb87aec2e),
	.w2(32'h39cf0eb0),
	.w3(32'hba0f58ca),
	.w4(32'h3969819e),
	.w5(32'h3a1e17cf),
	.w6(32'hba104f89),
	.w7(32'h3a8e02c7),
	.w8(32'h39b9d03f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbcb3a),
	.w1(32'hba4060b9),
	.w2(32'hb971ebfa),
	.w3(32'hba63567e),
	.w4(32'hb9b837cf),
	.w5(32'hbaa279c2),
	.w6(32'hbab5c9f0),
	.w7(32'hba0833d3),
	.w8(32'hbaf36d44),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db2c8),
	.w1(32'hbba7f963),
	.w2(32'hbab837bd),
	.w3(32'hba52764c),
	.w4(32'hbb2e116e),
	.w5(32'hba825549),
	.w6(32'hbb2e3171),
	.w7(32'hbb861233),
	.w8(32'hbb7afc92),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80d136),
	.w1(32'hbb3587e6),
	.w2(32'hba41dd97),
	.w3(32'hba673fde),
	.w4(32'hbb3b8b1d),
	.w5(32'hba93daa8),
	.w6(32'hba875cef),
	.w7(32'hbb80cfed),
	.w8(32'hbb5b86bb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadffe5),
	.w1(32'hbb15ecac),
	.w2(32'h3b051d06),
	.w3(32'h3b802156),
	.w4(32'hba8a6aca),
	.w5(32'h3ad61e4b),
	.w6(32'h3b5ce251),
	.w7(32'hb9070f12),
	.w8(32'h3b4deac3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac6cfa),
	.w1(32'h38a9c0d6),
	.w2(32'hb999d812),
	.w3(32'h39c66743),
	.w4(32'hb89adaa2),
	.w5(32'h3907c2ad),
	.w6(32'h3ab3b434),
	.w7(32'hb90dbce3),
	.w8(32'h38b1d790),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25ebd2),
	.w1(32'h3a8f82d6),
	.w2(32'h3a00d5e4),
	.w3(32'h39bdb874),
	.w4(32'h396c848e),
	.w5(32'h39e1e12a),
	.w6(32'h3a6c36cb),
	.w7(32'hb8c6ee37),
	.w8(32'hb999c919),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa59420),
	.w1(32'h3a505660),
	.w2(32'h3b3d7426),
	.w3(32'h3b2ecea4),
	.w4(32'h3a8bf14d),
	.w5(32'h3af8e126),
	.w6(32'h3b13e47e),
	.w7(32'h3a99c7fb),
	.w8(32'h3ae5e50a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e63ae),
	.w1(32'h39a96850),
	.w2(32'h3a57f0fc),
	.w3(32'h3b133180),
	.w4(32'hb8da5cb7),
	.w5(32'h3a9b49a1),
	.w6(32'h3b2ad5a7),
	.w7(32'h3ab5effa),
	.w8(32'h3ab78580),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7a60e),
	.w1(32'hb9321669),
	.w2(32'h399bbc0e),
	.w3(32'h3a9727ec),
	.w4(32'h3adff1e7),
	.w5(32'h39bf0b09),
	.w6(32'hb92d06b0),
	.w7(32'h3a33cc31),
	.w8(32'h37d87e01),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fd11d),
	.w1(32'h3988dc5a),
	.w2(32'h3ac1026a),
	.w3(32'h3a579040),
	.w4(32'h3a9d0ba3),
	.w5(32'h3ae32a33),
	.w6(32'h3a4af988),
	.w7(32'h3a092591),
	.w8(32'h385020ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef4a22),
	.w1(32'hbabafd1f),
	.w2(32'h3b6af5c8),
	.w3(32'h3abd7c83),
	.w4(32'h3697bc8d),
	.w5(32'h3b711306),
	.w6(32'hbb92d68f),
	.w7(32'hbb572613),
	.w8(32'h3b83b518),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86b76e),
	.w1(32'hbbd161de),
	.w2(32'h3a2719d2),
	.w3(32'h3b7ae888),
	.w4(32'hbbd1658d),
	.w5(32'hb86d1e80),
	.w6(32'h3bbd6f6f),
	.w7(32'hbbb3a663),
	.w8(32'h3a7b2430),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05e907),
	.w1(32'hbc37c79e),
	.w2(32'hbb6befc5),
	.w3(32'h3b2d9ae8),
	.w4(32'hbbbef93a),
	.w5(32'h3a818cec),
	.w6(32'h3bb121d1),
	.w7(32'hbb265518),
	.w8(32'h3b573cc8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7d510),
	.w1(32'hba2ffb24),
	.w2(32'h3969806f),
	.w3(32'h3a7546d0),
	.w4(32'hba437ba1),
	.w5(32'h397883c5),
	.w6(32'h3b10dc75),
	.w7(32'h3a1a4759),
	.w8(32'h3a944cab),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a968a2d),
	.w1(32'h3aa1b194),
	.w2(32'h3a1bd0dc),
	.w3(32'h3a98aab9),
	.w4(32'h3a639d25),
	.w5(32'h3a1c903c),
	.w6(32'h3a0da15c),
	.w7(32'h3a8b902d),
	.w8(32'h3969e438),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba687f5e),
	.w1(32'hba481a08),
	.w2(32'hb91cc6c9),
	.w3(32'hba5db926),
	.w4(32'hb9b27540),
	.w5(32'h3a2964fe),
	.w6(32'hba4e689a),
	.w7(32'hb758b3f1),
	.w8(32'h3a11be8f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d9d0e),
	.w1(32'h3a36edb7),
	.w2(32'h3a7c3637),
	.w3(32'h3a91cd97),
	.w4(32'h39ef1f73),
	.w5(32'h3a398ae0),
	.w6(32'h3a9f1f85),
	.w7(32'h3a9fe8d1),
	.w8(32'h380e39e1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beede8a),
	.w1(32'h3bd3697d),
	.w2(32'h3bc02a7b),
	.w3(32'h3bf0def1),
	.w4(32'h3ba6bc96),
	.w5(32'h3b011be8),
	.w6(32'h3be5c722),
	.w7(32'h3bd200ec),
	.w8(32'h3baad23c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b564287),
	.w1(32'hba8c2500),
	.w2(32'h3b97a830),
	.w3(32'h3b16071e),
	.w4(32'hbb322add),
	.w5(32'h3b7fba22),
	.w6(32'h3b14e7e1),
	.w7(32'hbac9eefc),
	.w8(32'h3bc2e790),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba82127),
	.w1(32'h3a9b5dc0),
	.w2(32'h3be28ca6),
	.w3(32'h3b14208e),
	.w4(32'hbad5edbe),
	.w5(32'h3b93f57b),
	.w6(32'h3bcf28a0),
	.w7(32'h3adfccb6),
	.w8(32'h3bca8826),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd66eab),
	.w1(32'h3b39683b),
	.w2(32'h3bf61e83),
	.w3(32'h3bcc4c2d),
	.w4(32'h3b03c72b),
	.w5(32'h3bc7cd98),
	.w6(32'h3bdd386b),
	.w7(32'h3b819de4),
	.w8(32'h3c01fbf6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af20371),
	.w1(32'h3b587dde),
	.w2(32'h3b6f117a),
	.w3(32'h3b94677a),
	.w4(32'h3bd1fe3b),
	.w5(32'h3bf0ae98),
	.w6(32'h3b7beb4c),
	.w7(32'h3bb94dfd),
	.w8(32'h3bf1f085),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52626f),
	.w1(32'h3a47a84e),
	.w2(32'h3a821279),
	.w3(32'h38a5b2a1),
	.w4(32'h3a1f26af),
	.w5(32'hba0aec48),
	.w6(32'h37a2a0cd),
	.w7(32'hb8d73db4),
	.w8(32'h3846c485),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa835b9),
	.w1(32'hb9cacc28),
	.w2(32'h3aa7e5ac),
	.w3(32'hba3b256f),
	.w4(32'h39eac4af),
	.w5(32'h3943bce5),
	.w6(32'h393649d8),
	.w7(32'h3ac72c73),
	.w8(32'h3ac8a845),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb180b42),
	.w1(32'hbaed3b5e),
	.w2(32'hb924f060),
	.w3(32'hbb5a4f02),
	.w4(32'hba166424),
	.w5(32'h3913f1aa),
	.w6(32'hbb359766),
	.w7(32'hba0e1b3f),
	.w8(32'h3a3fe3f4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27c97c),
	.w1(32'h3a974a6f),
	.w2(32'h3b510185),
	.w3(32'h3a95d39e),
	.w4(32'hba150b56),
	.w5(32'h3afe8b86),
	.w6(32'h3af31796),
	.w7(32'h3a03aff9),
	.w8(32'h3b2754f0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad667f8),
	.w1(32'h3abba1c2),
	.w2(32'h3a80ec64),
	.w3(32'h39ab904e),
	.w4(32'hb908a2ae),
	.w5(32'h3abda810),
	.w6(32'h3a904b1c),
	.w7(32'h3a4bc91a),
	.w8(32'h3a9ae8ec),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8de9d6),
	.w1(32'h3b0ed7d9),
	.w2(32'h3bb32f3b),
	.w3(32'h3b89a304),
	.w4(32'h3b5d3624),
	.w5(32'h3bc94456),
	.w6(32'h3a9c6007),
	.w7(32'h3ab08169),
	.w8(32'h3b90c16c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cea30d),
	.w1(32'hb983cee2),
	.w2(32'h3a4c5626),
	.w3(32'h3912bea9),
	.w4(32'hb9705adb),
	.w5(32'h3a283b78),
	.w6(32'hb81af0bc),
	.w7(32'hb9af4394),
	.w8(32'hb9146cd1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920f764),
	.w1(32'hb9efb193),
	.w2(32'h39eb982c),
	.w3(32'hb9c781eb),
	.w4(32'h3963f4c5),
	.w5(32'h3a04e37b),
	.w6(32'hba475b80),
	.w7(32'hb9c8f9f4),
	.w8(32'h39db5e08),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c9656),
	.w1(32'hb9685566),
	.w2(32'hb851b4b2),
	.w3(32'h39cdb0f6),
	.w4(32'h39c6d7c9),
	.w5(32'hb830b720),
	.w6(32'hb91ac25d),
	.w7(32'h3832a0d5),
	.w8(32'hba0eee78),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9278ac2),
	.w1(32'hb9e5aab2),
	.w2(32'hb8fd8dba),
	.w3(32'hb9afc477),
	.w4(32'hba4bb3f8),
	.w5(32'hb9b293f9),
	.w6(32'hba3da5a2),
	.w7(32'h387640e8),
	.w8(32'hb92fc6b5),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a28da),
	.w1(32'hbb096603),
	.w2(32'hba6dcdcc),
	.w3(32'hba1ee10c),
	.w4(32'hba885fb7),
	.w5(32'h3a05e3d4),
	.w6(32'h38df947a),
	.w7(32'hb98335ff),
	.w8(32'h3a7357e2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82a64f),
	.w1(32'h3ae3d3c0),
	.w2(32'h3ab956b9),
	.w3(32'h3ab1bc0e),
	.w4(32'h3aa5cd9a),
	.w5(32'h391e074f),
	.w6(32'h3b1a97e7),
	.w7(32'h3acc2cbb),
	.w8(32'h38c4ccc6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16104d),
	.w1(32'h3a3a0acd),
	.w2(32'h3ad2c4a5),
	.w3(32'h3ac1c04a),
	.w4(32'h3a056ec7),
	.w5(32'h3a62776b),
	.w6(32'h3b00cddf),
	.w7(32'h3a77ede0),
	.w8(32'h3a223b32),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0143b3),
	.w1(32'h3a29f526),
	.w2(32'h3a993456),
	.w3(32'h3ad29563),
	.w4(32'h3a9cfda2),
	.w5(32'h3a863697),
	.w6(32'h3af9da76),
	.w7(32'h3b0b7004),
	.w8(32'h3a4a746d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b60e55),
	.w1(32'hba21c339),
	.w2(32'hb91efcca),
	.w3(32'h3738f2c1),
	.w4(32'h3a089b36),
	.w5(32'h3a2aaf52),
	.w6(32'hb98612ff),
	.w7(32'hb8c0d3bd),
	.w8(32'h387a3796),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398776c0),
	.w1(32'hb9d261eb),
	.w2(32'h39524e5c),
	.w3(32'h39c660da),
	.w4(32'h3a549c8b),
	.w5(32'h399dee2c),
	.w6(32'hba124451),
	.w7(32'h3a00b6cb),
	.w8(32'hb8a7b892),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f616c),
	.w1(32'hb8dd5128),
	.w2(32'h395a3289),
	.w3(32'h3a4a4ff7),
	.w4(32'h3aad3728),
	.w5(32'hba07dfe9),
	.w6(32'hb7105567),
	.w7(32'h3a24f124),
	.w8(32'h395e524c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a417b81),
	.w1(32'h3a6ab799),
	.w2(32'h3a01763c),
	.w3(32'hba3cfaea),
	.w4(32'hb9b46591),
	.w5(32'hba19223d),
	.w6(32'h3a623c88),
	.w7(32'h39dfdd84),
	.w8(32'hba1d0d97),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a2b2a),
	.w1(32'h3aa010e2),
	.w2(32'h3b03bc29),
	.w3(32'h3b77e515),
	.w4(32'h3b4d7a84),
	.w5(32'h3b38560d),
	.w6(32'h3aa317a2),
	.w7(32'h3adea18d),
	.w8(32'h3a7a599f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40c302),
	.w1(32'hb9f4dfdc),
	.w2(32'h3bc606da),
	.w3(32'hba24ea57),
	.w4(32'hb9384e47),
	.w5(32'h3bc18c80),
	.w6(32'h3a650d6a),
	.w7(32'hba8cbfb1),
	.w8(32'h3ba9674f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff5d6b),
	.w1(32'hbb31998f),
	.w2(32'h3b7e6980),
	.w3(32'h38eb194a),
	.w4(32'hbb227a98),
	.w5(32'h3b5b7a97),
	.w6(32'h3a95a05a),
	.w7(32'hbae0b9d4),
	.w8(32'h3b3b76df),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b708935),
	.w1(32'hbb6c17fd),
	.w2(32'h3c16db55),
	.w3(32'h3b38aa29),
	.w4(32'hbbd3f288),
	.w5(32'h3b245255),
	.w6(32'h3bbd2832),
	.w7(32'hbb557d75),
	.w8(32'h3baf9a39),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982133e),
	.w1(32'hb9dea514),
	.w2(32'h3979719f),
	.w3(32'hb9c9a7df),
	.w4(32'hb9371366),
	.w5(32'hb90326db),
	.w6(32'hba4560b2),
	.w7(32'h399ff0fc),
	.w8(32'hba5f479f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3927dd3c),
	.w1(32'h39abec85),
	.w2(32'hb924411f),
	.w3(32'hb94509b5),
	.w4(32'h3970c284),
	.w5(32'hb9622711),
	.w6(32'h3a26be10),
	.w7(32'h3a0f9627),
	.w8(32'h3a892f8f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a989eec),
	.w1(32'h3ad25666),
	.w2(32'h3a35e072),
	.w3(32'hb9bb239f),
	.w4(32'h39b2c304),
	.w5(32'h399eb0bf),
	.w6(32'h3b31308e),
	.w7(32'h3b03399d),
	.w8(32'hb8c798b1),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c1a6e),
	.w1(32'hb967e3b8),
	.w2(32'hba771d1b),
	.w3(32'h3afe6c0b),
	.w4(32'h3a983f9a),
	.w5(32'h38a0e895),
	.w6(32'h3aeb8b30),
	.w7(32'h39cb6129),
	.w8(32'hba963f92),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47cff2),
	.w1(32'hba02c732),
	.w2(32'hb9373bd2),
	.w3(32'hb9b983d6),
	.w4(32'hb9b8d14c),
	.w5(32'h3a501309),
	.w6(32'hbaaec8cd),
	.w7(32'hba68f2d1),
	.w8(32'h3a0eae59),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6d57b),
	.w1(32'h38920472),
	.w2(32'h390b74cc),
	.w3(32'h3b599271),
	.w4(32'h3b08c6b8),
	.w5(32'h3af4fb2d),
	.w6(32'h3abaaf19),
	.w7(32'h39f54f52),
	.w8(32'h3aaffe77),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf82969),
	.w1(32'h3b5d6624),
	.w2(32'h3b143613),
	.w3(32'h3b980d53),
	.w4(32'h3afccf87),
	.w5(32'h3b430cdb),
	.w6(32'h3baa5784),
	.w7(32'h3b4ed5cb),
	.w8(32'h3ba4a29d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e8708),
	.w1(32'h3a8715f3),
	.w2(32'h3b121341),
	.w3(32'h3b566437),
	.w4(32'hba5a4771),
	.w5(32'h3aa4fde0),
	.w6(32'h3b68c432),
	.w7(32'h3a64a524),
	.w8(32'h3b10b5bb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4aa09),
	.w1(32'h3a19149d),
	.w2(32'h3af41065),
	.w3(32'h3ab3ed63),
	.w4(32'hb9cdedbd),
	.w5(32'h3a866b47),
	.w6(32'h3b17e8ed),
	.w7(32'hb99d2467),
	.w8(32'h3a86a050),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1db0c5),
	.w1(32'hb9e5797b),
	.w2(32'h3adfdb03),
	.w3(32'h391a9dac),
	.w4(32'h3a3670c9),
	.w5(32'h3b72ec0c),
	.w6(32'hba19b0e4),
	.w7(32'hb9c292f1),
	.w8(32'h3b200840),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ecbc3),
	.w1(32'h3a41eddc),
	.w2(32'h3b38a35e),
	.w3(32'h3afbea24),
	.w4(32'h38067868),
	.w5(32'h3ad3b051),
	.w6(32'h3b03dedf),
	.w7(32'h39d43921),
	.w8(32'h3af28a4a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8456c2),
	.w1(32'h3a563f3e),
	.w2(32'h3a9d5352),
	.w3(32'h3b3282b5),
	.w4(32'h3b1b6a5b),
	.w5(32'h3b49a881),
	.w6(32'h3b16d255),
	.w7(32'h3ac3da99),
	.w8(32'h3b2bea8f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c644b),
	.w1(32'h39ddd713),
	.w2(32'h39b80d2a),
	.w3(32'h38f295dd),
	.w4(32'h3a1f57ff),
	.w5(32'h3a5e9307),
	.w6(32'h399c31bf),
	.w7(32'h3966111d),
	.w8(32'h3a5c8289),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cd471),
	.w1(32'h3aa94b26),
	.w2(32'h3a7e037f),
	.w3(32'h3a56f70c),
	.w4(32'h3a19cab8),
	.w5(32'h39c09dbc),
	.w6(32'h3ab8a0e6),
	.w7(32'h3a102e11),
	.w8(32'h394af428),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a135083),
	.w1(32'h3a4d453b),
	.w2(32'h3a029b5e),
	.w3(32'h38cd6cd7),
	.w4(32'h39b114ad),
	.w5(32'hba097cf7),
	.w6(32'h393ca8f7),
	.w7(32'h381a8256),
	.w8(32'h390ba7da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bdd62),
	.w1(32'hb9fd3c32),
	.w2(32'h399915e8),
	.w3(32'hba2d8e46),
	.w4(32'hba0f00c2),
	.w5(32'h3a1c7022),
	.w6(32'h3a65e208),
	.w7(32'h39f3b62f),
	.w8(32'h394ea132),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b863336),
	.w1(32'hba88e1c4),
	.w2(32'h3add8464),
	.w3(32'h3b570869),
	.w4(32'hbaa8d22d),
	.w5(32'hb9e4d106),
	.w6(32'h3b451981),
	.w7(32'hb993e4c7),
	.w8(32'h3a9dbb69),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39309ada),
	.w1(32'hba329bc0),
	.w2(32'h38e59d9b),
	.w3(32'hba3bb5ae),
	.w4(32'hbabd94de),
	.w5(32'hba37df74),
	.w6(32'h3a865c5f),
	.w7(32'hb91334b8),
	.w8(32'hba4c6c9d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7bf46),
	.w1(32'h3a221f77),
	.w2(32'h3b34d107),
	.w3(32'h39947627),
	.w4(32'h395fdd0b),
	.w5(32'h3af9f464),
	.w6(32'h3a6513c0),
	.w7(32'h37bd6c3d),
	.w8(32'h3af814bb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9acc83),
	.w1(32'h3ad69ff2),
	.w2(32'h3a4fcea9),
	.w3(32'h3bb8172d),
	.w4(32'h3a3ece81),
	.w5(32'h3ae72841),
	.w6(32'h3bbfe1fb),
	.w7(32'h3b10894d),
	.w8(32'h3b26ada0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2589a6),
	.w1(32'hbb60f168),
	.w2(32'hba1e955d),
	.w3(32'h3972003f),
	.w4(32'hbb40684c),
	.w5(32'h38d92e80),
	.w6(32'h399ca8fc),
	.w7(32'hbb654728),
	.w8(32'hb92b25ef),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add96e4),
	.w1(32'h39726304),
	.w2(32'h3ac7c952),
	.w3(32'h3b743f59),
	.w4(32'h3ac8633e),
	.w5(32'h3b59b8ef),
	.w6(32'h3a838816),
	.w7(32'h3ab2ba58),
	.w8(32'h3b73b9c4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b9129),
	.w1(32'hbb587aec),
	.w2(32'h3ac0dd48),
	.w3(32'hba8ad8aa),
	.w4(32'hbace5b54),
	.w5(32'h3adaec7f),
	.w6(32'hbaffa121),
	.w7(32'hbb34537a),
	.w8(32'hba9f3900),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55dea9),
	.w1(32'h3ab2eead),
	.w2(32'h3b9c2708),
	.w3(32'h3b2d9d33),
	.w4(32'h350c9da4),
	.w5(32'h3b740661),
	.w6(32'h3b415576),
	.w7(32'h3a4b4ffa),
	.w8(32'h3b950784),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78bdb7),
	.w1(32'h392fe3f9),
	.w2(32'h3b47f9fe),
	.w3(32'h39c4ceb9),
	.w4(32'hba43eb5d),
	.w5(32'h3af9dfde),
	.w6(32'h3a3a3df9),
	.w7(32'h3a5ff6fc),
	.w8(32'h3afdbadc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44ec66),
	.w1(32'hba449706),
	.w2(32'h3b4d9af2),
	.w3(32'h3b030060),
	.w4(32'hbb08fdd1),
	.w5(32'h3b44423c),
	.w6(32'h3b44d258),
	.w7(32'hb8803d60),
	.w8(32'h3b4d01e6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e8196),
	.w1(32'hb93dfae1),
	.w2(32'hbadd10ee),
	.w3(32'hb9f1fac2),
	.w4(32'h38903bc7),
	.w5(32'hba2adb26),
	.w6(32'h398b975d),
	.w7(32'hba008b2b),
	.w8(32'h3a014c5f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab42c50),
	.w1(32'h39f1146b),
	.w2(32'h3ba3e901),
	.w3(32'h399f8505),
	.w4(32'h38e6d46f),
	.w5(32'h3b7c39e6),
	.w6(32'h3b4b2f61),
	.w7(32'h3b7c3b9f),
	.w8(32'h3be85139),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01df80),
	.w1(32'hbb3189a3),
	.w2(32'h3b30e33b),
	.w3(32'hba9a0252),
	.w4(32'hbaf854d8),
	.w5(32'h3a1b5a97),
	.w6(32'hbaa818ef),
	.w7(32'h3a7a324b),
	.w8(32'h3b862d07),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b616b96),
	.w1(32'hb9ef52c8),
	.w2(32'h3bcdb89c),
	.w3(32'hbaaee767),
	.w4(32'hbaa9a855),
	.w5(32'h3bae271a),
	.w6(32'hb9f10fcc),
	.w7(32'hba6b10d3),
	.w8(32'h3bb7ba59),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4945b),
	.w1(32'hbb34de37),
	.w2(32'h3b56bda5),
	.w3(32'h3b907994),
	.w4(32'hbbdae55e),
	.w5(32'h398761fb),
	.w6(32'h3c081068),
	.w7(32'h3a1e0e27),
	.w8(32'h3bd40291),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15da23),
	.w1(32'h3aba86cc),
	.w2(32'h3bb27ad3),
	.w3(32'h3ae5fe43),
	.w4(32'hbae2dc6a),
	.w5(32'h3b76d0ab),
	.w6(32'h3aaeb5cc),
	.w7(32'h3a900cba),
	.w8(32'h3bc5846f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84cde4),
	.w1(32'h39b30419),
	.w2(32'h3b9c2a85),
	.w3(32'h3b0bcb2b),
	.w4(32'h3b110c4e),
	.w5(32'h3b5f2279),
	.w6(32'hbadfb578),
	.w7(32'h39a47b39),
	.w8(32'h3bb3553d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b56bd),
	.w1(32'hba137a85),
	.w2(32'h3a4904df),
	.w3(32'hba158623),
	.w4(32'hbad0908a),
	.w5(32'h39ff9957),
	.w6(32'h39e24d44),
	.w7(32'h3b2737ad),
	.w8(32'h3ac3e92d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0b90d),
	.w1(32'h3ab62b3f),
	.w2(32'h3b46b3ca),
	.w3(32'h3bbb043c),
	.w4(32'h3a4c5c79),
	.w5(32'h3b768a83),
	.w6(32'h3a76bcc9),
	.w7(32'hbb86bb8e),
	.w8(32'hbafa8dfb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e28ae),
	.w1(32'h3b877c2d),
	.w2(32'h3bc4f6dd),
	.w3(32'hb9fd52db),
	.w4(32'h3a920074),
	.w5(32'h3b5a6b16),
	.w6(32'hb8d47580),
	.w7(32'h3b56cff4),
	.w8(32'h3b488bf7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f0c4f),
	.w1(32'hbb0c4481),
	.w2(32'h3a8fb39b),
	.w3(32'h3a29484f),
	.w4(32'h384e5a83),
	.w5(32'h3a65123e),
	.w6(32'hbad6cb1f),
	.w7(32'hbb16f189),
	.w8(32'h3a3439d7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af15fef),
	.w1(32'h39c7414d),
	.w2(32'h3a2950fe),
	.w3(32'h390b0e0a),
	.w4(32'h39216e47),
	.w5(32'h39b0de48),
	.w6(32'h392440fb),
	.w7(32'h391b3d0e),
	.w8(32'h3a9e68ef),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a161848),
	.w1(32'h39ee8837),
	.w2(32'hba631c1c),
	.w3(32'h3af391c0),
	.w4(32'h3a9eeedb),
	.w5(32'h3aa13258),
	.w6(32'h3b852f03),
	.w7(32'h3ba47d73),
	.w8(32'h3bc82807),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25a017),
	.w1(32'hbb1de6f7),
	.w2(32'h3abde2ef),
	.w3(32'hbb11ac34),
	.w4(32'hbb7c309e),
	.w5(32'h3b69364e),
	.w6(32'hba06758b),
	.w7(32'hbaeaf36f),
	.w8(32'h3b9e362f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b669ac0),
	.w1(32'h3b2b2edd),
	.w2(32'h3b92687c),
	.w3(32'h3b5e6f2b),
	.w4(32'h3aeebf6d),
	.w5(32'h3ae58f6f),
	.w6(32'h3b686859),
	.w7(32'h3b68092a),
	.w8(32'h3b9eaad5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a615a),
	.w1(32'h3a2e2163),
	.w2(32'h3b4e6aa2),
	.w3(32'h3b1ee3e2),
	.w4(32'hba5bc1ed),
	.w5(32'h3956f39a),
	.w6(32'h3b8f37ba),
	.w7(32'h3ac3fad6),
	.w8(32'h3b3f32be),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a566713),
	.w1(32'hbaccfe98),
	.w2(32'hb9af6425),
	.w3(32'h3a5a19ad),
	.w4(32'hbb5c4e07),
	.w5(32'h3aa8b059),
	.w6(32'h3a890b0f),
	.w7(32'hbb563676),
	.w8(32'h3983aa94),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30b56d),
	.w1(32'h3b44031e),
	.w2(32'h3b7ad702),
	.w3(32'h3af92ba7),
	.w4(32'h3ab1f5bb),
	.w5(32'h3abdf54f),
	.w6(32'h3b498193),
	.w7(32'h3b2243c6),
	.w8(32'hba8c6d21),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c1945),
	.w1(32'h3a5b3092),
	.w2(32'h3a6d92b2),
	.w3(32'h39d78c03),
	.w4(32'hb8f5888f),
	.w5(32'h3ad7b6bb),
	.w6(32'h3b00baee),
	.w7(32'hb97b3bb5),
	.w8(32'h3b37a93a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdb216),
	.w1(32'h3b2739e8),
	.w2(32'h3a2a2767),
	.w3(32'h3afbd97f),
	.w4(32'h3a004e47),
	.w5(32'h39ed09c8),
	.w6(32'h3a8d0e0f),
	.w7(32'h3a8462dd),
	.w8(32'h3a885d6e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a695708),
	.w1(32'h3a36dd0a),
	.w2(32'h38e3fadd),
	.w3(32'h39c13feb),
	.w4(32'hba287852),
	.w5(32'hb9e39757),
	.w6(32'h3a419d1d),
	.w7(32'hb9aa8019),
	.w8(32'hbae7a85c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdf77d),
	.w1(32'hbacfd6fe),
	.w2(32'hbad031d7),
	.w3(32'hba862c31),
	.w4(32'hbadcffce),
	.w5(32'hb91de0b3),
	.w6(32'hba31e9ee),
	.w7(32'hba5bb0ba),
	.w8(32'hb9a38166),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87dc1fa),
	.w1(32'hb94922d5),
	.w2(32'h3ab28656),
	.w3(32'hbabfd6e1),
	.w4(32'hb7b34ffc),
	.w5(32'hb8b474d4),
	.w6(32'hba54caa5),
	.w7(32'h3ae5887e),
	.w8(32'hba6b7e55),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa190d0),
	.w1(32'h39277b12),
	.w2(32'h3b6dc84e),
	.w3(32'h3a31067b),
	.w4(32'hba79c8a5),
	.w5(32'h39df4939),
	.w6(32'h39ce7560),
	.w7(32'h370f343f),
	.w8(32'h3aa4e6a9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd4150),
	.w1(32'h3a17d448),
	.w2(32'h3a757e68),
	.w3(32'h3a5a5809),
	.w4(32'hb83683b2),
	.w5(32'hb9b67e28),
	.w6(32'h38a722db),
	.w7(32'hba182da3),
	.w8(32'hbad530b6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d23023),
	.w1(32'h3b5a73c4),
	.w2(32'h3b84edc7),
	.w3(32'h3b57951a),
	.w4(32'h3b1fafbc),
	.w5(32'hb9db2fa6),
	.w6(32'h3aed1d53),
	.w7(32'h3b28d94c),
	.w8(32'h3aea0822),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac78f8f),
	.w1(32'hbb7cb600),
	.w2(32'hbad1b138),
	.w3(32'h3a013599),
	.w4(32'hba0b4ddf),
	.w5(32'hb9ec420f),
	.w6(32'h3b87dc3c),
	.w7(32'h3b4ea21d),
	.w8(32'h3a91bf8e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb134501),
	.w1(32'h3ae407c7),
	.w2(32'hb93fce68),
	.w3(32'hb98370db),
	.w4(32'hbb04ea73),
	.w5(32'hbb16b83b),
	.w6(32'hba7ccf3d),
	.w7(32'hbb4d20dc),
	.w8(32'h39cfd875),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad12f0d),
	.w1(32'hba70a9d4),
	.w2(32'hba4bc974),
	.w3(32'hbb775349),
	.w4(32'hbb094f3c),
	.w5(32'h3a3cbabf),
	.w6(32'h3aaefa17),
	.w7(32'h3b36b9ff),
	.w8(32'h385e2c1a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf9f89),
	.w1(32'hb903eb9f),
	.w2(32'hba4f93a9),
	.w3(32'hb9cc7662),
	.w4(32'hbad35e9a),
	.w5(32'hb8b31418),
	.w6(32'hba1de36c),
	.w7(32'hbab646f7),
	.w8(32'hba0b3f57),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c9518f),
	.w1(32'hb9d397d8),
	.w2(32'hb8432e32),
	.w3(32'hb8e4dd5f),
	.w4(32'hba1b145c),
	.w5(32'hbaa05924),
	.w6(32'h39b3d23f),
	.w7(32'h3a16b930),
	.w8(32'hba2dabac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b7c01),
	.w1(32'h3b5f0dfe),
	.w2(32'h3b6572a4),
	.w3(32'hb8b4c11a),
	.w4(32'h3b52cd84),
	.w5(32'h3b846a76),
	.w6(32'h3b01bb21),
	.w7(32'h3b43a1fa),
	.w8(32'h3ace1190),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b372619),
	.w1(32'h3b15a74e),
	.w2(32'h3bb71f45),
	.w3(32'h3a505469),
	.w4(32'h3a34f084),
	.w5(32'h3b7ea85b),
	.w6(32'hba027f24),
	.w7(32'h39bc598e),
	.w8(32'h3aeb6adf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202f7b),
	.w1(32'hbaf0d34e),
	.w2(32'hbad27fb0),
	.w3(32'hba275073),
	.w4(32'hba8f88dc),
	.w5(32'h39a04ecd),
	.w6(32'hbab6675a),
	.w7(32'hbab9c64e),
	.w8(32'h3afe36f2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b322589),
	.w1(32'h3ac0ec0a),
	.w2(32'h3a1e8e63),
	.w3(32'h3b97008a),
	.w4(32'h3aef82c1),
	.w5(32'h3ade62bb),
	.w6(32'h3b5d66bf),
	.w7(32'h3a7f0523),
	.w8(32'h3b1c0b6b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7110e8),
	.w1(32'hb9e0d1a0),
	.w2(32'h3a17914d),
	.w3(32'h3afe972a),
	.w4(32'h3a4381e1),
	.w5(32'hbb476033),
	.w6(32'h3b176a34),
	.w7(32'hb7ba5067),
	.w8(32'hbb0fb22b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bee70a),
	.w1(32'hba401c5e),
	.w2(32'h3b0e4cd2),
	.w3(32'hbba3e30a),
	.w4(32'hbb5a2a27),
	.w5(32'h3a8d9f26),
	.w6(32'hbb5a3e18),
	.w7(32'hbab8b4c8),
	.w8(32'h3ae89d11),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3047e5),
	.w1(32'h3a69c974),
	.w2(32'h3b44a725),
	.w3(32'h3a5bc88e),
	.w4(32'hba86500e),
	.w5(32'hb9c5fc42),
	.w6(32'h3b00e93e),
	.w7(32'h3a6ba5f4),
	.w8(32'hba87682f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25e26d),
	.w1(32'h3a9171ca),
	.w2(32'h3b8efd19),
	.w3(32'h3b356c53),
	.w4(32'h3b16506e),
	.w5(32'h3ba65e05),
	.w6(32'h3aef93aa),
	.w7(32'h3afe3309),
	.w8(32'h3ba666f7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b010b),
	.w1(32'h3a3dd5bb),
	.w2(32'h3adeb086),
	.w3(32'h38e65f93),
	.w4(32'hba9f36d2),
	.w5(32'h39f0e2d1),
	.w6(32'h3ab5c4ab),
	.w7(32'h3a2ce89b),
	.w8(32'h3b429bbc),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0359f3),
	.w1(32'h3aa0e31a),
	.w2(32'h3b6603d6),
	.w3(32'hba9ed7a5),
	.w4(32'hbb1af003),
	.w5(32'h3a0fb42a),
	.w6(32'hb887476a),
	.w7(32'hba261dd2),
	.w8(32'h3b0dc523),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ebb44),
	.w1(32'h3a624be5),
	.w2(32'h3b5e15d5),
	.w3(32'h3b1b7f98),
	.w4(32'h3abcacc1),
	.w5(32'h3b7299f9),
	.w6(32'h3b07c337),
	.w7(32'h3aaffa0f),
	.w8(32'h3b5509ba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5557cd),
	.w1(32'h3a3a82f8),
	.w2(32'h3b5169c2),
	.w3(32'h3a593b6a),
	.w4(32'h3989ced4),
	.w5(32'hb9d35930),
	.w6(32'h3b4599cf),
	.w7(32'h3b10e751),
	.w8(32'h3b2bc486),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d23e58),
	.w1(32'h3aa090a8),
	.w2(32'h3b291c03),
	.w3(32'h3a703f67),
	.w4(32'h3af1eaf7),
	.w5(32'h3b081a32),
	.w6(32'h3b0b9eeb),
	.w7(32'h3b62dfdb),
	.w8(32'h3b6d97ac),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba970db8),
	.w1(32'hba89237d),
	.w2(32'h3a4258c2),
	.w3(32'hbb2942bd),
	.w4(32'hbb329a16),
	.w5(32'h3a36cd8a),
	.w6(32'hba38b535),
	.w7(32'hb89d240a),
	.w8(32'h3a09dd0d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7608b),
	.w1(32'hbbed4c2f),
	.w2(32'h38f09e2b),
	.w3(32'h3ade906b),
	.w4(32'hbb5ea7b1),
	.w5(32'h3b85c5ef),
	.w6(32'h3a3aef28),
	.w7(32'hbae3426a),
	.w8(32'h3bcdfa46),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b403b56),
	.w1(32'h3ab73e34),
	.w2(32'h3ad50eba),
	.w3(32'h3b1911d5),
	.w4(32'h3a9d3517),
	.w5(32'h3a3d4156),
	.w6(32'h3b71e80a),
	.w7(32'h3b337e62),
	.w8(32'h3b0c4a2b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26fe7c),
	.w1(32'hbb1996ba),
	.w2(32'hba05f108),
	.w3(32'hb96a3431),
	.w4(32'h3a43632e),
	.w5(32'hb9574bdd),
	.w6(32'hb9c683e3),
	.w7(32'h3a3a2d18),
	.w8(32'h38c8385a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbb2d0),
	.w1(32'hba307e66),
	.w2(32'hba22475b),
	.w3(32'hb9f5b19f),
	.w4(32'h383b7e48),
	.w5(32'hba7ecd03),
	.w6(32'h3a52bceb),
	.w7(32'hb83e5a41),
	.w8(32'hbb072061),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3a4bb),
	.w1(32'h3b0fb8ad),
	.w2(32'h3b5458da),
	.w3(32'h39a65b00),
	.w4(32'hb89f27cf),
	.w5(32'hb9d8e1b2),
	.w6(32'h39d75e98),
	.w7(32'h3b0ea38e),
	.w8(32'hb99d2fde),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b935b40),
	.w1(32'h3ab0a1ea),
	.w2(32'h3b5b93b5),
	.w3(32'h3adbb001),
	.w4(32'hba83c8d8),
	.w5(32'h3a9ec641),
	.w6(32'h3b251c1f),
	.w7(32'h3a8a16c4),
	.w8(32'h3aaeba95),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c5d959),
	.w1(32'hbb00d1a3),
	.w2(32'hba55be96),
	.w3(32'h3aa81c3c),
	.w4(32'hbb47b1d5),
	.w5(32'hb8988186),
	.w6(32'h3b4ddd82),
	.w7(32'hba952951),
	.w8(32'h3b5f6d9a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba504e24),
	.w1(32'hbb27c279),
	.w2(32'hbab123c0),
	.w3(32'hbb189a1d),
	.w4(32'h3a67afce),
	.w5(32'h3b1a8aca),
	.w6(32'hba6ead98),
	.w7(32'h3aa005b4),
	.w8(32'h3b1c7cff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1038),
	.w1(32'h3b36a09c),
	.w2(32'h3b8580ae),
	.w3(32'h3b9f1944),
	.w4(32'h3b01d95f),
	.w5(32'h3b8c1e0b),
	.w6(32'h3baf3c10),
	.w7(32'h3b36e476),
	.w8(32'h3b9c5ad9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a299d),
	.w1(32'h37e3285f),
	.w2(32'h3b186800),
	.w3(32'hb87b5ce6),
	.w4(32'h39f068a8),
	.w5(32'h3a39f552),
	.w6(32'h3aa4b45c),
	.w7(32'h3ad24d63),
	.w8(32'h3b1e7121),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c431e),
	.w1(32'h3a26f111),
	.w2(32'h3c07ca8e),
	.w3(32'hba891c47),
	.w4(32'h3b432b65),
	.w5(32'h3bd50dee),
	.w6(32'hbb6bab75),
	.w7(32'h3b842f25),
	.w8(32'h3b7b7be5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a819d),
	.w1(32'hbacedb4a),
	.w2(32'h3b8dd11f),
	.w3(32'hba390543),
	.w4(32'hbbadbe37),
	.w5(32'h3b5843d3),
	.w6(32'h3a3aec66),
	.w7(32'hbb2fdfe3),
	.w8(32'h3af00a63),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c1574),
	.w1(32'hba0a3dc2),
	.w2(32'hba92fd23),
	.w3(32'h3a99e3a1),
	.w4(32'h3a08c63d),
	.w5(32'h3b69549e),
	.w6(32'h3b1112a2),
	.w7(32'h3a0d1f0f),
	.w8(32'h3ba691a0),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3811617e),
	.w1(32'hbb27d37d),
	.w2(32'hba88de71),
	.w3(32'hb9163b75),
	.w4(32'hbb3c1024),
	.w5(32'hbb61bb13),
	.w6(32'hbacc1863),
	.w7(32'hbb41aef9),
	.w8(32'hbb098f00),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b657e38),
	.w1(32'hb9cf876f),
	.w2(32'h3b30ecf1),
	.w3(32'h3afdc631),
	.w4(32'hbb232f03),
	.w5(32'h3b2e5e80),
	.w6(32'h3b5587cb),
	.w7(32'hb87c672f),
	.w8(32'h3b7614bb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b613b89),
	.w1(32'h3916780e),
	.w2(32'h3a38040b),
	.w3(32'h3abec8d4),
	.w4(32'hbb878177),
	.w5(32'h3b430502),
	.w6(32'h3a87cc6e),
	.w7(32'hbb16bba6),
	.w8(32'h3b838bca),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a925aa1),
	.w1(32'hba67aa44),
	.w2(32'hbaa116c3),
	.w3(32'h3b734c81),
	.w4(32'hbb09ee48),
	.w5(32'hbb0c78e5),
	.w6(32'h3a35d441),
	.w7(32'hbb5772d4),
	.w8(32'hbb56a632),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e3987),
	.w1(32'hb8f9255c),
	.w2(32'hbb0905c2),
	.w3(32'hba28dedb),
	.w4(32'h39ededf8),
	.w5(32'h3926032c),
	.w6(32'hba1bfce0),
	.w7(32'hb9555189),
	.w8(32'h39e14db8),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9d2cd),
	.w1(32'hba59d220),
	.w2(32'hba856790),
	.w3(32'hba3943ec),
	.w4(32'hbab4525c),
	.w5(32'h3ab88e46),
	.w6(32'h39a26760),
	.w7(32'h3920053d),
	.w8(32'h3963e798),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b62b6),
	.w1(32'h3b6ab56e),
	.w2(32'h3b8aae93),
	.w3(32'h3a951864),
	.w4(32'h3aeb51f0),
	.w5(32'h3a7e48e2),
	.w6(32'h3b309ee5),
	.w7(32'h3b2d62c2),
	.w8(32'h39c5a691),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fafcd),
	.w1(32'h3a0c1d43),
	.w2(32'h3b1f2f47),
	.w3(32'hbb36bd90),
	.w4(32'hba8d0bbe),
	.w5(32'hba32458e),
	.w6(32'hbaffd773),
	.w7(32'h3b1b9a93),
	.w8(32'h3a026b21),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12760d),
	.w1(32'h399b149c),
	.w2(32'h3b5814b7),
	.w3(32'hba655120),
	.w4(32'hbafcf6a0),
	.w5(32'hbaff69db),
	.w6(32'h3b15b657),
	.w7(32'h3a57241c),
	.w8(32'hbb4b768e),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cdf40),
	.w1(32'hb99303e2),
	.w2(32'h3a59161a),
	.w3(32'hbb80a27d),
	.w4(32'h3a7d6021),
	.w5(32'hbac72e68),
	.w6(32'hbae5039f),
	.w7(32'h3a47ccc7),
	.w8(32'hbb16e6ad),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac90fbc),
	.w1(32'hbb35808a),
	.w2(32'hba29873e),
	.w3(32'hbaf8e568),
	.w4(32'hbaaa517d),
	.w5(32'h3ba870be),
	.w6(32'hb83414ec),
	.w7(32'hba6397c8),
	.w8(32'h3b64ec93),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0761e9),
	.w1(32'h3aa7f279),
	.w2(32'h3a261bae),
	.w3(32'h3aa8177c),
	.w4(32'h3a0fa116),
	.w5(32'hbafab4ce),
	.w6(32'h3ad76093),
	.w7(32'hb73ca653),
	.w8(32'hbb5fda20),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba625a52),
	.w1(32'h3ae9519e),
	.w2(32'h3aec03b6),
	.w3(32'hbace6907),
	.w4(32'hbb1268ac),
	.w5(32'h3a7c175d),
	.w6(32'hbafd9ed4),
	.w7(32'hbb0a763f),
	.w8(32'h3ae01e3d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17adcd),
	.w1(32'h3af85ecb),
	.w2(32'h3b8243ea),
	.w3(32'h3b7e1535),
	.w4(32'h3b0752cc),
	.w5(32'h39922a9b),
	.w6(32'h3b808ae0),
	.w7(32'h3b896838),
	.w8(32'h3b2bac97),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d4c0b),
	.w1(32'h3ba54eff),
	.w2(32'h3bf9d660),
	.w3(32'h3b980442),
	.w4(32'h3b8ed1bf),
	.w5(32'h3c2c98f0),
	.w6(32'h3b9edbaa),
	.w7(32'h3b5b6bb8),
	.w8(32'h3c2025a7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5cd6c),
	.w1(32'hbae83408),
	.w2(32'hba5b9ea9),
	.w3(32'hb9c9816d),
	.w4(32'hbac2c724),
	.w5(32'hb89708e4),
	.w6(32'h3a97996b),
	.w7(32'hbb3aafbb),
	.w8(32'hbb2ab55c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef3c4a),
	.w1(32'hb94ea285),
	.w2(32'h3b280a29),
	.w3(32'h39ff7edb),
	.w4(32'hbaa909ca),
	.w5(32'h3b5ecdef),
	.w6(32'h3a83b2e9),
	.w7(32'h3a5b685a),
	.w8(32'h3b6a79b3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6352ab),
	.w1(32'hbb3ffa10),
	.w2(32'hbb068b00),
	.w3(32'hb92b3ed8),
	.w4(32'h391b74f5),
	.w5(32'h39f9f7ba),
	.w6(32'h3a3f970f),
	.w7(32'hba640273),
	.w8(32'hba47bbc3),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4731f),
	.w1(32'h3b3291fb),
	.w2(32'h3bc3a499),
	.w3(32'h3bb19ae4),
	.w4(32'h38ddffbf),
	.w5(32'h3b616bd7),
	.w6(32'h3bc47e82),
	.w7(32'h3a4b59b3),
	.w8(32'h3b9188f0),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2251bc),
	.w1(32'hbaa4e39e),
	.w2(32'h3b1b66b8),
	.w3(32'h3b027a9f),
	.w4(32'hbb1450a6),
	.w5(32'h3b6f2329),
	.w6(32'h3b30f23c),
	.w7(32'hbacb73c9),
	.w8(32'h3b85dd3b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8da961),
	.w1(32'h3b5f3a9f),
	.w2(32'h3bb8e518),
	.w3(32'h3baf302f),
	.w4(32'h3b35d269),
	.w5(32'h3be3c98f),
	.w6(32'h3b7ee041),
	.w7(32'h3ac53dd9),
	.w8(32'h3be84243),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39051157),
	.w1(32'h3a2f71c1),
	.w2(32'h3a41a340),
	.w3(32'h3a528e40),
	.w4(32'hba6c65ae),
	.w5(32'hba647f11),
	.w6(32'h3b00d8ad),
	.w7(32'hba8ed14f),
	.w8(32'hbb0f5176),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e8d7),
	.w1(32'h3b8d30f3),
	.w2(32'h3ba68dde),
	.w3(32'h3aa6d657),
	.w4(32'h3a9fa52c),
	.w5(32'h3b8c542f),
	.w6(32'h3b344846),
	.w7(32'h3b825d14),
	.w8(32'h3b8aa764),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c2c5a),
	.w1(32'h3a51e069),
	.w2(32'h38f203a4),
	.w3(32'h3acec0e3),
	.w4(32'h3a1661e5),
	.w5(32'hbabb2ea1),
	.w6(32'h3aacc729),
	.w7(32'h38a9310c),
	.w8(32'hb912d223),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3c509),
	.w1(32'h3b3e780a),
	.w2(32'h3b68f416),
	.w3(32'h37a2e994),
	.w4(32'hb93f9036),
	.w5(32'hba65fdd9),
	.w6(32'h3a113ea3),
	.w7(32'h3b1f95e7),
	.w8(32'hbade09ef),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23a949),
	.w1(32'hba9db1fe),
	.w2(32'hba4f736b),
	.w3(32'hba0c11c9),
	.w4(32'hba007005),
	.w5(32'hbadc2e89),
	.w6(32'hb9bee783),
	.w7(32'hb8ec89b5),
	.w8(32'h3a59ebd7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78fe04),
	.w1(32'h38e1cfe8),
	.w2(32'h3b185709),
	.w3(32'h3b755787),
	.w4(32'h39dfbfb2),
	.w5(32'h397ae839),
	.w6(32'h3b9edffa),
	.w7(32'h3a41c0e5),
	.w8(32'h3b04ad56),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01f8e8),
	.w1(32'h3b2b62d8),
	.w2(32'h3849a2dd),
	.w3(32'h3ae877a2),
	.w4(32'h39a7c68d),
	.w5(32'hbabceb54),
	.w6(32'h3a2efd45),
	.w7(32'h3aec3ce5),
	.w8(32'hbb3c709a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cdcf8),
	.w1(32'hbb4285f8),
	.w2(32'hbae7c936),
	.w3(32'hbb0567a3),
	.w4(32'hba50bcd8),
	.w5(32'h3a2677e9),
	.w6(32'hbadfc8ce),
	.w7(32'hba1c4d30),
	.w8(32'hb8c220ff),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d7ff),
	.w1(32'hbacfe05c),
	.w2(32'h39c164b0),
	.w3(32'hbb247534),
	.w4(32'hbb55271c),
	.w5(32'hba7e0184),
	.w6(32'hbaaacdde),
	.w7(32'hba7d27a4),
	.w8(32'hbad398ca),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39577e87),
	.w1(32'h39e3104a),
	.w2(32'h3a8362ef),
	.w3(32'hba3fbf31),
	.w4(32'hbafccd3d),
	.w5(32'h3aab7e74),
	.w6(32'h3968513a),
	.w7(32'hb8c315b3),
	.w8(32'h3ab52fd6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd851b),
	.w1(32'hbaa43834),
	.w2(32'hb9850767),
	.w3(32'h3ad66e38),
	.w4(32'hb9a7e4a0),
	.w5(32'h3b2c1775),
	.w6(32'hb9a865d6),
	.w7(32'hbae6a11d),
	.w8(32'h3b0d7e29),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01be59),
	.w1(32'h3a8229fb),
	.w2(32'h3a4acf2c),
	.w3(32'h3adcfd6a),
	.w4(32'h3a42a2b3),
	.w5(32'hba39737d),
	.w6(32'h3af7355c),
	.w7(32'h39f15ff9),
	.w8(32'h3ae8f60a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3716c),
	.w1(32'h3bc9d206),
	.w2(32'h3c2e68dc),
	.w3(32'h3b4c80c7),
	.w4(32'hbb2ff2f4),
	.w5(32'h3bd3fac4),
	.w6(32'h38749b35),
	.w7(32'hbb1a3b4d),
	.w8(32'h3b327633),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb20825),
	.w1(32'h3b0c6c3e),
	.w2(32'h3b6be187),
	.w3(32'h3bca26ff),
	.w4(32'hbab4d0d7),
	.w5(32'h3abc58a1),
	.w6(32'h3b8e90fd),
	.w7(32'hbab5d50c),
	.w8(32'h3b4cf329),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac87494),
	.w1(32'hbaa6fbfe),
	.w2(32'hba329cef),
	.w3(32'hb8ae655a),
	.w4(32'h3aa59a6a),
	.w5(32'hbaba2279),
	.w6(32'hba8d9cb1),
	.w7(32'hbaa80787),
	.w8(32'hba950f87),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883417c),
	.w1(32'hba0ae53f),
	.w2(32'hba57f270),
	.w3(32'hba773739),
	.w4(32'hb9ebc2bb),
	.w5(32'hb8922cfa),
	.w6(32'hb9909ecd),
	.w7(32'hba5eae0c),
	.w8(32'hba1fd23b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e17bb),
	.w1(32'h3a76e367),
	.w2(32'h3aa8bbcd),
	.w3(32'hba9ad5b6),
	.w4(32'hba47d53b),
	.w5(32'h398b0a91),
	.w6(32'hba1c3258),
	.w7(32'h3a6b4197),
	.w8(32'hb9d27130),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b20e84),
	.w1(32'hbb433261),
	.w2(32'hba47c018),
	.w3(32'hbb1c0275),
	.w4(32'hb9f2cc52),
	.w5(32'hba0ed902),
	.w6(32'hbb1c72c5),
	.w7(32'hb821adf2),
	.w8(32'hbac5f9aa),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340d98),
	.w1(32'hba775b91),
	.w2(32'h3a5ab1df),
	.w3(32'hba26ea0f),
	.w4(32'h3b208455),
	.w5(32'h3a48b917),
	.w6(32'hb984d2e3),
	.w7(32'h3b052429),
	.w8(32'h3ace6cef),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b650b10),
	.w1(32'h3ac76c56),
	.w2(32'h3b47b2ba),
	.w3(32'h3a86d86e),
	.w4(32'h39a59f25),
	.w5(32'h3addfb1e),
	.w6(32'h3b083274),
	.w7(32'h3aad76a4),
	.w8(32'h3b9064fd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63f313),
	.w1(32'h37f2c88f),
	.w2(32'h3a5dc98f),
	.w3(32'h3ab749a2),
	.w4(32'hbafb7d93),
	.w5(32'hb99f3bab),
	.w6(32'h3b9979a0),
	.w7(32'hba8b9c25),
	.w8(32'hb9e6cc9b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4a22),
	.w1(32'hbb837a92),
	.w2(32'hb65433f2),
	.w3(32'hbb8b8ac8),
	.w4(32'hba834a14),
	.w5(32'h3a5df162),
	.w6(32'hbb7c0b7f),
	.w7(32'hb9333ee8),
	.w8(32'hb325da38),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012bbf),
	.w1(32'h3b3f7541),
	.w2(32'h3bc4f61b),
	.w3(32'h3972fbda),
	.w4(32'h3afa05fe),
	.w5(32'h3b910816),
	.w6(32'h3b4fd6ac),
	.w7(32'h3b9ee8e8),
	.w8(32'h3b9ddb9d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b197651),
	.w1(32'h3ab9eeff),
	.w2(32'h3aa84cdc),
	.w3(32'h3b0ef971),
	.w4(32'h3b289081),
	.w5(32'h3b7f953c),
	.w6(32'h3b05241a),
	.w7(32'h3abb21da),
	.w8(32'h3b60615e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39286a),
	.w1(32'hbb2fdbf6),
	.w2(32'h3a6e32d7),
	.w3(32'h393ea10d),
	.w4(32'hba2dd135),
	.w5(32'h3a80c07f),
	.w6(32'hbac030e2),
	.w7(32'hbaf66362),
	.w8(32'hbab7bf25),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8c695),
	.w1(32'h3a464a4c),
	.w2(32'h39c1288d),
	.w3(32'h3b60f6d5),
	.w4(32'h3af889be),
	.w5(32'hbb117977),
	.w6(32'hbace95a6),
	.w7(32'hbb739743),
	.w8(32'hbb3d5c2d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b2251),
	.w1(32'h399e4d48),
	.w2(32'h3a8fd5ea),
	.w3(32'hbb32802e),
	.w4(32'hba5609f7),
	.w5(32'hba7bac28),
	.w6(32'hbb043ab2),
	.w7(32'h3ad32e21),
	.w8(32'hba25cd73),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396035a8),
	.w1(32'hbb0a83dd),
	.w2(32'hb8cd8cd6),
	.w3(32'hb99c8e9b),
	.w4(32'hb9c7b376),
	.w5(32'hbac2ee88),
	.w6(32'h3b2cddf0),
	.w7(32'h3af303da),
	.w8(32'hba83eae7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37ecb7),
	.w1(32'hba149780),
	.w2(32'h3b92ff9f),
	.w3(32'hbab0c6fc),
	.w4(32'hbb745915),
	.w5(32'h3a2ad560),
	.w6(32'h3ac2d9af),
	.w7(32'h3993d591),
	.w8(32'h396e0818),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c981e),
	.w1(32'hba8edcad),
	.w2(32'h3aed1b19),
	.w3(32'hba259b42),
	.w4(32'hbacc0e49),
	.w5(32'h3a020857),
	.w6(32'h3988e462),
	.w7(32'hb9dbc8e1),
	.w8(32'h3aeff25e),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc8c7c),
	.w1(32'hbb43d37b),
	.w2(32'hbac697b1),
	.w3(32'hbaab7706),
	.w4(32'hba92b699),
	.w5(32'hba47230c),
	.w6(32'hba941b9d),
	.w7(32'hba1cb204),
	.w8(32'hb99e7509),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b066946),
	.w1(32'h3a9f5ef1),
	.w2(32'h3b3e56ee),
	.w3(32'h3a79d5a3),
	.w4(32'hbab28ac7),
	.w5(32'hb88d17ea),
	.w6(32'h3b5b2952),
	.w7(32'h3b1975c9),
	.w8(32'h3b1714fb),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2dd8e6),
	.w1(32'h3a1005e8),
	.w2(32'h3b178038),
	.w3(32'hb8acf2f0),
	.w4(32'hba9e356c),
	.w5(32'h3adb695d),
	.w6(32'h3ae64ebb),
	.w7(32'h39eedf76),
	.w8(32'h3b5088eb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7bb49),
	.w1(32'h3b3a099c),
	.w2(32'h3bbc5ffa),
	.w3(32'h3bb6316e),
	.w4(32'hb97f92fa),
	.w5(32'h3b11faab),
	.w6(32'h3bb1e9ba),
	.w7(32'h3a90e8e7),
	.w8(32'h3b4825ed),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0ad4a),
	.w1(32'h3b148c0a),
	.w2(32'h3b0ffd0c),
	.w3(32'hbae6e60b),
	.w4(32'hb93bd224),
	.w5(32'h3ae0e9b9),
	.w6(32'hb9e59a5d),
	.w7(32'h3b3c6df3),
	.w8(32'h3a851d7f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f6cb8),
	.w1(32'hbb0ab83b),
	.w2(32'h3a6f29cd),
	.w3(32'hb9f74a47),
	.w4(32'hb9638f21),
	.w5(32'hba96864b),
	.w6(32'hbb55a9b7),
	.w7(32'hba74a941),
	.w8(32'h3a7a67a6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c7aff),
	.w1(32'hba618977),
	.w2(32'h3bc5c997),
	.w3(32'h3a801f28),
	.w4(32'h3a953389),
	.w5(32'h3bae06af),
	.w6(32'h3b340062),
	.w7(32'h3965be17),
	.w8(32'h3b983dae),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62d04f),
	.w1(32'h39b9a239),
	.w2(32'h3beb9cd0),
	.w3(32'h3b0af2f5),
	.w4(32'h3a9a945f),
	.w5(32'h3bcf222d),
	.w6(32'h3b101aca),
	.w7(32'h3a744660),
	.w8(32'h3b7b21bf),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57e9b9),
	.w1(32'h3a02c96a),
	.w2(32'h3b8bf70a),
	.w3(32'h3a850e41),
	.w4(32'hb9fc05ce),
	.w5(32'h3b4ae77d),
	.w6(32'h3b3b3043),
	.w7(32'h3a963127),
	.w8(32'h3bb62093),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96dc502),
	.w1(32'h3a0f46b5),
	.w2(32'hba919416),
	.w3(32'h3b9c849b),
	.w4(32'h3b6fcc55),
	.w5(32'h399bacfd),
	.w6(32'h3a56b77c),
	.w7(32'hb93ac5cf),
	.w8(32'hbb164beb),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a0aa6),
	.w1(32'hbac31500),
	.w2(32'hbad6603c),
	.w3(32'hbb03671f),
	.w4(32'hbaebdf73),
	.w5(32'h3959ba91),
	.w6(32'hbb407cfb),
	.w7(32'hbb2d3ced),
	.w8(32'hb9161dbc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d644a),
	.w1(32'h3a1fd4fb),
	.w2(32'h3a3a192d),
	.w3(32'h3a1c1c68),
	.w4(32'h3a00ac11),
	.w5(32'hba9a5c2e),
	.w6(32'h3a384a39),
	.w7(32'h3a9a7ad9),
	.w8(32'hbab6515f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e449c),
	.w1(32'h3b47f619),
	.w2(32'h3a06e886),
	.w3(32'h3b0a1202),
	.w4(32'h3abc6111),
	.w5(32'h3b2cd1aa),
	.w6(32'h3404aca0),
	.w7(32'hbaf78cb1),
	.w8(32'h3a9ba24c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb7d99),
	.w1(32'h3ba11c02),
	.w2(32'h3bd132c9),
	.w3(32'h3bb20b74),
	.w4(32'h3b98dcec),
	.w5(32'h3bed7a77),
	.w6(32'h3bccbd9e),
	.w7(32'h3b6a557e),
	.w8(32'h3bb2aa55),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab7e3),
	.w1(32'h3b1c7973),
	.w2(32'h3ba87303),
	.w3(32'h3b8df837),
	.w4(32'h3b435185),
	.w5(32'h3b801cf8),
	.w6(32'hb98045e3),
	.w7(32'h3b18e201),
	.w8(32'h3b133a27),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9912b6b),
	.w1(32'hbb48f655),
	.w2(32'hbb1d8884),
	.w3(32'h3a1bf4b9),
	.w4(32'hbafa8d9e),
	.w5(32'hb9c4b4f6),
	.w6(32'h3b0a51b2),
	.w7(32'hba874a7d),
	.w8(32'h3aa6ab05),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60e316),
	.w1(32'h3abd276a),
	.w2(32'h3b9199d4),
	.w3(32'h3b157681),
	.w4(32'hba9da590),
	.w5(32'h3b2a47ca),
	.w6(32'h3b4b0d54),
	.w7(32'h3959f2de),
	.w8(32'h3b979d5c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac2226),
	.w1(32'hb9a15c1c),
	.w2(32'hb841836f),
	.w3(32'hba36a69c),
	.w4(32'h37c51181),
	.w5(32'h3a87c526),
	.w6(32'hb9784296),
	.w7(32'hba69f6ee),
	.w8(32'h3af28229),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912dec5),
	.w1(32'hba7577a0),
	.w2(32'hba491a60),
	.w3(32'h3a558410),
	.w4(32'hb80b8072),
	.w5(32'hbafbc164),
	.w6(32'h3a200453),
	.w7(32'hb9974305),
	.w8(32'hba62c20c),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbd0f),
	.w1(32'hb9278d70),
	.w2(32'hb9da2dc9),
	.w3(32'hb7fe28ae),
	.w4(32'hb9d395e5),
	.w5(32'h3b1ce580),
	.w6(32'h3aaf3ff0),
	.w7(32'h3a75763b),
	.w8(32'hb97a3cdd),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a969da7),
	.w1(32'h39f6560d),
	.w2(32'h39e617dd),
	.w3(32'hbb350bed),
	.w4(32'h3a8e67b1),
	.w5(32'h3962892e),
	.w6(32'hbb5195fc),
	.w7(32'h39f57940),
	.w8(32'hba98e135),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f14afc),
	.w1(32'h3a6d34e5),
	.w2(32'h39b82e77),
	.w3(32'h3b30a151),
	.w4(32'h3b50d967),
	.w5(32'hbb4b3f4f),
	.w6(32'h39f63a0a),
	.w7(32'h3b1d31a7),
	.w8(32'h3b96e519),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0df4b5),
	.w1(32'h3b472458),
	.w2(32'h3b7f55c2),
	.w3(32'hba06797f),
	.w4(32'hbaddb248),
	.w5(32'h3b80072b),
	.w6(32'hba4936a9),
	.w7(32'hbacefe95),
	.w8(32'hbb59fe23),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b938a9f),
	.w1(32'h3a93dd8d),
	.w2(32'h3aea17ee),
	.w3(32'h3bb2b69f),
	.w4(32'h3b1f8783),
	.w5(32'h3c23527e),
	.w6(32'hbbe844ad),
	.w7(32'hbab580fc),
	.w8(32'h3c71db3c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e2e5d),
	.w1(32'h3bb386be),
	.w2(32'h3c051558),
	.w3(32'h3c3044ec),
	.w4(32'h3bb566dc),
	.w5(32'hbb75bb4e),
	.w6(32'h3c498d96),
	.w7(32'h3c8ecf5f),
	.w8(32'hbb2a0631),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1bfdd),
	.w1(32'h398b2d18),
	.w2(32'h3c0c314a),
	.w3(32'h39d3a72a),
	.w4(32'hb98bd2f6),
	.w5(32'hba858344),
	.w6(32'h3b61a961),
	.w7(32'h3bd633c4),
	.w8(32'h3b5eb011),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04c3d0),
	.w1(32'h3b665b3e),
	.w2(32'h380f885b),
	.w3(32'hbb80d1da),
	.w4(32'hbb10bc9b),
	.w5(32'hb7905e5b),
	.w6(32'h3b9cc2e8),
	.w7(32'hba61c69d),
	.w8(32'hbbe5e586),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a83ca),
	.w1(32'hbc0cfeac),
	.w2(32'hbb5dbde2),
	.w3(32'hb9caeabc),
	.w4(32'h3c0629bc),
	.w5(32'hbb5a36d9),
	.w6(32'hbb14dc20),
	.w7(32'h3a3b0b5e),
	.w8(32'hbb344204),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0cd7),
	.w1(32'h3b579c49),
	.w2(32'h3aaf593a),
	.w3(32'hba296d6b),
	.w4(32'hbb2244b1),
	.w5(32'hbb94dc89),
	.w6(32'hbbe86730),
	.w7(32'hbab5c326),
	.w8(32'h3b7d4f17),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6322f),
	.w1(32'hbbeae05f),
	.w2(32'hb891a9ff),
	.w3(32'hba958789),
	.w4(32'h39a70e25),
	.w5(32'hbb9cdc72),
	.w6(32'hbaf61149),
	.w7(32'h3b886626),
	.w8(32'hbb57cc1c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba782f37),
	.w1(32'hbae334c6),
	.w2(32'h39696fbe),
	.w3(32'hbb1dc265),
	.w4(32'h3acac9b1),
	.w5(32'h3b276a34),
	.w6(32'hbb9fc37e),
	.w7(32'hba6f00bb),
	.w8(32'h3abae039),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a1c91),
	.w1(32'h3a3c973e),
	.w2(32'h390f4c1a),
	.w3(32'h3bd94b4d),
	.w4(32'h3ae44a33),
	.w5(32'hbb1d0271),
	.w6(32'h3afb6456),
	.w7(32'h3b3dc3c0),
	.w8(32'h3bca5bb0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f27cc1),
	.w1(32'hb9ce6650),
	.w2(32'h3a887fe8),
	.w3(32'hbaf24995),
	.w4(32'hba9c8d30),
	.w5(32'hba67e303),
	.w6(32'h3b99eba4),
	.w7(32'h3bfe1d5e),
	.w8(32'hbb0b9e49),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c38ba),
	.w1(32'hbb901c08),
	.w2(32'hba84a1bf),
	.w3(32'hbb7f01c2),
	.w4(32'hba521ebe),
	.w5(32'hbab06dc5),
	.w6(32'hbb8e8213),
	.w7(32'h3b6082d9),
	.w8(32'hb8da1a05),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ce419),
	.w1(32'h3c79784b),
	.w2(32'h3c55b464),
	.w3(32'h3c433eb1),
	.w4(32'h3c1bb238),
	.w5(32'h3bb188f6),
	.w6(32'h3c9c62f1),
	.w7(32'h3be2df58),
	.w8(32'h3c3ae479),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f99a),
	.w1(32'h3b7916c1),
	.w2(32'h3c0a57e5),
	.w3(32'h3b4ad8b9),
	.w4(32'h3ac30b34),
	.w5(32'h3b8b5bd2),
	.w6(32'h3babf3c5),
	.w7(32'h3c00b49a),
	.w8(32'hbb39d3c8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed0e5f),
	.w1(32'h3bf3b3e4),
	.w2(32'h3c2ac970),
	.w3(32'h3b6bf28e),
	.w4(32'h37bc62e4),
	.w5(32'hbbca65c0),
	.w6(32'hbb3d9806),
	.w7(32'hba7f8947),
	.w8(32'hbb82cb85),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4f40),
	.w1(32'h3b43d057),
	.w2(32'hbbf4dd86),
	.w3(32'hbb834cd5),
	.w4(32'hbb708acc),
	.w5(32'hbb933626),
	.w6(32'hbc097ee2),
	.w7(32'hbbc3c4cf),
	.w8(32'h3ba21f4c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba7a47),
	.w1(32'h3c53056e),
	.w2(32'h3bc2c16d),
	.w3(32'h3c7058c8),
	.w4(32'h3c8db6a9),
	.w5(32'hb904b0e1),
	.w6(32'h3ca25e35),
	.w7(32'h3c73b0b8),
	.w8(32'hbb37f3c6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba7d68),
	.w1(32'hbaf95527),
	.w2(32'hba6e49b4),
	.w3(32'hbb2c46fe),
	.w4(32'hbb066158),
	.w5(32'h3b8dd94a),
	.w6(32'hbb64e31d),
	.w7(32'hbb63c9d8),
	.w8(32'h3b88ac0d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abf98),
	.w1(32'hb9f77a91),
	.w2(32'h3ae7704f),
	.w3(32'hbb29869d),
	.w4(32'hba9394c0),
	.w5(32'h3aafa224),
	.w6(32'h3b60fa0b),
	.w7(32'h3bf25561),
	.w8(32'h3aa64abc),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2de3),
	.w1(32'h37d61e72),
	.w2(32'h3b8264cc),
	.w3(32'h3902d0d9),
	.w4(32'h3aee3de1),
	.w5(32'h3b49a931),
	.w6(32'h3a696f24),
	.w7(32'h3bf6cf3b),
	.w8(32'h3bc83a96),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad489c),
	.w1(32'h3bd529b3),
	.w2(32'h3ba60357),
	.w3(32'h3b9ad82e),
	.w4(32'h3aad4356),
	.w5(32'hbb43b96d),
	.w6(32'h3be4eeb3),
	.w7(32'h3c225bc5),
	.w8(32'hbbfe56b3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729258),
	.w1(32'hbb158858),
	.w2(32'h3b9d612d),
	.w3(32'hbb885cae),
	.w4(32'hbbfc918e),
	.w5(32'hbc1e5604),
	.w6(32'hbb74c5da),
	.w7(32'hbb2c57fc),
	.w8(32'hbb830a85),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2b1aa),
	.w1(32'h3b027409),
	.w2(32'hbb448f34),
	.w3(32'hbb9cdd0d),
	.w4(32'hbb356b40),
	.w5(32'h3bb8d0c8),
	.w6(32'h3a9fb9b6),
	.w7(32'hbb07b0ab),
	.w8(32'h3bc2bd13),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b325),
	.w1(32'hbae49f68),
	.w2(32'h3abc1479),
	.w3(32'h3ba8e781),
	.w4(32'hbb3b2152),
	.w5(32'hbc0ce33b),
	.w6(32'h3b96f588),
	.w7(32'hbb40e7a9),
	.w8(32'hbb8a36e7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8b60),
	.w1(32'hb90346d7),
	.w2(32'hba98c4a5),
	.w3(32'hbb1550a2),
	.w4(32'hbaf06737),
	.w5(32'h3ac9751f),
	.w6(32'hbbd1df9b),
	.w7(32'hbba016c7),
	.w8(32'h3bfbb154),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a059279),
	.w1(32'hbbd57c2c),
	.w2(32'hbac9f9a3),
	.w3(32'hbb238794),
	.w4(32'hbb999c0c),
	.w5(32'hbba057ae),
	.w6(32'h3bb5557c),
	.w7(32'h3a676ddd),
	.w8(32'h3a40a5e1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4e3fb),
	.w1(32'h3b86cb8d),
	.w2(32'h3b54b795),
	.w3(32'hbbba5b33),
	.w4(32'hbb8baca3),
	.w5(32'h3aa3e615),
	.w6(32'h3bb50ee5),
	.w7(32'h3b0c90e5),
	.w8(32'h3afbacf6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f8d3d5),
	.w1(32'hb9ecf89b),
	.w2(32'hb9e0757b),
	.w3(32'h39a8b948),
	.w4(32'h3a942252),
	.w5(32'h3b277ca6),
	.w6(32'hb97a8fcb),
	.w7(32'h3b1c5553),
	.w8(32'hbb8779b1),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e31a12),
	.w1(32'hbb41e046),
	.w2(32'hbc095c1d),
	.w3(32'h3b783c67),
	.w4(32'hbbbc449c),
	.w5(32'hbb341667),
	.w6(32'h3b872c07),
	.w7(32'hbba3d8a1),
	.w8(32'h3bedb520),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule