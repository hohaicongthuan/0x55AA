module layer_8_featuremap_158(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f5103),
	.w1(32'hbbdcbce6),
	.w2(32'hbb8e580e),
	.w3(32'hbb8b4e4b),
	.w4(32'hbbd65407),
	.w5(32'hbbc62245),
	.w6(32'hbc1d19bf),
	.w7(32'h3aa3c750),
	.w8(32'hbb419f1c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0f4c3),
	.w1(32'h3a947a20),
	.w2(32'hb98e180e),
	.w3(32'hbb1cf11c),
	.w4(32'h3b65e4f6),
	.w5(32'h3b9ea4c1),
	.w6(32'hbb508706),
	.w7(32'hbb832591),
	.w8(32'h3ab76ddc),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9e3ed),
	.w1(32'hbc8604b1),
	.w2(32'hbca0de7c),
	.w3(32'h3b3b2b39),
	.w4(32'hbb8c3e86),
	.w5(32'hbc2ccc4a),
	.w6(32'h3bb8d5ed),
	.w7(32'h3c9c56be),
	.w8(32'h3c0a0c01),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce0b86),
	.w1(32'h3c8ca07d),
	.w2(32'h3d18b635),
	.w3(32'hbc5e6887),
	.w4(32'hbc838ca2),
	.w5(32'hbce0a72a),
	.w6(32'h3c9de168),
	.w7(32'h3d0e362b),
	.w8(32'h3cd5309d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d18d732),
	.w1(32'h3bac67e3),
	.w2(32'h3c26fbb3),
	.w3(32'hbc82017b),
	.w4(32'hbb8c4774),
	.w5(32'hbbf9445b),
	.w6(32'h3b9e564e),
	.w7(32'h3bab7877),
	.w8(32'h3bc835a3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c352cea),
	.w1(32'h39f10f72),
	.w2(32'hba32ca1f),
	.w3(32'hbb846c7b),
	.w4(32'hba3879de),
	.w5(32'hbc1de516),
	.w6(32'hba73e9d8),
	.w7(32'hbc4ddfa8),
	.w8(32'hbc5da220),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e5f1),
	.w1(32'hba1aff4a),
	.w2(32'h3b5212e9),
	.w3(32'hbbf9ce35),
	.w4(32'hbb78a0b9),
	.w5(32'hbbf7da85),
	.w6(32'h3ad239e3),
	.w7(32'h3b5dfb58),
	.w8(32'hba14d23b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21fe87),
	.w1(32'hbb874a03),
	.w2(32'hba5427f3),
	.w3(32'hbbf1e697),
	.w4(32'hbbf3cb18),
	.w5(32'h3986909e),
	.w6(32'hb9bb783e),
	.w7(32'hbae77907),
	.w8(32'h396474dc),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b8ca),
	.w1(32'h3b26fa08),
	.w2(32'h3bf01caa),
	.w3(32'hbb5577b8),
	.w4(32'hbc80466a),
	.w5(32'hbcd4785c),
	.w6(32'h3bd746db),
	.w7(32'h3c5f3f7a),
	.w8(32'h3c3c5aae),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966728),
	.w1(32'h3c22e1fe),
	.w2(32'h3cd81d14),
	.w3(32'hbc8c7419),
	.w4(32'hba5be406),
	.w5(32'h3bab443a),
	.w6(32'h3b7308fb),
	.w7(32'h3c5398c5),
	.w8(32'h3c1908f9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c704fce),
	.w1(32'h3c2d2f80),
	.w2(32'h3b9ab3da),
	.w3(32'h3bc02224),
	.w4(32'h3c42cd1d),
	.w5(32'h3c0803b4),
	.w6(32'hbc0b942e),
	.w7(32'hbc6a9666),
	.w8(32'hbbd12fdb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27ed80),
	.w1(32'hba81aa6f),
	.w2(32'hbc3507ee),
	.w3(32'h3bfddfec),
	.w4(32'h3a0fc0ce),
	.w5(32'h398410c5),
	.w6(32'hbb5c2169),
	.w7(32'hbc0eaa86),
	.w8(32'h3a562283),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f70988),
	.w1(32'h3c91dd76),
	.w2(32'h3d1f3022),
	.w3(32'hb9b2aefa),
	.w4(32'h3c84a674),
	.w5(32'h3cd388aa),
	.w6(32'hbb953772),
	.w7(32'hbb6902dc),
	.w8(32'hbc13f536),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caedafe),
	.w1(32'hbcbde603),
	.w2(32'hbd02eff5),
	.w3(32'h3ca8e1e5),
	.w4(32'hbb5838e4),
	.w5(32'hbb7c0135),
	.w6(32'hbc2ed431),
	.w7(32'hbbea37d6),
	.w8(32'hbc7caf6b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5ba8c),
	.w1(32'h3a421179),
	.w2(32'h3b0f6293),
	.w3(32'hbc267f02),
	.w4(32'hbc16ba70),
	.w5(32'hbc920538),
	.w6(32'h3c2bc694),
	.w7(32'h3c8b1656),
	.w8(32'h3c692c65),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7414e2),
	.w1(32'h3bcffe07),
	.w2(32'h3bccd3ba),
	.w3(32'hbc25ced9),
	.w4(32'h3bfbee13),
	.w5(32'h3b55d834),
	.w6(32'hbc176cdf),
	.w7(32'hbb503285),
	.w8(32'hbafbd25f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd79099),
	.w1(32'hbb36969a),
	.w2(32'h3b0f656e),
	.w3(32'hbb0f29ab),
	.w4(32'h3b9a6513),
	.w5(32'h3b8ec891),
	.w6(32'hbb7b0838),
	.w7(32'h3bb4c389),
	.w8(32'hbb3aedb2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8919aa),
	.w1(32'hbb0797d8),
	.w2(32'h3a545d70),
	.w3(32'h3bfd6c58),
	.w4(32'h3bc5086f),
	.w5(32'h3c80274f),
	.w6(32'h3a12e979),
	.w7(32'h3b9b87a8),
	.w8(32'h3b8ee3e6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc855179),
	.w1(32'hbbe876c9),
	.w2(32'h3c2566b2),
	.w3(32'h37d70c93),
	.w4(32'hba1c47e7),
	.w5(32'h3caa0e10),
	.w6(32'hbc4133e1),
	.w7(32'hbb9c0cfe),
	.w8(32'hbabc73ef),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20aee),
	.w1(32'hbb94755f),
	.w2(32'hbb6642df),
	.w3(32'h3c613bfc),
	.w4(32'hbb958b4f),
	.w5(32'hbc161142),
	.w6(32'h3b8eb737),
	.w7(32'h3c070b84),
	.w8(32'h3b9394db),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961231c),
	.w1(32'hbba37311),
	.w2(32'hb99f0c0b),
	.w3(32'hbbefa740),
	.w4(32'hbb975530),
	.w5(32'hbb45f119),
	.w6(32'hbbee6d05),
	.w7(32'hbc35e03b),
	.w8(32'hbc216b75),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc425d2b),
	.w1(32'h39d59e58),
	.w2(32'hbc1988bd),
	.w3(32'h3b43c7e3),
	.w4(32'hbc19d1b4),
	.w5(32'hbc19191a),
	.w6(32'hbbd93846),
	.w7(32'h3b228850),
	.w8(32'hbbd2c63f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cfcab),
	.w1(32'hbcb65c89),
	.w2(32'hbb5c3efb),
	.w3(32'hbb3383d0),
	.w4(32'h3c1d7135),
	.w5(32'h3d02c723),
	.w6(32'h3b16e5d1),
	.w7(32'h3c6cca0d),
	.w8(32'h3c102e44),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9de539),
	.w1(32'h3c25b9cb),
	.w2(32'h3b63289c),
	.w3(32'h3ca9bea1),
	.w4(32'hbb8a5d90),
	.w5(32'hba314891),
	.w6(32'h397b5ad1),
	.w7(32'h3bd6d5fc),
	.w8(32'h3b14697b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad23076),
	.w1(32'hbc3f84ad),
	.w2(32'hbcc75cce),
	.w3(32'h3beb815d),
	.w4(32'h3a91cf8b),
	.w5(32'h3b641ab6),
	.w6(32'h3c5152ae),
	.w7(32'h3c8f9192),
	.w8(32'h3c6127d9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc958445),
	.w1(32'hbb36d553),
	.w2(32'hbcdb0631),
	.w3(32'hba72a4e3),
	.w4(32'h3c7b47af),
	.w5(32'h3d091b84),
	.w6(32'h3906cc66),
	.w7(32'h3b350076),
	.w8(32'h3b0c8696),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89e728),
	.w1(32'h3b1b6dc0),
	.w2(32'h3b16b4b8),
	.w3(32'h3cee19da),
	.w4(32'hbc059d3a),
	.w5(32'hbc90eea1),
	.w6(32'hbaa6e99d),
	.w7(32'h3be2dad9),
	.w8(32'h3c409643),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c2c15),
	.w1(32'hbcbe7674),
	.w2(32'hbca52dd3),
	.w3(32'hbcdc8311),
	.w4(32'hbad551e0),
	.w5(32'hbc7221ef),
	.w6(32'hbccebf26),
	.w7(32'h3b43ca77),
	.w8(32'hbc39559a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc48b),
	.w1(32'hbb2147ff),
	.w2(32'h3b1b3ce2),
	.w3(32'hbbe25247),
	.w4(32'h3b3c5ad9),
	.w5(32'h3c182764),
	.w6(32'hbb9f7c96),
	.w7(32'hbba14fda),
	.w8(32'h3b4536e0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f292),
	.w1(32'h3a8590d2),
	.w2(32'h3bc46b21),
	.w3(32'h3b6a491b),
	.w4(32'h3c483f25),
	.w5(32'h3c01b285),
	.w6(32'hbad14bf2),
	.w7(32'h3af14168),
	.w8(32'h3b8bf848),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c060b3a),
	.w1(32'h3ca879d9),
	.w2(32'h3d2a782a),
	.w3(32'h3c52118e),
	.w4(32'h3c13dbcf),
	.w5(32'h3cc3d0a4),
	.w6(32'h39891a1c),
	.w7(32'hbc36b9c4),
	.w8(32'hbc11d6ce),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdcec7c),
	.w1(32'h3b1ab193),
	.w2(32'hbc482e30),
	.w3(32'h3c9cf4cf),
	.w4(32'h3c8de56e),
	.w5(32'h3cd31fb7),
	.w6(32'hba79be6a),
	.w7(32'hbcbdfe9d),
	.w8(32'hbc804b0d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc759ce5),
	.w1(32'h3a5ebb56),
	.w2(32'h3b8a4d79),
	.w3(32'h3cc29755),
	.w4(32'h3a81e819),
	.w5(32'hbc1634b6),
	.w6(32'h3ad9b9b2),
	.w7(32'h3bcddf43),
	.w8(32'h3bb51e13),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbd3c0),
	.w1(32'h3bbd0d3f),
	.w2(32'h3bca0d93),
	.w3(32'hbc11ca5d),
	.w4(32'h3bd64b12),
	.w5(32'h3b476e3a),
	.w6(32'hb9868777),
	.w7(32'hba9b44f0),
	.w8(32'hb85fd9cd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17aebe),
	.w1(32'h3c03f78c),
	.w2(32'h3c997fcd),
	.w3(32'h3bc19407),
	.w4(32'h3bac0743),
	.w5(32'h3c40af51),
	.w6(32'h3b7313e6),
	.w7(32'h3b0aea7d),
	.w8(32'hbb76898e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e53e7),
	.w1(32'h3ba0729c),
	.w2(32'h3afcf1d9),
	.w3(32'h3c13466d),
	.w4(32'h3a5bd92c),
	.w5(32'hbba449bd),
	.w6(32'hbbe47d4c),
	.w7(32'hbba04e1e),
	.w8(32'hbb6de9c2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af30de9),
	.w1(32'hbc4385ea),
	.w2(32'hbc73ece0),
	.w3(32'hbb4d9601),
	.w4(32'hbba6d709),
	.w5(32'hbc1c5d05),
	.w6(32'hbaa20eec),
	.w7(32'hba5eaff6),
	.w8(32'hbb2e4358),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a7ff4),
	.w1(32'h3ba9f5bb),
	.w2(32'h3bf27210),
	.w3(32'hbbf66777),
	.w4(32'hbc43b7ea),
	.w5(32'hbca54502),
	.w6(32'h3c12f75a),
	.w7(32'h3c80ca10),
	.w8(32'h3c36c8db),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3113),
	.w1(32'h3b3b3b11),
	.w2(32'h3a66da60),
	.w3(32'hbc656f48),
	.w4(32'hbb722f0e),
	.w5(32'hbab7a9ea),
	.w6(32'h3b284a71),
	.w7(32'h3bba9c3d),
	.w8(32'hbb91a175),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f70263),
	.w1(32'h3b9453cf),
	.w2(32'h3c3a3603),
	.w3(32'hbb7dbb0f),
	.w4(32'h3ab41a59),
	.w5(32'h3bf08af5),
	.w6(32'hbb59bfab),
	.w7(32'hbba59062),
	.w8(32'hbadd06a9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cdf85),
	.w1(32'hbb3220f1),
	.w2(32'hbbc810f0),
	.w3(32'h39317a34),
	.w4(32'h3b8a0e6b),
	.w5(32'h3b001cba),
	.w6(32'hbb17ebbd),
	.w7(32'hb98c56d1),
	.w8(32'hbae0aacb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e2199),
	.w1(32'h3c0c4429),
	.w2(32'h3c00c474),
	.w3(32'h3ab8a1db),
	.w4(32'hbbd848fa),
	.w5(32'h3c323f0f),
	.w6(32'h3c10351c),
	.w7(32'h3bd749b6),
	.w8(32'hbb26de1e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc4460),
	.w1(32'hbc91fd9f),
	.w2(32'hbce10357),
	.w3(32'h3c067fc2),
	.w4(32'h3b4bbe32),
	.w5(32'hbc4069b1),
	.w6(32'h3b0673ab),
	.w7(32'h3b8612cb),
	.w8(32'h3ba6d80a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b1753),
	.w1(32'h3aea70ec),
	.w2(32'h3af89e55),
	.w3(32'hbc571fe9),
	.w4(32'hbb913c90),
	.w5(32'hbba855e9),
	.w6(32'h3ba1ce91),
	.w7(32'h3ba609af),
	.w8(32'h3b261e8c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8c5b3),
	.w1(32'hba6ae214),
	.w2(32'h3b6924bb),
	.w3(32'hb9eff339),
	.w4(32'h3ad914a1),
	.w5(32'h3b5c03b6),
	.w6(32'h3aa94257),
	.w7(32'h3bdf081d),
	.w8(32'h3c429345),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21b776),
	.w1(32'h3bb7676f),
	.w2(32'h3b47efe2),
	.w3(32'h3ba6f4e1),
	.w4(32'h3ba6869a),
	.w5(32'h39d6939b),
	.w6(32'h3c0b022d),
	.w7(32'h3c010294),
	.w8(32'h3c388d9e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f0fe),
	.w1(32'h3a27e039),
	.w2(32'hbb62bbf1),
	.w3(32'h3b9bfba6),
	.w4(32'h3b9df7ff),
	.w5(32'hbb8e2384),
	.w6(32'h3ba65047),
	.w7(32'h3b9a4c25),
	.w8(32'h3a67c3bf),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903ffc2),
	.w1(32'h3b8f4637),
	.w2(32'h3b21e3d2),
	.w3(32'hb97ad834),
	.w4(32'hbb9d56e8),
	.w5(32'h3ad63d44),
	.w6(32'hb926b48d),
	.w7(32'h3a41caf4),
	.w8(32'h3c09cdf6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4a372),
	.w1(32'hbc0a513f),
	.w2(32'hbcfaab13),
	.w3(32'h3c25e951),
	.w4(32'hbc83a68d),
	.w5(32'hbc1983e3),
	.w6(32'hbbcc23db),
	.w7(32'hbb37f607),
	.w8(32'hbb982325),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce549c1),
	.w1(32'h3a33f9cc),
	.w2(32'hbbd1f25b),
	.w3(32'hbb6951ce),
	.w4(32'h3b8bc5bb),
	.w5(32'h3c95943b),
	.w6(32'hba97419f),
	.w7(32'h3b397e33),
	.w8(32'h3c1f7b66),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5369f),
	.w1(32'hbbc8b7fe),
	.w2(32'hbc92d54b),
	.w3(32'h3c46030b),
	.w4(32'h3b163472),
	.w5(32'hbbb2d29d),
	.w6(32'h3aeaa869),
	.w7(32'hbb6af8a1),
	.w8(32'h39e1257d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fb808),
	.w1(32'hbb7cae13),
	.w2(32'h3bb39c70),
	.w3(32'hbb081d0a),
	.w4(32'hbbf81100),
	.w5(32'h3bfde7c7),
	.w6(32'hbb9caa0b),
	.w7(32'hbb8357c2),
	.w8(32'h3b6adbe2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea3c35),
	.w1(32'h3b1c6ad4),
	.w2(32'hb9c38dc1),
	.w3(32'h3c48f853),
	.w4(32'h39ebccb9),
	.w5(32'hbb346b59),
	.w6(32'h3b4f3aee),
	.w7(32'h3acae62d),
	.w8(32'h3bbea42b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39070393),
	.w1(32'hbb8f5914),
	.w2(32'h3bb5e640),
	.w3(32'hba7770c2),
	.w4(32'h3b6203fe),
	.w5(32'h3c57f925),
	.w6(32'hba539b22),
	.w7(32'h3c191abb),
	.w8(32'h3b356fdf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dc004),
	.w1(32'hbac3ba26),
	.w2(32'hbac61728),
	.w3(32'h3c48f262),
	.w4(32'hbbe65924),
	.w5(32'hbbea040f),
	.w6(32'hbb9884c2),
	.w7(32'hbc0b8060),
	.w8(32'hbc09a560),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115115),
	.w1(32'hbb708e51),
	.w2(32'h3b55fec5),
	.w3(32'h39ef2b19),
	.w4(32'h3ad3dae2),
	.w5(32'h3aa5bb32),
	.w6(32'hbbe42dac),
	.w7(32'hb96605bc),
	.w8(32'h3c16b0fe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d2c9b),
	.w1(32'h3bc2a53a),
	.w2(32'hbaae2ecb),
	.w3(32'h3b4f7971),
	.w4(32'h3c78a94c),
	.w5(32'hbb964123),
	.w6(32'hbc197f2a),
	.w7(32'hbca104fc),
	.w8(32'hbbc35f89),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59376),
	.w1(32'hbb6db739),
	.w2(32'hbb5c067a),
	.w3(32'hbbdc4392),
	.w4(32'hbb83d275),
	.w5(32'hbc0edf96),
	.w6(32'hbbbba8a2),
	.w7(32'h3b1c833c),
	.w8(32'h3a790168),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8792aa),
	.w1(32'hbb9b08b9),
	.w2(32'hba8ab4a6),
	.w3(32'hbb350dd0),
	.w4(32'hbb01906c),
	.w5(32'hba1d5993),
	.w6(32'hba7a6d88),
	.w7(32'hbb4d7375),
	.w8(32'hba4acf8b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d4300),
	.w1(32'h3b06fdfc),
	.w2(32'h3bce82e5),
	.w3(32'hbae191a8),
	.w4(32'h3ad4ed4a),
	.w5(32'hbb988b7a),
	.w6(32'hbb6c8830),
	.w7(32'hbb82ff85),
	.w8(32'h3c170380),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8bbd3),
	.w1(32'hbc14f65b),
	.w2(32'hbcb53a59),
	.w3(32'hbb7a08c0),
	.w4(32'hbbbe9465),
	.w5(32'hbca51d20),
	.w6(32'h3bc850dd),
	.w7(32'h3c26aa43),
	.w8(32'h3c1e669a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc914e01),
	.w1(32'hbcac4093),
	.w2(32'hbd07d5d3),
	.w3(32'hbc63fb78),
	.w4(32'hbaf7259b),
	.w5(32'hbca7876f),
	.w6(32'h3c7cc537),
	.w7(32'h3cc976db),
	.w8(32'h3ca20e3d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbda368),
	.w1(32'hbaf8f1ad),
	.w2(32'hbc0c971b),
	.w3(32'hbc490340),
	.w4(32'h3c0163ef),
	.w5(32'h3c0f22f2),
	.w6(32'hbbbfd769),
	.w7(32'hbc78ffb2),
	.w8(32'hbc3873d5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f739),
	.w1(32'h3b29219d),
	.w2(32'hb9b67ae3),
	.w3(32'h3aac965b),
	.w4(32'h3aa9de47),
	.w5(32'hbb120d3e),
	.w6(32'h3ba34d02),
	.w7(32'h3b0a4536),
	.w8(32'h3ba9b7f1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaeb465),
	.w1(32'hb9db9ed7),
	.w2(32'hbbccb497),
	.w3(32'hbb82b5fb),
	.w4(32'h3bb69232),
	.w5(32'h3bf85c20),
	.w6(32'hba87ce6e),
	.w7(32'hbbf1923f),
	.w8(32'hbb4e5842),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c312),
	.w1(32'h3bf0d29a),
	.w2(32'h3b97561f),
	.w3(32'h3b44c86f),
	.w4(32'h3c067ad3),
	.w5(32'h3b4e8a16),
	.w6(32'h39bf4e83),
	.w7(32'h3ad020d6),
	.w8(32'h3b56de28),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f35e7),
	.w1(32'hbbbe8775),
	.w2(32'hbc8c263f),
	.w3(32'h3a69a637),
	.w4(32'hbb339bd9),
	.w5(32'hbc3ea2e2),
	.w6(32'hba42c9ec),
	.w7(32'hba95953c),
	.w8(32'h3b8d284c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a6d45),
	.w1(32'hbc43489b),
	.w2(32'hbc067af1),
	.w3(32'hbbb9efa4),
	.w4(32'hbbee1b6f),
	.w5(32'hbb8b6677),
	.w6(32'h3a21e840),
	.w7(32'h3bbddfaf),
	.w8(32'h3bbbe356),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef320a),
	.w1(32'h396cc6b7),
	.w2(32'hbbfba777),
	.w3(32'h3b451475),
	.w4(32'hba97e748),
	.w5(32'h3b34d86e),
	.w6(32'hbb8d942a),
	.w7(32'h3aa7acf7),
	.w8(32'h3b0334c4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bd108),
	.w1(32'hbbc7f891),
	.w2(32'hbc18e7ab),
	.w3(32'hbb3e5ce4),
	.w4(32'hbc4567fe),
	.w5(32'hbc23f016),
	.w6(32'hbba6fc79),
	.w7(32'h39512564),
	.w8(32'h3c2b90d6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1696bb),
	.w1(32'h3c4c5924),
	.w2(32'h3c8a1b15),
	.w3(32'hbc075763),
	.w4(32'hbba81fcd),
	.w5(32'hbbc737e8),
	.w6(32'h3be9130a),
	.w7(32'h3c491d84),
	.w8(32'hba080e91),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bec0f),
	.w1(32'hbc0db78e),
	.w2(32'hbcb753bc),
	.w3(32'hba9e7431),
	.w4(32'h3b47ccbe),
	.w5(32'hbb00ba65),
	.w6(32'h3a419503),
	.w7(32'hba7c086d),
	.w8(32'hbb1d56fa),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc0202),
	.w1(32'hbc1738af),
	.w2(32'hbca9cb49),
	.w3(32'hbc2529a4),
	.w4(32'hbc1e7acc),
	.w5(32'hbc32b9fc),
	.w6(32'hbb9c71b7),
	.w7(32'hbc0cbc42),
	.w8(32'hbb05707c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca22583),
	.w1(32'h3c5e0012),
	.w2(32'h3d0fbd5d),
	.w3(32'hbbd690f7),
	.w4(32'h3c244534),
	.w5(32'h3c3ad207),
	.w6(32'hbb317757),
	.w7(32'h3c21c3a5),
	.w8(32'hbaff0029),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb28cbb),
	.w1(32'hbcc716cf),
	.w2(32'hbcf56264),
	.w3(32'h3beec86a),
	.w4(32'hbb9c8b11),
	.w5(32'hbb72008b),
	.w6(32'hbc007cd5),
	.w7(32'hbb441e9f),
	.w8(32'h3b669666),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7e17f4),
	.w1(32'hbaa965dc),
	.w2(32'h3c5934da),
	.w3(32'h3bbeceb4),
	.w4(32'hbc411382),
	.w5(32'h3781f9b8),
	.w6(32'h3c1bbbfe),
	.w7(32'hbb8e1d33),
	.w8(32'h3b791058),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a2e2c),
	.w1(32'h3b1b1b6a),
	.w2(32'h3c0e93de),
	.w3(32'hbb18669a),
	.w4(32'h3c135567),
	.w5(32'h3c3b2645),
	.w6(32'hbbbfbe1d),
	.w7(32'h3b8001be),
	.w8(32'h3b1aea9c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c4206),
	.w1(32'hbb893adf),
	.w2(32'hbb52545d),
	.w3(32'h3b349f20),
	.w4(32'h3b4aa40b),
	.w5(32'hb9dc363a),
	.w6(32'hbc188d16),
	.w7(32'h3aeff7a6),
	.w8(32'h3aa4ef42),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e69d49),
	.w1(32'h3bd5dfb2),
	.w2(32'h3d08400f),
	.w3(32'hbae67274),
	.w4(32'hb8094b4e),
	.w5(32'h3c9167a1),
	.w6(32'hbb95d44b),
	.w7(32'h3c4f3688),
	.w8(32'h3b9ad68d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf15a9d),
	.w1(32'h3b96b849),
	.w2(32'hbb491843),
	.w3(32'h3c881a32),
	.w4(32'hbb4dce1d),
	.w5(32'hbbecf7ad),
	.w6(32'hbb5c8b39),
	.w7(32'hbbc728b9),
	.w8(32'hb9d1350e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855d31),
	.w1(32'hbc4d0a10),
	.w2(32'hbcf5eb8f),
	.w3(32'h3c113370),
	.w4(32'hbc169a5c),
	.w5(32'hbc3c9989),
	.w6(32'h3c3a47e3),
	.w7(32'h3c365824),
	.w8(32'h3b915637),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca02cbe),
	.w1(32'hbb859014),
	.w2(32'hbc017a58),
	.w3(32'hbc2a7309),
	.w4(32'h3bc887aa),
	.w5(32'hba14c498),
	.w6(32'hbaa1e820),
	.w7(32'h3ae0389a),
	.w8(32'hbb52b3db),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b8af1d),
	.w1(32'hbb21ca6a),
	.w2(32'h3a75aa9f),
	.w3(32'hbc4c711a),
	.w4(32'hbb4ae3d2),
	.w5(32'hbc3a7353),
	.w6(32'hb92ac8ca),
	.w7(32'h3c205347),
	.w8(32'h3beb0404),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb972c6bf),
	.w1(32'h3b28bb6c),
	.w2(32'h3b2b1bbe),
	.w3(32'hbb2b7552),
	.w4(32'hbb1b3a28),
	.w5(32'hbc0639ca),
	.w6(32'h3a9f1cb3),
	.w7(32'h3c8c2fae),
	.w8(32'hbb82fca3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33e068),
	.w1(32'hbc485f74),
	.w2(32'hbbd1efd8),
	.w3(32'h3b5e0fcd),
	.w4(32'hbc93ab7b),
	.w5(32'hbc79f217),
	.w6(32'hbbfbf127),
	.w7(32'h3ad517db),
	.w8(32'hbb9dfff6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadc9ad),
	.w1(32'h3c20791e),
	.w2(32'h3c1a50a2),
	.w3(32'hbc9a93f7),
	.w4(32'h3c45055d),
	.w5(32'h3ca674e8),
	.w6(32'hbb804c67),
	.w7(32'hbbf1f259),
	.w8(32'hbc049e94),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccfbf2),
	.w1(32'h3be7b261),
	.w2(32'h3c83ddbc),
	.w3(32'h3c53e9fb),
	.w4(32'hbc07d121),
	.w5(32'hbacb8ff3),
	.w6(32'hbb0736a0),
	.w7(32'hb9beb50a),
	.w8(32'hbbb488d1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09701c),
	.w1(32'hbca9c903),
	.w2(32'hbd296724),
	.w3(32'hba010aae),
	.w4(32'h3c4b5a24),
	.w5(32'h3c639fb2),
	.w6(32'h3c40a82b),
	.w7(32'h3c775fef),
	.w8(32'h3c9c05c9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8bb62),
	.w1(32'h3c22c7af),
	.w2(32'h3c8f30e2),
	.w3(32'h3c1713b3),
	.w4(32'h3bbc32a3),
	.w5(32'h3c4db062),
	.w6(32'hbc04abb3),
	.w7(32'hbc5f1c95),
	.w8(32'hbc8ddcef),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55f71f),
	.w1(32'hbb51fd0c),
	.w2(32'hbc93be72),
	.w3(32'h3c2b6261),
	.w4(32'hbc61d389),
	.w5(32'hbc573618),
	.w6(32'h3a9ef132),
	.w7(32'hbb071aa6),
	.w8(32'hbb0b35c6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c7e13),
	.w1(32'h382a0bda),
	.w2(32'hbc139c7e),
	.w3(32'hbbddd3eb),
	.w4(32'hbb3b2e13),
	.w5(32'hbbf23e06),
	.w6(32'h39e09349),
	.w7(32'h3bd5b2ae),
	.w8(32'hbb662649),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ab28),
	.w1(32'h3c8a9386),
	.w2(32'h3c2ed429),
	.w3(32'hbc385b69),
	.w4(32'h3c57d094),
	.w5(32'h3c074a19),
	.w6(32'h3b9d304e),
	.w7(32'h3a9c819a),
	.w8(32'hbba5d564),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4423fc),
	.w1(32'h3b53f3de),
	.w2(32'h3b7fa266),
	.w3(32'h3c0c0de9),
	.w4(32'h39345bb3),
	.w5(32'h3a81c51d),
	.w6(32'hbb969180),
	.w7(32'hbbc517ff),
	.w8(32'hbbc79d9e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a05b8),
	.w1(32'h3a34e534),
	.w2(32'hbb1a10e7),
	.w3(32'h3a39069a),
	.w4(32'h3bc1be0e),
	.w5(32'h3bed2b7b),
	.w6(32'h3b2d281c),
	.w7(32'hba58ac3b),
	.w8(32'h3b153b0b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd5ac),
	.w1(32'h3b5427b0),
	.w2(32'h3bc28878),
	.w3(32'h3b0285fe),
	.w4(32'h39d57369),
	.w5(32'hba977a02),
	.w6(32'hbb36cc5d),
	.w7(32'h3c417be9),
	.w8(32'h3c9dc511),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c443655),
	.w1(32'h3c85f9f8),
	.w2(32'h3c7205e7),
	.w3(32'hbc402bf2),
	.w4(32'h3c0c396e),
	.w5(32'h3bef8312),
	.w6(32'h3ab81250),
	.w7(32'hbb34b4b9),
	.w8(32'hbb47d2dd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb2458),
	.w1(32'hbbb78491),
	.w2(32'h3b50b836),
	.w3(32'h3ba9720f),
	.w4(32'h3b36a03e),
	.w5(32'h3c221993),
	.w6(32'h3a946427),
	.w7(32'h3c0439c9),
	.w8(32'h3b71cdbb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3f5c),
	.w1(32'hbb48c5aa),
	.w2(32'h3bef8a6a),
	.w3(32'hbab2e1a2),
	.w4(32'h3ad2cea8),
	.w5(32'hbbb3e8e6),
	.w6(32'h3b5e716d),
	.w7(32'h3b8ecf71),
	.w8(32'h3c0a9228),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37cbd6),
	.w1(32'h3bd93a4c),
	.w2(32'hbb3cd296),
	.w3(32'hbb87d622),
	.w4(32'h3a11a90a),
	.w5(32'hbbb8a250),
	.w6(32'h3b0c0592),
	.w7(32'hbb97513b),
	.w8(32'h3b374ae7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7506dd),
	.w1(32'hbc5bdf3d),
	.w2(32'hbc74d29c),
	.w3(32'hbb629a78),
	.w4(32'hbaeb91b1),
	.w5(32'hbbeb6825),
	.w6(32'hbab3ebe5),
	.w7(32'h3b69a4be),
	.w8(32'h3bd843ab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98bebc),
	.w1(32'h393d999c),
	.w2(32'h3b966d25),
	.w3(32'hbb166219),
	.w4(32'hbbc58a01),
	.w5(32'hbb6dffdf),
	.w6(32'hbbe877f4),
	.w7(32'h3c04e107),
	.w8(32'h3a2fa5dd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c4c64),
	.w1(32'h3b02866d),
	.w2(32'h3bbc7551),
	.w3(32'hbac05c15),
	.w4(32'hbc0275b3),
	.w5(32'hbc0dae66),
	.w6(32'hbb067221),
	.w7(32'hbbb8ccc3),
	.w8(32'hba3460a4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfce26),
	.w1(32'hbb856897),
	.w2(32'h3b84a33d),
	.w3(32'h38d5298f),
	.w4(32'h3ba7aafe),
	.w5(32'h3c56c09b),
	.w6(32'h3abcee89),
	.w7(32'h3b87bb1f),
	.w8(32'h3b2d9e86),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68659c),
	.w1(32'h3a51a7a4),
	.w2(32'hbb89c9de),
	.w3(32'h39bec4fa),
	.w4(32'hbb63f84f),
	.w5(32'hbc8bf80a),
	.w6(32'hbb48d41e),
	.w7(32'hbc36accb),
	.w8(32'hbbeee862),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5f2b0),
	.w1(32'h3b20ace3),
	.w2(32'h3b208d4e),
	.w3(32'hbc5c89d4),
	.w4(32'hba8095c6),
	.w5(32'h3c1bacec),
	.w6(32'h39700ec0),
	.w7(32'h3bad2170),
	.w8(32'h3b5948e9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b2543),
	.w1(32'h3b29692b),
	.w2(32'hba774d13),
	.w3(32'h3b6ef7aa),
	.w4(32'h3a146adf),
	.w5(32'hbb23f070),
	.w6(32'h3b4f13c1),
	.w7(32'h3b466f8f),
	.w8(32'h3bd4e111),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f020),
	.w1(32'h3c6d1da9),
	.w2(32'h3cc10a21),
	.w3(32'h3aa1ac9b),
	.w4(32'h3b928c0b),
	.w5(32'h3c05b488),
	.w6(32'h3ab236ca),
	.w7(32'hbb199af0),
	.w8(32'hbb8b61e6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d418e),
	.w1(32'hbcd97774),
	.w2(32'hbd18332b),
	.w3(32'h3c0de3e4),
	.w4(32'hbb9cc6ca),
	.w5(32'hbc945895),
	.w6(32'hbb06bbb5),
	.w7(32'h3c085847),
	.w8(32'h3c4bf27a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3455b8),
	.w1(32'hbbd09bea),
	.w2(32'hbc34450f),
	.w3(32'hbb3ecb77),
	.w4(32'hbbfaf66d),
	.w5(32'hbba50833),
	.w6(32'hbaf5ff44),
	.w7(32'hbc13d343),
	.w8(32'hbbe9aa4e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1715fb),
	.w1(32'h3aa8069e),
	.w2(32'hbad7b902),
	.w3(32'hba1e2e55),
	.w4(32'h3b64fad0),
	.w5(32'h3bdb0ee8),
	.w6(32'hbb8d978e),
	.w7(32'hbc0c94c6),
	.w8(32'hbbd4fd9b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba47e42),
	.w1(32'h3ba2e411),
	.w2(32'hbb94e5f6),
	.w3(32'h3af1e7f1),
	.w4(32'h3ad22abc),
	.w5(32'hba5a53d4),
	.w6(32'h3bff8146),
	.w7(32'h3b39dc76),
	.w8(32'h3b2c8997),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a57ed),
	.w1(32'h3aaffb65),
	.w2(32'hba978443),
	.w3(32'hbbf77fc6),
	.w4(32'h3c360039),
	.w5(32'h3c29d847),
	.w6(32'h3a9b8b5f),
	.w7(32'hbb0e10bd),
	.w8(32'h3aeeeb37),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a874a),
	.w1(32'hbb7072d3),
	.w2(32'hbc18a375),
	.w3(32'h3c0f6160),
	.w4(32'hbb0f1aa1),
	.w5(32'hbb9cf668),
	.w6(32'hbba5e110),
	.w7(32'hbc349222),
	.w8(32'hbbe28e45),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf31ff),
	.w1(32'hbb9b3e95),
	.w2(32'hbcbae0bb),
	.w3(32'hbc22d118),
	.w4(32'h3cffa5f9),
	.w5(32'h3d5796af),
	.w6(32'hbc016f7a),
	.w7(32'hbbf60542),
	.w8(32'hbc2f428c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff3209),
	.w1(32'h3c376dfb),
	.w2(32'h3ccc4a27),
	.w3(32'h3d1e2897),
	.w4(32'h3a8d0b45),
	.w5(32'h3c84cff7),
	.w6(32'hbc0a12c5),
	.w7(32'hbc4fe37a),
	.w8(32'hbc8c3b64),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86a74e),
	.w1(32'hb9c6033f),
	.w2(32'hbba08ef9),
	.w3(32'h3c80f692),
	.w4(32'h3bb0a526),
	.w5(32'h3bf0eaaa),
	.w6(32'hbb30a9da),
	.w7(32'hbc0f15d2),
	.w8(32'hbbcd6bf1),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b2409),
	.w1(32'hbc14e89e),
	.w2(32'hbc3f89a5),
	.w3(32'h3b2ca8c5),
	.w4(32'h3ba9acf8),
	.w5(32'hbb5417fc),
	.w6(32'hbaa47c80),
	.w7(32'hbabc3ea1),
	.w8(32'h3bf5af57),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc489569),
	.w1(32'hbc126961),
	.w2(32'hbbe0caac),
	.w3(32'h3b25d2bb),
	.w4(32'hbb9df8de),
	.w5(32'hbc11e63d),
	.w6(32'hbc212407),
	.w7(32'hbbcf1ab0),
	.w8(32'hbbb92c02),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc095d5b),
	.w1(32'hbc5530e5),
	.w2(32'hbcbf2c39),
	.w3(32'hbc18ad99),
	.w4(32'h3b2a8164),
	.w5(32'h3c3a81fd),
	.w6(32'hba1326cc),
	.w7(32'hbb3b8ef4),
	.w8(32'h39fd60cd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec8ae6),
	.w1(32'hbc322e9f),
	.w2(32'hbc9f444a),
	.w3(32'hbbad336f),
	.w4(32'hbbf705f0),
	.w5(32'hbc436b96),
	.w6(32'h3b3f4e8a),
	.w7(32'h3a613b4c),
	.w8(32'h3b7ceae6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e4a46),
	.w1(32'h3bca821d),
	.w2(32'hbbb8ad47),
	.w3(32'h39ab5797),
	.w4(32'h3a90d144),
	.w5(32'h3ba294d3),
	.w6(32'h3ad9a601),
	.w7(32'h3b131ac6),
	.w8(32'h3b09e4b3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe47ba),
	.w1(32'h3aa87837),
	.w2(32'hbb6297b2),
	.w3(32'h3a57ba35),
	.w4(32'h3add9eb2),
	.w5(32'hbc56c8e4),
	.w6(32'hba5bfb51),
	.w7(32'hbc1993dd),
	.w8(32'hbb812f88),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc411765),
	.w1(32'h3a20ef72),
	.w2(32'hbb0dfcf1),
	.w3(32'hbc62e526),
	.w4(32'h3af7cabb),
	.w5(32'h3b2cf257),
	.w6(32'h3a1b3fb3),
	.w7(32'hbba54d56),
	.w8(32'h397ec6fa),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02f94d),
	.w1(32'h3ac97149),
	.w2(32'hbb78df4d),
	.w3(32'hba9eb669),
	.w4(32'h3a132f75),
	.w5(32'hbb1643a6),
	.w6(32'hbbd90ba3),
	.w7(32'hbb5bc321),
	.w8(32'hbb642d36),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f97c0),
	.w1(32'hbc4b0a22),
	.w2(32'hbccf4503),
	.w3(32'hbba9263d),
	.w4(32'h3b8a176c),
	.w5(32'hbb5ae4fe),
	.w6(32'hbb90cfe7),
	.w7(32'hbc8afb63),
	.w8(32'hbba4215e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf54225),
	.w1(32'h3b8adc63),
	.w2(32'h3a0edbdd),
	.w3(32'h3b103573),
	.w4(32'hbc2f946b),
	.w5(32'hb914d502),
	.w6(32'h3a8ef55d),
	.w7(32'hba84c7dc),
	.w8(32'h3bcd9218),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc459fc1),
	.w1(32'h39bf98a8),
	.w2(32'h3ab179aa),
	.w3(32'h3ba170c1),
	.w4(32'h3ab300e7),
	.w5(32'h3a7e22bd),
	.w6(32'h39115d84),
	.w7(32'h3a8902f3),
	.w8(32'h3a8feab7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1a97b),
	.w1(32'hbb498709),
	.w2(32'hba30b590),
	.w3(32'hba289745),
	.w4(32'hbb32bf01),
	.w5(32'h3a0705ca),
	.w6(32'hbb040baf),
	.w7(32'hbab48591),
	.w8(32'hb939cb8c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule