module layer_8_featuremap_139(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d1e45),
	.w1(32'hbc8045a8),
	.w2(32'hbbe071b2),
	.w3(32'hbb52428b),
	.w4(32'h3bb5e8d1),
	.w5(32'h3bc4af5b),
	.w6(32'h3b85d53c),
	.w7(32'hbc280eaa),
	.w8(32'h3c3442e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cc10c),
	.w1(32'h3c0575a8),
	.w2(32'h3c0acc0b),
	.w3(32'hb9a60be1),
	.w4(32'h3b3c326e),
	.w5(32'h3b689e29),
	.w6(32'h3b66526e),
	.w7(32'h3ba2ce1d),
	.w8(32'hbbaf4bd3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a949d),
	.w1(32'h3c842f88),
	.w2(32'hbb724cd8),
	.w3(32'hb9453604),
	.w4(32'hbb70268f),
	.w5(32'h3c0c34f6),
	.w6(32'hbabde578),
	.w7(32'h3c450944),
	.w8(32'hbca6fb3c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b013a63),
	.w1(32'h3bb67aba),
	.w2(32'h3bb200d6),
	.w3(32'h3be60f7d),
	.w4(32'hbcbd2a0d),
	.w5(32'hbc8db1bb),
	.w6(32'hbc3e8308),
	.w7(32'hbd0463ed),
	.w8(32'hbaa7b3bc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6feb2d),
	.w1(32'hbbee5a09),
	.w2(32'hbbe21995),
	.w3(32'hbc22e5d2),
	.w4(32'hbc20c64a),
	.w5(32'hba7da5a5),
	.w6(32'h3c7b485a),
	.w7(32'h3b0a4a29),
	.w8(32'hbc410b27),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca518e7),
	.w1(32'h3957aa07),
	.w2(32'hbb9d6ff5),
	.w3(32'hbbf482aa),
	.w4(32'hbb961ed7),
	.w5(32'hbbf6af1c),
	.w6(32'hbc55112a),
	.w7(32'hbc5bcb35),
	.w8(32'hbc114459),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43238b),
	.w1(32'hbae2e71f),
	.w2(32'hbc6a70a6),
	.w3(32'hbc25b562),
	.w4(32'h3c26fd66),
	.w5(32'hbc312589),
	.w6(32'h3bba55c1),
	.w7(32'hbcdba29b),
	.w8(32'h3c4178d6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8d511),
	.w1(32'hbb58d377),
	.w2(32'h3bcf5fc2),
	.w3(32'hbc9aee42),
	.w4(32'hbbf88ae9),
	.w5(32'h3ba44d51),
	.w6(32'hbc54470a),
	.w7(32'h3c149c94),
	.w8(32'hbc164e3a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885fbb3),
	.w1(32'h3c995ca3),
	.w2(32'hbcbf09d5),
	.w3(32'h3b34f2f1),
	.w4(32'hbc26d457),
	.w5(32'h3a9aae91),
	.w6(32'hbc070e2b),
	.w7(32'hbbdc7f1a),
	.w8(32'h3d2b888b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf170e),
	.w1(32'hbcd297bf),
	.w2(32'hbb209239),
	.w3(32'hba84b506),
	.w4(32'h3bf1e19b),
	.w5(32'hbc2d976e),
	.w6(32'h3ca20ad5),
	.w7(32'h3c8c4a31),
	.w8(32'h3ccb9f6a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85a4b3),
	.w1(32'h3bfbe781),
	.w2(32'hbb84e7ee),
	.w3(32'hbbc81c0c),
	.w4(32'hbc8c1205),
	.w5(32'hbc8676ff),
	.w6(32'h3aac0904),
	.w7(32'h3bea64b0),
	.w8(32'hbad98f2e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85b745),
	.w1(32'h3c01b752),
	.w2(32'hbba5a223),
	.w3(32'hbb87a672),
	.w4(32'hbc7f3654),
	.w5(32'hbb4fe85a),
	.w6(32'hbb3fc245),
	.w7(32'h3c26a070),
	.w8(32'hbc017dff),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e8cf3),
	.w1(32'h3c5d62ae),
	.w2(32'h3b1aa883),
	.w3(32'hbc2ebca5),
	.w4(32'h3b095a0e),
	.w5(32'h3c037c65),
	.w6(32'h3b2c09ca),
	.w7(32'h3bec2157),
	.w8(32'h3c216631),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc9d6f),
	.w1(32'h3b831198),
	.w2(32'hbab1f698),
	.w3(32'h3be925d3),
	.w4(32'hbb2ff2f5),
	.w5(32'hbafc8068),
	.w6(32'h3b903360),
	.w7(32'hb922d1a1),
	.w8(32'h3b45816a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4abb),
	.w1(32'hb80dfee9),
	.w2(32'hba8e70e1),
	.w3(32'h3b6d5008),
	.w4(32'hbb4ebd97),
	.w5(32'hba67e888),
	.w6(32'h3c3ebb97),
	.w7(32'h393c0f42),
	.w8(32'h3b35088c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba965a77),
	.w1(32'hbac6d499),
	.w2(32'hb9d85a4f),
	.w3(32'hb98fce93),
	.w4(32'hba986717),
	.w5(32'hba6fe54d),
	.w6(32'h3b801eec),
	.w7(32'hba91e21c),
	.w8(32'hbbaa0014),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d579),
	.w1(32'hbc866981),
	.w2(32'hba35ab88),
	.w3(32'hbba012ec),
	.w4(32'h3bc46e43),
	.w5(32'hbba014d8),
	.w6(32'hbbe3b3d2),
	.w7(32'h3a9810ca),
	.w8(32'h399fe429),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19453c),
	.w1(32'h37edc29c),
	.w2(32'h39999790),
	.w3(32'hbb4da5ce),
	.w4(32'hbbb9f5df),
	.w5(32'hbc1ffc57),
	.w6(32'h3c0a1ee3),
	.w7(32'hbc248325),
	.w8(32'hbcd39c4b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83b966),
	.w1(32'hbae6d4a4),
	.w2(32'h3abd1e46),
	.w3(32'hbc9e541f),
	.w4(32'hbba4b2c2),
	.w5(32'hbb3aec48),
	.w6(32'hbc41ecbd),
	.w7(32'h381586c9),
	.w8(32'hbc1aa1fc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6975),
	.w1(32'hbc4ea440),
	.w2(32'hbc824962),
	.w3(32'hbbfe7f61),
	.w4(32'hbc10496d),
	.w5(32'hbc80dd56),
	.w6(32'hbbe93597),
	.w7(32'h3c122838),
	.w8(32'h3d16d3db),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8acb25),
	.w1(32'hba84f518),
	.w2(32'h3ae9ca18),
	.w3(32'hbbb5309c),
	.w4(32'h3c007340),
	.w5(32'h3b369d53),
	.w6(32'h3cba8fc5),
	.w7(32'hbc9d2a82),
	.w8(32'h3b97e5f5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46520),
	.w1(32'hbc31da37),
	.w2(32'hb8eb707d),
	.w3(32'hbbe3d969),
	.w4(32'hbc061590),
	.w5(32'hbb701492),
	.w6(32'h3c987329),
	.w7(32'h3ba732ef),
	.w8(32'h3b496f1e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82a777),
	.w1(32'hbbf5b9b7),
	.w2(32'hbc429dbe),
	.w3(32'hbbbbd22f),
	.w4(32'hbbe6d73f),
	.w5(32'h3acd1401),
	.w6(32'h3bf30e2e),
	.w7(32'h3bf6f6fa),
	.w8(32'h3c9d58fb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc256604),
	.w1(32'hbc57bfac),
	.w2(32'h3c260889),
	.w3(32'hbbb568ec),
	.w4(32'h3b2b68b8),
	.w5(32'hbb683947),
	.w6(32'h3c05f499),
	.w7(32'h3c27e280),
	.w8(32'hbb25a6db),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba21c6b),
	.w1(32'h3bc7b7d2),
	.w2(32'h3a8dcce6),
	.w3(32'h3b579ef1),
	.w4(32'h3b78e78b),
	.w5(32'hbb2a5d2e),
	.w6(32'h37a1ebe3),
	.w7(32'h3b3f9d6f),
	.w8(32'hba29f96a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6c4bf),
	.w1(32'hbba8e9ae),
	.w2(32'h3b78c00c),
	.w3(32'hbb90893e),
	.w4(32'h3c480ed5),
	.w5(32'hbb8e02de),
	.w6(32'h3a95f78c),
	.w7(32'hbb40bb31),
	.w8(32'h3bdaba45),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5703ca),
	.w1(32'h3c66056e),
	.w2(32'hbc031609),
	.w3(32'hbbc4d789),
	.w4(32'hbaf5e8fd),
	.w5(32'hbc30530c),
	.w6(32'h3c6a31c0),
	.w7(32'h3c8f59ff),
	.w8(32'h3bdf1887),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2de30),
	.w1(32'hbcc6feff),
	.w2(32'hbd28765d),
	.w3(32'hbc32d6e9),
	.w4(32'hbce60c57),
	.w5(32'hbcf489a2),
	.w6(32'h3d0101f5),
	.w7(32'h3cd7a40f),
	.w8(32'h3d5734e1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd357f8),
	.w1(32'hbd0e4c07),
	.w2(32'hbb797c8a),
	.w3(32'hbcacf51b),
	.w4(32'hbb525fcb),
	.w5(32'hbbd4cde7),
	.w6(32'h3ce011ad),
	.w7(32'h3c32eec5),
	.w8(32'hbbfc0e6b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a80ef),
	.w1(32'hbc417adb),
	.w2(32'hbc9e83e3),
	.w3(32'h39050424),
	.w4(32'hbba93538),
	.w5(32'h3c0bb4ba),
	.w6(32'hbb6c0799),
	.w7(32'h3c69a223),
	.w8(32'h3d3debe2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabb638),
	.w1(32'hbc8ec05a),
	.w2(32'h3b996d4d),
	.w3(32'h3bcc10ba),
	.w4(32'h3b1e64b1),
	.w5(32'h3b5b1188),
	.w6(32'h3c8c9afd),
	.w7(32'h3c0eaaaa),
	.w8(32'h3c2f3a52),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8bc5),
	.w1(32'h3b3d0126),
	.w2(32'hbc5718d7),
	.w3(32'h3996fb25),
	.w4(32'hbc50c606),
	.w5(32'hba753d0e),
	.w6(32'h3be6e236),
	.w7(32'hbc88a7d7),
	.w8(32'hbb8d090e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbed086),
	.w1(32'hbce2d9d2),
	.w2(32'h3b05f7a1),
	.w3(32'hbc6d46d1),
	.w4(32'h398f6588),
	.w5(32'h3be685c6),
	.w6(32'hbc322320),
	.w7(32'h3c892511),
	.w8(32'h3cbc8e59),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b6e8b),
	.w1(32'hba86f25f),
	.w2(32'h3b8643b6),
	.w3(32'h3c3e0e50),
	.w4(32'h3bca4cfa),
	.w5(32'h3c081fd7),
	.w6(32'h3c1b2051),
	.w7(32'hbc8dd11e),
	.w8(32'hbcbd7844),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348a82),
	.w1(32'h3c5733cc),
	.w2(32'h3b978f49),
	.w3(32'h3a17a3b4),
	.w4(32'h3c7b8818),
	.w5(32'h3c453f14),
	.w6(32'hbc95d667),
	.w7(32'h3c00dcf4),
	.w8(32'h3b05f36a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2666),
	.w1(32'hbbd66004),
	.w2(32'h3b2309f1),
	.w3(32'h3bd52da7),
	.w4(32'hbc3cfb01),
	.w5(32'hba509a39),
	.w6(32'h3c0373e7),
	.w7(32'h3c3bbf4c),
	.w8(32'hbc0d8ad8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee06a0),
	.w1(32'h3c5029c4),
	.w2(32'hbbe73862),
	.w3(32'h3c23485c),
	.w4(32'hbc8fa4c9),
	.w5(32'hbc2b588c),
	.w6(32'hbcbcda3d),
	.w7(32'hbbe7194c),
	.w8(32'hbadc5020),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3082a0),
	.w1(32'hbb86f9f5),
	.w2(32'h3b073ba1),
	.w3(32'hbc6069de),
	.w4(32'h3bad6fdc),
	.w5(32'hb98b4ce8),
	.w6(32'hbc2f5c16),
	.w7(32'hbb40c6ba),
	.w8(32'hba94491c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad181f9),
	.w1(32'h3aa24d38),
	.w2(32'hbc439b4b),
	.w3(32'hbb817cbd),
	.w4(32'hbacff17e),
	.w5(32'hbb0cef08),
	.w6(32'hbb7fe061),
	.w7(32'hbc4d0ea6),
	.w8(32'hbcae7172),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f35e9),
	.w1(32'hbca29b39),
	.w2(32'hbb512fba),
	.w3(32'hbacd5c66),
	.w4(32'hb9f14887),
	.w5(32'hba9390b6),
	.w6(32'hbc84aa94),
	.w7(32'h3c7d0e3c),
	.w8(32'h3c8a81ec),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81142a),
	.w1(32'hbc5b3fd8),
	.w2(32'hbc5a2afe),
	.w3(32'hbbf8f8fd),
	.w4(32'h3c399256),
	.w5(32'hbbb6b42f),
	.w6(32'h3c4764e7),
	.w7(32'hbb3be759),
	.w8(32'hbc8d7f98),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48235d),
	.w1(32'hbc80efe2),
	.w2(32'hbbbc247a),
	.w3(32'hbbaa0a04),
	.w4(32'hbc85ac6e),
	.w5(32'hbc86c85f),
	.w6(32'hbc9004f3),
	.w7(32'h3d0ad13c),
	.w8(32'h3d726901),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97e69a),
	.w1(32'hbc08efd8),
	.w2(32'h3ab930b9),
	.w3(32'hbc73aa27),
	.w4(32'h3c23c451),
	.w5(32'h3c3c74f6),
	.w6(32'h3cc1fc83),
	.w7(32'hbb8eeac1),
	.w8(32'hbd1d0bfa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e8e3b),
	.w1(32'hb9161163),
	.w2(32'h3afac48c),
	.w3(32'h3c4f6736),
	.w4(32'hbae771d4),
	.w5(32'h3bd8d48b),
	.w6(32'hbd2137c8),
	.w7(32'h3c60b11c),
	.w8(32'h3c725039),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8adc8),
	.w1(32'hb94e0914),
	.w2(32'hbc081cf4),
	.w3(32'h3ba4ce9b),
	.w4(32'h39eff08b),
	.w5(32'hbb25f8d4),
	.w6(32'h3c215597),
	.w7(32'h3c629c29),
	.w8(32'hbbdd1cb6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93f782),
	.w1(32'hbbc030e6),
	.w2(32'h3baeedbd),
	.w3(32'h3c13ee16),
	.w4(32'hbc2b2ebb),
	.w5(32'h3b4e3d05),
	.w6(32'h3c0de76a),
	.w7(32'h3b95a7d8),
	.w8(32'h3bcdada1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c303848),
	.w1(32'h3c7a5fb3),
	.w2(32'h3bac6684),
	.w3(32'h3c7c5cd2),
	.w4(32'hbb07221c),
	.w5(32'h3aa9cfa8),
	.w6(32'hbc884f68),
	.w7(32'hbb9e7594),
	.w8(32'h3c9d6690),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37474),
	.w1(32'hbc1120e2),
	.w2(32'h3ba5b3ec),
	.w3(32'h3b5d2680),
	.w4(32'hbbfe53a0),
	.w5(32'h39acbbf2),
	.w6(32'h3a1a75d9),
	.w7(32'hbb7a4e71),
	.w8(32'hbc2afc3c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb39691),
	.w1(32'h3b22c828),
	.w2(32'h3bcd9643),
	.w3(32'h3b69fe70),
	.w4(32'hbb3af8e3),
	.w5(32'h3accb656),
	.w6(32'h3b9e6b75),
	.w7(32'h3bea956f),
	.w8(32'h3cf02237),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c323d6d),
	.w1(32'h3c4d12f9),
	.w2(32'hbc46a149),
	.w3(32'hbc38d5e1),
	.w4(32'hbc9d19b4),
	.w5(32'hbca58896),
	.w6(32'h3ca334e3),
	.w7(32'hbc9bc0ea),
	.w8(32'hbcc9b791),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952f690),
	.w1(32'hba740bbe),
	.w2(32'h3ab7bf9d),
	.w3(32'hbc6390a3),
	.w4(32'hbb92c1ae),
	.w5(32'hbc27da0f),
	.w6(32'hbc57813e),
	.w7(32'hba53c06d),
	.w8(32'h3bae5b89),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb9c24),
	.w1(32'h3ab3a412),
	.w2(32'hbbd5f3fc),
	.w3(32'hbcbf6dfe),
	.w4(32'hbbb3c8cf),
	.w5(32'hbc53eef5),
	.w6(32'h3a0449dc),
	.w7(32'hbc9d6d50),
	.w8(32'hbc127c05),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0a990),
	.w1(32'hba8d9408),
	.w2(32'hbb3b177f),
	.w3(32'hbb806cd7),
	.w4(32'h3a4b8e4a),
	.w5(32'hbbfca488),
	.w6(32'h3c286df8),
	.w7(32'hbc0f9811),
	.w8(32'hbc96c5b9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc547aaa),
	.w1(32'hbb6fbcdc),
	.w2(32'hbb3cea04),
	.w3(32'h3aca75f7),
	.w4(32'h3a7a96ee),
	.w5(32'h3bb5b11d),
	.w6(32'hbbfddbb9),
	.w7(32'h3c299389),
	.w8(32'h3c479e7d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01369e),
	.w1(32'h3b11cc3e),
	.w2(32'hbc467d81),
	.w3(32'h3b958065),
	.w4(32'hbc559c37),
	.w5(32'hbcf2f3e7),
	.w6(32'h3c12e2b7),
	.w7(32'h3b904c64),
	.w8(32'hbca3af34),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6053d6),
	.w1(32'hbb2c2aff),
	.w2(32'hbb9039ee),
	.w3(32'hbc94b58d),
	.w4(32'hba82ecc6),
	.w5(32'hbb8f239d),
	.w6(32'h3b903efc),
	.w7(32'hbc13794a),
	.w8(32'hbc84e5e0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd11221),
	.w1(32'h3bc88e2b),
	.w2(32'hbb392e86),
	.w3(32'h3b6f64cd),
	.w4(32'hbc14bf02),
	.w5(32'hbc0cf42e),
	.w6(32'hbbed88fd),
	.w7(32'h3ae246f2),
	.w8(32'h3c1acf7a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6e4e5),
	.w1(32'h39a9d7a0),
	.w2(32'hbb968698),
	.w3(32'hbbaaa393),
	.w4(32'hbb8ebf0e),
	.w5(32'h3c11c3c1),
	.w6(32'h3c5a976f),
	.w7(32'h3c959b16),
	.w8(32'h3bafcb03),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fc644),
	.w1(32'hbc6c046b),
	.w2(32'h3b0ffd82),
	.w3(32'h3bba18e3),
	.w4(32'hb9fee59e),
	.w5(32'h3bba06d3),
	.w6(32'hbaeccf35),
	.w7(32'h3c6dfc54),
	.w8(32'h3c7d49f6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3686f2),
	.w1(32'h3ab2c6ac),
	.w2(32'h3c4ea1ab),
	.w3(32'h3b98ab80),
	.w4(32'h3c9e3e59),
	.w5(32'h3c045a59),
	.w6(32'h3bee7c3b),
	.w7(32'hbd4bcfe0),
	.w8(32'hbda181a7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2bb57),
	.w1(32'h3cc122ff),
	.w2(32'hbbe46930),
	.w3(32'h3c7db989),
	.w4(32'hbb43affd),
	.w5(32'h39a5e3cf),
	.w6(32'hbd7f3ccb),
	.w7(32'hbba711dc),
	.w8(32'hbcd91bb6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f20c2),
	.w1(32'hbb4d0b8f),
	.w2(32'hbbf5fcb9),
	.w3(32'h3c654c7c),
	.w4(32'h3ba89322),
	.w5(32'h3a8bb252),
	.w6(32'hbc6f335e),
	.w7(32'hba737746),
	.w8(32'h39c1ba9a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81c249),
	.w1(32'hbc04fb74),
	.w2(32'h3a2aa221),
	.w3(32'h3b88e75a),
	.w4(32'h3aec5662),
	.w5(32'hbb51ccfc),
	.w6(32'h3b9e27e2),
	.w7(32'hbc6bebdc),
	.w8(32'hbcad02ae),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05b564),
	.w1(32'h3b9d755e),
	.w2(32'hbb77d2a3),
	.w3(32'h3abec62a),
	.w4(32'hbabcf106),
	.w5(32'h3c5c72d4),
	.w6(32'hbbe49472),
	.w7(32'h3ba0d885),
	.w8(32'h3c9f11b3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17433d),
	.w1(32'hbba485d0),
	.w2(32'hbae4032e),
	.w3(32'h3b6da89d),
	.w4(32'hbc2f8c87),
	.w5(32'hbc389169),
	.w6(32'h3c1a68d1),
	.w7(32'hb9ac6395),
	.w8(32'h3cad1a04),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c39e6),
	.w1(32'hbb1a6ec9),
	.w2(32'h3b60f7ef),
	.w3(32'hbca56c08),
	.w4(32'h3c3353b2),
	.w5(32'h3b951c72),
	.w6(32'h3c03d4c0),
	.w7(32'hba4c630e),
	.w8(32'hbbde58d2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a529c),
	.w1(32'h3c38cd80),
	.w2(32'hbb18092f),
	.w3(32'h3c211b48),
	.w4(32'h3b71ba87),
	.w5(32'hbbf9f3c1),
	.w6(32'hbb56a576),
	.w7(32'hba076acb),
	.w8(32'hbc025cbf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe363a7),
	.w1(32'hbc318461),
	.w2(32'h3bd6b718),
	.w3(32'h3b22b91e),
	.w4(32'hba807656),
	.w5(32'hbba97e5d),
	.w6(32'hba8804e9),
	.w7(32'hbc8cb8db),
	.w8(32'hbca4c563),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd31fb),
	.w1(32'hbafe34f1),
	.w2(32'hbc74c7d9),
	.w3(32'hbc019ae8),
	.w4(32'hbc54028c),
	.w5(32'hbcfa5c4e),
	.w6(32'hbc581a69),
	.w7(32'hbb66df6b),
	.w8(32'hbc812832),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc869161),
	.w1(32'hbc71321f),
	.w2(32'h3b9c3beb),
	.w3(32'hbce018ab),
	.w4(32'hbbcdb3ba),
	.w5(32'hbc26c00a),
	.w6(32'hbc9aaafd),
	.w7(32'h3be66b65),
	.w8(32'hbbc9b900),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9428cb),
	.w1(32'h3c19d41b),
	.w2(32'hba8816a0),
	.w3(32'hbb55aad4),
	.w4(32'hbafad9ae),
	.w5(32'hbbc0446a),
	.w6(32'hba8fc2c7),
	.w7(32'hbc41b000),
	.w8(32'hbc4bdd89),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5162f0),
	.w1(32'hba8b5ae7),
	.w2(32'h3b83bc2a),
	.w3(32'hbace882e),
	.w4(32'hb9a7c272),
	.w5(32'h3c546617),
	.w6(32'hba9f0bd0),
	.w7(32'hbc2508c0),
	.w8(32'hbc81f48e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3af737),
	.w1(32'h3b9c01c7),
	.w2(32'h3b6c5355),
	.w3(32'h3af89f80),
	.w4(32'hb9929c68),
	.w5(32'h3bdc77ee),
	.w6(32'hbc8121c2),
	.w7(32'hbb8fb302),
	.w8(32'h3c8cbd18),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80fd3f),
	.w1(32'hbc1ce55e),
	.w2(32'h3c18b4a9),
	.w3(32'hbbc8ceae),
	.w4(32'h3c047aa5),
	.w5(32'h3bb23450),
	.w6(32'h3bd8b024),
	.w7(32'hbc249cd3),
	.w8(32'hbcde47cf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc91890),
	.w1(32'h3c53969e),
	.w2(32'hb853a155),
	.w3(32'h3b3fff77),
	.w4(32'hbc81537a),
	.w5(32'hbadd1f0e),
	.w6(32'hbcfd8d10),
	.w7(32'h3bab2efb),
	.w8(32'h3c531d7d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f027),
	.w1(32'hbba597f8),
	.w2(32'hb9166856),
	.w3(32'hbbb7d898),
	.w4(32'hbb94371a),
	.w5(32'hbbc0cb26),
	.w6(32'hbc197a2b),
	.w7(32'hbc2696cb),
	.w8(32'hbc8b25e9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b829da3),
	.w1(32'h3c09e791),
	.w2(32'h393f85cb),
	.w3(32'h3adc24ba),
	.w4(32'hb6cac55b),
	.w5(32'h3752b320),
	.w6(32'hbbdf3924),
	.w7(32'hb901dfaf),
	.w8(32'hb8de751f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb33290),
	.w1(32'hbb9fb785),
	.w2(32'hbb2a461b),
	.w3(32'hbb8fdf50),
	.w4(32'hbba81d10),
	.w5(32'hbb8c1e8e),
	.w6(32'h3ab0b097),
	.w7(32'h3a6095e9),
	.w8(32'hbace5616),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb867649),
	.w1(32'hbb607bc4),
	.w2(32'hba8dcc02),
	.w3(32'hbabffdbf),
	.w4(32'hba27bade),
	.w5(32'h3acd6107),
	.w6(32'hba60a71f),
	.w7(32'h3928954b),
	.w8(32'h39af3a90),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab02e4b),
	.w1(32'hbaa1f61e),
	.w2(32'hbad0aade),
	.w3(32'hba1d6f32),
	.w4(32'hb9d0d9d7),
	.w5(32'hbaa39012),
	.w6(32'hbaa366eb),
	.w7(32'hbade2285),
	.w8(32'hbb1f186c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcfe1c),
	.w1(32'hbaa74c1c),
	.w2(32'hba1128f7),
	.w3(32'hba514161),
	.w4(32'h39e6f676),
	.w5(32'h3a639beb),
	.w6(32'hbaa689b6),
	.w7(32'hb98897c0),
	.w8(32'hb99d8958),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb222431),
	.w1(32'hb9163305),
	.w2(32'hbac8c664),
	.w3(32'h3902d1b7),
	.w4(32'hbb420aa5),
	.w5(32'hbac7b437),
	.w6(32'hbb2d5a15),
	.w7(32'hbbabe563),
	.w8(32'hbacb6e0d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbed96b),
	.w1(32'hbb835030),
	.w2(32'hbb53f019),
	.w3(32'hbb8ec512),
	.w4(32'hbba18717),
	.w5(32'hbaf6ceae),
	.w6(32'h3b01089c),
	.w7(32'hb95445af),
	.w8(32'hba8e03c8),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc810517),
	.w1(32'hbc0db636),
	.w2(32'hbc2d8c75),
	.w3(32'hbc15045f),
	.w4(32'hbb49af04),
	.w5(32'hbbb62721),
	.w6(32'hbb374b1b),
	.w7(32'hbab6d2c3),
	.w8(32'hbbff0319),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a9d9b),
	.w1(32'hbc430679),
	.w2(32'h37dc5768),
	.w3(32'hbc2ad0e1),
	.w4(32'hbc01969f),
	.w5(32'h3a287251),
	.w6(32'h37d09821),
	.w7(32'h3b3cc959),
	.w8(32'h3b8f1481),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9310cc),
	.w1(32'hbb4ca061),
	.w2(32'hb9f647a4),
	.w3(32'hbb9980db),
	.w4(32'hbb4fa883),
	.w5(32'hbb186f41),
	.w6(32'hbb8397fd),
	.w7(32'hbb82f01b),
	.w8(32'hbb201403),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b5bb7),
	.w1(32'hb63b311b),
	.w2(32'hba6b21b3),
	.w3(32'h3a5fc843),
	.w4(32'hba48938d),
	.w5(32'hbafbac92),
	.w6(32'hb9a84d22),
	.w7(32'hbb1904d3),
	.w8(32'hbb86dd84),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb179c5a),
	.w1(32'hbaef476d),
	.w2(32'hb86230b7),
	.w3(32'hbab1337e),
	.w4(32'hb99405b3),
	.w5(32'hb997a131),
	.w6(32'hbb5a703e),
	.w7(32'hb9db6f3f),
	.w8(32'hba11e743),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d7a70a),
	.w1(32'h399dffe1),
	.w2(32'hba51a388),
	.w3(32'h38737e63),
	.w4(32'hba0edd46),
	.w5(32'hba364cf8),
	.w6(32'hb95156f0),
	.w7(32'hba3bf908),
	.w8(32'hba71b32e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e66bb),
	.w1(32'h384282e9),
	.w2(32'h3b11f43e),
	.w3(32'h3a10d24f),
	.w4(32'h3a96e21c),
	.w5(32'h3ad64a29),
	.w6(32'h39c88570),
	.w7(32'h3b079cbe),
	.w8(32'h3b23ca47),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace49ff),
	.w1(32'h3b05158a),
	.w2(32'hbaf07448),
	.w3(32'h3b17eabf),
	.w4(32'hba2dee0d),
	.w5(32'hbabb6012),
	.w6(32'h3b297b80),
	.w7(32'hbb3bf806),
	.w8(32'hbb6e13fc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff80b8),
	.w1(32'hba3b3816),
	.w2(32'h3aeeb071),
	.w3(32'h3a2f1dc7),
	.w4(32'h3a9d4834),
	.w5(32'h390d0cef),
	.w6(32'hb9b6fe11),
	.w7(32'h3a43e5b3),
	.w8(32'hb966d748),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac90d79),
	.w1(32'h3b22787d),
	.w2(32'h3b212fb3),
	.w3(32'hbabe7c9a),
	.w4(32'h3a68d385),
	.w5(32'h3ae4f161),
	.w6(32'hbb80ca20),
	.w7(32'h3a1f6845),
	.w8(32'h3b10dbf0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4b62f),
	.w1(32'hbae7fa46),
	.w2(32'hbb68c2a9),
	.w3(32'hbb546d25),
	.w4(32'hbb9240f6),
	.w5(32'hbb3e3c36),
	.w6(32'h3af8ed5c),
	.w7(32'hbb0bbc74),
	.w8(32'hbb301b3f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28b960),
	.w1(32'hbb730682),
	.w2(32'hbb2d3e1b),
	.w3(32'h3aa1e666),
	.w4(32'h3902164b),
	.w5(32'hbad183c7),
	.w6(32'hbb1407ac),
	.w7(32'hbae863f2),
	.w8(32'hbb0ecdfe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e529d),
	.w1(32'hbb47be9e),
	.w2(32'hbb359f70),
	.w3(32'hba235838),
	.w4(32'hbb314b1e),
	.w5(32'hbb013346),
	.w6(32'hb778eb88),
	.w7(32'hbae74273),
	.w8(32'hbad7cf41),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95c69),
	.w1(32'hbb6403a6),
	.w2(32'h39f3a882),
	.w3(32'hbbb2f133),
	.w4(32'hbabd5417),
	.w5(32'h3a84a304),
	.w6(32'h37638bf2),
	.w7(32'h3acc28be),
	.w8(32'h3b0d09bb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17072d),
	.w1(32'h39873102),
	.w2(32'hb9c7a743),
	.w3(32'h3abb5c19),
	.w4(32'h38bd9cdd),
	.w5(32'h396cefcd),
	.w6(32'h3a94a897),
	.w7(32'hba235017),
	.w8(32'hba49b40e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b143e),
	.w1(32'h39f2f0ff),
	.w2(32'hb955a84b),
	.w3(32'h3a9d856d),
	.w4(32'h398aca8e),
	.w5(32'h382a6ca8),
	.w6(32'h3a0cafa0),
	.w7(32'hb834aec7),
	.w8(32'hb9a4af54),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba079b0e),
	.w1(32'hbaaa6ca8),
	.w2(32'h3b02d5f5),
	.w3(32'hba709a29),
	.w4(32'h3a544863),
	.w5(32'h3a631d2f),
	.w6(32'hba994b1b),
	.w7(32'h3ac64dc9),
	.w8(32'h3abf7509),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af1dd11),
	.w1(32'h3a7d1006),
	.w2(32'hba34a112),
	.w3(32'hba45159c),
	.w4(32'h3a398122),
	.w5(32'h3995409d),
	.w6(32'h392777f7),
	.w7(32'hb97e08ed),
	.w8(32'hba08379b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97428a),
	.w1(32'hbb066993),
	.w2(32'hbb181168),
	.w3(32'hb9c57f3c),
	.w4(32'hbab04952),
	.w5(32'hbb008a0c),
	.w6(32'hbacdfe5c),
	.w7(32'hbb311854),
	.w8(32'hbb2d2dab),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82d7c0),
	.w1(32'h3abfa43d),
	.w2(32'h3a85f13d),
	.w3(32'hba17dc13),
	.w4(32'h396c6580),
	.w5(32'h3af38eb9),
	.w6(32'hba066d72),
	.w7(32'h386b4c6d),
	.w8(32'h3ac66dcf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23d136),
	.w1(32'h3a88d5e7),
	.w2(32'h3ad6a1a7),
	.w3(32'hb9abf595),
	.w4(32'h3a7913ba),
	.w5(32'h3aaec7f8),
	.w6(32'hbb3d65de),
	.w7(32'hbb14ae7d),
	.w8(32'hba0401db),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afce1d3),
	.w1(32'h3af04aa8),
	.w2(32'h3a5db785),
	.w3(32'h3abc5b03),
	.w4(32'h3b24a29b),
	.w5(32'h3ab08425),
	.w6(32'hb8e59e63),
	.w7(32'h3a12e739),
	.w8(32'hba049ea4),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67db03),
	.w1(32'hbb115824),
	.w2(32'h3b22e0f6),
	.w3(32'hbbb060cb),
	.w4(32'hbbb8a88c),
	.w5(32'hbad7c766),
	.w6(32'hbacdd337),
	.w7(32'hbb597195),
	.w8(32'hbb28ab2e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57d015),
	.w1(32'hbb87c6e1),
	.w2(32'hba5cbd74),
	.w3(32'hbb8a1445),
	.w4(32'hbaad61e0),
	.w5(32'h3a80fa63),
	.w6(32'hbb8829b6),
	.w7(32'h391ad3ce),
	.w8(32'h39ac8c2d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f42ef),
	.w1(32'hba2db1bc),
	.w2(32'hb9fe7dd0),
	.w3(32'hb7fb0918),
	.w4(32'hb9bc0044),
	.w5(32'hb9927a46),
	.w6(32'hbaa628a9),
	.w7(32'hba85dbc9),
	.w8(32'hba15c12f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9ca05),
	.w1(32'h3a461b74),
	.w2(32'h3a6a8856),
	.w3(32'h3a4b2e13),
	.w4(32'h3b079a94),
	.w5(32'h3a4a18cb),
	.w6(32'hba63e306),
	.w7(32'h3ab7d561),
	.w8(32'h36012110),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf0b15),
	.w1(32'hba0ef5a9),
	.w2(32'h3a941e91),
	.w3(32'h395d7f31),
	.w4(32'hba74c9ab),
	.w5(32'h3a64bce5),
	.w6(32'h3a358ea4),
	.w7(32'h39861da4),
	.w8(32'h3b4308a0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b6b29c),
	.w1(32'h395b2949),
	.w2(32'h388a50af),
	.w3(32'hb853ffa8),
	.w4(32'h3aef6fed),
	.w5(32'h3a8767c3),
	.w6(32'hb9dcc065),
	.w7(32'h3b7ad6b6),
	.w8(32'h3bbf40e3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381947a3),
	.w1(32'h39aa3bc7),
	.w2(32'hb9721846),
	.w3(32'hbb340720),
	.w4(32'hba744461),
	.w5(32'hbb150efc),
	.w6(32'hb9f44f1a),
	.w7(32'h3a37427d),
	.w8(32'hba9b9e6d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b519e8d),
	.w1(32'h3b8c116c),
	.w2(32'h3b25bae8),
	.w3(32'h3ad78fbf),
	.w4(32'h3adf9c85),
	.w5(32'h3b0d407c),
	.w6(32'hba8bc68a),
	.w7(32'hbaa1dcf0),
	.w8(32'h394e9e69),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9512d66),
	.w1(32'hba1ad49f),
	.w2(32'hba12eb35),
	.w3(32'hba7741ad),
	.w4(32'h385ded2a),
	.w5(32'hb922f814),
	.w6(32'hb9cf7351),
	.w7(32'hb98bab2c),
	.w8(32'hb99eaf0e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f16a13),
	.w1(32'h36480186),
	.w2(32'hb9e1c2d6),
	.w3(32'hb9bc9b85),
	.w4(32'hbaa0b370),
	.w5(32'hbacdbcdc),
	.w6(32'h3a224d3b),
	.w7(32'hba4a2049),
	.w8(32'hbb0c49f1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915f45b),
	.w1(32'h39c3ce90),
	.w2(32'h3a614479),
	.w3(32'hb8bec865),
	.w4(32'h39bba851),
	.w5(32'h389c30be),
	.w6(32'hba3315c8),
	.w7(32'h3a904c3b),
	.w8(32'h3a47ccc2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a8bbd),
	.w1(32'h3aa519cb),
	.w2(32'hbb039f53),
	.w3(32'h3b0db7d4),
	.w4(32'h3901041c),
	.w5(32'hba9c563f),
	.w6(32'h3a498fbe),
	.w7(32'hbaacd238),
	.w8(32'hbae3e026),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53d313),
	.w1(32'hbb04062d),
	.w2(32'hbae4fb0b),
	.w3(32'hbb7ee95a),
	.w4(32'hbb0295ac),
	.w5(32'hbb043d00),
	.w6(32'hb9e363ab),
	.w7(32'h384d3a3d),
	.w8(32'hba871a4e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99564fb),
	.w1(32'hb9c9cb6a),
	.w2(32'h3a4ea059),
	.w3(32'hb98f2742),
	.w4(32'h3a52bf56),
	.w5(32'hb953fe17),
	.w6(32'hba0169bd),
	.w7(32'h3b0679b7),
	.w8(32'hb9d55e0e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab19000),
	.w1(32'h3a770acf),
	.w2(32'hb7f03477),
	.w3(32'h38b81e3b),
	.w4(32'hb8bea8e1),
	.w5(32'hb919a2e5),
	.w6(32'h3ad9a0c2),
	.w7(32'h39e5782e),
	.w8(32'h39168e8e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61f145),
	.w1(32'hbac9924f),
	.w2(32'hbaf49b1f),
	.w3(32'h3781061b),
	.w4(32'h39318924),
	.w5(32'hb914b807),
	.w6(32'hbb7cd2cc),
	.w7(32'hbb7a645b),
	.w8(32'hbb1cbd83),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198b6d),
	.w1(32'hbb1cd09b),
	.w2(32'hbabcf123),
	.w3(32'hba389f00),
	.w4(32'hb9b64671),
	.w5(32'hb95efea9),
	.w6(32'hba325da6),
	.w7(32'hba357e29),
	.w8(32'hbb08bad0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9bf67),
	.w1(32'hba66f803),
	.w2(32'hba2f659b),
	.w3(32'hb9611aff),
	.w4(32'h39f47723),
	.w5(32'h391fd5a8),
	.w6(32'hbab6ebb4),
	.w7(32'hba1289f5),
	.w8(32'hba5f91de),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cb2ec),
	.w1(32'h3aad33a9),
	.w2(32'h3a879932),
	.w3(32'h3a96b893),
	.w4(32'h3b2b5172),
	.w5(32'h3ae9258c),
	.w6(32'hba38ff09),
	.w7(32'h3ad04e3b),
	.w8(32'h3a0aa452),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad708a1),
	.w1(32'h3aa81ca7),
	.w2(32'h3a21d803),
	.w3(32'hba7e15ee),
	.w4(32'h3a39f863),
	.w5(32'h38dd3b68),
	.w6(32'h3ac7a448),
	.w7(32'h3a37d9ce),
	.w8(32'hb9b72bbf),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb682),
	.w1(32'hbb0ea85f),
	.w2(32'hba03cdb4),
	.w3(32'hbaaf98de),
	.w4(32'hb948a259),
	.w5(32'hb8b94324),
	.w6(32'hbb4a80e3),
	.w7(32'h3a552ae9),
	.w8(32'h3adb3278),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf06f0f),
	.w1(32'hb907f23b),
	.w2(32'hba38c934),
	.w3(32'hb9b06e1c),
	.w4(32'h39c411a2),
	.w5(32'h38b95401),
	.w6(32'h392f86af),
	.w7(32'h3a5828a0),
	.w8(32'h39eb951e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa0737),
	.w1(32'hbac5f883),
	.w2(32'hbb092a9b),
	.w3(32'h390fdf24),
	.w4(32'hbb171f43),
	.w5(32'hbb2921bf),
	.w6(32'h38f69c70),
	.w7(32'hbac3f7a3),
	.w8(32'hbab6ab70),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule