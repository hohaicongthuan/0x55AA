module layer_10_featuremap_77(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92578fc),
	.w1(32'hb9bfd893),
	.w2(32'hbacf5894),
	.w3(32'hbb18eeaa),
	.w4(32'hbb35d4b1),
	.w5(32'hbbae7396),
	.w6(32'hbbd19f51),
	.w7(32'hbb0f3efe),
	.w8(32'hbc0564cd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6e427),
	.w1(32'h3c2202b2),
	.w2(32'h39c8a04a),
	.w3(32'h3a23be1c),
	.w4(32'h3b5c90d0),
	.w5(32'hba45f1a1),
	.w6(32'h3aa54160),
	.w7(32'h3ba0136d),
	.w8(32'hb99a18e1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5570a),
	.w1(32'hb97634e0),
	.w2(32'hbb9ced91),
	.w3(32'hbb227a79),
	.w4(32'h3b4cd8dd),
	.w5(32'hbb31086f),
	.w6(32'hbbd65211),
	.w7(32'h3bafa0ee),
	.w8(32'hbb4c10e7),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba073871),
	.w1(32'h3b1471d8),
	.w2(32'hbc204c16),
	.w3(32'h39730c8f),
	.w4(32'hbad77684),
	.w5(32'hbb962fa7),
	.w6(32'hbb56b1ee),
	.w7(32'hbbef0324),
	.w8(32'hbb44a591),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60f3c7),
	.w1(32'h3aa08883),
	.w2(32'hbb461304),
	.w3(32'hba747814),
	.w4(32'hbb65bc42),
	.w5(32'h3a9fb183),
	.w6(32'hbb93d7d3),
	.w7(32'hbb6adb28),
	.w8(32'h3a71c537),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c6010),
	.w1(32'hbb566276),
	.w2(32'h3bf838d1),
	.w3(32'h3b940908),
	.w4(32'h3aa44c36),
	.w5(32'h3b18df68),
	.w6(32'h3a94a03a),
	.w7(32'h3b06a3b1),
	.w8(32'hbbdbcb0e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5ea94a),
	.w1(32'h3c7d927c),
	.w2(32'hbbac105e),
	.w3(32'h3c06c31f),
	.w4(32'h3bfeedaa),
	.w5(32'hbbbc8aca),
	.w6(32'hbb844314),
	.w7(32'hbb9e69ce),
	.w8(32'hbbf598c8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17d117),
	.w1(32'hbb333df7),
	.w2(32'hbbfb9044),
	.w3(32'hbc65bd28),
	.w4(32'hbbf2917f),
	.w5(32'hbb8a8f26),
	.w6(32'hbc829f15),
	.w7(32'hbc69ec99),
	.w8(32'hbc3b0688),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2e71b),
	.w1(32'h3b2904f3),
	.w2(32'h3abca43c),
	.w3(32'h3a0a1ec4),
	.w4(32'hbae090b9),
	.w5(32'hba988a2b),
	.w6(32'hba45d044),
	.w7(32'h395c507f),
	.w8(32'hbb9dfa8f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a062e9e),
	.w1(32'hbb808829),
	.w2(32'h3b589be1),
	.w3(32'h3aa618c8),
	.w4(32'hbb8bda16),
	.w5(32'h3b2e001e),
	.w6(32'hbb66b157),
	.w7(32'hbb84bbd6),
	.w8(32'h3b095570),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36634d),
	.w1(32'h3b149b1b),
	.w2(32'h39f9473e),
	.w3(32'h3b146d31),
	.w4(32'h3b3aed1f),
	.w5(32'hbace661d),
	.w6(32'h3b176e95),
	.w7(32'h3b09363d),
	.w8(32'hbb65e10b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8addc2),
	.w1(32'h3bbf6254),
	.w2(32'h3a50bea4),
	.w3(32'hba623f17),
	.w4(32'hbacf68f7),
	.w5(32'hba743caa),
	.w6(32'hbb1b1343),
	.w7(32'hbbd8c70a),
	.w8(32'hbb9c2d8c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa24c69),
	.w1(32'hbb9d6b28),
	.w2(32'hba95594a),
	.w3(32'hba69c148),
	.w4(32'hbb9e5f47),
	.w5(32'hbb9d7374),
	.w6(32'hbb6a5444),
	.w7(32'hbbbfd43b),
	.w8(32'hbb8ef65d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e8b54),
	.w1(32'hbb46b6ab),
	.w2(32'hbbf58a2b),
	.w3(32'hbbf4fd96),
	.w4(32'hbafee030),
	.w5(32'hbc1851bb),
	.w6(32'hbbb65e90),
	.w7(32'hbad15e84),
	.w8(32'hba9700e9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8adb09),
	.w1(32'hbc0b5342),
	.w2(32'hbbdb02fc),
	.w3(32'h3a30f4cc),
	.w4(32'h3a615aad),
	.w5(32'hbb3dbbf3),
	.w6(32'h3bbdfed4),
	.w7(32'h3ab181ae),
	.w8(32'hba650790),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9047b5),
	.w1(32'h39a6bc82),
	.w2(32'h3bbf57fa),
	.w3(32'hbb0dfc27),
	.w4(32'hba59e20b),
	.w5(32'h3bad13c9),
	.w6(32'hbb2e6c3a),
	.w7(32'hba5f5419),
	.w8(32'hba610857),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7dc14),
	.w1(32'h3bde8e6c),
	.w2(32'h3b989728),
	.w3(32'h3b9cd3da),
	.w4(32'h3bcf9ddd),
	.w5(32'h3b8f9252),
	.w6(32'h3b26ab93),
	.w7(32'h3b3afdd3),
	.w8(32'h3b8a49b5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0359f5),
	.w1(32'hbc525669),
	.w2(32'hbc790686),
	.w3(32'hbbebfbb4),
	.w4(32'hbc518125),
	.w5(32'hbc084328),
	.w6(32'hbc0b0963),
	.w7(32'hbc7a731c),
	.w8(32'hbc50588d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9d2a),
	.w1(32'hbb696a03),
	.w2(32'hbb8b61e8),
	.w3(32'hbb841a53),
	.w4(32'hb9e426da),
	.w5(32'hbbc8212f),
	.w6(32'hbbb01a37),
	.w7(32'hbbc8383c),
	.w8(32'hbbd0700c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b2af4),
	.w1(32'hbaa93263),
	.w2(32'h38a97fa3),
	.w3(32'hbac8b4bf),
	.w4(32'hbb5a8e7f),
	.w5(32'h3b08861d),
	.w6(32'hbb000f60),
	.w7(32'hbb8c02fa),
	.w8(32'h3b3ee048),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29c791),
	.w1(32'h3b28c6bf),
	.w2(32'hbb311d06),
	.w3(32'h3b463e2a),
	.w4(32'h3a34fe4a),
	.w5(32'h3a9b983d),
	.w6(32'h3ad5d4fe),
	.w7(32'hbaa2fc18),
	.w8(32'h39a13a43),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea52b),
	.w1(32'h3b267088),
	.w2(32'h3aeaaf04),
	.w3(32'h3a88362d),
	.w4(32'h3bc3c054),
	.w5(32'hb9cdbe77),
	.w6(32'h3b2b4128),
	.w7(32'hbb057e45),
	.w8(32'h3af3f261),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc675244),
	.w1(32'hbc91f291),
	.w2(32'hbcb0119e),
	.w3(32'hbc4e5f1a),
	.w4(32'hbbf25135),
	.w5(32'hbc70965b),
	.w6(32'hbc8e8270),
	.w7(32'hbc86ff3a),
	.w8(32'hbc8d4893),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f3191),
	.w1(32'hbb96c9d4),
	.w2(32'h3af9f7d7),
	.w3(32'h3b75ffc1),
	.w4(32'h3aa280bc),
	.w5(32'h3b50e9fd),
	.w6(32'h3b9adf42),
	.w7(32'h3b57bebe),
	.w8(32'h3aa497f6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b576433),
	.w1(32'h3bf6aa77),
	.w2(32'hbaf100a9),
	.w3(32'h3bc85281),
	.w4(32'h3bfe6617),
	.w5(32'h3b169f0f),
	.w6(32'h3b7073af),
	.w7(32'h3a48e0c8),
	.w8(32'hbb8528f2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea3f2e),
	.w1(32'hbbfe9284),
	.w2(32'hbaf16b6a),
	.w3(32'hbb31b516),
	.w4(32'h3a944f39),
	.w5(32'hbb88c821),
	.w6(32'hbb1a503f),
	.w7(32'h39816390),
	.w8(32'hbbbe7236),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e1d8c),
	.w1(32'h3b149032),
	.w2(32'h38014fad),
	.w3(32'hbb2290fd),
	.w4(32'hbb8f6f9c),
	.w5(32'hbab0d208),
	.w6(32'hbb868515),
	.w7(32'hbb6dfd41),
	.w8(32'h3aa34b14),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02231a),
	.w1(32'h3b13f331),
	.w2(32'h392a5265),
	.w3(32'h3b17d82f),
	.w4(32'h3a1d11d0),
	.w5(32'hba408c4a),
	.w6(32'h3b975b71),
	.w7(32'h3b13d092),
	.w8(32'h3b78f169),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f7ce5),
	.w1(32'h3ca13e1b),
	.w2(32'hbbe69a76),
	.w3(32'hbae98eb6),
	.w4(32'h3aa2535a),
	.w5(32'h3cd6a667),
	.w6(32'h3bc4f81d),
	.w7(32'h3c42ea2c),
	.w8(32'hbca734fd),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805a2e),
	.w1(32'hbbf704c3),
	.w2(32'hbb6cd0f1),
	.w3(32'h3d0d98a3),
	.w4(32'h3c13798d),
	.w5(32'hba57133f),
	.w6(32'hbab8084e),
	.w7(32'h3c6e79b4),
	.w8(32'hba4ed820),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37702),
	.w1(32'hbbb2c1e8),
	.w2(32'hbc0f1e81),
	.w3(32'hbb72e12e),
	.w4(32'hbbb9296f),
	.w5(32'h3c1418dc),
	.w6(32'hbb3f6cb8),
	.w7(32'hbb07651e),
	.w8(32'hbc0403fa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6deaed),
	.w1(32'hbb4e21e5),
	.w2(32'hbc8bb438),
	.w3(32'h3c825d54),
	.w4(32'h3b1fae14),
	.w5(32'h3c1738cc),
	.w6(32'h3b67d402),
	.w7(32'h3c005938),
	.w8(32'h385820bb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb636a42),
	.w1(32'h3b0edf21),
	.w2(32'hba10b3d4),
	.w3(32'h3bc86c8e),
	.w4(32'hbb4ffdeb),
	.w5(32'hbadde503),
	.w6(32'h3c2f65ec),
	.w7(32'h3b956c3a),
	.w8(32'h3b18c490),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d04e),
	.w1(32'h3b2c71c9),
	.w2(32'h3ba87b4a),
	.w3(32'hbb39f55b),
	.w4(32'hbb01e9aa),
	.w5(32'h3b3da8f2),
	.w6(32'h3bedf934),
	.w7(32'h3b54da86),
	.w8(32'hb9d991dd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a14f6),
	.w1(32'h3c1df298),
	.w2(32'h3b2fcea4),
	.w3(32'h3ad752a7),
	.w4(32'hbc26eb79),
	.w5(32'h39dca3a3),
	.w6(32'h3ca6921d),
	.w7(32'h3c883a99),
	.w8(32'h3b346ca3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab07b1),
	.w1(32'h3b0f9ebc),
	.w2(32'hbc108031),
	.w3(32'hbaf8b1ca),
	.w4(32'hba9624e5),
	.w5(32'h3be300e3),
	.w6(32'h3b94de0e),
	.w7(32'h3b1e9936),
	.w8(32'hbb1342cb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df754),
	.w1(32'hbc477635),
	.w2(32'hbb9b2d2a),
	.w3(32'h3af0b082),
	.w4(32'hbbb0416e),
	.w5(32'hbc06e678),
	.w6(32'h3b9e9faa),
	.w7(32'h3c26e944),
	.w8(32'hbbe5acb0),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25588b),
	.w1(32'h3c47f9ef),
	.w2(32'h3c064c1a),
	.w3(32'h3b65f4e7),
	.w4(32'h3b72f041),
	.w5(32'hbbef2baa),
	.w6(32'h3c427a2e),
	.w7(32'h3c0ccfec),
	.w8(32'h3d29bd28),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3231e5),
	.w1(32'h3d13b308),
	.w2(32'hba1343f4),
	.w3(32'hbcb67cdf),
	.w4(32'hbb8560c6),
	.w5(32'h3c13dc41),
	.w6(32'h3d421962),
	.w7(32'h3aa5ff95),
	.w8(32'hbb506dd9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69fb7d),
	.w1(32'hbc491668),
	.w2(32'hbb48f7df),
	.w3(32'h3c5eac79),
	.w4(32'h3c460f97),
	.w5(32'hbb009c21),
	.w6(32'hbcd0fc3c),
	.w7(32'h3ac58b26),
	.w8(32'h3bcb37cd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4c352),
	.w1(32'h3a4b052c),
	.w2(32'h3ba3616b),
	.w3(32'h39fcd7ea),
	.w4(32'hb9593598),
	.w5(32'hbc7e3480),
	.w6(32'h3ba8f338),
	.w7(32'h3b8101b0),
	.w8(32'hb9498f02),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a344e),
	.w1(32'h3c4e80a8),
	.w2(32'h3c9a1698),
	.w3(32'hbca5252f),
	.w4(32'hb9f0570e),
	.w5(32'h3b905e7e),
	.w6(32'hbc03b4ce),
	.w7(32'hbc81ec1a),
	.w8(32'hbaa86613),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586939),
	.w1(32'hba28611a),
	.w2(32'h3aa19cfc),
	.w3(32'h3ccb28a4),
	.w4(32'h3cdbf58a),
	.w5(32'hbb165aa0),
	.w6(32'hbb367601),
	.w7(32'hbc09c0d4),
	.w8(32'hbb635eaa),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cfbd5),
	.w1(32'hbb2e7e4a),
	.w2(32'h3b433afd),
	.w3(32'hbbd8cac5),
	.w4(32'hbb811e19),
	.w5(32'h3ba49b3b),
	.w6(32'hbb5b9ccb),
	.w7(32'hbbae101f),
	.w8(32'hbc99388b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7590ad),
	.w1(32'hbadda93b),
	.w2(32'hbc336f98),
	.w3(32'h3bed2825),
	.w4(32'h3c66434d),
	.w5(32'h3ca38d0b),
	.w6(32'hbc08ae91),
	.w7(32'h3b6b83d7),
	.w8(32'hbaa9c83c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52491d),
	.w1(32'h3bc872ed),
	.w2(32'h3b2f54d7),
	.w3(32'h3bce2b02),
	.w4(32'hbc9b39f8),
	.w5(32'hbc07ea3c),
	.w6(32'h3cc266fd),
	.w7(32'h3cc792bb),
	.w8(32'h3af1dd1f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38ef57),
	.w1(32'hbba24e9f),
	.w2(32'h3cadb023),
	.w3(32'hbba8f3e8),
	.w4(32'hbba6a212),
	.w5(32'hb7354632),
	.w6(32'hbbd8dbc7),
	.w7(32'hbc030f0a),
	.w8(32'h3a70d3dc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03cb38),
	.w1(32'hbc356ab8),
	.w2(32'hbc803d7f),
	.w3(32'hbc40b0fc),
	.w4(32'hbb233b3b),
	.w5(32'hbc39bd26),
	.w6(32'hbc8597c8),
	.w7(32'hbcade7b2),
	.w8(32'hbcb223f3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba210dfe),
	.w1(32'hbad80cd7),
	.w2(32'hbc13676b),
	.w3(32'hbae5d8e1),
	.w4(32'hbb7ac7c5),
	.w5(32'hbb5fd08a),
	.w6(32'hbb82712f),
	.w7(32'hbba4c6ee),
	.w8(32'h3c86667c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46fe0c),
	.w1(32'h3b091ca8),
	.w2(32'hbc089073),
	.w3(32'hbbcbbfeb),
	.w4(32'h3b88bb6b),
	.w5(32'h3c1cabd1),
	.w6(32'h3ccc2032),
	.w7(32'h3bedfc78),
	.w8(32'hba5500f2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ca44),
	.w1(32'h3c34f41a),
	.w2(32'hbc0d8e00),
	.w3(32'h3a1d88f5),
	.w4(32'hbba5654d),
	.w5(32'h3ca1b964),
	.w6(32'h3c1bb586),
	.w7(32'h3bc938b8),
	.w8(32'h3b92bfea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefd01b),
	.w1(32'h3bbd8e83),
	.w2(32'hbc3496ab),
	.w3(32'h3becfbbf),
	.w4(32'h3b09dec8),
	.w5(32'hbb238546),
	.w6(32'hba529504),
	.w7(32'h3aba03bc),
	.w8(32'hba940d1d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b2e07),
	.w1(32'h3b9e2d24),
	.w2(32'hbad8ecc7),
	.w3(32'hbc2a83cd),
	.w4(32'hbc9dc36b),
	.w5(32'h3a02c1e1),
	.w6(32'h3b617184),
	.w7(32'hbb3f0d14),
	.w8(32'hbc3cda6b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fdad1),
	.w1(32'hbcbb6054),
	.w2(32'h3ba8afe4),
	.w3(32'h3ba75f7f),
	.w4(32'h3a0faa9c),
	.w5(32'hbbad2692),
	.w6(32'hbc568c69),
	.w7(32'hbba3b48a),
	.w8(32'hbc9b0185),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb3cd),
	.w1(32'hbc2da2ea),
	.w2(32'hbca4ba2f),
	.w3(32'h3caa96ac),
	.w4(32'h3cdfaf57),
	.w5(32'h3cf6d49a),
	.w6(32'hbc39a694),
	.w7(32'h3b33d5e5),
	.w8(32'hbc86e0dd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b29d1),
	.w1(32'hbb8d1ff8),
	.w2(32'hbc4d44dc),
	.w3(32'h3d08ea17),
	.w4(32'h3bd21527),
	.w5(32'h3c07a3fe),
	.w6(32'h3c0bb640),
	.w7(32'h3caf2d36),
	.w8(32'hbc2a25fe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58c0fa),
	.w1(32'h3bb3abf0),
	.w2(32'h3bc4a749),
	.w3(32'hbbb1cbb4),
	.w4(32'hbcb6e5e3),
	.w5(32'h3b20886f),
	.w6(32'h3c7a1060),
	.w7(32'h3c5ce29c),
	.w8(32'h3bdfe6ff),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab0d3),
	.w1(32'hbbfbd29e),
	.w2(32'h3ac336d5),
	.w3(32'hbac74c08),
	.w4(32'hbb08d40f),
	.w5(32'h3affa73d),
	.w6(32'hbbb9c9ae),
	.w7(32'hbb7c75ab),
	.w8(32'h3acac97a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386c1394),
	.w1(32'h3b9dee3a),
	.w2(32'h3c6c87c7),
	.w3(32'hbb489920),
	.w4(32'h3b926b82),
	.w5(32'hbb2e3397),
	.w6(32'h3a7ce53c),
	.w7(32'h3bf731d3),
	.w8(32'h3bf20b80),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c2619),
	.w1(32'hbaa4937d),
	.w2(32'h3ae55880),
	.w3(32'hb913d00b),
	.w4(32'h3baa48cd),
	.w5(32'h3a6d5721),
	.w6(32'hbb2e9c61),
	.w7(32'hbc003a9a),
	.w8(32'hbb801096),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53debd),
	.w1(32'hbc2196d3),
	.w2(32'hbb60ca05),
	.w3(32'h39abc37c),
	.w4(32'h3bc240fd),
	.w5(32'h3bb634e6),
	.w6(32'hbc139ad1),
	.w7(32'hbc17c16a),
	.w8(32'hbab41c1a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb551c40),
	.w1(32'hbb60da26),
	.w2(32'h3bec007a),
	.w3(32'h3bc92964),
	.w4(32'h3c8487ad),
	.w5(32'hbc3a013a),
	.w6(32'h39d5b6f6),
	.w7(32'h3c038f00),
	.w8(32'h3a3ad3a6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a285dc5),
	.w1(32'hbb78a09e),
	.w2(32'h3c1140e8),
	.w3(32'hbbebb7db),
	.w4(32'h3ba05a8d),
	.w5(32'hbba69618),
	.w6(32'hbc25ee6b),
	.w7(32'hbc012a2f),
	.w8(32'h3bae280b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd555df),
	.w1(32'h3b0f7827),
	.w2(32'hbc1265a3),
	.w3(32'hbc2a1b8e),
	.w4(32'hbbc90ad5),
	.w5(32'hbbd5aecf),
	.w6(32'hbb05606c),
	.w7(32'hbbabb737),
	.w8(32'hbb788c08),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5375be),
	.w1(32'hbc76e775),
	.w2(32'hbb5114f6),
	.w3(32'hbcf81068),
	.w4(32'hbc89421e),
	.w5(32'h3b3e50e3),
	.w6(32'hbc515009),
	.w7(32'hbc2baaa7),
	.w8(32'h3c29c542),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b22c5),
	.w1(32'h3ad01b66),
	.w2(32'hbafbbafc),
	.w3(32'hba1a5551),
	.w4(32'hbb2c3b08),
	.w5(32'hbb005977),
	.w6(32'h3c42663f),
	.w7(32'h3c1890ce),
	.w8(32'hba6f2654),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998d174),
	.w1(32'h3b0c6ed2),
	.w2(32'hbbe46843),
	.w3(32'hbb88b8b1),
	.w4(32'hbac9b049),
	.w5(32'hbb0b704b),
	.w6(32'h3a6090f6),
	.w7(32'hb9e0f7e8),
	.w8(32'hbc167383),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59b7d),
	.w1(32'h398e1b09),
	.w2(32'hbaf88a37),
	.w3(32'hbc094c15),
	.w4(32'hbc6fbbfc),
	.w5(32'h3b9f0285),
	.w6(32'h3b5ac1db),
	.w7(32'hb92d03c8),
	.w8(32'h39790fb6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69cb57),
	.w1(32'h3c17f8ae),
	.w2(32'hbbd8d948),
	.w3(32'hbc0cb034),
	.w4(32'hbb2945ba),
	.w5(32'hbc0df13c),
	.w6(32'hb82f1445),
	.w7(32'h3b76e38b),
	.w8(32'hbc561205),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b907ad5),
	.w1(32'h3b2d70c5),
	.w2(32'h3b861840),
	.w3(32'h3bcf71c7),
	.w4(32'h3ab0a07f),
	.w5(32'h3b96e469),
	.w6(32'h3a913874),
	.w7(32'hba11facb),
	.w8(32'h3bae0d16),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7e5b6),
	.w1(32'h3af8657e),
	.w2(32'hbab69834),
	.w3(32'hbb93d5e2),
	.w4(32'hbb1eeb2f),
	.w5(32'h3c354bbb),
	.w6(32'hbb1e1f9f),
	.w7(32'hbc185b79),
	.w8(32'hbbaf5dd8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfde6df),
	.w1(32'hbb21a613),
	.w2(32'h3c02a6e3),
	.w3(32'h3bf9f997),
	.w4(32'hbbc4f522),
	.w5(32'h3c148bbb),
	.w6(32'hbc129892),
	.w7(32'h38f5affc),
	.w8(32'h3c29b08c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a77ed),
	.w1(32'h3c6ba78b),
	.w2(32'h3ba2b55e),
	.w3(32'hbbdeb6be),
	.w4(32'hba8b4244),
	.w5(32'hbc1e88da),
	.w6(32'h3c13525d),
	.w7(32'h3c0d3a9e),
	.w8(32'hbc205866),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54aba7),
	.w1(32'hbc9863a3),
	.w2(32'h3ade89b0),
	.w3(32'h3c00c3cb),
	.w4(32'h3bd79dbb),
	.w5(32'h3b803c7f),
	.w6(32'hbc883de7),
	.w7(32'hbc66a4af),
	.w8(32'hbaf93c33),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2105e),
	.w1(32'hb9e25789),
	.w2(32'h3b800907),
	.w3(32'h3aa4932a),
	.w4(32'hbb219114),
	.w5(32'h3bd3e55f),
	.w6(32'hbb24fa3b),
	.w7(32'h3a132fc5),
	.w8(32'h3a292d18),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61773f),
	.w1(32'hbad68528),
	.w2(32'hbc27dc68),
	.w3(32'hbbeff7e3),
	.w4(32'hbbe06b1d),
	.w5(32'hbc01dfa2),
	.w6(32'h3b446e7b),
	.w7(32'h3b765614),
	.w8(32'hbc0a62ae),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc580a94),
	.w1(32'hbc01ea5f),
	.w2(32'hbc2f9436),
	.w3(32'hbccee752),
	.w4(32'hbca412f9),
	.w5(32'hbc46665e),
	.w6(32'hbc69943d),
	.w7(32'hbc157e7b),
	.w8(32'hbc43894e),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044b53),
	.w1(32'h39aecdeb),
	.w2(32'h3a4e648f),
	.w3(32'hbc34f3c2),
	.w4(32'hbba7607b),
	.w5(32'h3b9f1861),
	.w6(32'h3b58df9c),
	.w7(32'h3ba8d45a),
	.w8(32'hbb7378d6),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89703d),
	.w1(32'hbc5a63df),
	.w2(32'hba9c31ae),
	.w3(32'h3c2ddac8),
	.w4(32'h3c0ae94b),
	.w5(32'hbbbb61f4),
	.w6(32'hbb78afb5),
	.w7(32'hbbd9f345),
	.w8(32'hba802a5d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91279c),
	.w1(32'hba17d708),
	.w2(32'h3abfea5a),
	.w3(32'h3b8fef58),
	.w4(32'h398233ae),
	.w5(32'h3b034734),
	.w6(32'hb9d94466),
	.w7(32'hbb2e800a),
	.w8(32'h39d1253a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac0f30),
	.w1(32'h3b8e1a57),
	.w2(32'hba89b0e5),
	.w3(32'hbb9ee0c7),
	.w4(32'hbb77de35),
	.w5(32'h39730b81),
	.w6(32'h3ba84716),
	.w7(32'h3ab99bc6),
	.w8(32'h3bbbe0b7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eeb8b),
	.w1(32'hbaf21f44),
	.w2(32'hbc310c21),
	.w3(32'hbc119518),
	.w4(32'hbbf785da),
	.w5(32'hbc5816ea),
	.w6(32'hb96155d7),
	.w7(32'h381b7f83),
	.w8(32'hbbcfdfda),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9761b7),
	.w1(32'hbc09977a),
	.w2(32'hbc86b7f6),
	.w3(32'hbc3e8d69),
	.w4(32'hbc180c5c),
	.w5(32'hbc988380),
	.w6(32'h3bce137e),
	.w7(32'h3c40b16a),
	.w8(32'hbc2ec88b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15a836),
	.w1(32'hbb6d6ba5),
	.w2(32'h3b19bd55),
	.w3(32'hbc4be8f8),
	.w4(32'hbb062fac),
	.w5(32'h3a5f5149),
	.w6(32'hbb41d43a),
	.w7(32'hbc2222e6),
	.w8(32'h3b649b70),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7515ad),
	.w1(32'h3b22ad4d),
	.w2(32'h3c17602f),
	.w3(32'hbb48827e),
	.w4(32'h3c038e87),
	.w5(32'h3b0519fd),
	.w6(32'h3ae6b691),
	.w7(32'h3af3b3eb),
	.w8(32'hbbb2f57f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b563bf2),
	.w1(32'h3bdcbc78),
	.w2(32'h3b6ab936),
	.w3(32'hbc60bf89),
	.w4(32'h3aa8c636),
	.w5(32'h3b9eb876),
	.w6(32'h3b73e643),
	.w7(32'h3b13d9d8),
	.w8(32'h3ba41f3a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ae26c),
	.w1(32'h3bb9e6c4),
	.w2(32'h3bbe3334),
	.w3(32'h3a58a590),
	.w4(32'h3be564f4),
	.w5(32'h3b9e703c),
	.w6(32'h3a8295a6),
	.w7(32'h3ba5c583),
	.w8(32'h3b7aa351),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5a374),
	.w1(32'h3b42f565),
	.w2(32'hbc148301),
	.w3(32'h3b009bdd),
	.w4(32'h3ade0d46),
	.w5(32'hbbacebca),
	.w6(32'h3b135017),
	.w7(32'h3ba18c50),
	.w8(32'hbc296d80),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcef8ce),
	.w1(32'hbbff2f52),
	.w2(32'hbcbf588a),
	.w3(32'hbc854315),
	.w4(32'hbc95010a),
	.w5(32'h3b8b0491),
	.w6(32'h3b1c9f4a),
	.w7(32'hbc088865),
	.w8(32'hbbe5b2f0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd3bdb8),
	.w1(32'hbc09dd9c),
	.w2(32'hbc99b4d6),
	.w3(32'hbc866bdb),
	.w4(32'hbca89404),
	.w5(32'hbc827e97),
	.w6(32'hbc8996ed),
	.w7(32'hbc34897e),
	.w8(32'hbcd83155),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b7a7),
	.w1(32'h3bca954e),
	.w2(32'h3ba3933b),
	.w3(32'hbb0433b4),
	.w4(32'hbbad32a3),
	.w5(32'h3a84d55a),
	.w6(32'h3acb979c),
	.w7(32'h3a827485),
	.w8(32'h3c0fbfc2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a594d69),
	.w1(32'hbb131dc7),
	.w2(32'hbb32426f),
	.w3(32'hbb8d5dcb),
	.w4(32'h3a08a631),
	.w5(32'hbb45b72f),
	.w6(32'hbbbe19b6),
	.w7(32'hbbd11fb2),
	.w8(32'hbb82b5f3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a09e2),
	.w1(32'h3a1d70d2),
	.w2(32'h3b6ad498),
	.w3(32'h3a92020c),
	.w4(32'h3b83f089),
	.w5(32'h3aafcc3e),
	.w6(32'hb9be0a95),
	.w7(32'h3aeb257a),
	.w8(32'h3b60c605),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb941b63),
	.w1(32'hbba2c9de),
	.w2(32'h3b40abe6),
	.w3(32'hbb2a0c3c),
	.w4(32'hbb1d8b34),
	.w5(32'h3ba34677),
	.w6(32'hbbd8be22),
	.w7(32'hbc2167a7),
	.w8(32'h3b406b96),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3b89c),
	.w1(32'h3b9aef58),
	.w2(32'h3b7fc00d),
	.w3(32'hba2e1ac1),
	.w4(32'hb8a55f02),
	.w5(32'hbc205aaa),
	.w6(32'h3c883509),
	.w7(32'h3c208b03),
	.w8(32'h3b8b436d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c0475),
	.w1(32'h3b73c980),
	.w2(32'hbbf6a4e3),
	.w3(32'hbc3d8eaf),
	.w4(32'hb94835ec),
	.w5(32'hbb7eb52c),
	.w6(32'h3bade54f),
	.w7(32'hbbbd351b),
	.w8(32'hbc95a657),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd26b4a),
	.w1(32'hbaf53e20),
	.w2(32'h3a82126e),
	.w3(32'hbbd9fb30),
	.w4(32'hbc188d91),
	.w5(32'hbcb1984a),
	.w6(32'hbb78f72f),
	.w7(32'h39dd314b),
	.w8(32'hbba83586),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc407509),
	.w1(32'hbcc02cef),
	.w2(32'hbb4e4ac2),
	.w3(32'hbbffe9c0),
	.w4(32'hbb4ebe87),
	.w5(32'h3a092dc5),
	.w6(32'hbcf53350),
	.w7(32'hbc819c25),
	.w8(32'hbc8d9b53),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36a3c0),
	.w1(32'hbc71d8b0),
	.w2(32'h3b6f9952),
	.w3(32'h38c858b3),
	.w4(32'hbc4bb015),
	.w5(32'h3b2b9af4),
	.w6(32'h3c0f1ec7),
	.w7(32'hbb34d93f),
	.w8(32'h3913de0d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4410),
	.w1(32'hbc0a985a),
	.w2(32'h3be0d02b),
	.w3(32'hbca58af8),
	.w4(32'hbc85ed7f),
	.w5(32'h3b5b86f7),
	.w6(32'hbba1dc2c),
	.w7(32'hbbd8305e),
	.w8(32'hbc4ec512),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c007961),
	.w1(32'h3adeb575),
	.w2(32'h3a2d453a),
	.w3(32'h3d170816),
	.w4(32'h3d200e39),
	.w5(32'hbaec5be8),
	.w6(32'h3bc09c1a),
	.w7(32'h3a88a542),
	.w8(32'h399d7d77),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6599c9),
	.w1(32'hbc57abf8),
	.w2(32'h3b7979fd),
	.w3(32'h3bf7f783),
	.w4(32'h3b91d4cf),
	.w5(32'hbb48e056),
	.w6(32'hba9f254d),
	.w7(32'h3b1c133b),
	.w8(32'h3a889f78),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd6cc4),
	.w1(32'h3a863739),
	.w2(32'hbb902851),
	.w3(32'hbc9c115b),
	.w4(32'hbbb4de1d),
	.w5(32'h3aa39a97),
	.w6(32'hbb6e2305),
	.w7(32'hb9b6b63f),
	.w8(32'hbb1a027e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3da35b),
	.w1(32'hba5f4292),
	.w2(32'hbc03fbf8),
	.w3(32'h3c079d95),
	.w4(32'h3be3c69e),
	.w5(32'h3b127094),
	.w6(32'h3c2d2b88),
	.w7(32'h3c144cd6),
	.w8(32'h3c916076),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc3181d),
	.w1(32'hbc95929e),
	.w2(32'hbcc6865f),
	.w3(32'hbd05b28a),
	.w4(32'hbcf0ed35),
	.w5(32'hbc1f00d0),
	.w6(32'h3a27967c),
	.w7(32'hbb415c69),
	.w8(32'hbb9133f6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30e98b),
	.w1(32'h3b0b742e),
	.w2(32'hbc07f663),
	.w3(32'h37c39b74),
	.w4(32'hbaad6168),
	.w5(32'h3a40113d),
	.w6(32'h3c54b13b),
	.w7(32'h3b82e55f),
	.w8(32'h3b782ee4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ff0eb),
	.w1(32'h3b25eead),
	.w2(32'h3bf397df),
	.w3(32'h3a4230ef),
	.w4(32'h3b07fc81),
	.w5(32'hbc2eb196),
	.w6(32'h3b89078b),
	.w7(32'h3ac36587),
	.w8(32'h3a2b0a90),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5aa85f),
	.w1(32'h3c40d390),
	.w2(32'h3bfbc46c),
	.w3(32'hbb4275c9),
	.w4(32'h3c051481),
	.w5(32'hba49483f),
	.w6(32'hbba3d52b),
	.w7(32'hbc10f9d1),
	.w8(32'h3c3a3dfd),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af778cd),
	.w1(32'h3bcf1837),
	.w2(32'h3cbc020b),
	.w3(32'h3b8f8bc9),
	.w4(32'h3c407a8f),
	.w5(32'h3ccd20ea),
	.w6(32'h3af39736),
	.w7(32'h3bba5d3f),
	.w8(32'hba468c56),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb5f9ce),
	.w1(32'h394d225b),
	.w2(32'h3b9cc85a),
	.w3(32'h3d62b651),
	.w4(32'h3d1c54b3),
	.w5(32'hbc819216),
	.w6(32'h3c5370ba),
	.w7(32'h3caa0ae8),
	.w8(32'hbc5c07ca),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805096),
	.w1(32'hbc79d3ad),
	.w2(32'hbb5b1d1a),
	.w3(32'h3b9b0146),
	.w4(32'h3b8c7303),
	.w5(32'h3c311a2d),
	.w6(32'hbca9cc2a),
	.w7(32'hbc49aece),
	.w8(32'h3bf58760),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c9808),
	.w1(32'h3c95bc2c),
	.w2(32'h3c3e5c65),
	.w3(32'hbc25002c),
	.w4(32'hbc88e931),
	.w5(32'hba2d4fac),
	.w6(32'h3c965924),
	.w7(32'h3c272ebc),
	.w8(32'h3beab2fb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d8bd1),
	.w1(32'h3c2fb265),
	.w2(32'h3b7036ce),
	.w3(32'hbb957692),
	.w4(32'hbadfe8b0),
	.w5(32'h3c125b64),
	.w6(32'h3c88706e),
	.w7(32'h3c42fde5),
	.w8(32'hbc5e67fb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac67c49),
	.w1(32'hbca11a1e),
	.w2(32'h3bc7d49e),
	.w3(32'h3d1d6282),
	.w4(32'h3d1cb6e9),
	.w5(32'hbc15d527),
	.w6(32'hbbe2ead6),
	.w7(32'h3b847b14),
	.w8(32'hbc2eea15),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8788b),
	.w1(32'h3a4e0ea9),
	.w2(32'hbaf2ce8f),
	.w3(32'hbc288db2),
	.w4(32'h3b1a05f6),
	.w5(32'hbbb3e84d),
	.w6(32'hbc8e87c5),
	.w7(32'hbc5a1d9d),
	.w8(32'h39fb9de7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b265dd8),
	.w1(32'h3ba9f053),
	.w2(32'hbc2f9f9f),
	.w3(32'hbc0fa192),
	.w4(32'hbc2577ac),
	.w5(32'h3b913e82),
	.w6(32'hbb8a5afa),
	.w7(32'hbb407f74),
	.w8(32'hbb8bb8ed),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6792e8),
	.w1(32'hbb420298),
	.w2(32'hbb3d8b28),
	.w3(32'h3b329963),
	.w4(32'hbb8bc6df),
	.w5(32'hbc2904a1),
	.w6(32'hbbd6e034),
	.w7(32'h3ac7aceb),
	.w8(32'h3bbaea2c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92906f4),
	.w1(32'hbb2dc9da),
	.w2(32'hbbdfc670),
	.w3(32'hbbd8631e),
	.w4(32'hbb16a87f),
	.w5(32'hbb19c6a9),
	.w6(32'h3b57a5f6),
	.w7(32'h3a2ca4da),
	.w8(32'hb9f921ec),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f539d),
	.w1(32'hbc341111),
	.w2(32'hbc0c0a59),
	.w3(32'hbb46e5bf),
	.w4(32'hb91c28ab),
	.w5(32'h3b02487f),
	.w6(32'h37a4c296),
	.w7(32'hbbad1883),
	.w8(32'h398bf86b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a0c93),
	.w1(32'hbcb6feb9),
	.w2(32'h3c1c33f5),
	.w3(32'h3c9ae13e),
	.w4(32'h3c0389eb),
	.w5(32'hbaead54b),
	.w6(32'hbc0b633f),
	.w7(32'h3a53d327),
	.w8(32'h3baddff7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd66b71),
	.w1(32'hbb957c08),
	.w2(32'hbb1734c1),
	.w3(32'h3b939f12),
	.w4(32'h3b181507),
	.w5(32'hba16dd15),
	.w6(32'hbc7e7b7a),
	.w7(32'hbc570eb3),
	.w8(32'h3ab19140),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba2a7c),
	.w1(32'hbbb1691d),
	.w2(32'hbb4ce083),
	.w3(32'hbb8f3258),
	.w4(32'hbb97feba),
	.w5(32'h3b2e4409),
	.w6(32'hbb4f994e),
	.w7(32'hbb1dfcef),
	.w8(32'hbb40de2c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c196e),
	.w1(32'h3ba21b7f),
	.w2(32'hbc0b99a7),
	.w3(32'h3c006047),
	.w4(32'h3b46b047),
	.w5(32'h3c90ed77),
	.w6(32'h3bed582e),
	.w7(32'h3b95164f),
	.w8(32'hbb8e424d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc60bfe),
	.w1(32'hbbee31d6),
	.w2(32'h3a8ef69f),
	.w3(32'hbb230746),
	.w4(32'hbc801710),
	.w5(32'hbb4fa9a9),
	.w6(32'h3bea5f1f),
	.w7(32'h3c4e10a7),
	.w8(32'hba98f3cc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb87d63),
	.w1(32'h3b9f4733),
	.w2(32'hbc71efa1),
	.w3(32'hbac3a2e1),
	.w4(32'h3abcd2e3),
	.w5(32'h3b99c4cc),
	.w6(32'hbb1113ed),
	.w7(32'hbb43fb2b),
	.w8(32'h3b217838),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec72ef),
	.w1(32'h3a0f9262),
	.w2(32'hbc6f15c9),
	.w3(32'hbc703c20),
	.w4(32'hbc9191fb),
	.w5(32'h3b0e74e7),
	.w6(32'h3bfbfe80),
	.w7(32'h3bfcb67c),
	.w8(32'h3b2c84a7),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba247be9),
	.w1(32'h3b12be19),
	.w2(32'hbb3a285b),
	.w3(32'h3b10d2e2),
	.w4(32'hbc233108),
	.w5(32'h3b50fea5),
	.w6(32'h3cce33cb),
	.w7(32'h3c6f18ff),
	.w8(32'hb8d248e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2acb7f),
	.w1(32'h3ac24fef),
	.w2(32'hbc1bab77),
	.w3(32'hbbede66b),
	.w4(32'hbc6900e0),
	.w5(32'h3cf59fa7),
	.w6(32'h3c14186f),
	.w7(32'h3be4701d),
	.w8(32'hbbfe5806),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaaace7),
	.w1(32'hbbf957d7),
	.w2(32'h3c7bf5ba),
	.w3(32'h3c7449aa),
	.w4(32'hba93643f),
	.w5(32'hbcb706d3),
	.w6(32'h3b9441bd),
	.w7(32'h3c7c7192),
	.w8(32'h3cb676d1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6dbd30),
	.w1(32'h3ba93c9d),
	.w2(32'h3c121ace),
	.w3(32'hbc734a38),
	.w4(32'h3c20fa03),
	.w5(32'hbbbd515c),
	.w6(32'h3c099949),
	.w7(32'hbc0b8936),
	.w8(32'hbc28a236),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac4626),
	.w1(32'hbc07a5fd),
	.w2(32'h3ca154c1),
	.w3(32'hb9c3bd9c),
	.w4(32'h3b739d76),
	.w5(32'h3bceaf41),
	.w6(32'hbc863e6c),
	.w7(32'hbc9c8005),
	.w8(32'hbbd65b7a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8288ba),
	.w1(32'hbbaf7512),
	.w2(32'hbc9a947d),
	.w3(32'h3d28c82a),
	.w4(32'h3d033681),
	.w5(32'hbca18c78),
	.w6(32'hbbbb800c),
	.w7(32'hbabb0ea5),
	.w8(32'hbc1246f9),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcda1a10),
	.w1(32'hbc7dda68),
	.w2(32'h3af984b6),
	.w3(32'hbcdf4e31),
	.w4(32'hbcb99041),
	.w5(32'hbba8509b),
	.w6(32'hbc0afa18),
	.w7(32'hbc9951e5),
	.w8(32'h3c340357),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaf6b6),
	.w1(32'h3c1859ba),
	.w2(32'h3b7d4ba7),
	.w3(32'hbc9e88c4),
	.w4(32'h3c030a5b),
	.w5(32'h3baeae87),
	.w6(32'h3be9198c),
	.w7(32'h3c1e174d),
	.w8(32'h3b7074f7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3976a6),
	.w1(32'hbc34783c),
	.w2(32'h3b5301ec),
	.w3(32'hbc553288),
	.w4(32'hbbff6f23),
	.w5(32'hbc666a3e),
	.w6(32'hbc4bfe7b),
	.w7(32'hbbf18dc7),
	.w8(32'hbc7549d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7598d6),
	.w1(32'h3b04be83),
	.w2(32'h3affc7d2),
	.w3(32'hba4fa161),
	.w4(32'hbaa01bc9),
	.w5(32'h3c262c97),
	.w6(32'hbb648f14),
	.w7(32'hbb864b76),
	.w8(32'hbc1f458c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a2bde),
	.w1(32'h39d33844),
	.w2(32'h3c0505af),
	.w3(32'h3bf4eba5),
	.w4(32'h3a8d0982),
	.w5(32'hbad928cd),
	.w6(32'hbbda1783),
	.w7(32'hba713df7),
	.w8(32'h3af8d173),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4529f4),
	.w1(32'h3b143176),
	.w2(32'hbb428021),
	.w3(32'hbba2f6b4),
	.w4(32'h3b104c57),
	.w5(32'hb79850dd),
	.w6(32'hbbeabf2b),
	.w7(32'hbab32e26),
	.w8(32'hb9c7d4c9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20290d),
	.w1(32'h3b2b7606),
	.w2(32'hbbfaf424),
	.w3(32'h3bbabe6e),
	.w4(32'h3ba59f81),
	.w5(32'h3cbf9e85),
	.w6(32'h3aa96df4),
	.w7(32'h3b948f12),
	.w8(32'hbc88ccd9),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cf1cb),
	.w1(32'hbcab6fc4),
	.w2(32'hb9975592),
	.w3(32'h3d15d182),
	.w4(32'h3c7dba40),
	.w5(32'h392f3e1c),
	.w6(32'hbc20e051),
	.w7(32'h3ac1e21a),
	.w8(32'h3a9a56d8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9076a6f),
	.w1(32'h39775336),
	.w2(32'hbb93dada),
	.w3(32'h3aa78a65),
	.w4(32'h3a7aa654),
	.w5(32'h3ba6e556),
	.w6(32'hbb4c4bb1),
	.w7(32'hbadd2c00),
	.w8(32'h3ab7c88b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87e4ac),
	.w1(32'h3b9f10ff),
	.w2(32'h3cb3285b),
	.w3(32'h3cedc829),
	.w4(32'h3bdb479d),
	.w5(32'hbc96b41a),
	.w6(32'h3cb6f647),
	.w7(32'h3c295e2a),
	.w8(32'h3adc02a3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ade4d),
	.w1(32'hbc0b52d7),
	.w2(32'hbbf793fa),
	.w3(32'h3c45044e),
	.w4(32'h3cca7412),
	.w5(32'hbc0c36da),
	.w6(32'hbc37498a),
	.w7(32'hbc8096ae),
	.w8(32'h3a364143),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a6f7a),
	.w1(32'h3b245961),
	.w2(32'h3aa9b268),
	.w3(32'hbbb4ed6d),
	.w4(32'h3b8fbb38),
	.w5(32'h3adeb0ad),
	.w6(32'hbb15314f),
	.w7(32'hbb7cc53d),
	.w8(32'h3b7bb68f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa19d93),
	.w1(32'h3b053c49),
	.w2(32'hba7c0722),
	.w3(32'h3af2ee8f),
	.w4(32'h3b02b6ef),
	.w5(32'h3b1668c9),
	.w6(32'h3a2c8271),
	.w7(32'hb9da8673),
	.w8(32'hbbf18407),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd175fb),
	.w1(32'h3b20a3f7),
	.w2(32'h3b28dba2),
	.w3(32'h3c5fb9d6),
	.w4(32'h3bd5f79b),
	.w5(32'h3b5d0510),
	.w6(32'h3c06ae32),
	.w7(32'h3c805d1b),
	.w8(32'h39d67249),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb88b1),
	.w1(32'h3b2d4f11),
	.w2(32'h3cb93495),
	.w3(32'h3c7eb266),
	.w4(32'h3b86d6e7),
	.w5(32'h3a13d123),
	.w6(32'h3c05a39c),
	.w7(32'h3bc7786f),
	.w8(32'h3c045639),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e0ca),
	.w1(32'h3b445f89),
	.w2(32'h399eda6b),
	.w3(32'h3d1102b1),
	.w4(32'h3d230de4),
	.w5(32'h3c328082),
	.w6(32'hbc20c3b6),
	.w7(32'hbc32df88),
	.w8(32'h3bd24594),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb661bd),
	.w1(32'hbb3d7b4c),
	.w2(32'h3b7aee2b),
	.w3(32'h3b8193a9),
	.w4(32'h38197a6e),
	.w5(32'hbc3c7530),
	.w6(32'h3c24bdec),
	.w7(32'h3bea927f),
	.w8(32'hbb5d6dc1),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205852),
	.w1(32'hbc1b2f0a),
	.w2(32'h3b95ea65),
	.w3(32'hbb706a76),
	.w4(32'h3b82aa4c),
	.w5(32'hba2b599e),
	.w6(32'hbc90dc9c),
	.w7(32'hbcaf4cab),
	.w8(32'hba2b90a5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c014483),
	.w1(32'h39775116),
	.w2(32'h3b050b10),
	.w3(32'h3b7a7150),
	.w4(32'h3a0c971d),
	.w5(32'hbafa97b2),
	.w6(32'hbbd44917),
	.w7(32'hbbc5160b),
	.w8(32'h3b524345),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17dfa4),
	.w1(32'hbc42b5a1),
	.w2(32'hbb99a697),
	.w3(32'hbc010725),
	.w4(32'hbbe280ff),
	.w5(32'hba595dca),
	.w6(32'hbbfccaa7),
	.w7(32'hbbfad8de),
	.w8(32'hbb90f402),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1accb1),
	.w1(32'h3c09f366),
	.w2(32'h3c51d528),
	.w3(32'h3c8c9fac),
	.w4(32'h3bf68ec4),
	.w5(32'hbc62d8d0),
	.w6(32'h3c86cc09),
	.w7(32'h3a915cfb),
	.w8(32'hbc4079f7),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf355d),
	.w1(32'h3c8793fb),
	.w2(32'hbadbf0fb),
	.w3(32'hbc75a190),
	.w4(32'h3a88f2bf),
	.w5(32'h3b96cec4),
	.w6(32'hbbbfc135),
	.w7(32'hbc9b7ecb),
	.w8(32'h3b754eda),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0830b8),
	.w1(32'h3bbc227d),
	.w2(32'h3b2976f7),
	.w3(32'hbb73b685),
	.w4(32'hbba442df),
	.w5(32'h3b2fe2d0),
	.w6(32'h3c5a9bdd),
	.w7(32'h3bed2469),
	.w8(32'h3acda2ed),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb483b13),
	.w1(32'hbb3c71dd),
	.w2(32'hbc084f17),
	.w3(32'hb8bc4d3d),
	.w4(32'h398560f3),
	.w5(32'hbb5987dc),
	.w6(32'hb99ad81c),
	.w7(32'hb84168d9),
	.w8(32'hbbd52537),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb111fda),
	.w1(32'h38643c9a),
	.w2(32'h3a6bf510),
	.w3(32'h3b226f9b),
	.w4(32'hbab78fc6),
	.w5(32'h3a909df7),
	.w6(32'hba28645e),
	.w7(32'hbb403e17),
	.w8(32'hbb7865b2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75692b),
	.w1(32'hbc118a50),
	.w2(32'h3b8a745c),
	.w3(32'hbbb819f1),
	.w4(32'h3ab48718),
	.w5(32'h3b07afba),
	.w6(32'hbb897453),
	.w7(32'h3a31a354),
	.w8(32'hb94f4421),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47ad1c),
	.w1(32'hbb978059),
	.w2(32'h3ad7ed90),
	.w3(32'hbb896cb7),
	.w4(32'hbaa151e2),
	.w5(32'hbc5f30ae),
	.w6(32'hbb82c69b),
	.w7(32'hba830424),
	.w8(32'hbc976c48),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30e363),
	.w1(32'hbc82b659),
	.w2(32'h3bcc1094),
	.w3(32'hbd268f41),
	.w4(32'hbcabce47),
	.w5(32'hbb5bba63),
	.w6(32'hbc98e014),
	.w7(32'hbb8eca49),
	.w8(32'hbc629164),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08995a),
	.w1(32'hbbe1b726),
	.w2(32'hbbb87278),
	.w3(32'hbcb7b52f),
	.w4(32'hbc846f8f),
	.w5(32'hbb93b54f),
	.w6(32'hbcb68e29),
	.w7(32'h3b041766),
	.w8(32'hbc00e197),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eaf1d),
	.w1(32'hbb49cedf),
	.w2(32'hb9c4eeec),
	.w3(32'hbb278765),
	.w4(32'hba6258c1),
	.w5(32'h3c00a7a9),
	.w6(32'hbb09570c),
	.w7(32'h3a2006fe),
	.w8(32'hbbeb48ab),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c567abd),
	.w1(32'h3bd017aa),
	.w2(32'h39bce668),
	.w3(32'h3c69e78a),
	.w4(32'h3aed4381),
	.w5(32'h3b82ca5c),
	.w6(32'hbbdd4d91),
	.w7(32'hba884b4e),
	.w8(32'h3b39cbd5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abab759),
	.w1(32'h3ab8c7f0),
	.w2(32'hbc5135d7),
	.w3(32'h3ab0491b),
	.w4(32'hba37e033),
	.w5(32'hbbf893bf),
	.w6(32'h39871a35),
	.w7(32'h3acc9ccc),
	.w8(32'hbbc9854f),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58203a),
	.w1(32'h3b9a3b55),
	.w2(32'h3b815461),
	.w3(32'h3ba33a98),
	.w4(32'h3bb83d08),
	.w5(32'h3bd71a90),
	.w6(32'h3ba252d2),
	.w7(32'h3c02d75e),
	.w8(32'h3b402619),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb94202),
	.w1(32'h3b3f2160),
	.w2(32'h398a7af8),
	.w3(32'h3bdc5def),
	.w4(32'h3bb50ed1),
	.w5(32'hbc3516aa),
	.w6(32'h3b6257d8),
	.w7(32'h3b4d41fe),
	.w8(32'hbc3d547b),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f06be),
	.w1(32'hbb5afe25),
	.w2(32'hbbfe0fe0),
	.w3(32'hbc0c46d8),
	.w4(32'h3a9e66b4),
	.w5(32'hba81d0ad),
	.w6(32'hb9f9eb28),
	.w7(32'h3be5e4b3),
	.w8(32'h3ab19987),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce55dd),
	.w1(32'h3af45af0),
	.w2(32'hbb875653),
	.w3(32'hba2adba7),
	.w4(32'h3ab7fc01),
	.w5(32'h3a89d030),
	.w6(32'hb8922645),
	.w7(32'hbb5bb31e),
	.w8(32'h3b7d64ba),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4cbf4),
	.w1(32'hbb9e17b0),
	.w2(32'h3a8b5dbc),
	.w3(32'hbbb93dd2),
	.w4(32'hbbb1b8ca),
	.w5(32'hb9852560),
	.w6(32'hbc5ce433),
	.w7(32'hbc166b2a),
	.w8(32'hbc630fe6),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad82b73),
	.w1(32'hbac9e7cf),
	.w2(32'hbbe0b0e1),
	.w3(32'h3a7e3198),
	.w4(32'hb9ed9754),
	.w5(32'hbc8deb2a),
	.w6(32'h3b278fb3),
	.w7(32'h3c269f45),
	.w8(32'hbcb2673e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad36d4),
	.w1(32'hbcc85bfd),
	.w2(32'hbb467e7f),
	.w3(32'hbd04b8f1),
	.w4(32'hbca5dbd3),
	.w5(32'hba08313b),
	.w6(32'hbccca1bf),
	.w7(32'hbbc5943c),
	.w8(32'h3a3c6fe0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba132e62),
	.w1(32'hb9d8c96c),
	.w2(32'h3bd52852),
	.w3(32'hbace9ddf),
	.w4(32'hbab04949),
	.w5(32'h3c30bd35),
	.w6(32'hba0b82e3),
	.w7(32'hba860bf4),
	.w8(32'hb980c2db),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd852f),
	.w1(32'hbc314243),
	.w2(32'h3b8a2d43),
	.w3(32'hbb18f862),
	.w4(32'hbc2129d6),
	.w5(32'hbbe867b8),
	.w6(32'hbbfea647),
	.w7(32'hbba337d6),
	.w8(32'h3a65d6c1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2af49d),
	.w1(32'hba337164),
	.w2(32'h3be2283e),
	.w3(32'hbc13934d),
	.w4(32'hbab49935),
	.w5(32'h3b1880f9),
	.w6(32'hbba92e57),
	.w7(32'hbb83bc05),
	.w8(32'hbb81ce15),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0d245),
	.w1(32'hbcdded05),
	.w2(32'h3c1e9bb3),
	.w3(32'hbcd5db04),
	.w4(32'hbcb7a206),
	.w5(32'h3c24f88c),
	.w6(32'hbce86bab),
	.w7(32'hbc2a0570),
	.w8(32'h3b9e74fc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cb4c8),
	.w1(32'h3a44b440),
	.w2(32'h3b5aa518),
	.w3(32'hba76ec0d),
	.w4(32'hbba8a6dd),
	.w5(32'h3b31f55b),
	.w6(32'hbbc81d4c),
	.w7(32'hbb88157c),
	.w8(32'h3b888d84),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8039dce),
	.w1(32'hb9cb0459),
	.w2(32'h39c27048),
	.w3(32'h3ad8fbe8),
	.w4(32'hbad7099b),
	.w5(32'h38f9cfe2),
	.w6(32'hb8ba6778),
	.w7(32'hb98ebb29),
	.w8(32'hbc3018e3),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d1432),
	.w1(32'hbc1937df),
	.w2(32'hbb622d1b),
	.w3(32'h3b3c6a04),
	.w4(32'h393188c4),
	.w5(32'hb9b7473e),
	.w6(32'hbaa860ac),
	.w7(32'hbb229e27),
	.w8(32'hbb0aad13),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1057d5),
	.w1(32'h3be64a3c),
	.w2(32'h3b58406f),
	.w3(32'h3c236df8),
	.w4(32'h3c278e4a),
	.w5(32'h3b2052ed),
	.w6(32'hbbbe4ff6),
	.w7(32'h3b100910),
	.w8(32'hbaafbfc0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ebe04),
	.w1(32'h3c032afb),
	.w2(32'hbb989d3b),
	.w3(32'hba2ba364),
	.w4(32'h3c689347),
	.w5(32'h3bccf0d4),
	.w6(32'h3c4f09ce),
	.w7(32'h3bf17abe),
	.w8(32'hb9b40ce9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f63c8),
	.w1(32'h3c25855a),
	.w2(32'h3b98bb4a),
	.w3(32'h3c84ed26),
	.w4(32'h3c48e42d),
	.w5(32'h3ad3f68a),
	.w6(32'h3b2b1f6f),
	.w7(32'hbae521e7),
	.w8(32'hb9f0369b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea6188),
	.w1(32'h3b8f9119),
	.w2(32'h3b0ba47d),
	.w3(32'hba6236bb),
	.w4(32'h3babea20),
	.w5(32'hbb038b3d),
	.w6(32'h3be55678),
	.w7(32'h3c6539cf),
	.w8(32'hbbbd94ae),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32f779),
	.w1(32'h3bf852da),
	.w2(32'h3b818d2d),
	.w3(32'hbb346c71),
	.w4(32'h3c34e053),
	.w5(32'h3b8978e8),
	.w6(32'h3b538834),
	.w7(32'h3c5d632b),
	.w8(32'hbb7ee0a1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5da03),
	.w1(32'h3b98d786),
	.w2(32'hbb6819c7),
	.w3(32'hbbd2debd),
	.w4(32'hbc9d841e),
	.w5(32'hbc2ca317),
	.w6(32'hbc65dbb9),
	.w7(32'h3a94a764),
	.w8(32'hbc37e0ad),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0bfb3),
	.w1(32'hbc3ce170),
	.w2(32'h3985673a),
	.w3(32'hbc9ff6e5),
	.w4(32'hbbb9d8dd),
	.w5(32'h3b0e18ea),
	.w6(32'hbc526c42),
	.w7(32'hbbda252a),
	.w8(32'hbacf56d5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b671e82),
	.w1(32'h396f8583),
	.w2(32'h3a5935de),
	.w3(32'h3a9cf9e1),
	.w4(32'h399f3df6),
	.w5(32'h3b855a8c),
	.w6(32'hbb31b9a3),
	.w7(32'hbb0aec5b),
	.w8(32'h3b9f6ba2),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff3106),
	.w1(32'hbb26dab1),
	.w2(32'hbb7e5fd4),
	.w3(32'h3b43f130),
	.w4(32'hb9d0c2f7),
	.w5(32'hbb8017e7),
	.w6(32'h3ba70084),
	.w7(32'hba40a388),
	.w8(32'hbbafede8),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63fb4e),
	.w1(32'hbc2052c3),
	.w2(32'h3b0e9817),
	.w3(32'hbba0b0a6),
	.w4(32'hbbd272aa),
	.w5(32'hbad4e6c2),
	.w6(32'hbbc0fde8),
	.w7(32'hbb6d5a4d),
	.w8(32'h3ab86a88),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c142d90),
	.w1(32'h3c2206ac),
	.w2(32'h3c1f863b),
	.w3(32'h3c8e4a63),
	.w4(32'h3c0ed424),
	.w5(32'hbb01e37b),
	.w6(32'h3c3ffdc1),
	.w7(32'h3b98893f),
	.w8(32'hbbb59953),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc458dfe),
	.w1(32'hbc7ccea4),
	.w2(32'h3c1499ef),
	.w3(32'hbcc9a916),
	.w4(32'hbca36f68),
	.w5(32'h3c1dd00f),
	.w6(32'hbca240c4),
	.w7(32'hbc3249c2),
	.w8(32'h3b40cb5b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f552b),
	.w1(32'h3c17b0f5),
	.w2(32'h3b010e3a),
	.w3(32'h3c578c14),
	.w4(32'h3c5a6d88),
	.w5(32'h3c0eb62e),
	.w6(32'h3c1189de),
	.w7(32'h3c0069b3),
	.w8(32'h3bc0529c),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2dcc),
	.w1(32'h3bbe09f4),
	.w2(32'h3c02b61c),
	.w3(32'h3bf803e8),
	.w4(32'h3bd8af32),
	.w5(32'h3c22f8e4),
	.w6(32'h3c0c0037),
	.w7(32'h3bc6bcdc),
	.w8(32'h3be2b571),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9248be),
	.w1(32'hba3a14cd),
	.w2(32'h3bed7b93),
	.w3(32'h3ac8b6d0),
	.w4(32'hbb3a91b1),
	.w5(32'h3bba0e7d),
	.w6(32'h3b30cb37),
	.w7(32'h3aa2b9e6),
	.w8(32'h3b9444e6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbf79f),
	.w1(32'h3c1bb684),
	.w2(32'h3b2edad3),
	.w3(32'h3bbbee47),
	.w4(32'h3bd59c6b),
	.w5(32'h3b776f52),
	.w6(32'h3b39aafe),
	.w7(32'h3c03d341),
	.w8(32'h3a2d1e81),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3333a7),
	.w1(32'h3aa0fd7d),
	.w2(32'h3b9c597f),
	.w3(32'h3b8d681a),
	.w4(32'h3bbaa288),
	.w5(32'h3c43006a),
	.w6(32'h3b255a26),
	.w7(32'hb9fd1a20),
	.w8(32'h3a3c1d66),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963a9c3),
	.w1(32'hbb1d0854),
	.w2(32'h3c006ac5),
	.w3(32'h3b8bc204),
	.w4(32'hbb183427),
	.w5(32'h3bfb881a),
	.w6(32'h3b7baa58),
	.w7(32'h3b2d6ffa),
	.w8(32'h3c680c4a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8edfae),
	.w1(32'h3c1ce78a),
	.w2(32'h3b645f19),
	.w3(32'h3ba126e5),
	.w4(32'h3b84f44d),
	.w5(32'h3b87e7d8),
	.w6(32'hbb13db37),
	.w7(32'hbbdf3780),
	.w8(32'h3b96ea50),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9db9f9),
	.w1(32'h3b8ffc78),
	.w2(32'h3b70ef46),
	.w3(32'h3b9c0103),
	.w4(32'h3b686b34),
	.w5(32'h3b187c2d),
	.w6(32'h3b3dd732),
	.w7(32'h3ac5ac63),
	.w8(32'h3aa1f6d5),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d199b),
	.w1(32'h3ba143b2),
	.w2(32'h3bb94bfb),
	.w3(32'h3a32602a),
	.w4(32'h3b69f5ea),
	.w5(32'hb8dfec25),
	.w6(32'h3a989cf2),
	.w7(32'h3b702799),
	.w8(32'h3a091ed0),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefe036),
	.w1(32'hbb04d426),
	.w2(32'h3c008fcf),
	.w3(32'hbb98a7a5),
	.w4(32'hbb44f804),
	.w5(32'h3b69f03c),
	.w6(32'hbacede28),
	.w7(32'h3b04a44c),
	.w8(32'h3bce6730),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0df9c5),
	.w1(32'hbc4f70dd),
	.w2(32'h3b74b9b1),
	.w3(32'hbca87ed7),
	.w4(32'hbc42ad1e),
	.w5(32'hbbaf75bb),
	.w6(32'hbc140985),
	.w7(32'hbae7e2e7),
	.w8(32'hbcad3d75),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a411319),
	.w1(32'hb99b6f09),
	.w2(32'h3b775966),
	.w3(32'hba443c07),
	.w4(32'h39434434),
	.w5(32'h388d7b08),
	.w6(32'hbc579a5e),
	.w7(32'hbad1e828),
	.w8(32'h3af381b9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1be927),
	.w1(32'hba0cdacd),
	.w2(32'hbc328f55),
	.w3(32'hbb012688),
	.w4(32'hba92ad5a),
	.w5(32'hbc2080b1),
	.w6(32'hbb01251c),
	.w7(32'hba88576b),
	.w8(32'hbc249a96),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27917b),
	.w1(32'hbb0cdaf1),
	.w2(32'h3c55f07f),
	.w3(32'hbb82045f),
	.w4(32'hbb2c2198),
	.w5(32'h3b448e36),
	.w6(32'hbbc9e31d),
	.w7(32'hbae4ad66),
	.w8(32'h3b92611b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab57cee),
	.w1(32'h3bee9f76),
	.w2(32'hbab1469e),
	.w3(32'h3c06a5f8),
	.w4(32'h3c4b9e45),
	.w5(32'hbbb08364),
	.w6(32'h3c047d17),
	.w7(32'h3bff6969),
	.w8(32'hbc21aea3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf21497),
	.w1(32'hbb992679),
	.w2(32'h3b1fc92e),
	.w3(32'hbc9ccf56),
	.w4(32'hbb8a263c),
	.w5(32'h3a20a189),
	.w6(32'h3b34d2e5),
	.w7(32'h3c3236d9),
	.w8(32'hbb93f90b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10dfbb),
	.w1(32'hbb719a9d),
	.w2(32'h3a84cb6c),
	.w3(32'hbbea4353),
	.w4(32'hbbb1d79b),
	.w5(32'h3b328f51),
	.w6(32'hbbd1a7d7),
	.w7(32'hba94c116),
	.w8(32'h3b38bce8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98432e),
	.w1(32'hbb2897b3),
	.w2(32'h3bba11be),
	.w3(32'hbb98ed88),
	.w4(32'hba13d392),
	.w5(32'h3c2d33a5),
	.w6(32'hbb395480),
	.w7(32'h3a0d2a2f),
	.w8(32'h3be421f5),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64528d),
	.w1(32'h3c0121d7),
	.w2(32'h3b20b8e1),
	.w3(32'h3c04dff4),
	.w4(32'h3b454b5e),
	.w5(32'h39011823),
	.w6(32'h3c16b8f6),
	.w7(32'h3b863cf3),
	.w8(32'hbb0c190b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945d801),
	.w1(32'hba8a2d10),
	.w2(32'h3c244daa),
	.w3(32'hba1e8603),
	.w4(32'h3b219bc3),
	.w5(32'h3beb9e80),
	.w6(32'h3aadd8a1),
	.w7(32'h3b814721),
	.w8(32'h3bee17c6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffab3d),
	.w1(32'hbb2735db),
	.w2(32'h3b3f1e9a),
	.w3(32'h3beea80e),
	.w4(32'h3a55d4a0),
	.w5(32'hba846217),
	.w6(32'h3c0e8bb5),
	.w7(32'h3bef4ea7),
	.w8(32'hb8b8b465),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd92e33),
	.w1(32'hbc94efb1),
	.w2(32'h3bae7360),
	.w3(32'hbcc166c2),
	.w4(32'hbc9cfe40),
	.w5(32'h3b82ca18),
	.w6(32'hbce6385d),
	.w7(32'hbc82c543),
	.w8(32'h3b1e0109),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3e09d),
	.w1(32'hbbeca55b),
	.w2(32'h3b66143d),
	.w3(32'hbbe2487d),
	.w4(32'hbb3fed57),
	.w5(32'h3c041784),
	.w6(32'hbc700467),
	.w7(32'hbbdb08af),
	.w8(32'hbc444160),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cbea7),
	.w1(32'h3bbbf7cb),
	.w2(32'h3b94533d),
	.w3(32'h3c5ad611),
	.w4(32'h3c0f22a4),
	.w5(32'h3b91b366),
	.w6(32'h3c5580be),
	.w7(32'h3bdfbb53),
	.w8(32'h3b8209f1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fde2d0),
	.w1(32'h389e2da0),
	.w2(32'hbb253b0d),
	.w3(32'hba86eaf5),
	.w4(32'hba0f8f3e),
	.w5(32'hbad5c1cf),
	.w6(32'hb9c45f6e),
	.w7(32'h3b82d623),
	.w8(32'hbb99d7c8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb317981),
	.w1(32'hba6785b2),
	.w2(32'h3b51781d),
	.w3(32'hbb28354b),
	.w4(32'hbac0e6f5),
	.w5(32'h3bc3ba0c),
	.w6(32'hbb4a5604),
	.w7(32'hbb11dd5d),
	.w8(32'h398cc41b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b598c9c),
	.w1(32'h3c24d93d),
	.w2(32'hbae38993),
	.w3(32'h3c12be38),
	.w4(32'h3c235acd),
	.w5(32'hba26ca76),
	.w6(32'h3b377cdc),
	.w7(32'h3c0b2a6e),
	.w8(32'hbc437689),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4458b2),
	.w1(32'h3b475d6d),
	.w2(32'hba3703f1),
	.w3(32'hbc5f27e1),
	.w4(32'hb94db8d0),
	.w5(32'hba5cbfe8),
	.w6(32'hbc700265),
	.w7(32'h3b41b4bb),
	.w8(32'hbb63cf7b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ebfba),
	.w1(32'hbbffb375),
	.w2(32'hbc437a14),
	.w3(32'hbbc45d1f),
	.w4(32'hbb517123),
	.w5(32'hb9391d29),
	.w6(32'hbbd1bab6),
	.w7(32'hbc19f91d),
	.w8(32'hbbd6c3d1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f9bee),
	.w1(32'hbb8ae5f3),
	.w2(32'hbba61d58),
	.w3(32'h3bb88c35),
	.w4(32'hbb21351d),
	.w5(32'hbba9b89b),
	.w6(32'hbb9be35e),
	.w7(32'hbc45abba),
	.w8(32'hbb93500b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94c811),
	.w1(32'h39ed5c97),
	.w2(32'h3a04753f),
	.w3(32'hba867c9a),
	.w4(32'h3aaa5589),
	.w5(32'h3b2d90ee),
	.w6(32'hbaa0c869),
	.w7(32'hb9bf3822),
	.w8(32'h3b56d9ba),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd1f57),
	.w1(32'h3a93cb2e),
	.w2(32'h3ac9f2a1),
	.w3(32'h3b94d50c),
	.w4(32'h3b726215),
	.w5(32'h3be9893d),
	.w6(32'h3b17fff8),
	.w7(32'hbb0fc735),
	.w8(32'h3b2f05ec),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f77f),
	.w1(32'h3b703cc2),
	.w2(32'h3c6bc2f3),
	.w3(32'h3c235d77),
	.w4(32'h3bfa039a),
	.w5(32'h3bcbfc18),
	.w6(32'h3b70a5aa),
	.w7(32'h3bdb360b),
	.w8(32'hbaa61996),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0886b6),
	.w1(32'hbb514318),
	.w2(32'hbb9fff6a),
	.w3(32'h39ecbc36),
	.w4(32'h39f6307c),
	.w5(32'hbbb19810),
	.w6(32'hbbbf7d9a),
	.w7(32'hb99a97be),
	.w8(32'hbb641004),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b090992),
	.w1(32'h3bf825bf),
	.w2(32'hbb909b6f),
	.w3(32'h3b9b6e84),
	.w4(32'hbac3f6e3),
	.w5(32'hbba2d2b9),
	.w6(32'h3b885891),
	.w7(32'h3b44af33),
	.w8(32'hbc0f2650),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda409f),
	.w1(32'hbba0cf7e),
	.w2(32'hbb0bd2bc),
	.w3(32'hbc9ab01d),
	.w4(32'hbb8da71d),
	.w5(32'hbab256dd),
	.w6(32'hbc1b2f85),
	.w7(32'h37d87bc6),
	.w8(32'hbb57fba0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49e774),
	.w1(32'h3bc9ccb8),
	.w2(32'hbbc36b6d),
	.w3(32'hbbe71c38),
	.w4(32'h3be1eec4),
	.w5(32'hbb461902),
	.w6(32'h3b3508af),
	.w7(32'h3be04bf9),
	.w8(32'hbb5e3935),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6529c1),
	.w1(32'hbb7b0bd2),
	.w2(32'h38fe785c),
	.w3(32'h3b9fae4f),
	.w4(32'h3b2c4c2f),
	.w5(32'hbb87ff1f),
	.w6(32'h3b4f84f5),
	.w7(32'hbb124b71),
	.w8(32'hbafb866e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04fc2a),
	.w1(32'hbc409dfd),
	.w2(32'h3b8b818b),
	.w3(32'hbb5daef1),
	.w4(32'hbb648063),
	.w5(32'h3bb255ff),
	.w6(32'h3b1b4688),
	.w7(32'h3b49cfc7),
	.w8(32'hbc15fd89),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35afe7),
	.w1(32'hbc015154),
	.w2(32'hbb1985d5),
	.w3(32'hbc377d8c),
	.w4(32'hbbb899f7),
	.w5(32'hb9b8bd2d),
	.w6(32'hbc1767ae),
	.w7(32'h3b12da67),
	.w8(32'hbb68889a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ab30),
	.w1(32'hbbcd1768),
	.w2(32'hbb553e5c),
	.w3(32'hbbc5a739),
	.w4(32'hbbab8666),
	.w5(32'hb9b8c84e),
	.w6(32'hbc650731),
	.w7(32'hbbc20858),
	.w8(32'hbc1c676a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c175a54),
	.w1(32'h3b250aa8),
	.w2(32'h3c92022f),
	.w3(32'h3b4473d1),
	.w4(32'h3ae89cb9),
	.w5(32'h3c301fbc),
	.w6(32'h3b3fa3e0),
	.w7(32'h3be0a379),
	.w8(32'h3bf9cddc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3c9b2),
	.w1(32'h39cc0420),
	.w2(32'h3b9da19c),
	.w3(32'h3c2bd6a6),
	.w4(32'h3c17ccda),
	.w5(32'h3c218c9c),
	.w6(32'h3bdc6690),
	.w7(32'h3bcd7cef),
	.w8(32'h3bf29911),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43518c),
	.w1(32'h3b8d0319),
	.w2(32'hb89143fb),
	.w3(32'h3b86fc65),
	.w4(32'h3be4b22b),
	.w5(32'h3ac5d7f6),
	.w6(32'h3c06226d),
	.w7(32'h3c00d2f7),
	.w8(32'hba324705),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6fc03),
	.w1(32'h3a91627d),
	.w2(32'h3a1e5db1),
	.w3(32'h3b431bf2),
	.w4(32'h3b410062),
	.w5(32'hbaef8947),
	.w6(32'h3b034def),
	.w7(32'h3bf025af),
	.w8(32'hbac15b40),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f44f),
	.w1(32'hbaa21448),
	.w2(32'h3a3dbdec),
	.w3(32'hbc1804fa),
	.w4(32'hbb787c8c),
	.w5(32'hbbb94277),
	.w6(32'hbbafa2a3),
	.w7(32'h3bde3228),
	.w8(32'hb9d8196b),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09e44d),
	.w1(32'h3bb271eb),
	.w2(32'hba18a794),
	.w3(32'hbbd8f6bf),
	.w4(32'hbb30c4ab),
	.w5(32'hbc46bba0),
	.w6(32'hba027655),
	.w7(32'h3b8fb4b6),
	.w8(32'hbc5078e7),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc703d02),
	.w1(32'hbcb609c1),
	.w2(32'h3b9adccf),
	.w3(32'hbcfefe41),
	.w4(32'hbca98c86),
	.w5(32'hbac7ac8a),
	.w6(32'hbc944201),
	.w7(32'hbafbcc79),
	.w8(32'hbc077fcc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec1bc3),
	.w1(32'hb971081c),
	.w2(32'h3be3700a),
	.w3(32'h3a3da580),
	.w4(32'h3b459bd0),
	.w5(32'h3b15ff5b),
	.w6(32'hbbba81f1),
	.w7(32'h3b10fcca),
	.w8(32'h3b3e91b6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc023ae3),
	.w1(32'hbc2020c0),
	.w2(32'hb8827e84),
	.w3(32'hbc14e5fc),
	.w4(32'hbbcb55d0),
	.w5(32'hba98d285),
	.w6(32'hbbb5042b),
	.w7(32'hba8ff152),
	.w8(32'hbbb024f4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab10ae8),
	.w1(32'hbb92e612),
	.w2(32'hbbf30b88),
	.w3(32'h3bb572cd),
	.w4(32'hbbb3d6f3),
	.w5(32'hbce2ef3f),
	.w6(32'h3b049c24),
	.w7(32'hb5395ddd),
	.w8(32'hbcf8079e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd053c88),
	.w1(32'hbce97d91),
	.w2(32'h3b8615ce),
	.w3(32'hbd505860),
	.w4(32'hbd1aeee5),
	.w5(32'h3c1fb732),
	.w6(32'hbd19800a),
	.w7(32'hbcafabd8),
	.w8(32'hbb36554d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf7ff0),
	.w1(32'hbb42afca),
	.w2(32'h39cccac5),
	.w3(32'h39900c0b),
	.w4(32'hbbbb1f67),
	.w5(32'h3b0afd28),
	.w6(32'hbbe834b6),
	.w7(32'hbb3920c5),
	.w8(32'h3b0e5906),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459f37),
	.w1(32'h3ba6a4d6),
	.w2(32'h38f15208),
	.w3(32'h3ba4c96e),
	.w4(32'h3c009cd6),
	.w5(32'h3b50a8cb),
	.w6(32'h3bb18e82),
	.w7(32'h3bc2d8eb),
	.w8(32'h3bd395b0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b63f),
	.w1(32'h3aeb4b49),
	.w2(32'h3aafcfc3),
	.w3(32'hbab0a2ef),
	.w4(32'hbaeea4a9),
	.w5(32'hb9d37aaa),
	.w6(32'h3b07a4d9),
	.w7(32'hbb57386c),
	.w8(32'h3abeb05a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe63fa),
	.w1(32'hba045ed7),
	.w2(32'hba1ff7cd),
	.w3(32'hb9597e22),
	.w4(32'h3aa3adef),
	.w5(32'hbc36019b),
	.w6(32'h3b00f43a),
	.w7(32'h3bc8876e),
	.w8(32'hbc6c4b1a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc512ec2),
	.w1(32'hbc7cd7e0),
	.w2(32'h3bbeab16),
	.w3(32'hbca38ea4),
	.w4(32'hbc5ca9fa),
	.w5(32'h379d6cc7),
	.w6(32'hbc5bc783),
	.w7(32'h3b55668e),
	.w8(32'h3bad477f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd85a8),
	.w1(32'hbc0327cd),
	.w2(32'h3bb30294),
	.w3(32'hbb17321e),
	.w4(32'hbb6d75e9),
	.w5(32'h3c0ea62c),
	.w6(32'h3b04c44f),
	.w7(32'h3b850b30),
	.w8(32'h3c09a5fc),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c156498),
	.w1(32'h3c5466ac),
	.w2(32'hba8e55f4),
	.w3(32'h3c4ac9c3),
	.w4(32'h3c7da848),
	.w5(32'hb9ada499),
	.w6(32'h3c4a61c4),
	.w7(32'h3c5b9990),
	.w8(32'h3af40d46),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac98bb4),
	.w1(32'h3aa6f04e),
	.w2(32'h3aadafb5),
	.w3(32'h3b066fc7),
	.w4(32'h3ab69028),
	.w5(32'hba007b86),
	.w6(32'h3afb2091),
	.w7(32'h3b436f7e),
	.w8(32'hb9ceebaf),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710c463),
	.w1(32'h39437cd9),
	.w2(32'h3bb277f6),
	.w3(32'h3a672033),
	.w4(32'h3b1a055c),
	.w5(32'h3c8008d1),
	.w6(32'h3a307bb0),
	.w7(32'h3b3527bd),
	.w8(32'h3c6172f0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36ac04),
	.w1(32'hbb7c6883),
	.w2(32'hbb21954b),
	.w3(32'h3b658ee0),
	.w4(32'hbbd41b2c),
	.w5(32'h3a4c9bd6),
	.w6(32'hba77ec09),
	.w7(32'hbc19d40e),
	.w8(32'h3b462804),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e9582),
	.w1(32'h39296def),
	.w2(32'h3bc1043b),
	.w3(32'h38bc1025),
	.w4(32'h39892783),
	.w5(32'h3c098f7f),
	.w6(32'h39cb8d8f),
	.w7(32'h3b3997df),
	.w8(32'h3c0062e3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55a618),
	.w1(32'hbb87570a),
	.w2(32'hbb74a366),
	.w3(32'h3be1379b),
	.w4(32'h3b2c993c),
	.w5(32'hba942066),
	.w6(32'hbbb62231),
	.w7(32'hbb851fa1),
	.w8(32'hba63d4a8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada0e96),
	.w1(32'hbc92108b),
	.w2(32'h3c011cc9),
	.w3(32'hbbc8cbe6),
	.w4(32'hbbd6d8f1),
	.w5(32'h3b92eb25),
	.w6(32'hbc11014f),
	.w7(32'hbbc65b3e),
	.w8(32'h3c1dcb40),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80710),
	.w1(32'hbbba8910),
	.w2(32'h3966996d),
	.w3(32'hbbacfc81),
	.w4(32'hbc121753),
	.w5(32'hbc1d4d12),
	.w6(32'hbc1d639d),
	.w7(32'hbbbf9a01),
	.w8(32'hbc54afa9),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule