module layer_10_featuremap_257(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88374d),
	.w1(32'h3a9c7121),
	.w2(32'h3b298dde),
	.w3(32'h39896d66),
	.w4(32'h3ac84279),
	.w5(32'hbb05dd78),
	.w6(32'h3b4b4313),
	.w7(32'h3a5b1a6e),
	.w8(32'hba3a3455),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e099),
	.w1(32'hbab67ae4),
	.w2(32'hbad9c2cf),
	.w3(32'h3b063dcc),
	.w4(32'hb8dcfb3a),
	.w5(32'h3934b485),
	.w6(32'h3b4b4f61),
	.w7(32'hbaaf6031),
	.w8(32'h3a1a7342),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9222b),
	.w1(32'hb9d475ba),
	.w2(32'hbaf14cc8),
	.w3(32'hbb5bc04d),
	.w4(32'hb841052b),
	.w5(32'h3b93b072),
	.w6(32'hbad04737),
	.w7(32'h3b880c33),
	.w8(32'h3b2b8c29),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274065),
	.w1(32'h3b341cc2),
	.w2(32'h37b7b8cd),
	.w3(32'h3bd3e252),
	.w4(32'h3ad2a04a),
	.w5(32'hbb4830ca),
	.w6(32'h3bbef47b),
	.w7(32'h3a5ad13e),
	.w8(32'hbbd7ecdd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2dc31),
	.w1(32'h3aa1ee45),
	.w2(32'h3b3a2dae),
	.w3(32'h3a711661),
	.w4(32'h3b6903bb),
	.w5(32'h3b083148),
	.w6(32'h3af22d2c),
	.w7(32'h3bcf8dd3),
	.w8(32'h3b07e414),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9720b),
	.w1(32'h39d9f37e),
	.w2(32'hbb002ab6),
	.w3(32'h3b8f388f),
	.w4(32'hba052ef6),
	.w5(32'h3b646e34),
	.w6(32'h3b4ba2a9),
	.w7(32'hbb0c565a),
	.w8(32'h3b448d65),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b1724),
	.w1(32'hbb14f425),
	.w2(32'hbacb6462),
	.w3(32'hba13f656),
	.w4(32'h38737b69),
	.w5(32'hba5ecfac),
	.w6(32'h38250fa2),
	.w7(32'h3b004698),
	.w8(32'hbb98ce49),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3474c7),
	.w1(32'h39c77a32),
	.w2(32'h357be846),
	.w3(32'hbba4e778),
	.w4(32'hbab8df4e),
	.w5(32'h3b7d04ce),
	.w6(32'h3aeb1526),
	.w7(32'hb9ec475a),
	.w8(32'h3ae16d01),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a584e),
	.w1(32'h3afd556f),
	.w2(32'h3ac21e00),
	.w3(32'h3abf4872),
	.w4(32'h3b65a535),
	.w5(32'h3ab75e98),
	.w6(32'h3a490977),
	.w7(32'h3aaaf22a),
	.w8(32'h3b1de282),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0450cb),
	.w1(32'h39d00702),
	.w2(32'hbbc19847),
	.w3(32'h3b91d4b1),
	.w4(32'hbb1d725a),
	.w5(32'hba364dc4),
	.w6(32'h3b9bde15),
	.w7(32'hbae83802),
	.w8(32'hbaaa0200),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fc954),
	.w1(32'hbb01d9a6),
	.w2(32'hbb4a142a),
	.w3(32'h3b02aa86),
	.w4(32'hba315ad7),
	.w5(32'h3b94becb),
	.w6(32'h3b423aa1),
	.w7(32'hbb46e806),
	.w8(32'h3b6fc63a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c68215),
	.w1(32'h3ac7e6cd),
	.w2(32'h3a57cc4e),
	.w3(32'hb996a4f9),
	.w4(32'hbb1329f9),
	.w5(32'hbb84f493),
	.w6(32'hba9e0e6e),
	.w7(32'h3b8b34ea),
	.w8(32'hbb5e49be),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10e822),
	.w1(32'hbb37ceaf),
	.w2(32'hbb66cbb0),
	.w3(32'hba73832c),
	.w4(32'hbb001df8),
	.w5(32'hbb8dfea3),
	.w6(32'h3aa3d96b),
	.w7(32'hbaa3193e),
	.w8(32'hbb81eb6c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c433e),
	.w1(32'h3b4c4e3f),
	.w2(32'h39b55077),
	.w3(32'h38524b99),
	.w4(32'h3b119ddc),
	.w5(32'h3aaccbed),
	.w6(32'h3b5d2ff8),
	.w7(32'hbaacf550),
	.w8(32'h3ab2d11d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f44d3),
	.w1(32'hbb44f9bc),
	.w2(32'hbb2a67c1),
	.w3(32'h3a00c543),
	.w4(32'hba078b9d),
	.w5(32'hbb475797),
	.w6(32'hba7e04d0),
	.w7(32'hba9b148e),
	.w8(32'hbb1fb3fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d9814),
	.w1(32'h3b981b14),
	.w2(32'hbc285129),
	.w3(32'h3bab22b9),
	.w4(32'hbaf93db5),
	.w5(32'h3aee9b16),
	.w6(32'h3c45a451),
	.w7(32'hbba50225),
	.w8(32'h395cfd97),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5494bc),
	.w1(32'h3ae93bab),
	.w2(32'h3a45d811),
	.w3(32'h3b923ae5),
	.w4(32'h3abf91ad),
	.w5(32'hba877de2),
	.w6(32'h3bb1c606),
	.w7(32'h3aa30410),
	.w8(32'hba83a240),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b8aad),
	.w1(32'hbb15133c),
	.w2(32'h3939dd04),
	.w3(32'hbb09c61a),
	.w4(32'hba6ecec8),
	.w5(32'hb90efe67),
	.w6(32'hbb07cf69),
	.w7(32'hbab07807),
	.w8(32'h3ac4190d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fb642),
	.w1(32'hb9df7a1c),
	.w2(32'h3b9e3742),
	.w3(32'hba1e156e),
	.w4(32'h3b01f7b3),
	.w5(32'h39fd19f1),
	.w6(32'h3aadccd5),
	.w7(32'h3b21699e),
	.w8(32'hba4b52ca),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba869be2),
	.w1(32'hbb2190e5),
	.w2(32'hbabbbe09),
	.w3(32'hba8b4231),
	.w4(32'hb938be42),
	.w5(32'hbb68b183),
	.w6(32'hba9c3fdd),
	.w7(32'hba0f2d51),
	.w8(32'hbb5e03a4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae63852),
	.w1(32'h3c508bfe),
	.w2(32'hbbbe50bb),
	.w3(32'h3c2d4d9f),
	.w4(32'h3b6384ac),
	.w5(32'h3af2c305),
	.w6(32'h3ca4794e),
	.w7(32'hbb0cf65c),
	.w8(32'hbabc2834),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a326838),
	.w1(32'hb953bad3),
	.w2(32'h397e61f1),
	.w3(32'h3a17f4ff),
	.w4(32'h3b257998),
	.w5(32'h389fc81a),
	.w6(32'hbb292b9e),
	.w7(32'hba4f78a9),
	.w8(32'hbaeac7c0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d661),
	.w1(32'hbad5b431),
	.w2(32'hbae22d14),
	.w3(32'hbbc9ad4c),
	.w4(32'hba4e4cd5),
	.w5(32'hba6bdfd5),
	.w6(32'hbb0ce8f1),
	.w7(32'h3b075ade),
	.w8(32'hb95ef8e6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba892403),
	.w1(32'h3c44f74b),
	.w2(32'hbc36e1f6),
	.w3(32'h3c5a5902),
	.w4(32'hbc008925),
	.w5(32'hbac9dc63),
	.w6(32'h3cf101f9),
	.w7(32'hbc250b6f),
	.w8(32'hb9ca0fce),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0938fb),
	.w1(32'hbb26f8a8),
	.w2(32'h3a9769aa),
	.w3(32'hbaf85a7d),
	.w4(32'hbabdb2df),
	.w5(32'h3a82976d),
	.w6(32'hbbac76b3),
	.w7(32'hbae14b13),
	.w8(32'h3943b5bb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6b099),
	.w1(32'hbb91c40d),
	.w2(32'hba46f8d7),
	.w3(32'hbb7604c2),
	.w4(32'h39662217),
	.w5(32'h3a97ff20),
	.w6(32'hbb24b2d9),
	.w7(32'h3a8272fa),
	.w8(32'hb9d632f6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5eb3c),
	.w1(32'hba71e4bb),
	.w2(32'hba8e10e7),
	.w3(32'hbb1c564a),
	.w4(32'hba799141),
	.w5(32'h3aa8f574),
	.w6(32'hbb3e7147),
	.w7(32'h3a036a1d),
	.w8(32'h3a51d5eb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a698fd),
	.w1(32'h3b71484e),
	.w2(32'h3ac82f01),
	.w3(32'h3abe5bf6),
	.w4(32'h3a310fe5),
	.w5(32'h3ab85e22),
	.w6(32'hb8040bbd),
	.w7(32'h3a1b356a),
	.w8(32'hba03edcf),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29468f),
	.w1(32'h39f49942),
	.w2(32'hb9c3d19b),
	.w3(32'hbb4bb3a4),
	.w4(32'hbb11e11d),
	.w5(32'h3adb64c2),
	.w6(32'hbb03bb55),
	.w7(32'hbb2b212e),
	.w8(32'hba10ac54),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb358461),
	.w1(32'hbbef235b),
	.w2(32'hbbce5a58),
	.w3(32'hbbde9018),
	.w4(32'hbba5b019),
	.w5(32'hbb1ca40c),
	.w6(32'hbafb9aa0),
	.w7(32'hbb19fdbb),
	.w8(32'h3b321f1d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bc198),
	.w1(32'h3b9bdff9),
	.w2(32'h3ba0cbf5),
	.w3(32'hbb4dc08e),
	.w4(32'hba0e810a),
	.w5(32'h3b9479d2),
	.w6(32'h3a158de0),
	.w7(32'hbacc8792),
	.w8(32'h3abfc831),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a437a3c),
	.w1(32'hb9aeae26),
	.w2(32'hbb558476),
	.w3(32'h396c46f8),
	.w4(32'hbb82d4e9),
	.w5(32'hbb07afe1),
	.w6(32'hbb8630b7),
	.w7(32'h3a86b38f),
	.w8(32'h390876a0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badf8ac),
	.w1(32'h3b1b43d9),
	.w2(32'h3bc8a52e),
	.w3(32'h38a8def1),
	.w4(32'h3ac8c619),
	.w5(32'hba8b4cd3),
	.w6(32'h3ab96bb7),
	.w7(32'h3ad7ad56),
	.w8(32'h3932e3dc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05f019),
	.w1(32'hbaffb3e6),
	.w2(32'hbaa9b85b),
	.w3(32'hbb380426),
	.w4(32'hbab8301a),
	.w5(32'h3ac869f9),
	.w6(32'hbb054e7e),
	.w7(32'hbba09d65),
	.w8(32'h39bf692e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e95b),
	.w1(32'hbb285c31),
	.w2(32'hbace9bbb),
	.w3(32'h3b77d92d),
	.w4(32'h3b22e017),
	.w5(32'hbba364f8),
	.w6(32'h3acd55c6),
	.w7(32'h3abb4193),
	.w8(32'hbb5bbed3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97750f0),
	.w1(32'h3be62255),
	.w2(32'h3ba8f6fd),
	.w3(32'hbad5963d),
	.w4(32'h3bca0737),
	.w5(32'h3af46b51),
	.w6(32'h3c0ac4e5),
	.w7(32'h3bcfc103),
	.w8(32'h3b5805dc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79cfad),
	.w1(32'h3a9927d8),
	.w2(32'h3aba2eda),
	.w3(32'hbaac8f75),
	.w4(32'hb91e7e2a),
	.w5(32'hbad65cc7),
	.w6(32'hbba6f34f),
	.w7(32'h3b0fcbf9),
	.w8(32'hbac55772),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9853968),
	.w1(32'hbb4a5fd6),
	.w2(32'h3aa83b1a),
	.w3(32'hbafe610b),
	.w4(32'h3b154e03),
	.w5(32'hbb900ddc),
	.w6(32'hbb8c6146),
	.w7(32'hb8d66c6a),
	.w8(32'hbb8656c7),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60bb4d),
	.w1(32'h3a4b157c),
	.w2(32'hba97a07b),
	.w3(32'hbb85cc93),
	.w4(32'hbaab3729),
	.w5(32'hba726ece),
	.w6(32'hba76030f),
	.w7(32'hbb4fac27),
	.w8(32'hbb045529),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186fd0),
	.w1(32'h3af4e5bc),
	.w2(32'h3a69f5ea),
	.w3(32'h3bd23a53),
	.w4(32'h3b1e3f83),
	.w5(32'h3aeaa375),
	.w6(32'h3b5f793d),
	.w7(32'h3a8689f8),
	.w8(32'h39b9f94c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23433b),
	.w1(32'hbaf9f17a),
	.w2(32'h3acc338b),
	.w3(32'hbbba0115),
	.w4(32'hba6bbd92),
	.w5(32'h3af99ffe),
	.w6(32'hbb39c49a),
	.w7(32'hb96ca4b7),
	.w8(32'h3a0e6aa3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7e833),
	.w1(32'hbae56350),
	.w2(32'hba1b3541),
	.w3(32'hb99a54f0),
	.w4(32'hba86b79c),
	.w5(32'hbb3d076d),
	.w6(32'hba81006a),
	.w7(32'h3b128466),
	.w8(32'hbaff53cf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5e93),
	.w1(32'h3ab404a2),
	.w2(32'h3b2caf81),
	.w3(32'hba7e8cd5),
	.w4(32'h3ad3faa5),
	.w5(32'hbba12635),
	.w6(32'h3b0a7820),
	.w7(32'h3a8edd31),
	.w8(32'hbab12100),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d6e4c),
	.w1(32'hbb976575),
	.w2(32'hbab9d3c3),
	.w3(32'hba2487d1),
	.w4(32'hb993c541),
	.w5(32'hba4bb2e8),
	.w6(32'h3b076ec7),
	.w7(32'h39d19588),
	.w8(32'h3aa1a299),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf007d9),
	.w1(32'hbb554154),
	.w2(32'h37f4307e),
	.w3(32'hbb0deec8),
	.w4(32'hb91b0a01),
	.w5(32'h394d1597),
	.w6(32'hbb4d18bc),
	.w7(32'h3ab224bb),
	.w8(32'hb9983932),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9171d9),
	.w1(32'h3ba826b6),
	.w2(32'h3b10fe2b),
	.w3(32'h38a0cfc4),
	.w4(32'hbb2bd037),
	.w5(32'h3b5b1fff),
	.w6(32'h3b135fe1),
	.w7(32'h3aa7aff8),
	.w8(32'h3ad6058d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17cdf8),
	.w1(32'hbbb0b7f0),
	.w2(32'h3aec1d47),
	.w3(32'hbbd1c85e),
	.w4(32'hbb0ca45c),
	.w5(32'h3b84359d),
	.w6(32'hbbedaa1b),
	.w7(32'h3a663c39),
	.w8(32'h3b035eac),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8d04),
	.w1(32'h39fd44fd),
	.w2(32'hb9def880),
	.w3(32'h3ba2a390),
	.w4(32'h3b6c6b9b),
	.w5(32'hbb91671b),
	.w6(32'h3b65abe8),
	.w7(32'hb93b4af2),
	.w8(32'hbb54d156),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b0331),
	.w1(32'h3ab09512),
	.w2(32'h3b2aa027),
	.w3(32'hb9729a80),
	.w4(32'hb978f038),
	.w5(32'h39f29d84),
	.w6(32'h3b20e420),
	.w7(32'hbb37a688),
	.w8(32'hbb12bf79),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5cd1),
	.w1(32'hbbaa4370),
	.w2(32'hbb0adc17),
	.w3(32'hbb945d64),
	.w4(32'h3a956e28),
	.w5(32'hbafc3219),
	.w6(32'hbb940f2c),
	.w7(32'hba01a679),
	.w8(32'hbb4ec772),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaedbb0),
	.w1(32'hbb840b57),
	.w2(32'hbae37526),
	.w3(32'hbbef1d4d),
	.w4(32'hbb5c657f),
	.w5(32'hba49b090),
	.w6(32'hbbbb12c6),
	.w7(32'hbb0ce23d),
	.w8(32'h39975719),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82983d),
	.w1(32'hbb153b64),
	.w2(32'hb9b8a65a),
	.w3(32'h3aaf3734),
	.w4(32'h3b42135e),
	.w5(32'h3b20c9a4),
	.w6(32'hba6d6449),
	.w7(32'h392d718d),
	.w8(32'hba525f88),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf0262),
	.w1(32'hbb83c769),
	.w2(32'hbba7f8a0),
	.w3(32'hbb4d9293),
	.w4(32'hba5a81e7),
	.w5(32'h3c2fca7e),
	.w6(32'hba644268),
	.w7(32'hb9641762),
	.w8(32'h3c1ec964),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd71227),
	.w1(32'hbaade0f8),
	.w2(32'h3924912a),
	.w3(32'hbb4541d5),
	.w4(32'h3a1325ce),
	.w5(32'h3b12a62b),
	.w6(32'h39c15ea4),
	.w7(32'hba01f0e1),
	.w8(32'h39c3d3ab),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba271348),
	.w1(32'h38e1913f),
	.w2(32'hbae8b312),
	.w3(32'h3b1229a3),
	.w4(32'hb9f3a338),
	.w5(32'hbab022c3),
	.w6(32'h3b246eaf),
	.w7(32'hb9b992f6),
	.w8(32'hbb099242),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9146b30),
	.w1(32'hbb18f4f7),
	.w2(32'hbb43e114),
	.w3(32'h3ae43465),
	.w4(32'h3a8cc5ff),
	.w5(32'h3b9e4c20),
	.w6(32'hba615a76),
	.w7(32'hb9c22349),
	.w8(32'h3a9248d0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f15b5),
	.w1(32'hba088c76),
	.w2(32'h3a4fa5d2),
	.w3(32'hb86f32de),
	.w4(32'h3a537e18),
	.w5(32'h3b07ec5a),
	.w6(32'hbb1504b8),
	.w7(32'hba2c5898),
	.w8(32'h3b1a62b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0b618),
	.w1(32'hbb1c41e4),
	.w2(32'hbb7d670b),
	.w3(32'hbb88da48),
	.w4(32'h3b6dc248),
	.w5(32'h3ab147ed),
	.w6(32'hb9be9975),
	.w7(32'h39b7cdeb),
	.w8(32'hba7777f6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade8217),
	.w1(32'hbbc019dd),
	.w2(32'hbb2625c2),
	.w3(32'hbba0261c),
	.w4(32'hb86ea222),
	.w5(32'h3b58ce3e),
	.w6(32'hbbbf754b),
	.w7(32'h3a595be7),
	.w8(32'hbbb15569),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c04f5),
	.w1(32'hbc13277d),
	.w2(32'h3b7b85d6),
	.w3(32'hbbe17fba),
	.w4(32'hbb5aac56),
	.w5(32'hbb8a8a97),
	.w6(32'hbc7b8044),
	.w7(32'hbaef2d65),
	.w8(32'hbb6479e6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb541f25),
	.w1(32'hba256b68),
	.w2(32'hb974b3d7),
	.w3(32'hbb885e56),
	.w4(32'hb9d21ed9),
	.w5(32'hbb1b4d7a),
	.w6(32'h3ac5f869),
	.w7(32'h3ab73a0c),
	.w8(32'hbb7ff08e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44ba33),
	.w1(32'hbb5e5373),
	.w2(32'hbbd64565),
	.w3(32'hbb83354c),
	.w4(32'hbbd1ca44),
	.w5(32'hbb08927f),
	.w6(32'hb9c1a4bb),
	.w7(32'hbb4b671e),
	.w8(32'hb9fc8ec6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf20660),
	.w1(32'hbb903660),
	.w2(32'hbb0c5541),
	.w3(32'hba1ee0e2),
	.w4(32'hbb27de86),
	.w5(32'h3a0a3dd3),
	.w6(32'hba47b7a9),
	.w7(32'hba229f71),
	.w8(32'h39c1f488),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7993),
	.w1(32'hba7b07b0),
	.w2(32'h3afaf185),
	.w3(32'hb99a7ec8),
	.w4(32'h3b138ec8),
	.w5(32'h3aa5653d),
	.w6(32'h39f23156),
	.w7(32'hb969d45c),
	.w8(32'hbab68110),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8727c8),
	.w1(32'hba12f981),
	.w2(32'hbba1c772),
	.w3(32'h3a967cfc),
	.w4(32'hbba63f67),
	.w5(32'hbab9543f),
	.w6(32'h3b21e72c),
	.w7(32'hbb99ae5f),
	.w8(32'hbb548abb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af0dc),
	.w1(32'hbb8ef56e),
	.w2(32'hbabe02a3),
	.w3(32'hbb25d9d6),
	.w4(32'hbb7c1035),
	.w5(32'hbac47ab9),
	.w6(32'hbb8c43d4),
	.w7(32'hb8c6e630),
	.w8(32'hbaafa943),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93429b2),
	.w1(32'h3ae4accc),
	.w2(32'hb990db0b),
	.w3(32'h39b42d3a),
	.w4(32'h3a273362),
	.w5(32'h3b82cf87),
	.w6(32'h3b643c0c),
	.w7(32'h3a9553c5),
	.w8(32'h3bdc0952),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431b72),
	.w1(32'hb922c26e),
	.w2(32'hbb82e40a),
	.w3(32'h3c031f28),
	.w4(32'hba8096b8),
	.w5(32'hbb0306a2),
	.w6(32'h3b7ea2e3),
	.w7(32'hbc0316ca),
	.w8(32'hbb8fcd08),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fa6b3),
	.w1(32'h3bd0a1e1),
	.w2(32'hbb612235),
	.w3(32'h3bc7533e),
	.w4(32'hba313cf9),
	.w5(32'h3a4b6c56),
	.w6(32'h3c064091),
	.w7(32'hbac5fbad),
	.w8(32'h3b53edde),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ac99c),
	.w1(32'h3a8ca0db),
	.w2(32'h3baf4f7e),
	.w3(32'hbba49f70),
	.w4(32'h3b0c856f),
	.w5(32'hbad490a0),
	.w6(32'hba8e4853),
	.w7(32'h3b5f33bf),
	.w8(32'hba55d38d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015ac1),
	.w1(32'hbb2d78d6),
	.w2(32'h3b7f0cb7),
	.w3(32'hbb36f0e6),
	.w4(32'h3a4af8ca),
	.w5(32'hba35e7a9),
	.w6(32'hbb406651),
	.w7(32'h3b799542),
	.w8(32'hbbb1ae8c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f702),
	.w1(32'h3cac1922),
	.w2(32'hbb05721b),
	.w3(32'h3bde88b4),
	.w4(32'h3baa3846),
	.w5(32'hb84e7588),
	.w6(32'h3cb297e3),
	.w7(32'h3c1ca37a),
	.w8(32'hbb625c0e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb564cf4),
	.w1(32'h39da8fa7),
	.w2(32'hbb9c93be),
	.w3(32'h3b47320d),
	.w4(32'hbadc9d9c),
	.w5(32'hba820681),
	.w6(32'h3b30a18f),
	.w7(32'h3a9d637b),
	.w8(32'hb994c4d2),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f92c6d),
	.w1(32'hbbe7da4e),
	.w2(32'hbb0bc815),
	.w3(32'hbba7e9a6),
	.w4(32'h38d93752),
	.w5(32'h39d7e55f),
	.w6(32'hbb7ff2b5),
	.w7(32'hbaf7ac6d),
	.w8(32'h3a1146a8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92817e4),
	.w1(32'h3b1bd9f4),
	.w2(32'hb82df428),
	.w3(32'h3b762d64),
	.w4(32'h3a9495b8),
	.w5(32'hba87688a),
	.w6(32'h3b21e4d5),
	.w7(32'hba8ac39f),
	.w8(32'hb7575b15),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4b0e5),
	.w1(32'h3b6d833f),
	.w2(32'h3b51c29a),
	.w3(32'h3af1263c),
	.w4(32'h3a3a356a),
	.w5(32'hbad494b8),
	.w6(32'h3ae01513),
	.w7(32'hba8516b9),
	.w8(32'hba9dfd1d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ed667),
	.w1(32'hbaecaaeb),
	.w2(32'h388719e0),
	.w3(32'hbb95a670),
	.w4(32'hba0c1ed8),
	.w5(32'hba94b693),
	.w6(32'hbae840ea),
	.w7(32'h3b0c54fb),
	.w8(32'h3a09fc40),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b504d0b),
	.w1(32'h3a5aa222),
	.w2(32'h3ba68663),
	.w3(32'hb9b682df),
	.w4(32'h3b356386),
	.w5(32'hbb4bde9a),
	.w6(32'h39a1ba6d),
	.w7(32'h3b53c46e),
	.w8(32'hbb21ea59),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe0a89),
	.w1(32'hba813857),
	.w2(32'hbaac499d),
	.w3(32'h3a86d0f8),
	.w4(32'hbb1a9485),
	.w5(32'h3ad1a5f9),
	.w6(32'hbb106eb9),
	.w7(32'hbb394882),
	.w8(32'h3afea794),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb638),
	.w1(32'h3b006c33),
	.w2(32'hba923de0),
	.w3(32'h3b284e3c),
	.w4(32'h3a9ae390),
	.w5(32'hba90e99a),
	.w6(32'h3b8ee7e3),
	.w7(32'hbb1c3d72),
	.w8(32'hbb91d81a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8de6ff),
	.w1(32'h3b06ae26),
	.w2(32'hbb07e740),
	.w3(32'h39145f3d),
	.w4(32'h3a36df00),
	.w5(32'hbb6d6e56),
	.w6(32'h3b01b565),
	.w7(32'hba6d0b36),
	.w8(32'hbaadf84c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb4746),
	.w1(32'hb9a2531e),
	.w2(32'h3b9855b2),
	.w3(32'hbb53cbc3),
	.w4(32'h3b0382a2),
	.w5(32'hbb2b639d),
	.w6(32'hb9d0b4c0),
	.w7(32'h3b463de2),
	.w8(32'hbb86df90),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa30dc4),
	.w1(32'h3b52601c),
	.w2(32'hbaee619b),
	.w3(32'hbb2cc2de),
	.w4(32'hba84efad),
	.w5(32'hba43e7f1),
	.w6(32'h3ac6d22b),
	.w7(32'h3af522b5),
	.w8(32'h3a365e87),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa440e2),
	.w1(32'h3c01cc32),
	.w2(32'hbc1d495b),
	.w3(32'h3c66ed3f),
	.w4(32'hbb8e2301),
	.w5(32'h3a8cd8a5),
	.w6(32'h3c8db8e4),
	.w7(32'hbc24c57c),
	.w8(32'hba2cf650),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c61a81),
	.w1(32'h3b45c373),
	.w2(32'h3b2476c8),
	.w3(32'hba937974),
	.w4(32'h3b683d32),
	.w5(32'hbb9d9dd3),
	.w6(32'hb988c41c),
	.w7(32'h3bc35277),
	.w8(32'hbb916cc8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b9398),
	.w1(32'hbb69399b),
	.w2(32'hbad11bf0),
	.w3(32'h38ea5f6e),
	.w4(32'hbb71a918),
	.w5(32'h3ac6cb67),
	.w6(32'hbab34ed2),
	.w7(32'hba91e32d),
	.w8(32'h3af4f422),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2caf66),
	.w1(32'hbb07e0a4),
	.w2(32'hbb0f84b0),
	.w3(32'hbbdfffc6),
	.w4(32'hb9c44ac4),
	.w5(32'h3a2016b1),
	.w6(32'hbb8e4d81),
	.w7(32'h3bc1efe3),
	.w8(32'h397281e8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3c28d),
	.w1(32'hb9917ada),
	.w2(32'hb9af510b),
	.w3(32'hba9d21b7),
	.w4(32'hbaea4823),
	.w5(32'h3b2d74e2),
	.w6(32'hbacbdd2c),
	.w7(32'h3774da18),
	.w8(32'h39e8b80a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7c0f3),
	.w1(32'hbb3ec543),
	.w2(32'hba85c9c5),
	.w3(32'hbb1095d1),
	.w4(32'h3a4be18e),
	.w5(32'h3b66f8a6),
	.w6(32'h39c5a6eb),
	.w7(32'hba85a29e),
	.w8(32'h3c0ad952),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb7073),
	.w1(32'hbbd4823a),
	.w2(32'h3c07a471),
	.w3(32'hbbf5c87e),
	.w4(32'h3b13327b),
	.w5(32'h3b1cfeb9),
	.w6(32'hbba5acb1),
	.w7(32'h3ba8fd51),
	.w8(32'h3bad6270),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba51f42),
	.w1(32'h3c29eef2),
	.w2(32'hbb46f08b),
	.w3(32'h3c30c61b),
	.w4(32'hbbbdb3dc),
	.w5(32'h3bb8e55d),
	.w6(32'h3c1e48ac),
	.w7(32'hbb6de0d6),
	.w8(32'h3baefd5c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78d8fb),
	.w1(32'hbb113c80),
	.w2(32'h37a2daa6),
	.w3(32'hba885459),
	.w4(32'hba6d6200),
	.w5(32'h39ff3335),
	.w6(32'h3a941264),
	.w7(32'h3ae85703),
	.w8(32'h39bd5cc4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b390b86),
	.w1(32'hba972856),
	.w2(32'h3a2b2b41),
	.w3(32'h3a41f2f0),
	.w4(32'h3a98f8bd),
	.w5(32'h3b1f1b73),
	.w6(32'hbb67b8e0),
	.w7(32'h3b97e0c3),
	.w8(32'h3ae85b9d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaf100),
	.w1(32'hbaac43c3),
	.w2(32'hbb2f6521),
	.w3(32'hb91732bc),
	.w4(32'hba92e2f5),
	.w5(32'hb997519f),
	.w6(32'h38bd5d3c),
	.w7(32'hbac5351d),
	.w8(32'hbb0f633a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0f4a0),
	.w1(32'h3b8362da),
	.w2(32'h3a9a3707),
	.w3(32'h3ab82b12),
	.w4(32'h3af7d372),
	.w5(32'hba506c3f),
	.w6(32'h3be95c50),
	.w7(32'h3b7ff050),
	.w8(32'hbaa48ccd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6668e4),
	.w1(32'hbaebea1c),
	.w2(32'hbb8dc26f),
	.w3(32'hba52f23c),
	.w4(32'h3b955aff),
	.w5(32'hba4f00f2),
	.w6(32'hbb682540),
	.w7(32'h3b810a1a),
	.w8(32'hba84376a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb500097),
	.w1(32'hbab8cbf3),
	.w2(32'h3ac30cfc),
	.w3(32'h3b585ef5),
	.w4(32'h3a18e28b),
	.w5(32'h3b7c2cd2),
	.w6(32'hbba0935c),
	.w7(32'h3a702171),
	.w8(32'h39c6101e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfd022),
	.w1(32'hbb8cd1b8),
	.w2(32'h3b988fb5),
	.w3(32'h3b7ca5bb),
	.w4(32'hba840b7e),
	.w5(32'hbb51ee25),
	.w6(32'h3a1d5f2d),
	.w7(32'h3ab0d7fc),
	.w8(32'hbbb9eb51),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc026d4e),
	.w1(32'hbb80e3fc),
	.w2(32'h3a834af7),
	.w3(32'hbb3ae186),
	.w4(32'h39d254b9),
	.w5(32'h3b68de75),
	.w6(32'hbaf404e1),
	.w7(32'h3a66c354),
	.w8(32'h3bab7b27),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093a70),
	.w1(32'h3ce2573b),
	.w2(32'h3c21d676),
	.w3(32'hbc49787c),
	.w4(32'h3b21a743),
	.w5(32'h38acebc3),
	.w6(32'hbac8f322),
	.w7(32'h3bbee329),
	.w8(32'hbbebe25f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44a5bd),
	.w1(32'hbb63ac9b),
	.w2(32'h3bf44d5e),
	.w3(32'hbaf32387),
	.w4(32'hb810e30e),
	.w5(32'hbbdccc2d),
	.w6(32'h3c8818e9),
	.w7(32'h3c06b2c6),
	.w8(32'hba6524b6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28ba4c),
	.w1(32'h3bd9c609),
	.w2(32'h3b8308f9),
	.w3(32'hbc18bc00),
	.w4(32'hbc10b8c1),
	.w5(32'hb98107fc),
	.w6(32'hbbc9048f),
	.w7(32'hb9dbe983),
	.w8(32'h3952e198),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4415f0),
	.w1(32'h3b32172a),
	.w2(32'h3b8fc35d),
	.w3(32'h3b8a947a),
	.w4(32'h39392295),
	.w5(32'hbbc36576),
	.w6(32'h3b84ae32),
	.w7(32'h3a008fe6),
	.w8(32'h3a9d43e0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccde13a),
	.w1(32'h3d1afbad),
	.w2(32'h3ccd0a62),
	.w3(32'hbccc3e48),
	.w4(32'hbc3bfd46),
	.w5(32'h3b208b72),
	.w6(32'hbc192ca9),
	.w7(32'hbbdb9cae),
	.w8(32'hbbdd474c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb506901),
	.w1(32'hbc38a3a3),
	.w2(32'hba0be2af),
	.w3(32'h3a45fbd0),
	.w4(32'hbb206c30),
	.w5(32'hbc096f9d),
	.w6(32'hbc568970),
	.w7(32'hbbf4d182),
	.w8(32'h3b98cfe9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c677e35),
	.w1(32'h3cb2f01c),
	.w2(32'h3b9804e8),
	.w3(32'hbca478af),
	.w4(32'hbcaa8d5d),
	.w5(32'hbbb4b97e),
	.w6(32'hbb85236e),
	.w7(32'hbbbc1e7b),
	.w8(32'hbc0685e3),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f41c),
	.w1(32'h3cd0f129),
	.w2(32'h3c216503),
	.w3(32'hbc3ea657),
	.w4(32'hbc4a56f7),
	.w5(32'hbb5c713e),
	.w6(32'hbb3725ef),
	.w7(32'h3abdd828),
	.w8(32'hbb8b26da),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc665b1e),
	.w1(32'hbc105fa3),
	.w2(32'hbb6992b5),
	.w3(32'h392ab4cd),
	.w4(32'h3b1d8f8c),
	.w5(32'hbc15620a),
	.w6(32'h3af25a64),
	.w7(32'h3bd2787a),
	.w8(32'hbc38dac9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4242ff),
	.w1(32'hb9abb87d),
	.w2(32'h3ad3015d),
	.w3(32'hbbd3761d),
	.w4(32'hbabc51fa),
	.w5(32'h3b8f6864),
	.w6(32'hbb0c5708),
	.w7(32'hba3e2e83),
	.w8(32'hbc9366b7),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfff48c),
	.w1(32'hbce586d4),
	.w2(32'hbca1d6d2),
	.w3(32'h3c5e5868),
	.w4(32'h3c8770a8),
	.w5(32'hbbdb0455),
	.w6(32'hbc0bcf8a),
	.w7(32'hbb8a199f),
	.w8(32'hbb318b2e),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a488e),
	.w1(32'h3c6cf1d0),
	.w2(32'h3c1389ba),
	.w3(32'hb9ae4eb5),
	.w4(32'hbb39e2b6),
	.w5(32'h3c35ae6d),
	.w6(32'h3bf29e9e),
	.w7(32'h3b26f023),
	.w8(32'h3bc0bea1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41a687),
	.w1(32'h3a4303b7),
	.w2(32'h3a602daf),
	.w3(32'h3bdb0f60),
	.w4(32'h3aba7c52),
	.w5(32'h3c7fafbb),
	.w6(32'h3bd775da),
	.w7(32'h3bdc650a),
	.w8(32'hbb273a4d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e91a),
	.w1(32'hbc222085),
	.w2(32'hbab3ed78),
	.w3(32'h3ca0d3ee),
	.w4(32'h3c64718f),
	.w5(32'h3a9d0adf),
	.w6(32'hbb7c3570),
	.w7(32'hba80a54d),
	.w8(32'hbc11aee1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc1fec),
	.w1(32'hbb2ada67),
	.w2(32'hbad441f4),
	.w3(32'h3ae47b49),
	.w4(32'hbbacce78),
	.w5(32'hbbeecf88),
	.w6(32'hbc958a35),
	.w7(32'hbbde9871),
	.w8(32'h3b2650c1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe7f73),
	.w1(32'h3c5d3a0f),
	.w2(32'hbc16fe39),
	.w3(32'hbc2f60ea),
	.w4(32'hbc876f91),
	.w5(32'hb9875541),
	.w6(32'h3aebbbcb),
	.w7(32'hbb015a40),
	.w8(32'hba52dd33),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e10d7),
	.w1(32'h3bf93145),
	.w2(32'h3bf10d46),
	.w3(32'hbb788f36),
	.w4(32'hbba3501d),
	.w5(32'h3bf52273),
	.w6(32'hbb1c078a),
	.w7(32'hbab1c03e),
	.w8(32'hbb9b92a9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a7882),
	.w1(32'hbc9028a8),
	.w2(32'hbbe30118),
	.w3(32'h3c80689f),
	.w4(32'h3c77f898),
	.w5(32'hbc3ead1f),
	.w6(32'h3bbfb688),
	.w7(32'h3c0f78f8),
	.w8(32'h3bef8d5c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010e29),
	.w1(32'h3c459f9e),
	.w2(32'h3c52c368),
	.w3(32'hbc2c0f5c),
	.w4(32'hbbaa70e2),
	.w5(32'hbc165b86),
	.w6(32'hbceeec3f),
	.w7(32'hbca1b9fe),
	.w8(32'hbc9d2170),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca47604),
	.w1(32'hbbead233),
	.w2(32'hbc011a81),
	.w3(32'hbbd70eed),
	.w4(32'h39bfaf75),
	.w5(32'hbca7bfc4),
	.w6(32'hbc45907b),
	.w7(32'hbc0ec16b),
	.w8(32'hbc2b7358),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6d9bf),
	.w1(32'h3cd05fa0),
	.w2(32'h3c960177),
	.w3(32'hbd078942),
	.w4(32'hbca66903),
	.w5(32'hbab4a432),
	.w6(32'hbc526805),
	.w7(32'hbc043d3d),
	.w8(32'hbbaf74a8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa22acf),
	.w1(32'h3c360bc4),
	.w2(32'h3bba563d),
	.w3(32'h3acd69cc),
	.w4(32'hbaf0557c),
	.w5(32'h3bb6c1c6),
	.w6(32'hbbc076f5),
	.w7(32'h39fc90e7),
	.w8(32'h3bb31320),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc71993),
	.w1(32'h3bd512d3),
	.w2(32'h3c3164dd),
	.w3(32'h3ba0f0d7),
	.w4(32'h3b0e68ba),
	.w5(32'h3c07d51b),
	.w6(32'h3aee4a2b),
	.w7(32'h3b0e2cdf),
	.w8(32'h3c435056),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3a0f4),
	.w1(32'h3c541780),
	.w2(32'h3bb4bfdc),
	.w3(32'h3c6ee40b),
	.w4(32'h3aa62093),
	.w5(32'h3bded1c4),
	.w6(32'h3900aa75),
	.w7(32'h3bc90731),
	.w8(32'h3bb70981),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdabd82),
	.w1(32'hbbb4f261),
	.w2(32'h3bb5a9e3),
	.w3(32'h3bc722e8),
	.w4(32'hbb53b254),
	.w5(32'h3ac6af3b),
	.w6(32'h3ac867b4),
	.w7(32'h367bc964),
	.w8(32'h3c296010),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c151cd9),
	.w1(32'h3bcffc66),
	.w2(32'h3b957a56),
	.w3(32'h3bc04d0e),
	.w4(32'hbb93f91d),
	.w5(32'h3b72e543),
	.w6(32'h3c0a7f65),
	.w7(32'h3bc7c6b1),
	.w8(32'h3b6f5293),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c646c2a),
	.w1(32'h3c382f9b),
	.w2(32'hbabbe5f2),
	.w3(32'hbb7ca7f5),
	.w4(32'hbb8ab32b),
	.w5(32'h3a807597),
	.w6(32'hbc36942f),
	.w7(32'hbc09acb5),
	.w8(32'hbc3aaf42),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcabe4a4),
	.w1(32'hbcb1964d),
	.w2(32'hbbdf8e40),
	.w3(32'h3c357500),
	.w4(32'h3bdaa58d),
	.w5(32'hbbfef612),
	.w6(32'h3bd99d4e),
	.w7(32'h3c19d703),
	.w8(32'hbb3b107b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4714e),
	.w1(32'hbb513ac0),
	.w2(32'hba0ad7cd),
	.w3(32'hbbc96426),
	.w4(32'hbc1be88f),
	.w5(32'h3c3d1297),
	.w6(32'hbbac8b99),
	.w7(32'hbb80242b),
	.w8(32'h3a12ac13),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85a3c7),
	.w1(32'hbc08cd77),
	.w2(32'hbc29ec40),
	.w3(32'h3c1b0887),
	.w4(32'h3c507d68),
	.w5(32'h3c02c2e2),
	.w6(32'h3b17bd50),
	.w7(32'h3b310a9f),
	.w8(32'h3be3837c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c328db3),
	.w1(32'h3b8fd72c),
	.w2(32'h3b8c2422),
	.w3(32'h3b3ef2bc),
	.w4(32'hbc0338f0),
	.w5(32'hbbc372df),
	.w6(32'h3bea84d9),
	.w7(32'h3b89a23b),
	.w8(32'hbc113957),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb57628),
	.w1(32'h3c705d2b),
	.w2(32'h3b0d711d),
	.w3(32'hbbc96058),
	.w4(32'hbbf13e51),
	.w5(32'hbb805d13),
	.w6(32'h3aefa53f),
	.w7(32'hbbc912af),
	.w8(32'hbb161fe9),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038be3),
	.w1(32'hbbbcc15a),
	.w2(32'h38a82029),
	.w3(32'h3bdb3a69),
	.w4(32'h3b80f521),
	.w5(32'h3b621017),
	.w6(32'h3c1686ad),
	.w7(32'h3c029a57),
	.w8(32'hbcaf7214),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6588),
	.w1(32'h3c8f9a51),
	.w2(32'h3c18acde),
	.w3(32'h39c55132),
	.w4(32'h3be5895f),
	.w5(32'h3aa5a798),
	.w6(32'hbcda191a),
	.w7(32'hbc9f98f6),
	.w8(32'hbc26523a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd2010c),
	.w1(32'hbcce591a),
	.w2(32'hbc5d1f2c),
	.w3(32'h3c394258),
	.w4(32'h3c47f8f9),
	.w5(32'h3b7e147b),
	.w6(32'hb9b1da81),
	.w7(32'h3b63871a),
	.w8(32'hbb2fcfd3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a0fea),
	.w1(32'hbca64774),
	.w2(32'hbbe6f432),
	.w3(32'h3c3fcf1c),
	.w4(32'h3bfb3894),
	.w5(32'h3c17b277),
	.w6(32'h3c2cdb96),
	.w7(32'h3c597bcd),
	.w8(32'hbbe7bea9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf881fd),
	.w1(32'hbc67ed20),
	.w2(32'hbc4062d6),
	.w3(32'h3c1dc10a),
	.w4(32'h3c065743),
	.w5(32'h3c6529e3),
	.w6(32'h3bbbfdb1),
	.w7(32'hbb1ef4f0),
	.w8(32'hbb4368b3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19ae6b),
	.w1(32'hbc81c78a),
	.w2(32'hbbab4e5a),
	.w3(32'h3cae39e0),
	.w4(32'h3c99e2a7),
	.w5(32'hbab7099b),
	.w6(32'h3b77aa45),
	.w7(32'h3ba90e98),
	.w8(32'hbc4a983a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccef1f8),
	.w1(32'hbcd1063a),
	.w2(32'hbc5c0263),
	.w3(32'h3c0b95f1),
	.w4(32'h3c3926a2),
	.w5(32'hbbbc22a6),
	.w6(32'hb9fde1e3),
	.w7(32'h3b90e56f),
	.w8(32'hbc12bb63),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a4a84),
	.w1(32'hbc8c4f36),
	.w2(32'hbb70a84b),
	.w3(32'h3baa3388),
	.w4(32'h3bae1b2e),
	.w5(32'hbb5b9eeb),
	.w6(32'h3b55333a),
	.w7(32'h3baaa7dd),
	.w8(32'hbbbbfef5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f20d9),
	.w1(32'h39cdd6a9),
	.w2(32'h3bf5fd53),
	.w3(32'hbb8435a8),
	.w4(32'hbc3420b4),
	.w5(32'h392ce711),
	.w6(32'hbbde0056),
	.w7(32'hbbc4beb4),
	.w8(32'h3bb6c81e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e40ca),
	.w1(32'h3ca68a4d),
	.w2(32'h36e1e134),
	.w3(32'hbc118338),
	.w4(32'hbc9ae2f2),
	.w5(32'h3bb281f5),
	.w6(32'hbc05ee81),
	.w7(32'hbc0f215b),
	.w8(32'h3bd67dec),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baec02a),
	.w1(32'h3ba9dde2),
	.w2(32'h3a7cdb7c),
	.w3(32'h3ae7ff9b),
	.w4(32'hbabb6ec4),
	.w5(32'hbc24b627),
	.w6(32'h3b87e7b0),
	.w7(32'hb90efe40),
	.w8(32'hbbdc40e3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb218e),
	.w1(32'hbb1253d3),
	.w2(32'h3bbb1985),
	.w3(32'h3a398d79),
	.w4(32'hb96218a6),
	.w5(32'hbaf25284),
	.w6(32'h3b887de8),
	.w7(32'h3b0aa6e6),
	.w8(32'hba4252e6),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22aa09),
	.w1(32'hbb04b31f),
	.w2(32'hbadb032a),
	.w3(32'h3c018dad),
	.w4(32'h3c3f9533),
	.w5(32'h3c1b7283),
	.w6(32'hbba140a8),
	.w7(32'h3baa4555),
	.w8(32'hbc236289),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc709f01),
	.w1(32'hbcb70190),
	.w2(32'hbc423a0a),
	.w3(32'h3c83c82b),
	.w4(32'h3c244e96),
	.w5(32'hbbf7dbbe),
	.w6(32'hbb820bb9),
	.w7(32'h3a9f91c1),
	.w8(32'h3aa48a3e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c494248),
	.w1(32'h3c751fcd),
	.w2(32'h3c0794ac),
	.w3(32'hbc6b892e),
	.w4(32'hbc8a840c),
	.w5(32'hbc014d0c),
	.w6(32'hbc1708c1),
	.w7(32'hbc118ae5),
	.w8(32'hbb642453),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ae79c),
	.w1(32'h3cb446f2),
	.w2(32'h3c1d109c),
	.w3(32'hbc2c55d5),
	.w4(32'hbc2534ed),
	.w5(32'h3bbe2506),
	.w6(32'hbc5aa10e),
	.w7(32'hbc357e55),
	.w8(32'h3bbbb069),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8457bd),
	.w1(32'h3c0c2521),
	.w2(32'hbb95e6ab),
	.w3(32'h3b8284bb),
	.w4(32'hb9a3ceea),
	.w5(32'h3b8b3fce),
	.w6(32'hbc1721fa),
	.w7(32'h3a4a111d),
	.w8(32'h3b9a05e9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e286f),
	.w1(32'h3bd08479),
	.w2(32'hbb412d0e),
	.w3(32'hbb073d86),
	.w4(32'h3c26af21),
	.w5(32'h3c2b191e),
	.w6(32'hbb226332),
	.w7(32'h3be69476),
	.w8(32'hbb2a5728),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd64e22),
	.w1(32'hbc857800),
	.w2(32'hbbbb01ff),
	.w3(32'h3cb8056f),
	.w4(32'h3cf98160),
	.w5(32'h3b8b93c0),
	.w6(32'h3c47f668),
	.w7(32'h3c861133),
	.w8(32'hba156cbe),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a80e0),
	.w1(32'h3bd3f23c),
	.w2(32'h3bc8d6ec),
	.w3(32'h3a8e826c),
	.w4(32'hbb5a9058),
	.w5(32'hbb343c4a),
	.w6(32'h3b25aceb),
	.w7(32'hba630bfa),
	.w8(32'h3bfe1fd6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0626cd),
	.w1(32'h3b27ac23),
	.w2(32'h3babfe9b),
	.w3(32'h3b96a3c6),
	.w4(32'hba18ad23),
	.w5(32'hbba5d591),
	.w6(32'h3b848080),
	.w7(32'h3c308c31),
	.w8(32'hbc0d5db0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01ebc0),
	.w1(32'h3c2463be),
	.w2(32'h3b4d2db3),
	.w3(32'hbc288d95),
	.w4(32'hbbf3e78a),
	.w5(32'hbbb4050b),
	.w6(32'hbccbe62b),
	.w7(32'hbc9f4946),
	.w8(32'hbb8ab497),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734837),
	.w1(32'hbc529c69),
	.w2(32'hb95ad6e7),
	.w3(32'h3b3718a6),
	.w4(32'h39e4c9ef),
	.w5(32'hbad496fb),
	.w6(32'h3c375a0f),
	.w7(32'h3c0e3842),
	.w8(32'hbc18d99c),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc706a4e),
	.w1(32'hbba5c30d),
	.w2(32'h3899dd66),
	.w3(32'h3bbfd6b0),
	.w4(32'h3ba9c31f),
	.w5(32'h3c32a5b1),
	.w6(32'h3c18b4e1),
	.w7(32'h3baee655),
	.w8(32'hbc3b5fc2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85d493),
	.w1(32'hbc89cb52),
	.w2(32'hbc5c63fd),
	.w3(32'h3c6209d2),
	.w4(32'h3ca791c8),
	.w5(32'h39582067),
	.w6(32'hbc2878ad),
	.w7(32'hbb6afe0f),
	.w8(32'h3c62df74),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87625c),
	.w1(32'h3c0dbe2d),
	.w2(32'h3af97fd1),
	.w3(32'hbb1a0f05),
	.w4(32'hbb4051ab),
	.w5(32'h3b4f704f),
	.w6(32'hba9e4f97),
	.w7(32'hbadf419b),
	.w8(32'h39f85a1b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb033772),
	.w1(32'hbb0c07ca),
	.w2(32'h386dafef),
	.w3(32'h3ac9a078),
	.w4(32'h3ace0c53),
	.w5(32'hbbd22108),
	.w6(32'hbb40bca7),
	.w7(32'hb97fe8ae),
	.w8(32'h390e2931),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42bc85),
	.w1(32'h3c4d41a7),
	.w2(32'h3c9636f7),
	.w3(32'hbb018286),
	.w4(32'hbbbf0d1a),
	.w5(32'hbbb815aa),
	.w6(32'hbcc8d065),
	.w7(32'hbc92ea74),
	.w8(32'hbcc2c85c),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e7804),
	.w1(32'hbc9a50e5),
	.w2(32'hbc202851),
	.w3(32'hbc08ca33),
	.w4(32'hbc8c08f3),
	.w5(32'h3aef280c),
	.w6(32'hbc442c24),
	.w7(32'hbc25e561),
	.w8(32'h3b32f13d),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c213cb6),
	.w1(32'h3bbbd941),
	.w2(32'h3c640660),
	.w3(32'hbb46aa48),
	.w4(32'hbb8b302e),
	.w5(32'hbb085f5b),
	.w6(32'h3a93ae87),
	.w7(32'h3c3bdcdd),
	.w8(32'h3bb75270),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c5d9e),
	.w1(32'h3c83148d),
	.w2(32'h3c13e598),
	.w3(32'hbc679043),
	.w4(32'hbc5c0c4b),
	.w5(32'hbb483526),
	.w6(32'hbc6bfeb8),
	.w7(32'hbc055d41),
	.w8(32'h3b5b6ab9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4b871),
	.w1(32'hbaf63d66),
	.w2(32'hbbd2b3c7),
	.w3(32'hbbaee58f),
	.w4(32'hb9de4aa9),
	.w5(32'hbb6a878e),
	.w6(32'hbbd1cd91),
	.w7(32'hbb6ff65f),
	.w8(32'h3a4d92e8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c903a33),
	.w1(32'h3ca48da5),
	.w2(32'h3c3f140d),
	.w3(32'hbc252d71),
	.w4(32'hbc077e27),
	.w5(32'hbbc02e0f),
	.w6(32'hbb58de03),
	.w7(32'hbba9d193),
	.w8(32'h3b54da88),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6aca63),
	.w1(32'h3c476023),
	.w2(32'h3c95a6b7),
	.w3(32'hbc8d8c8c),
	.w4(32'hbbf5be03),
	.w5(32'hbb2a35bf),
	.w6(32'hbcb70c30),
	.w7(32'hbcacaf85),
	.w8(32'h3b675a32),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc710c3a),
	.w1(32'hbc685252),
	.w2(32'hbc832052),
	.w3(32'h3c088369),
	.w4(32'h3c3ab895),
	.w5(32'h3c26f3de),
	.w6(32'h3ca16604),
	.w7(32'h3c09ef51),
	.w8(32'h3c911e3e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c20d1),
	.w1(32'h3b3283a9),
	.w2(32'h3b8bc199),
	.w3(32'h3bc83b67),
	.w4(32'h3ba1c721),
	.w5(32'h3c7a6c40),
	.w6(32'h3baa8b57),
	.w7(32'h3c06c576),
	.w8(32'h3a160aa5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc37c09),
	.w1(32'hbc844e01),
	.w2(32'hbba22705),
	.w3(32'h3c5fc4e3),
	.w4(32'h3ce49d65),
	.w5(32'h3a99f1e0),
	.w6(32'h3c0b71ac),
	.w7(32'h3c31d58e),
	.w8(32'h3bfd0602),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb866ce),
	.w1(32'h3c0f30fd),
	.w2(32'h3bf56626),
	.w3(32'hbb3bf100),
	.w4(32'hbc1fde07),
	.w5(32'hbbdd3afe),
	.w6(32'hbb8fc79f),
	.w7(32'hbbd36561),
	.w8(32'hbc4a21db),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc99fb8),
	.w1(32'hbc8e745c),
	.w2(32'hbb02ee7d),
	.w3(32'h3c06cace),
	.w4(32'h3bf7a63d),
	.w5(32'hbc9f598b),
	.w6(32'h3c5e8dce),
	.w7(32'h3c49b795),
	.w8(32'h3afd963b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd91a27),
	.w1(32'h3cc91430),
	.w2(32'h3c36ca2a),
	.w3(32'hbc4b93d4),
	.w4(32'hbc609dd1),
	.w5(32'hb967c5a8),
	.w6(32'h3a09f80b),
	.w7(32'hbb970f88),
	.w8(32'hbb03aa70),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29dbf5),
	.w1(32'h3b5b9b9f),
	.w2(32'h3b058fc5),
	.w3(32'h3bc177ec),
	.w4(32'hbc2a5f47),
	.w5(32'hbbbcc09c),
	.w6(32'h3b081d9d),
	.w7(32'hbb907fe6),
	.w8(32'hbc2483f7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc315fea),
	.w1(32'h3b50626a),
	.w2(32'h3c8a83d8),
	.w3(32'hbc1da8f2),
	.w4(32'hba842a14),
	.w5(32'h3b06a2f1),
	.w6(32'hb8c940da),
	.w7(32'h3bcaf322),
	.w8(32'hbaf459a7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c299e),
	.w1(32'h3bfd9e8b),
	.w2(32'h3bdd59e3),
	.w3(32'h3b20719a),
	.w4(32'hbb273bab),
	.w5(32'h3b476fda),
	.w6(32'h3bfbaec1),
	.w7(32'h3a39f3ed),
	.w8(32'hbad11860),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad609e),
	.w1(32'h3be86708),
	.w2(32'h3c0b0eab),
	.w3(32'hbac271d8),
	.w4(32'h3b6f994e),
	.w5(32'h3c1ad363),
	.w6(32'h3c15ae80),
	.w7(32'h3c1c94f3),
	.w8(32'hbb6e46dc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1a50a),
	.w1(32'hbce00372),
	.w2(32'hbc41971c),
	.w3(32'h3cdd59a1),
	.w4(32'h3cbed66d),
	.w5(32'h3a50f772),
	.w6(32'h3bca15db),
	.w7(32'h3bea3326),
	.w8(32'h3c0ba0d8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b8416),
	.w1(32'h3bd01fb3),
	.w2(32'hbb5223c0),
	.w3(32'hba33378a),
	.w4(32'hbc8635d5),
	.w5(32'h3bbaf64b),
	.w6(32'h3ac1dffc),
	.w7(32'hbb582761),
	.w8(32'hbc44d2df),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05d829),
	.w1(32'hbc9e4cd2),
	.w2(32'hbbeb57cf),
	.w3(32'h3cb78901),
	.w4(32'h3cf13ff5),
	.w5(32'hba7c3aa6),
	.w6(32'h3c4de565),
	.w7(32'h3c3c3a4e),
	.w8(32'hbaf5da40),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002197),
	.w1(32'h3c5079e0),
	.w2(32'h3c2b12fa),
	.w3(32'h3b6dc2b7),
	.w4(32'hb90cb3b0),
	.w5(32'hbc9075f9),
	.w6(32'hba9b4b8c),
	.w7(32'h3b1dfac1),
	.w8(32'h3ae25a60),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d3d5e),
	.w1(32'h3cb7e5d2),
	.w2(32'hbb09b44d),
	.w3(32'hbc8b6c9d),
	.w4(32'hbc6c9aa4),
	.w5(32'h3b21cfcd),
	.w6(32'hbc1e1e3c),
	.w7(32'hbc59eadc),
	.w8(32'hbb84c2c5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f4cd8),
	.w1(32'h3c4fc985),
	.w2(32'h3c172775),
	.w3(32'h3b355af5),
	.w4(32'hb85bc1b5),
	.w5(32'h3b61f67d),
	.w6(32'h3b879e46),
	.w7(32'h3bdaa5c2),
	.w8(32'h3b6ca800),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58579c),
	.w1(32'h3b89194c),
	.w2(32'h3c1eb41b),
	.w3(32'hbb2e3a6d),
	.w4(32'hbbef8656),
	.w5(32'h3b018aa1),
	.w6(32'h3a798658),
	.w7(32'hbb302533),
	.w8(32'h3b79d555),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c689b06),
	.w1(32'h3c29cd1a),
	.w2(32'hbb764fbf),
	.w3(32'hbbcea692),
	.w4(32'hbc517471),
	.w5(32'hbc07a4cb),
	.w6(32'hbc5abf27),
	.w7(32'hbb9b2933),
	.w8(32'h3b23c464),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd774f1),
	.w1(32'h3b8c181f),
	.w2(32'hbb17e260),
	.w3(32'hbb885434),
	.w4(32'hbbece651),
	.w5(32'h3a60e7d3),
	.w6(32'hbc2b9e16),
	.w7(32'hbbe2848a),
	.w8(32'h3b64789b),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08600a),
	.w1(32'h3b21d979),
	.w2(32'hba181b8b),
	.w3(32'hbb06440c),
	.w4(32'hbb8231c9),
	.w5(32'h3b9b48a3),
	.w6(32'hbb9af953),
	.w7(32'hbba3427e),
	.w8(32'h3b501c03),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf67dcb),
	.w1(32'h3bdca8ad),
	.w2(32'hbb0a27c9),
	.w3(32'hbb378258),
	.w4(32'h3b5bd1fd),
	.w5(32'h3b8e488e),
	.w6(32'hbb808162),
	.w7(32'h3968fdcf),
	.w8(32'hbc732b3f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfe23d3),
	.w1(32'hbcbe0e98),
	.w2(32'hbc0a4396),
	.w3(32'h3c8cdcac),
	.w4(32'h3c9aaad8),
	.w5(32'h3aa3a71f),
	.w6(32'h3c1173f2),
	.w7(32'h3bd3802a),
	.w8(32'hbbe3795e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6b669),
	.w1(32'h39c08f36),
	.w2(32'hbb436f01),
	.w3(32'h3c18276e),
	.w4(32'h3bc0ccfa),
	.w5(32'h3c408de8),
	.w6(32'h3c95d349),
	.w7(32'h3b1c7c28),
	.w8(32'h3b3e89ee),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91fb9a),
	.w1(32'hbb1c417e),
	.w2(32'h38bdbb1e),
	.w3(32'h3c4664b1),
	.w4(32'h3c2b23c7),
	.w5(32'h3b4c4089),
	.w6(32'h3ac0bb12),
	.w7(32'h3b84ecce),
	.w8(32'hbc39bd32),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64f6b1),
	.w1(32'hbc34f051),
	.w2(32'h3a11f140),
	.w3(32'h3c484cd4),
	.w4(32'h3bd4ca40),
	.w5(32'hbb24b072),
	.w6(32'h3bdc10d7),
	.w7(32'h3c3b28e5),
	.w8(32'hbba61a1d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eba5b),
	.w1(32'h3c4d5554),
	.w2(32'h39052889),
	.w3(32'hbc46075e),
	.w4(32'hbbfa65ba),
	.w5(32'h3940156a),
	.w6(32'hbca14dbd),
	.w7(32'hbc609159),
	.w8(32'h3bfd0000),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24471),
	.w1(32'h3c15307f),
	.w2(32'hb9538280),
	.w3(32'hba9e39ef),
	.w4(32'hbb81fc16),
	.w5(32'h3bb0c50c),
	.w6(32'hbb148c87),
	.w7(32'hbc00bb68),
	.w8(32'h3c08994d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5201b1),
	.w1(32'h3b4d6ec2),
	.w2(32'hbb69c775),
	.w3(32'h3aec52a7),
	.w4(32'h3a462935),
	.w5(32'hbaf64bb5),
	.w6(32'hbc005bd9),
	.w7(32'hbae24818),
	.w8(32'hbb5da4d0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b685dbc),
	.w1(32'h3c1f412a),
	.w2(32'h3ab5f49a),
	.w3(32'hbb947bfa),
	.w4(32'hbbbbd169),
	.w5(32'h3b949b1a),
	.w6(32'hbc9c87f3),
	.w7(32'hbafdad00),
	.w8(32'hbb0d4274),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d236a),
	.w1(32'h3a402dec),
	.w2(32'hbbb4f7a9),
	.w3(32'h3c29cb8b),
	.w4(32'h3c123d60),
	.w5(32'h3b8b6509),
	.w6(32'h3b15b936),
	.w7(32'hbb1eeaa3),
	.w8(32'h396d74de),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dc458),
	.w1(32'hbba810ff),
	.w2(32'h3b3528ed),
	.w3(32'h3bfa1353),
	.w4(32'hbb0b1d2e),
	.w5(32'h3b2a8da0),
	.w6(32'h3bca552f),
	.w7(32'h3b3a9e4e),
	.w8(32'h3b413316),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8459dd),
	.w1(32'hbbcda695),
	.w2(32'h3843015d),
	.w3(32'h3ab41729),
	.w4(32'hba7a31c8),
	.w5(32'hbbad268f),
	.w6(32'h3a7919d2),
	.w7(32'h3c3c540a),
	.w8(32'hbb5045ab),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba2444),
	.w1(32'h3c23fd20),
	.w2(32'hba722a54),
	.w3(32'hbb737a42),
	.w4(32'hbc4d7e8b),
	.w5(32'hbc2d4b45),
	.w6(32'h3bac30b8),
	.w7(32'hbc23b7b7),
	.w8(32'h3a895dce),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2973dc),
	.w1(32'h3c0e0842),
	.w2(32'h3bfc5cfe),
	.w3(32'hbc0c9f2d),
	.w4(32'hbbe9c370),
	.w5(32'h3bb32bde),
	.w6(32'h3be885d8),
	.w7(32'hb97b5082),
	.w8(32'h3c023edf),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba858d4),
	.w1(32'hba9a87e5),
	.w2(32'hbbbf7b4f),
	.w3(32'hbb720009),
	.w4(32'h3ac63ff9),
	.w5(32'h3a36c342),
	.w6(32'h3a859126),
	.w7(32'h3b0d16fc),
	.w8(32'h3c63d786),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0bf02),
	.w1(32'h3b840869),
	.w2(32'h3b187458),
	.w3(32'h3a55145b),
	.w4(32'h3acbdf4c),
	.w5(32'hbbcc5514),
	.w6(32'h3c15775f),
	.w7(32'h3ac6bc61),
	.w8(32'h3b808187),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266f68),
	.w1(32'h3c538123),
	.w2(32'h3b17a3fc),
	.w3(32'hbcb23a87),
	.w4(32'hbc886e49),
	.w5(32'h3c12a99c),
	.w6(32'hbc945cbf),
	.w7(32'hbc7d4b7b),
	.w8(32'h3a9ad300),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e22f),
	.w1(32'hbbad2b5f),
	.w2(32'hbb88f080),
	.w3(32'h3c80fc89),
	.w4(32'h3c2125c7),
	.w5(32'hbc1cbe8e),
	.w6(32'hbaea2276),
	.w7(32'hbb27429d),
	.w8(32'h3c1947db),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1cb897),
	.w1(32'h3d00750c),
	.w2(32'h3c37524f),
	.w3(32'hbce5720c),
	.w4(32'hbd18c9fe),
	.w5(32'h390b6db0),
	.w6(32'hbc624a54),
	.w7(32'hbca094de),
	.w8(32'hbb3bc5b7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7602e6),
	.w1(32'h3c1670ab),
	.w2(32'h3c4d7993),
	.w3(32'h3a472842),
	.w4(32'hbb73dc99),
	.w5(32'hbc3b3056),
	.w6(32'hbbd3d122),
	.w7(32'hba95d454),
	.w8(32'hbc0c4204),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fdfc0),
	.w1(32'h3c8681e4),
	.w2(32'h3c54df04),
	.w3(32'hbc7e1ec3),
	.w4(32'hbc2688f9),
	.w5(32'h3b17fc26),
	.w6(32'hbc84e5b0),
	.w7(32'hbbf0f11e),
	.w8(32'hbb1ae371),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdca7bc),
	.w1(32'hbb809238),
	.w2(32'hbb9c81af),
	.w3(32'h3b3cc4b8),
	.w4(32'h3b41d434),
	.w5(32'h3c64d959),
	.w6(32'hba8ccc91),
	.w7(32'hba3ece7a),
	.w8(32'hbb625a8b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f828c),
	.w1(32'hbc63a20e),
	.w2(32'hbb95c9dd),
	.w3(32'h3c950728),
	.w4(32'h3c6f14e8),
	.w5(32'h3b17e2b7),
	.w6(32'h3b1ba785),
	.w7(32'h3b9a22c0),
	.w8(32'h3c408c1c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98d8b5),
	.w1(32'h3bd1bf9c),
	.w2(32'h3a7826b6),
	.w3(32'hbb1a232b),
	.w4(32'hbbb8fc5f),
	.w5(32'hbc37c31c),
	.w6(32'h3c5cab9b),
	.w7(32'h3b2d443f),
	.w8(32'h3b84ed37),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cae62),
	.w1(32'h3caae434),
	.w2(32'h3b977f57),
	.w3(32'hbc915db3),
	.w4(32'hbc9ec645),
	.w5(32'hba814f0b),
	.w6(32'hbc64846b),
	.w7(32'hbc8a2120),
	.w8(32'h393b6bb8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be40373),
	.w1(32'h3c07ac81),
	.w2(32'h3c30a517),
	.w3(32'hbb0cd5f4),
	.w4(32'hbb2dc8b8),
	.w5(32'hbba73737),
	.w6(32'h3baae20d),
	.w7(32'h3b8b5b88),
	.w8(32'hbc0b1ad2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ff8bf),
	.w1(32'hbc17a259),
	.w2(32'h3b47147c),
	.w3(32'h3aa8324b),
	.w4(32'hbaeb9765),
	.w5(32'h3b3fc576),
	.w6(32'hba88f306),
	.w7(32'h3b0cc1f6),
	.w8(32'hbbd26bcc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adedde6),
	.w1(32'h3b37563c),
	.w2(32'h3aaf3bf0),
	.w3(32'hbb56c1ab),
	.w4(32'hbbde740b),
	.w5(32'h3ba7f5d2),
	.w6(32'hbbeb7990),
	.w7(32'hbbe39ad6),
	.w8(32'h3a09995c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c09a9),
	.w1(32'hbc8e2ef4),
	.w2(32'hbc080510),
	.w3(32'h3b8c4b10),
	.w4(32'h3a02e58d),
	.w5(32'h3a02a52c),
	.w6(32'hbb134281),
	.w7(32'h3c63981e),
	.w8(32'hbc2fe0b3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74ead7),
	.w1(32'h3b26e282),
	.w2(32'hbacf5adf),
	.w3(32'h3b96e261),
	.w4(32'h3aef6e37),
	.w5(32'hbbcd5059),
	.w6(32'h3baf6348),
	.w7(32'hba811d9b),
	.w8(32'hbbcee944),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880de9),
	.w1(32'h3c3ad9b3),
	.w2(32'h3ad663fe),
	.w3(32'hbc082809),
	.w4(32'hbb7ebb58),
	.w5(32'h3bb0fd45),
	.w6(32'hbc93ba4f),
	.w7(32'hbbf20119),
	.w8(32'hbc519583),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fb19f),
	.w1(32'hbcb1b119),
	.w2(32'hbbe4bfdc),
	.w3(32'h3c8ce56d),
	.w4(32'h3c65cd12),
	.w5(32'h394b1ba5),
	.w6(32'h3b57e1e2),
	.w7(32'h3bff594a),
	.w8(32'hbb8e4d43),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b34bb8),
	.w1(32'hbb4191c4),
	.w2(32'h3be35e5b),
	.w3(32'h3bb49e45),
	.w4(32'hbb5f5baa),
	.w5(32'hb989d6fc),
	.w6(32'h39c8ae51),
	.w7(32'hb6319128),
	.w8(32'hbab3d7bd),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d1116),
	.w1(32'hbaaac199),
	.w2(32'h3bc24576),
	.w3(32'h3b83f5b2),
	.w4(32'hbbf6bcfe),
	.w5(32'h3b0fe8f0),
	.w6(32'hbafbdfcd),
	.w7(32'h3aee105f),
	.w8(32'h3c1a85a0),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b45eb),
	.w1(32'hbb56616d),
	.w2(32'h3c170807),
	.w3(32'hbb23b61c),
	.w4(32'h3b5bf9d6),
	.w5(32'hbc173f35),
	.w6(32'h3b8a53a3),
	.w7(32'h3c7bd842),
	.w8(32'hbcb4f0b8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b197c69),
	.w1(32'hbc538a7c),
	.w2(32'h3bd7ca5f),
	.w3(32'hbb1290b4),
	.w4(32'hbbaca6b9),
	.w5(32'h3a568de7),
	.w6(32'hbb434244),
	.w7(32'h3b852b1f),
	.w8(32'hbbdd9c8b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8fc03c),
	.w1(32'hbb7a6c26),
	.w2(32'hbbb1a4dd),
	.w3(32'h3a8208d8),
	.w4(32'h3bc9e8b8),
	.w5(32'h3a55be80),
	.w6(32'hba6f06e7),
	.w7(32'h3a436c18),
	.w8(32'h3b3921cc),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebfcac),
	.w1(32'hbbfd3e2e),
	.w2(32'hbbc59bd0),
	.w3(32'hba8d17fd),
	.w4(32'h3c1b2908),
	.w5(32'hbc331310),
	.w6(32'h3c055ecd),
	.w7(32'h3bfb0a68),
	.w8(32'hbc867f2d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3964b5),
	.w1(32'h3c397bb5),
	.w2(32'hbc151dd2),
	.w3(32'hbaf4fb55),
	.w4(32'hbc11bfc8),
	.w5(32'h3a71b760),
	.w6(32'hbaa0686e),
	.w7(32'hbbe0d803),
	.w8(32'hbb9d5ed2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ecfe7),
	.w1(32'h3960597c),
	.w2(32'hba9a7b57),
	.w3(32'h3b918f32),
	.w4(32'h3ba43fb6),
	.w5(32'hbb8fea07),
	.w6(32'h3aaa1878),
	.w7(32'hbb5006b5),
	.w8(32'h3a1146cc),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d1d74),
	.w1(32'hbbf3837a),
	.w2(32'h3c2b43a7),
	.w3(32'h3abaf41a),
	.w4(32'hbbb768af),
	.w5(32'h3a61a392),
	.w6(32'h3aa19dde),
	.w7(32'h3c044254),
	.w8(32'h39b44e3f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976bdf),
	.w1(32'h3af5dfa4),
	.w2(32'h3ae1b2cd),
	.w3(32'h3a5dd934),
	.w4(32'h3902d453),
	.w5(32'hbafecf1a),
	.w6(32'h3a568147),
	.w7(32'h3aaf7bf3),
	.w8(32'hbb1571a0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc8da),
	.w1(32'hbaabb2f7),
	.w2(32'hbb3b88ad),
	.w3(32'hbadd58a7),
	.w4(32'hbbd9a1e3),
	.w5(32'hbbd68f30),
	.w6(32'hbb1cceb7),
	.w7(32'hbb165690),
	.w8(32'h3a6d63cc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b3a66),
	.w1(32'h3a9c1cf0),
	.w2(32'h3a5656d7),
	.w3(32'hbbf724a2),
	.w4(32'hbb6b7584),
	.w5(32'h3b142b7b),
	.w6(32'h3b2164d4),
	.w7(32'h3b2f333e),
	.w8(32'hbc07501e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb366b6b),
	.w1(32'h391d9b5d),
	.w2(32'h3a5c215b),
	.w3(32'hba06d9a4),
	.w4(32'hbb8e4233),
	.w5(32'hbb670529),
	.w6(32'hbc26d265),
	.w7(32'hbbc8068a),
	.w8(32'hba9bd4e4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee5f44),
	.w1(32'h3b1410b1),
	.w2(32'h3b23db7f),
	.w3(32'hbb9829d4),
	.w4(32'h3ac7c822),
	.w5(32'h3a159347),
	.w6(32'h3a0d03b8),
	.w7(32'h3a02d205),
	.w8(32'h3953d820),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf87e1c),
	.w1(32'hbbb9ed3f),
	.w2(32'hbb8aef38),
	.w3(32'hb60519ea),
	.w4(32'hbb1a828b),
	.w5(32'hbb483fc9),
	.w6(32'hb8e1586d),
	.w7(32'hbae78d35),
	.w8(32'hbbcddd4e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8be847),
	.w1(32'hbb7643ef),
	.w2(32'hbb1de844),
	.w3(32'hbb4439a2),
	.w4(32'hb9b1bf2a),
	.w5(32'hbb94fef7),
	.w6(32'hbbcadb72),
	.w7(32'hbb84ac34),
	.w8(32'hbad1bbac),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cfeaf),
	.w1(32'hbae7ed13),
	.w2(32'hbb05e016),
	.w3(32'hbb0935c5),
	.w4(32'hbb898a0e),
	.w5(32'h3a119a7f),
	.w6(32'h37bdbf2e),
	.w7(32'hba1f3037),
	.w8(32'h3b69e4b1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cf847),
	.w1(32'hbbb3f810),
	.w2(32'hbb811417),
	.w3(32'h3b2ff276),
	.w4(32'hba278030),
	.w5(32'h3b056dc5),
	.w6(32'hbb15b370),
	.w7(32'hbb9d34fe),
	.w8(32'h3ac21386),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd221e),
	.w1(32'h3a83186f),
	.w2(32'h3b021a45),
	.w3(32'hbb0a2f1f),
	.w4(32'h3b99f57a),
	.w5(32'h3a34ab46),
	.w6(32'h3a50f547),
	.w7(32'h3b708df1),
	.w8(32'h39690f6c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5feca),
	.w1(32'h3a85d6d7),
	.w2(32'h3b2b799b),
	.w3(32'h3b210ca2),
	.w4(32'h3a9ff3bc),
	.w5(32'h3b122c2b),
	.w6(32'h3b236bcb),
	.w7(32'h3b7a32c2),
	.w8(32'h3aa17c24),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0491b1),
	.w1(32'h3b899100),
	.w2(32'h3bb9e613),
	.w3(32'h3b5b67b3),
	.w4(32'h3c214b1c),
	.w5(32'h39c70896),
	.w6(32'hb9cff348),
	.w7(32'h3bed6697),
	.w8(32'h3ac266f8),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c3af8),
	.w1(32'h3a204341),
	.w2(32'hba6bf554),
	.w3(32'hbb4ae799),
	.w4(32'hbb1f4989),
	.w5(32'hbb994ade),
	.w6(32'hbb7eed90),
	.w7(32'hbb50b382),
	.w8(32'hbbaa092b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e5bce),
	.w1(32'h3b09cac2),
	.w2(32'h3abaa8d1),
	.w3(32'hbb459ded),
	.w4(32'hbbfe4e61),
	.w5(32'h3a92bdc3),
	.w6(32'hbac242af),
	.w7(32'hbb22420a),
	.w8(32'h3a2b9bbf),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b777377),
	.w1(32'hba06dff6),
	.w2(32'h3ac374f4),
	.w3(32'hbb13aeff),
	.w4(32'h3b0fe27d),
	.w5(32'h39767694),
	.w6(32'hbb062a8a),
	.w7(32'h3b3f2699),
	.w8(32'h3a943e47),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76f25a),
	.w1(32'hb99c272a),
	.w2(32'hba0bd269),
	.w3(32'hba841449),
	.w4(32'h3b1a892c),
	.w5(32'hbba9c811),
	.w6(32'h3b3e4d4e),
	.w7(32'h3b039d17),
	.w8(32'hbb76d6af),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97c9d4),
	.w1(32'h39564e2b),
	.w2(32'hba772edf),
	.w3(32'hbb005cca),
	.w4(32'hbb5e338e),
	.w5(32'hb9d60028),
	.w6(32'h39ee66b3),
	.w7(32'h3909906e),
	.w8(32'hbb82e6df),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b3bee),
	.w1(32'h3bdef8cf),
	.w2(32'h3b8a8eca),
	.w3(32'hba8f4324),
	.w4(32'hbb914518),
	.w5(32'hb8b953c6),
	.w6(32'hba7747ee),
	.w7(32'hba8ffb84),
	.w8(32'hb91b58c9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9ef9c),
	.w1(32'h39199405),
	.w2(32'h3af21ab2),
	.w3(32'hb8975e2a),
	.w4(32'hbb07f213),
	.w5(32'hbb37c473),
	.w6(32'hba846b8d),
	.w7(32'h3af37be3),
	.w8(32'hbb38dc31),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27e54e),
	.w1(32'hbba411cd),
	.w2(32'hbb11e076),
	.w3(32'h3b047e6d),
	.w4(32'hbaad7746),
	.w5(32'h3a4913a2),
	.w6(32'hba5a8505),
	.w7(32'hba196aab),
	.w8(32'h3a046f10),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93de67),
	.w1(32'hba2633e4),
	.w2(32'hb93a8ba4),
	.w3(32'h394c1ee3),
	.w4(32'hbabad72b),
	.w5(32'hbb2bb9ab),
	.w6(32'h397ef91a),
	.w7(32'h3a94fc57),
	.w8(32'hbba1b895),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895566),
	.w1(32'hbb630686),
	.w2(32'hbb3ab416),
	.w3(32'h3a2cbe36),
	.w4(32'hbaf1684d),
	.w5(32'h3a026096),
	.w6(32'hbb6e50df),
	.w7(32'hbb5305da),
	.w8(32'hbb560724),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db3d63),
	.w1(32'h3a8b9a93),
	.w2(32'h3b0743f5),
	.w3(32'h3a4d8123),
	.w4(32'hbb310e40),
	.w5(32'h3b29811b),
	.w6(32'hbbd2dc86),
	.w7(32'hbb82a2fe),
	.w8(32'hbad91235),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39db65b7),
	.w1(32'h3bcc0304),
	.w2(32'hbbe296ba),
	.w3(32'hbba6122f),
	.w4(32'h39d00245),
	.w5(32'hbbdb5d55),
	.w6(32'h3abb7f9d),
	.w7(32'hbac7da25),
	.w8(32'hbbf13ccc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7eb636),
	.w1(32'hbcba0852),
	.w2(32'hbc5f8bcf),
	.w3(32'hbc5f3a28),
	.w4(32'hbbf17a2a),
	.w5(32'h3bbe577b),
	.w6(32'h3abace5d),
	.w7(32'hbbad373c),
	.w8(32'hba903cde),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fffff),
	.w1(32'h3cac9191),
	.w2(32'h3a83b491),
	.w3(32'h3c678b7d),
	.w4(32'h3bbe9e9d),
	.w5(32'hbc2905da),
	.w6(32'hbbfff7db),
	.w7(32'h3962de1c),
	.w8(32'hbb009bb4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6cfd6),
	.w1(32'hbbf52152),
	.w2(32'hbbbf317f),
	.w3(32'hbcbe75e8),
	.w4(32'hbc7b6e23),
	.w5(32'hb9a93f5e),
	.w6(32'h3aadff1b),
	.w7(32'hbc20656c),
	.w8(32'hbacf5fff),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4ab9b),
	.w1(32'h3b5c5f6a),
	.w2(32'h3b2ee7df),
	.w3(32'h3b386652),
	.w4(32'h398386e4),
	.w5(32'h39460d94),
	.w6(32'hbabafa73),
	.w7(32'hba95d3cb),
	.w8(32'h3a59dd40),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d35d1),
	.w1(32'h3633aac6),
	.w2(32'hbb0caddb),
	.w3(32'hbb15bc2b),
	.w4(32'hba9ff414),
	.w5(32'hbb226bdb),
	.w6(32'hbb0ea18b),
	.w7(32'hbb358ca9),
	.w8(32'hbadf186f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb537f5d),
	.w1(32'hbb1a9780),
	.w2(32'hbb7e59fa),
	.w3(32'hbb0a3d21),
	.w4(32'hbaaac75a),
	.w5(32'h3937d1a3),
	.w6(32'h39582a9c),
	.w7(32'h3a138f2c),
	.w8(32'h3a1b72b4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule