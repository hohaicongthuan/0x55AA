module layer_10_featuremap_355(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a8064),
	.w1(32'hbb106341),
	.w2(32'hbb83d700),
	.w3(32'hb9e9663b),
	.w4(32'hbb10e4fa),
	.w5(32'hb9d8898d),
	.w6(32'h3a15fefd),
	.w7(32'hbaf586c5),
	.w8(32'h3bca2372),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad054f3),
	.w1(32'hb974c222),
	.w2(32'hba3c4cee),
	.w3(32'h3b8fb5f1),
	.w4(32'h3959dedb),
	.w5(32'hb9fd36ee),
	.w6(32'h3c029d05),
	.w7(32'hbb54ac77),
	.w8(32'hbb5ee475),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb094cd7),
	.w1(32'hbb5b009c),
	.w2(32'hbb726e44),
	.w3(32'h3b46a72e),
	.w4(32'hbbb4fb4d),
	.w5(32'hbb240969),
	.w6(32'hbc1e136e),
	.w7(32'hbaa4929f),
	.w8(32'h3a67bf3c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adc863),
	.w1(32'h3b1bfe37),
	.w2(32'h3b653bf1),
	.w3(32'hba234f40),
	.w4(32'h3986d2ba),
	.w5(32'hbc0d950b),
	.w6(32'h3b362560),
	.w7(32'h3b0e0c4e),
	.w8(32'hbc2c3791),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a126a),
	.w1(32'hbc887a41),
	.w2(32'hbc446002),
	.w3(32'hbbbe7356),
	.w4(32'hbc1521fe),
	.w5(32'hbb904fb1),
	.w6(32'hbca36d75),
	.w7(32'hbc6df5c8),
	.w8(32'hbaa93f7b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4ba92),
	.w1(32'h3b0c366c),
	.w2(32'h3b1174b0),
	.w3(32'hbb1fbed2),
	.w4(32'hbb17e40f),
	.w5(32'hbba3ba03),
	.w6(32'h3b9e9a9f),
	.w7(32'h3aeedccd),
	.w8(32'h397da2f4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c55b7),
	.w1(32'hbab98fe8),
	.w2(32'h3a97e2d8),
	.w3(32'hbb9dd636),
	.w4(32'hbb8d195d),
	.w5(32'h3a10241e),
	.w6(32'hbaaeb91b),
	.w7(32'hbb6fccdb),
	.w8(32'hbb64f7da),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc708114),
	.w1(32'hbc38f964),
	.w2(32'hbbcfbd84),
	.w3(32'hbc5543ea),
	.w4(32'hbbb1e456),
	.w5(32'hbacc71c9),
	.w6(32'hbc34d4ed),
	.w7(32'hba5aea7e),
	.w8(32'hbaf2da0b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf595),
	.w1(32'h3a884954),
	.w2(32'hb8bb693a),
	.w3(32'hbb46aa90),
	.w4(32'hbab553d5),
	.w5(32'hbb8b747b),
	.w6(32'h3ab894a4),
	.w7(32'hb95a8998),
	.w8(32'hbaab28a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b719),
	.w1(32'hb93ce955),
	.w2(32'h3afcebf0),
	.w3(32'hbbaefa27),
	.w4(32'hbb4805ae),
	.w5(32'hbb3331ee),
	.w6(32'h3aed55e4),
	.w7(32'h3aaacf0e),
	.w8(32'h3a65ce29),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc62a),
	.w1(32'h38e11f7b),
	.w2(32'h3aab6160),
	.w3(32'hbab45372),
	.w4(32'hbb17efd0),
	.w5(32'h3bad229d),
	.w6(32'h3b5b7a01),
	.w7(32'h3815646d),
	.w8(32'hbb0318f3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3009),
	.w1(32'h38a92471),
	.w2(32'hbb5086a3),
	.w3(32'h39f812cd),
	.w4(32'hba5d290c),
	.w5(32'h3ba01d9a),
	.w6(32'hbc4cdfc0),
	.w7(32'h3b1a36f0),
	.w8(32'h3c0a1126),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ca2d7),
	.w1(32'hb98a0ce0),
	.w2(32'hbb94e2e3),
	.w3(32'hbb814cb8),
	.w4(32'h3ac51939),
	.w5(32'h3bc9bd59),
	.w6(32'h3b0e28fc),
	.w7(32'hba5added),
	.w8(32'h3bdface1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cae6a4),
	.w1(32'hba4fdb72),
	.w2(32'hbabe79e3),
	.w3(32'h3b720f9e),
	.w4(32'hbadc7678),
	.w5(32'hbb75164a),
	.w6(32'hb9b99642),
	.w7(32'h3a91c2db),
	.w8(32'hba9a806d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ae4a1),
	.w1(32'h3b955535),
	.w2(32'h3b8ea627),
	.w3(32'hbb88e103),
	.w4(32'hbb38f717),
	.w5(32'hba8e050d),
	.w6(32'h3ac466e6),
	.w7(32'h3ac97785),
	.w8(32'hbb76db93),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba91f34),
	.w1(32'h3b0e1130),
	.w2(32'hbb2a4063),
	.w3(32'h3b3286b4),
	.w4(32'h3ba52109),
	.w5(32'hbb2518e0),
	.w6(32'h3bff3894),
	.w7(32'h3b674e51),
	.w8(32'h3bc4f28d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e2610),
	.w1(32'h3b079e84),
	.w2(32'hba6ce5c9),
	.w3(32'hbbb170a8),
	.w4(32'hbb48f5c1),
	.w5(32'hba643d0b),
	.w6(32'h3b6e87f5),
	.w7(32'hba75e3c4),
	.w8(32'hbb7e9ab5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17f128),
	.w1(32'hbb70a75a),
	.w2(32'hb9694bb6),
	.w3(32'hbb73183d),
	.w4(32'h3b64d58d),
	.w5(32'h3c54d280),
	.w6(32'hbbba22af),
	.w7(32'h3b0bc079),
	.w8(32'hbb230cc3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0467ee),
	.w1(32'hbafc20ca),
	.w2(32'h3a59f75b),
	.w3(32'hbb49fd54),
	.w4(32'hbba6d629),
	.w5(32'h3b7fb833),
	.w6(32'h3ace4e90),
	.w7(32'h3a0d218c),
	.w8(32'h3afa63d9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83139d),
	.w1(32'hbb61593a),
	.w2(32'hbb877c27),
	.w3(32'h3b9fba36),
	.w4(32'h3a964350),
	.w5(32'hbb565cba),
	.w6(32'hbb1b6153),
	.w7(32'h3b6a5c3d),
	.w8(32'hbab319e4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8234a7),
	.w1(32'h3b36cc46),
	.w2(32'h3937fa07),
	.w3(32'hb8a79709),
	.w4(32'hbb19d995),
	.w5(32'hbb12e9da),
	.w6(32'h3c314bd7),
	.w7(32'h3b3f2d5c),
	.w8(32'h396affd1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc5d87),
	.w1(32'h399d8f87),
	.w2(32'h3b52b037),
	.w3(32'h3aadc1e0),
	.w4(32'hb9f4c4b7),
	.w5(32'hbaef7712),
	.w6(32'h3ac6591f),
	.w7(32'h3b03eefe),
	.w8(32'h3bb7cb33),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77b907),
	.w1(32'hbc2c3499),
	.w2(32'hb905ce60),
	.w3(32'hbba32298),
	.w4(32'hbb894c51),
	.w5(32'h3a200f85),
	.w6(32'hbb0edc0d),
	.w7(32'h39fd73e2),
	.w8(32'h3c01f981),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2506),
	.w1(32'h3a313dd9),
	.w2(32'hb9cca4e3),
	.w3(32'hbb8e8e47),
	.w4(32'hbb5006f6),
	.w5(32'h3b5564a6),
	.w6(32'h38bedd74),
	.w7(32'h3af06041),
	.w8(32'hbc6cb480),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372f86ee),
	.w1(32'hbb655462),
	.w2(32'hbb415f5e),
	.w3(32'h3c325176),
	.w4(32'hbb5c8ff3),
	.w5(32'hbb938bf1),
	.w6(32'hbbdb47aa),
	.w7(32'hbbb8dba9),
	.w8(32'h38b573b1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b853a24),
	.w1(32'h3af8d914),
	.w2(32'h3b3fe0a0),
	.w3(32'hbb598db9),
	.w4(32'hba7753d7),
	.w5(32'hbac83ce1),
	.w6(32'h3b71de4e),
	.w7(32'h3a7d240e),
	.w8(32'hbaa8ece4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7b8d5),
	.w1(32'h3ab7a0ed),
	.w2(32'h3b05b514),
	.w3(32'hba61b3bf),
	.w4(32'hbaceb09d),
	.w5(32'hba593f27),
	.w6(32'h3b2b259e),
	.w7(32'hba879018),
	.w8(32'hba81c6ff),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a895cd2),
	.w1(32'hbbd07a11),
	.w2(32'hba7499db),
	.w3(32'hbaafe44a),
	.w4(32'hbaf70063),
	.w5(32'h3bf80fa8),
	.w6(32'h3b08a953),
	.w7(32'hbbde37fb),
	.w8(32'hbb5b5c2b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4767),
	.w1(32'hbac2b2aa),
	.w2(32'hba0ef99e),
	.w3(32'h3b8c318f),
	.w4(32'hbb72d792),
	.w5(32'h3aca2eb6),
	.w6(32'hbb159592),
	.w7(32'h3b2cc029),
	.w8(32'hbb501b0c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b508079),
	.w1(32'hbb2e3226),
	.w2(32'hbb14c64f),
	.w3(32'h3b8a2f4e),
	.w4(32'hbb9fb08f),
	.w5(32'h3c11d83b),
	.w6(32'h3b712e81),
	.w7(32'hbab49d0d),
	.w8(32'hbbd61930),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36c2a),
	.w1(32'hba3e0889),
	.w2(32'hb9f01d49),
	.w3(32'h3c191866),
	.w4(32'h3bfc3036),
	.w5(32'h3bc6af0c),
	.w6(32'hbb08aa7d),
	.w7(32'hbb7d1af4),
	.w8(32'hbc04ab4f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45f1cf),
	.w1(32'hbb3ae423),
	.w2(32'hbb606799),
	.w3(32'h3c1098fb),
	.w4(32'hbaad1164),
	.w5(32'hbc3229c4),
	.w6(32'hbc42f236),
	.w7(32'hbb26ac32),
	.w8(32'hbbbaa296),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e707a),
	.w1(32'h3ac230f7),
	.w2(32'h3bbf4a5d),
	.w3(32'hbc38944b),
	.w4(32'hbba9b16e),
	.w5(32'h3baeb05d),
	.w6(32'h3b2c5aac),
	.w7(32'hba0ff908),
	.w8(32'h3b90c49b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64277e),
	.w1(32'h3b721840),
	.w2(32'hbae11629),
	.w3(32'hbb9da0f8),
	.w4(32'h3b512d82),
	.w5(32'h3b1bc1e3),
	.w6(32'hbbc0eebb),
	.w7(32'hb9e104e2),
	.w8(32'hbb4a4ead),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57537),
	.w1(32'hbb8c0e28),
	.w2(32'hbb0358a6),
	.w3(32'hba8dfc70),
	.w4(32'h39f67536),
	.w5(32'h3c1ce964),
	.w6(32'hbb81a908),
	.w7(32'hbb840480),
	.w8(32'hbbe9e1a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194da6),
	.w1(32'hbc21a188),
	.w2(32'hbb9bc201),
	.w3(32'hbb913e29),
	.w4(32'hbbb9d51a),
	.w5(32'h3b7b2e56),
	.w6(32'hbbfb1cd9),
	.w7(32'hbbe8e227),
	.w8(32'hbb471b85),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fa988),
	.w1(32'hbbe5c519),
	.w2(32'hbba48cc9),
	.w3(32'hbac69be9),
	.w4(32'hbb7cc2a0),
	.w5(32'h3b312017),
	.w6(32'hbb80cdc3),
	.w7(32'hbb95e9fd),
	.w8(32'hbaebaa30),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ac8a1),
	.w1(32'h3b625861),
	.w2(32'h3b9fbf9b),
	.w3(32'h3bb77e9e),
	.w4(32'hbb8021b6),
	.w5(32'h39fc0768),
	.w6(32'h3c1557ca),
	.w7(32'hbb6d3219),
	.w8(32'hbbbed16c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43698d),
	.w1(32'hba851c01),
	.w2(32'hba21473b),
	.w3(32'h3c0dbfb3),
	.w4(32'hba4c2b68),
	.w5(32'hbc8cdbd1),
	.w6(32'h3ac38f82),
	.w7(32'hbc02dca0),
	.w8(32'hbbda3f2a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9059652),
	.w1(32'h3b38ba18),
	.w2(32'h3bfaf54a),
	.w3(32'hbb00d479),
	.w4(32'hbb5a5bc6),
	.w5(32'h3b7f202a),
	.w6(32'h3b4a2602),
	.w7(32'h3b2a75db),
	.w8(32'h3bc835ac),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d5ebc),
	.w1(32'hbaf6a5bd),
	.w2(32'hbbcdc0e2),
	.w3(32'h3b7e7ce3),
	.w4(32'h3b271e99),
	.w5(32'hbbafa115),
	.w6(32'hbbc7df42),
	.w7(32'hbc108c19),
	.w8(32'hbae75e02),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b8378),
	.w1(32'h398bba84),
	.w2(32'hba9f5069),
	.w3(32'hbaa6dd08),
	.w4(32'hbb141bde),
	.w5(32'h3c3d454a),
	.w6(32'h3af10aca),
	.w7(32'hba893d6a),
	.w8(32'h3b21d9a7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5429),
	.w1(32'hbbbba002),
	.w2(32'hb99334be),
	.w3(32'h3c66f432),
	.w4(32'h3c6aa278),
	.w5(32'h394d1683),
	.w6(32'h3b3d34a9),
	.w7(32'h3be3dff4),
	.w8(32'hb9881c48),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ccd7a),
	.w1(32'hbc11e6bf),
	.w2(32'h3b04c006),
	.w3(32'hbbfc36d3),
	.w4(32'h385f32d4),
	.w5(32'h3a9c6d6f),
	.w6(32'h3a3b61af),
	.w7(32'h39c21b46),
	.w8(32'h3c217725),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba355b09),
	.w1(32'h3b5b467a),
	.w2(32'h3b8cac2e),
	.w3(32'hbb5c4549),
	.w4(32'hbbab0451),
	.w5(32'hba134fa9),
	.w6(32'h3b114231),
	.w7(32'h3b37a175),
	.w8(32'h3b9fec56),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd92d2b),
	.w1(32'h3be27c6a),
	.w2(32'h3bcd1904),
	.w3(32'hbb397a8f),
	.w4(32'h3abeadd3),
	.w5(32'hba54ccf1),
	.w6(32'h3c3180ec),
	.w7(32'h3b8c725c),
	.w8(32'h3c0fc9e0),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1508a7),
	.w1(32'h3bbd998a),
	.w2(32'h3bf1646a),
	.w3(32'hbc0fe6ed),
	.w4(32'hbb2e00c1),
	.w5(32'hbbd100c7),
	.w6(32'h3b563c91),
	.w7(32'h3b7bba95),
	.w8(32'hbb33fa35),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f355),
	.w1(32'hba3c5343),
	.w2(32'h3b6bbb8d),
	.w3(32'hbc3538ad),
	.w4(32'hbb87c027),
	.w5(32'h3b0a2d2e),
	.w6(32'h3b9b5a1b),
	.w7(32'h3bcdbfac),
	.w8(32'h3b983d13),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaf994),
	.w1(32'h3a37c959),
	.w2(32'hba48e335),
	.w3(32'hbba949a8),
	.w4(32'hbb229671),
	.w5(32'hbb2493ec),
	.w6(32'h3b676f5e),
	.w7(32'hba24ce1d),
	.w8(32'hbb39c244),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba692bea),
	.w1(32'hbb0b03df),
	.w2(32'h3b0bf989),
	.w3(32'hba87a847),
	.w4(32'hba3cd984),
	.w5(32'h3aa6e394),
	.w6(32'hbacc2aad),
	.w7(32'h3a781042),
	.w8(32'hba13c3fd),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6fc8a),
	.w1(32'hbaf23248),
	.w2(32'hbb9cf39f),
	.w3(32'hbaa943de),
	.w4(32'h390b2263),
	.w5(32'h39b98b43),
	.w6(32'hbb9ee4e7),
	.w7(32'hbbf5ac13),
	.w8(32'hbb9263a8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6055a5),
	.w1(32'hbc09a549),
	.w2(32'hb9ed7cb7),
	.w3(32'h3bb9f866),
	.w4(32'h3b8a8d4a),
	.w5(32'h3baf8b67),
	.w6(32'hbbc649f9),
	.w7(32'h3adc10ce),
	.w8(32'h3b7ba471),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8525b57),
	.w1(32'hbbbab2d3),
	.w2(32'hbbd8fca2),
	.w3(32'h3c39b0ca),
	.w4(32'h3b233384),
	.w5(32'hbb2eda6b),
	.w6(32'hbb880cd7),
	.w7(32'hbc183223),
	.w8(32'hba617074),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42f94f),
	.w1(32'h3ad31952),
	.w2(32'h3b65d670),
	.w3(32'hbc016c13),
	.w4(32'hbbf4e54f),
	.w5(32'h3c3f5f7b),
	.w6(32'h3bac0040),
	.w7(32'h3885e4c6),
	.w8(32'h3bb9e2ff),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1db504),
	.w1(32'hbb89f63a),
	.w2(32'hbb8ff5bb),
	.w3(32'h3c0a3ef7),
	.w4(32'h3c3f2c81),
	.w5(32'h3b203e6a),
	.w6(32'hbb5ccadb),
	.w7(32'h3bb4c52b),
	.w8(32'h3adae1d5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb501a9a),
	.w1(32'hba8d7781),
	.w2(32'hbb3e244f),
	.w3(32'h3afb84e4),
	.w4(32'h3bdc4d9d),
	.w5(32'h3a0d593f),
	.w6(32'hbb8f6758),
	.w7(32'hbb85b732),
	.w8(32'hbaae2669),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69f0c7),
	.w1(32'h3b3f7645),
	.w2(32'hbb837cad),
	.w3(32'hbaa2ebde),
	.w4(32'h3b7cc0b7),
	.w5(32'hba769a55),
	.w6(32'hbb85932a),
	.w7(32'hbac5a798),
	.w8(32'h3b80e716),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d2f8c),
	.w1(32'h3bb54128),
	.w2(32'hbacbc1c2),
	.w3(32'h3adaba9e),
	.w4(32'hbb54b9fe),
	.w5(32'hbb6288ad),
	.w6(32'h3c0ac88a),
	.w7(32'hbb53aa1a),
	.w8(32'hbb48e48d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397800c4),
	.w1(32'hbb2f1249),
	.w2(32'h3a8db69a),
	.w3(32'hba2dffdd),
	.w4(32'hbab21143),
	.w5(32'hbbea32b9),
	.w6(32'hbb827568),
	.w7(32'hbaa89706),
	.w8(32'hbc10a0cd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba816c47),
	.w1(32'hbba87f1a),
	.w2(32'hbbd7d922),
	.w3(32'hbbd55898),
	.w4(32'hbc3c294b),
	.w5(32'hbab06dbb),
	.w6(32'hbabe37bd),
	.w7(32'hbb6e7a73),
	.w8(32'h3afa049f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ab007),
	.w1(32'hba4e453f),
	.w2(32'h3ae2d3d6),
	.w3(32'hbb84fed8),
	.w4(32'hbababe07),
	.w5(32'hba4931d9),
	.w6(32'h3ae713b6),
	.w7(32'h3b2f0d68),
	.w8(32'h3bb714d3),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ba831),
	.w1(32'h3b832820),
	.w2(32'h3a5f2e2f),
	.w3(32'hbb956ffe),
	.w4(32'h3a4803c2),
	.w5(32'h3bdd0dbd),
	.w6(32'h3c0615fa),
	.w7(32'h377ee6f0),
	.w8(32'h3a8c00e0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9681a),
	.w1(32'hbc133560),
	.w2(32'hbbae9b75),
	.w3(32'h3c02e68a),
	.w4(32'h3c017600),
	.w5(32'h3b1acd53),
	.w6(32'hbaa533c9),
	.w7(32'hba33ec84),
	.w8(32'h3b807027),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b422fc),
	.w1(32'h3b1e9079),
	.w2(32'hba886ec7),
	.w3(32'hbba47f27),
	.w4(32'h38c576e1),
	.w5(32'h3baaf8ab),
	.w6(32'hbba61a8e),
	.w7(32'hbbace803),
	.w8(32'h3c30491e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bb85c),
	.w1(32'h3b90a075),
	.w2(32'h3a2f48d6),
	.w3(32'hbba82dc5),
	.w4(32'hba6067e1),
	.w5(32'h3c36f02e),
	.w6(32'hbbb58779),
	.w7(32'hbaacf3df),
	.w8(32'h3a9ed9c8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9a68),
	.w1(32'hbc36ffd2),
	.w2(32'hbc0d8c57),
	.w3(32'h3ce0cb38),
	.w4(32'h3c89b690),
	.w5(32'hbb771f0a),
	.w6(32'hbbe71d9b),
	.w7(32'hbae679ed),
	.w8(32'hbb82f643),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98fb8d),
	.w1(32'h3aff8612),
	.w2(32'h3b729d8e),
	.w3(32'hbc06c40a),
	.w4(32'h39078509),
	.w5(32'h39bdb58f),
	.w6(32'hbbd8b83b),
	.w7(32'h39c1de4e),
	.w8(32'h3be02989),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2357a5),
	.w1(32'h3c0ebc81),
	.w2(32'h3be89838),
	.w3(32'hbc181a39),
	.w4(32'hbb5ddcee),
	.w5(32'hba9ac983),
	.w6(32'h3c9df0a2),
	.w7(32'h3bd35dbf),
	.w8(32'h3c0b1a95),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9fc65),
	.w1(32'hbb8f59bd),
	.w2(32'hbb1a69b4),
	.w3(32'hbc1791c2),
	.w4(32'h3b3ac29f),
	.w5(32'h3b79f5f7),
	.w6(32'hbb8cf9aa),
	.w7(32'h3c12ebc4),
	.w8(32'h3b59bd9f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b054d),
	.w1(32'h3bc3b18d),
	.w2(32'h3ba9b597),
	.w3(32'hbb35cd2f),
	.w4(32'h3a0a154d),
	.w5(32'h3b839ff8),
	.w6(32'h3c3b6d06),
	.w7(32'h3b514f0f),
	.w8(32'hba59c082),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15c413),
	.w1(32'h3b3006f2),
	.w2(32'h399039d5),
	.w3(32'h3b3f8c29),
	.w4(32'hbaa54fe8),
	.w5(32'hba453ed4),
	.w6(32'h3b48746a),
	.w7(32'hb9ee495b),
	.w8(32'hbb9ce1e3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadae33f),
	.w1(32'h3c10ed4d),
	.w2(32'h3bb93b25),
	.w3(32'h3b28f7d8),
	.w4(32'hba874bc2),
	.w5(32'h3a9a941a),
	.w6(32'h3bae1119),
	.w7(32'h3b66c821),
	.w8(32'hbbdc9e9f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd45f14),
	.w1(32'h3bc6b5c2),
	.w2(32'h3bbe48d5),
	.w3(32'hbb089012),
	.w4(32'h3b66450f),
	.w5(32'h398a32bb),
	.w6(32'hbb8dbe45),
	.w7(32'h3a7addf3),
	.w8(32'h3b6bbeae),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bbcb4),
	.w1(32'hbb129ffb),
	.w2(32'h3a22e176),
	.w3(32'hbc11d06a),
	.w4(32'hbc0c545e),
	.w5(32'hb8caeca8),
	.w6(32'h3b16a2df),
	.w7(32'hbb8e49fa),
	.w8(32'h395ace80),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40367e),
	.w1(32'h3b3d841e),
	.w2(32'h3b22b1bf),
	.w3(32'hbaf22ce1),
	.w4(32'h3b4bc62e),
	.w5(32'h3b3bd3aa),
	.w6(32'h3b20b027),
	.w7(32'hb9f749bd),
	.w8(32'h3a1c38d2),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf71d),
	.w1(32'hbb1afcba),
	.w2(32'hbadedf05),
	.w3(32'hba99aa05),
	.w4(32'h39a7de85),
	.w5(32'h3bea14e0),
	.w6(32'hbb7af80a),
	.w7(32'hbb634251),
	.w8(32'h3c153399),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd02e2d),
	.w1(32'hbba01a8f),
	.w2(32'hb9cf53f0),
	.w3(32'h3c35d997),
	.w4(32'h39b563ef),
	.w5(32'h3b0cc268),
	.w6(32'hbb49d583),
	.w7(32'hbb6103a2),
	.w8(32'h3b9e4223),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ef83),
	.w1(32'h3b5239ad),
	.w2(32'h3ba0f5d9),
	.w3(32'h3b4dea34),
	.w4(32'h3be984a0),
	.w5(32'hbb0b929d),
	.w6(32'hbac69dba),
	.w7(32'h3b7e8188),
	.w8(32'hba672f29),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed081d),
	.w1(32'h3999a32b),
	.w2(32'h3a764416),
	.w3(32'hbbb6e917),
	.w4(32'hbb578143),
	.w5(32'hbbc1909b),
	.w6(32'h3b6c6d6a),
	.w7(32'h3b8bc6f7),
	.w8(32'hb916522f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ccbc),
	.w1(32'h3b3b78d4),
	.w2(32'h3b439ff2),
	.w3(32'hbbbf9086),
	.w4(32'hbb7661e8),
	.w5(32'hba9466b9),
	.w6(32'h3ba6b3df),
	.w7(32'hbb22c014),
	.w8(32'hbb3ac23e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d59a9),
	.w1(32'hbb2a5865),
	.w2(32'hbb3ecf70),
	.w3(32'hbb1b79e1),
	.w4(32'hbbb0ddd3),
	.w5(32'h3c15ab41),
	.w6(32'h3b3d7088),
	.w7(32'h3b6be36d),
	.w8(32'h3a5f1ca6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5bf4a),
	.w1(32'hbb92250b),
	.w2(32'hbb102192),
	.w3(32'h3aef079a),
	.w4(32'h3b551a9e),
	.w5(32'h3c26f2e7),
	.w6(32'hbaa4a776),
	.w7(32'h3b0bca78),
	.w8(32'h3c966fa7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c02c),
	.w1(32'hbb926294),
	.w2(32'h3a3fe176),
	.w3(32'h3c38c964),
	.w4(32'h3b05c8f8),
	.w5(32'hbbfc00b6),
	.w6(32'h39c71f2e),
	.w7(32'hba92827d),
	.w8(32'h3a6ac766),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ac7d8),
	.w1(32'h3c103a41),
	.w2(32'h3baec08a),
	.w3(32'hbb150057),
	.w4(32'hbb0f2735),
	.w5(32'h3c5e8bcf),
	.w6(32'h3c80819b),
	.w7(32'h3ac08ccc),
	.w8(32'h3c88afb1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf3568),
	.w1(32'hbc00dd9b),
	.w2(32'h37b916ad),
	.w3(32'h3c8c4f3a),
	.w4(32'h3b8cbeec),
	.w5(32'hbb5ad5e7),
	.w6(32'h3c03cd19),
	.w7(32'h3ab17ebe),
	.w8(32'h3b993674),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea2ab5),
	.w1(32'h3b099e40),
	.w2(32'h3a7b89a5),
	.w3(32'hbabd2e41),
	.w4(32'hbbcd43da),
	.w5(32'h3b1f67e3),
	.w6(32'h3bc66ab2),
	.w7(32'hba66deb5),
	.w8(32'h3acaa497),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51a81a),
	.w1(32'h3bf81524),
	.w2(32'hbacd70ff),
	.w3(32'h3b6c8f48),
	.w4(32'hbb4f0c66),
	.w5(32'h3c24a9c8),
	.w6(32'h3b42b40c),
	.w7(32'h3af30acf),
	.w8(32'hba105193),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa8de9),
	.w1(32'hbb994a79),
	.w2(32'h3a910a96),
	.w3(32'h3c94f298),
	.w4(32'h3bda7976),
	.w5(32'hbbb0d913),
	.w6(32'hbad1b360),
	.w7(32'h3bce5c6b),
	.w8(32'hbb17a403),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a378c14),
	.w1(32'h3ac38838),
	.w2(32'hba8b6f90),
	.w3(32'hbb8f1669),
	.w4(32'hbaa06b51),
	.w5(32'h3a0e08b1),
	.w6(32'h3b252bd7),
	.w7(32'hb9c53773),
	.w8(32'h3bf02013),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6b012),
	.w1(32'hbb8054da),
	.w2(32'h3af3756d),
	.w3(32'h3b85baa5),
	.w4(32'h3c1ad3a3),
	.w5(32'h3b0ffdc4),
	.w6(32'h3b23039f),
	.w7(32'h3b48c279),
	.w8(32'h3babd383),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b9762),
	.w1(32'hba72b13b),
	.w2(32'h3c0087be),
	.w3(32'hbafbf781),
	.w4(32'hba3f393b),
	.w5(32'hbb203970),
	.w6(32'hba9a281b),
	.w7(32'h3b565a6e),
	.w8(32'h3bbd3e8b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997c247),
	.w1(32'hbbcade05),
	.w2(32'h3b43031a),
	.w3(32'hbb997138),
	.w4(32'hbb29d361),
	.w5(32'h3bcdf9bd),
	.w6(32'hbc5fefdb),
	.w7(32'hbb253d32),
	.w8(32'h3c434392),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4038),
	.w1(32'hba12d82a),
	.w2(32'hbb003707),
	.w3(32'h3a2c74d2),
	.w4(32'h3af133a0),
	.w5(32'hbbd60126),
	.w6(32'h3b1055d8),
	.w7(32'hbb416ccb),
	.w8(32'h3b305ab6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77130e),
	.w1(32'h3b808583),
	.w2(32'h3bc5247b),
	.w3(32'hbbe17f0c),
	.w4(32'hbb66d1dd),
	.w5(32'h3ba4a650),
	.w6(32'h3a0b7f53),
	.w7(32'h3baf4e19),
	.w8(32'h3bf4bc92),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b608c7e),
	.w1(32'h3b22e488),
	.w2(32'h3a2a198d),
	.w3(32'h3bbe5739),
	.w4(32'h3b7a0368),
	.w5(32'h3c02c3c0),
	.w6(32'h3baee9c6),
	.w7(32'h3b094a80),
	.w8(32'hbb9f0bb6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e8730),
	.w1(32'hbb0e9596),
	.w2(32'hba66f9ac),
	.w3(32'h3cb313bb),
	.w4(32'h3c3498ef),
	.w5(32'hbbb6b700),
	.w6(32'hbb995004),
	.w7(32'h3bcc5985),
	.w8(32'hba237c6e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a644cc2),
	.w1(32'h3bca4eed),
	.w2(32'h3ae22c5e),
	.w3(32'hbbc83028),
	.w4(32'hbbddd5c1),
	.w5(32'h39ddc663),
	.w6(32'h3b9f0cec),
	.w7(32'h3a95dd52),
	.w8(32'h3b7785f9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf9d39),
	.w1(32'hbb0339b5),
	.w2(32'hba01c901),
	.w3(32'h3a230631),
	.w4(32'h3bc987b2),
	.w5(32'h3bc0f929),
	.w6(32'hbb93a306),
	.w7(32'hbac945cd),
	.w8(32'h3bb086a4),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e99ee),
	.w1(32'hbb182e4f),
	.w2(32'h3b15443b),
	.w3(32'hbad0810c),
	.w4(32'h3a789804),
	.w5(32'h3bcf8edb),
	.w6(32'hbb7f41d8),
	.w7(32'hbaca654b),
	.w8(32'h3b37ff6a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3464b),
	.w1(32'hbbfbc4f5),
	.w2(32'hbba6f3fe),
	.w3(32'hbbb1e778),
	.w4(32'hbb4b41e2),
	.w5(32'h3a06cd21),
	.w6(32'hbbb2268d),
	.w7(32'h3b9a2013),
	.w8(32'h3bdd7d1d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b611b2d),
	.w1(32'hbb3771bd),
	.w2(32'hbb1820a1),
	.w3(32'h39bdfc93),
	.w4(32'hbb845d37),
	.w5(32'hbbe76dfb),
	.w6(32'hbb859d90),
	.w7(32'hbc056c13),
	.w8(32'hbba64761),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90fa1c),
	.w1(32'h3b01eeca),
	.w2(32'h3aee3b55),
	.w3(32'h362f4dcc),
	.w4(32'h3b1180f3),
	.w5(32'h3acf4d5f),
	.w6(32'h3b205c72),
	.w7(32'h3c049b31),
	.w8(32'h3aa61033),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecc8cd),
	.w1(32'hbb1adf11),
	.w2(32'hbaefabaa),
	.w3(32'hb917c221),
	.w4(32'h3a98fd0e),
	.w5(32'h3b91d2b6),
	.w6(32'hb9761fdf),
	.w7(32'h3ab68716),
	.w8(32'h3bc76771),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398028c5),
	.w1(32'hbacfc824),
	.w2(32'hbb9c6cdc),
	.w3(32'h3a87aa19),
	.w4(32'hba81a226),
	.w5(32'hbb3994e7),
	.w6(32'hbb58b9cc),
	.w7(32'hbb422277),
	.w8(32'h3a7dc82d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359087),
	.w1(32'hbb4cf683),
	.w2(32'hbb31b8b7),
	.w3(32'hbb91e14d),
	.w4(32'hbadfff0a),
	.w5(32'h3a7540f2),
	.w6(32'hbb489a90),
	.w7(32'h3b819d94),
	.w8(32'hbaa063a5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda777),
	.w1(32'hb9c00e5d),
	.w2(32'h3ad2023a),
	.w3(32'hbb5f191b),
	.w4(32'hbabc5a88),
	.w5(32'hba45ab7f),
	.w6(32'hbb4e286c),
	.w7(32'h38978ca8),
	.w8(32'h3965644f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80836c6),
	.w1(32'hba173bb5),
	.w2(32'hbab4d325),
	.w3(32'hbaca0943),
	.w4(32'h3a213965),
	.w5(32'h3a8bf4eb),
	.w6(32'hb8268ded),
	.w7(32'hbb7f35e3),
	.w8(32'h39fc1b6a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b295c5d),
	.w1(32'h39f0524a),
	.w2(32'hbb10f2d3),
	.w3(32'h3a5041e5),
	.w4(32'hb9ec937b),
	.w5(32'h3b7699ab),
	.w6(32'hbb98a926),
	.w7(32'hb9fe34f2),
	.w8(32'h3b93c27d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da9b9a),
	.w1(32'hb9215114),
	.w2(32'h3a0b0758),
	.w3(32'h3951d453),
	.w4(32'hba5d3ed8),
	.w5(32'h3b13a4b7),
	.w6(32'h39814664),
	.w7(32'h36c7c834),
	.w8(32'h3a683a54),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadba1b),
	.w1(32'h3bcf33c8),
	.w2(32'h3beaabe6),
	.w3(32'h3bc6faa5),
	.w4(32'h3b1a3b3f),
	.w5(32'h3aabb0c1),
	.w6(32'h3be32c58),
	.w7(32'h3ba858cf),
	.w8(32'h3a5c00c2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc065),
	.w1(32'h3a968b43),
	.w2(32'h3b19638d),
	.w3(32'h3af340a9),
	.w4(32'h3ad72dfc),
	.w5(32'hba233895),
	.w6(32'h3aeb3d92),
	.w7(32'hbaa0b5bb),
	.w8(32'h3ab0675c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f752d),
	.w1(32'h3b1ef8a0),
	.w2(32'hbad3797b),
	.w3(32'h3ba5d5d9),
	.w4(32'h3afb094e),
	.w5(32'hbabaa7d2),
	.w6(32'h3bf2f6a0),
	.w7(32'hbad2f7fe),
	.w8(32'hbb0a22ca),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a261a05),
	.w1(32'h3b1b8c7a),
	.w2(32'h3c0c6bb8),
	.w3(32'hb97ea4db),
	.w4(32'hba27835d),
	.w5(32'h3ba73921),
	.w6(32'h3bd707ec),
	.w7(32'h3bbd5041),
	.w8(32'h3c00b72e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42f809),
	.w1(32'h3b75f883),
	.w2(32'h3947ba97),
	.w3(32'hba63390d),
	.w4(32'h3b882344),
	.w5(32'h3b69a704),
	.w6(32'hba8f6d64),
	.w7(32'h3b472030),
	.w8(32'h3b203bc9),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a840e25),
	.w1(32'h398e8979),
	.w2(32'h39662f77),
	.w3(32'hbb676db6),
	.w4(32'hbb40b0c1),
	.w5(32'hbb4b294c),
	.w6(32'hbb266cfd),
	.w7(32'hbb840dbb),
	.w8(32'h39de923d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac66614),
	.w1(32'h394253ce),
	.w2(32'hbb1c8c07),
	.w3(32'hb9a63eec),
	.w4(32'h392b6b1f),
	.w5(32'h3c09b09c),
	.w6(32'h3aaf41d2),
	.w7(32'hbab1bcc6),
	.w8(32'h3c27679a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a804f),
	.w1(32'h3bf3e954),
	.w2(32'h3b4c2f8f),
	.w3(32'h3bba284f),
	.w4(32'h3b9805f6),
	.w5(32'hbb8fb4ab),
	.w6(32'h3bc04bd9),
	.w7(32'h3b0c33c4),
	.w8(32'h39b01396),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecbbeb),
	.w1(32'hbb2a2f04),
	.w2(32'hbb7202fe),
	.w3(32'hbb83c70b),
	.w4(32'hbb184d6b),
	.w5(32'h3b1ffc28),
	.w6(32'h3a0a6579),
	.w7(32'h3b072a77),
	.w8(32'h3b432572),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b512c96),
	.w1(32'h39da7d5e),
	.w2(32'h3ab51303),
	.w3(32'hb9e88f68),
	.w4(32'h3ae3a2ea),
	.w5(32'hba01ef4b),
	.w6(32'hbaa70d39),
	.w7(32'h39dcde40),
	.w8(32'hbab8bcd6),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a140cfb),
	.w1(32'hbb118003),
	.w2(32'hbb76e46f),
	.w3(32'hbaa59dbf),
	.w4(32'hbb5a540c),
	.w5(32'hb684e7d2),
	.w6(32'hba52e666),
	.w7(32'hbb64b55f),
	.w8(32'h38e3f18d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ae858),
	.w1(32'hbac1c707),
	.w2(32'hbb061ac9),
	.w3(32'hba29e7f1),
	.w4(32'h3b057d82),
	.w5(32'h3ad4375a),
	.w6(32'h3a553d00),
	.w7(32'h3ac56948),
	.w8(32'h3a7b00d8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4c82f),
	.w1(32'hbb8fabd1),
	.w2(32'h3b652959),
	.w3(32'hbb040df1),
	.w4(32'hbbacdd0d),
	.w5(32'hbbbe5a53),
	.w6(32'hb5caf6cb),
	.w7(32'h3ad48c19),
	.w8(32'hbc022ac4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc1c24),
	.w1(32'hbb9d81e8),
	.w2(32'h3b37ae1e),
	.w3(32'h3ab68587),
	.w4(32'h3b4cb64c),
	.w5(32'hbb69c0b7),
	.w6(32'hbb32f4a7),
	.w7(32'h3b51c416),
	.w8(32'hbba3f728),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8616ae),
	.w1(32'h3b6377a8),
	.w2(32'h3be06814),
	.w3(32'hbaf99082),
	.w4(32'hbb46ad99),
	.w5(32'hbb2e3830),
	.w6(32'h3bca7b9b),
	.w7(32'h3b4e742d),
	.w8(32'hbc1b0115),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82e2e),
	.w1(32'hbb660bfd),
	.w2(32'h3afa0abb),
	.w3(32'h39d390ab),
	.w4(32'h3bc8be16),
	.w5(32'h399bf5c7),
	.w6(32'hbaafd392),
	.w7(32'h3b6e2d60),
	.w8(32'hba09ea02),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68b4bc),
	.w1(32'h39940ed0),
	.w2(32'h3b2a2b45),
	.w3(32'h3af51dbf),
	.w4(32'hba49e1d6),
	.w5(32'hbad4c324),
	.w6(32'h3b46e7b6),
	.w7(32'h3b5a5d4e),
	.w8(32'hbb15e8a3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39742c),
	.w1(32'h3aad84fa),
	.w2(32'h3b75c307),
	.w3(32'hbb719b18),
	.w4(32'hbbab5623),
	.w5(32'h39b0c572),
	.w6(32'hba794374),
	.w7(32'h3b03c632),
	.w8(32'hb9ac3fe8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980a896),
	.w1(32'hbb115c7a),
	.w2(32'hbac3f23e),
	.w3(32'hbaf36635),
	.w4(32'hbbc0012d),
	.w5(32'h3ac752d6),
	.w6(32'h3b12dc5b),
	.w7(32'h3ab13d5f),
	.w8(32'h3ae15f23),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc267637),
	.w1(32'hbb85e3de),
	.w2(32'h3ab66f69),
	.w3(32'h3a833a03),
	.w4(32'h3b50e27e),
	.w5(32'h3a8ed3fc),
	.w6(32'h3b8e4691),
	.w7(32'h3addc9af),
	.w8(32'h38842cc2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b1f1),
	.w1(32'h389ecaae),
	.w2(32'h3bb121fa),
	.w3(32'hbb0406d1),
	.w4(32'hbaa54a3f),
	.w5(32'h3b01d4d1),
	.w6(32'h3833124c),
	.w7(32'h3b020579),
	.w8(32'h3b888428),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb398dd9),
	.w1(32'hbb15781a),
	.w2(32'hbb5e5f8a),
	.w3(32'hba3c3e08),
	.w4(32'h3ae8db91),
	.w5(32'hb9f29825),
	.w6(32'h3b3dfc83),
	.w7(32'h3b155c2c),
	.w8(32'hba832121),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd95cc),
	.w1(32'hbb1579fe),
	.w2(32'hbaa834e9),
	.w3(32'hbb1bbcb2),
	.w4(32'hbae0fd85),
	.w5(32'hbb826162),
	.w6(32'hbb2d8a2a),
	.w7(32'hbac68167),
	.w8(32'h3b0f60fa),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bf7f1),
	.w1(32'hb7d09b97),
	.w2(32'h3bb127c1),
	.w3(32'hbc0c72b8),
	.w4(32'hbbb426ac),
	.w5(32'hb9d291f4),
	.w6(32'h3b00c96d),
	.w7(32'h3b1edb30),
	.w8(32'hbb072662),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08ff21),
	.w1(32'h3b84b72f),
	.w2(32'h3a6fdd26),
	.w3(32'h3b419807),
	.w4(32'h3a8175a7),
	.w5(32'h3a886416),
	.w6(32'h3b686854),
	.w7(32'h3934f0c6),
	.w8(32'h3a5639a8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbce6a),
	.w1(32'hbae0f79c),
	.w2(32'h3b187146),
	.w3(32'hbbeadf99),
	.w4(32'hbb48f1af),
	.w5(32'h3c3c9d26),
	.w6(32'hba316081),
	.w7(32'h3b067d8b),
	.w8(32'h3c4255ea),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bd2a1),
	.w1(32'hb9f1fbbc),
	.w2(32'hbb919404),
	.w3(32'h3c100063),
	.w4(32'h3b8e9d5c),
	.w5(32'h3b1f2461),
	.w6(32'h3b0d13b3),
	.w7(32'hbb1a92bf),
	.w8(32'h3ac0de70),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba741981),
	.w1(32'h3b8a69eb),
	.w2(32'h3c01baa3),
	.w3(32'h3ad92e8b),
	.w4(32'h3b8fe3b8),
	.w5(32'hbae88e35),
	.w6(32'h3b82781f),
	.w7(32'h3ba0c288),
	.w8(32'hbb140180),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bb61a),
	.w1(32'hb9b9937e),
	.w2(32'h3b3e97fc),
	.w3(32'hbb303fd7),
	.w4(32'hbb9f51f1),
	.w5(32'h3a77a6ba),
	.w6(32'h3adb9bec),
	.w7(32'h39b75102),
	.w8(32'h3b0297a7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb648c91),
	.w1(32'h3984f900),
	.w2(32'hbb0e1b99),
	.w3(32'hb9fa1c4b),
	.w4(32'hbb0857ab),
	.w5(32'h389d715f),
	.w6(32'h395068a3),
	.w7(32'hb8fd8812),
	.w8(32'h3b143631),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb550934),
	.w1(32'hbb800690),
	.w2(32'hbadbad4e),
	.w3(32'hbb88215a),
	.w4(32'hb9ee8deb),
	.w5(32'hbac229b8),
	.w6(32'hbb49eb88),
	.w7(32'hb851f908),
	.w8(32'hbb7031be),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cb40a),
	.w1(32'hbb758c6d),
	.w2(32'hb95e3d37),
	.w3(32'hbb5c97b7),
	.w4(32'hbaa2e970),
	.w5(32'h3aa76695),
	.w6(32'hbba67c25),
	.w7(32'hbb04801e),
	.w8(32'h39bf9d7d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9aab),
	.w1(32'h3a236af0),
	.w2(32'h3ac5276b),
	.w3(32'h3c07b57e),
	.w4(32'hbafeeda1),
	.w5(32'hbb713f53),
	.w6(32'h3c31fc5b),
	.w7(32'hbbd9b399),
	.w8(32'hbbe3cc77),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac76059),
	.w1(32'h3a3cb76a),
	.w2(32'hba0806fb),
	.w3(32'hbb0933ae),
	.w4(32'hba09ccb9),
	.w5(32'hba07d5c8),
	.w6(32'hbab17072),
	.w7(32'h3a0d7cb5),
	.w8(32'hbaeb5fe0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e2861),
	.w1(32'hbabe5b84),
	.w2(32'hbad5ec20),
	.w3(32'hba1e09bf),
	.w4(32'hbb4bc26c),
	.w5(32'hba937427),
	.w6(32'h3aa7edb6),
	.w7(32'hbafa4563),
	.w8(32'hbb388544),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919c2c1),
	.w1(32'h3a9aec58),
	.w2(32'h3af6627a),
	.w3(32'hba8b8476),
	.w4(32'hb8c08f3c),
	.w5(32'h3a4a782a),
	.w6(32'hbb9b2566),
	.w7(32'hb8c7e153),
	.w8(32'hb90d1145),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bc58e),
	.w1(32'h3ae2d28a),
	.w2(32'h3ba41cc7),
	.w3(32'h399e046f),
	.w4(32'h3b0f99d1),
	.w5(32'hba86213c),
	.w6(32'h3a5c72ba),
	.w7(32'h3b7b2bde),
	.w8(32'hba4340e6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a33e2),
	.w1(32'hba87afdb),
	.w2(32'hb9850e59),
	.w3(32'h39250d7b),
	.w4(32'h3a805b1d),
	.w5(32'h399da5d4),
	.w6(32'hba843e14),
	.w7(32'h3a16f83d),
	.w8(32'hbabd8835),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2039a),
	.w1(32'h3b19f49d),
	.w2(32'h3bde65e8),
	.w3(32'hbb039237),
	.w4(32'hbb4be721),
	.w5(32'hba55c563),
	.w6(32'h3b99aeed),
	.w7(32'h3b6808f7),
	.w8(32'h3a1f2ee2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d425ea),
	.w1(32'hbacac8aa),
	.w2(32'hbaa137fe),
	.w3(32'hbb211f69),
	.w4(32'hbb91cadd),
	.w5(32'h3ba23327),
	.w6(32'hbb285620),
	.w7(32'hbb4f2f7b),
	.w8(32'h3bb5019c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ac921),
	.w1(32'h397952f8),
	.w2(32'hbb23b291),
	.w3(32'h3999ce5c),
	.w4(32'h39031466),
	.w5(32'h3b159b02),
	.w6(32'hba468758),
	.w7(32'hbb17b526),
	.w8(32'h3b292080),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b18ec),
	.w1(32'h3a5bea7f),
	.w2(32'hb99a2317),
	.w3(32'h3a1bcfae),
	.w4(32'h3b6cbb94),
	.w5(32'hbb0a2d54),
	.w6(32'h3a592bc8),
	.w7(32'h3b18ec14),
	.w8(32'hba25a487),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb602d0),
	.w1(32'hbb6c8b1a),
	.w2(32'hbb1946cb),
	.w3(32'hbb26d63e),
	.w4(32'hbb9ecb2f),
	.w5(32'hba8536f1),
	.w6(32'h3b256600),
	.w7(32'hbbd0014a),
	.w8(32'h3b728a8b),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b558d83),
	.w1(32'hba386c9b),
	.w2(32'h3ad9b0f3),
	.w3(32'h3a6e3660),
	.w4(32'hba192e00),
	.w5(32'hbb0b59e3),
	.w6(32'h3aa74ce7),
	.w7(32'hbaa0795c),
	.w8(32'hbb9720e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb8117),
	.w1(32'hbaa37741),
	.w2(32'hbb8ea202),
	.w3(32'hbb368ec8),
	.w4(32'hba803abb),
	.w5(32'h3b091881),
	.w6(32'hbb48dbee),
	.w7(32'h3a020ae3),
	.w8(32'h3b746121),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b410741),
	.w1(32'h3b24eda0),
	.w2(32'h39e8d6f4),
	.w3(32'h3b63791c),
	.w4(32'h3a5973d9),
	.w5(32'h3b5ec0ab),
	.w6(32'h3b98cccb),
	.w7(32'h3a7212f6),
	.w8(32'h3b2581a4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b369a),
	.w1(32'h3c014af1),
	.w2(32'h3c3f9d4f),
	.w3(32'h3bd843f4),
	.w4(32'h3b00e92b),
	.w5(32'hbb0f5f11),
	.w6(32'h3c29b198),
	.w7(32'h3bca1579),
	.w8(32'hbafdf252),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bccaa),
	.w1(32'hbb2e5868),
	.w2(32'h3afef08f),
	.w3(32'h3a65d2a6),
	.w4(32'hba97de44),
	.w5(32'hba1a4c7f),
	.w6(32'h3af0d97a),
	.w7(32'h3a087478),
	.w8(32'hba3e8d0c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42f91d),
	.w1(32'hb976e573),
	.w2(32'h3aac8a8b),
	.w3(32'hb9256376),
	.w4(32'hbb568400),
	.w5(32'hbb0e8b53),
	.w6(32'h3bbe739b),
	.w7(32'hba917beb),
	.w8(32'h3b851915),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab28d5c),
	.w1(32'hbb55355f),
	.w2(32'hbb2ba8a6),
	.w3(32'hbb246d84),
	.w4(32'hbb2a882e),
	.w5(32'h3b5c2ddc),
	.w6(32'h3a773a5b),
	.w7(32'h3bc08065),
	.w8(32'h3bd33435),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1e8f),
	.w1(32'h3b168b14),
	.w2(32'h3ada99f4),
	.w3(32'hba220a3f),
	.w4(32'h3b5b09e5),
	.w5(32'hb9cca54a),
	.w6(32'h3b58eb96),
	.w7(32'h3973e737),
	.w8(32'h39cae16e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8cda8),
	.w1(32'hbb21d08a),
	.w2(32'hbb13e2e0),
	.w3(32'hbba2c828),
	.w4(32'h3967c6dc),
	.w5(32'h3b25a61b),
	.w6(32'hbb6da702),
	.w7(32'hb94b9e64),
	.w8(32'h3b19e444),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f7622),
	.w1(32'h3a5027f4),
	.w2(32'h3ba0c7e3),
	.w3(32'hba8da1bc),
	.w4(32'h39de49fd),
	.w5(32'hb9d1352f),
	.w6(32'h39b09d13),
	.w7(32'h3af5b704),
	.w8(32'hb9d025ac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b230acc),
	.w1(32'hbb11a691),
	.w2(32'h3ab71f8c),
	.w3(32'h3a21527b),
	.w4(32'h3aa9174e),
	.w5(32'hb9f3da58),
	.w6(32'h3b5cd452),
	.w7(32'h3b5d19ca),
	.w8(32'h3a454844),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c07e7),
	.w1(32'h3a1d6c54),
	.w2(32'hba39a6b2),
	.w3(32'hbaca085c),
	.w4(32'hbb3a07bb),
	.w5(32'hbb317525),
	.w6(32'hbab0b26a),
	.w7(32'hbb039073),
	.w8(32'h3aaf65af),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e26e3),
	.w1(32'hbb47f901),
	.w2(32'hbb156d52),
	.w3(32'hbb7a828b),
	.w4(32'hbbb2a377),
	.w5(32'hbbe4678b),
	.w6(32'hb9794428),
	.w7(32'h3b6ba902),
	.w8(32'hbc0312fb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff4ea0),
	.w1(32'h3b173885),
	.w2(32'hbb21385c),
	.w3(32'h3b7ba633),
	.w4(32'hbaa1eb6f),
	.w5(32'hbb737c4d),
	.w6(32'h3bf8961a),
	.w7(32'hbab040e0),
	.w8(32'hbbc247f7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb43f),
	.w1(32'hb97f3ec7),
	.w2(32'h3c0ea6c9),
	.w3(32'hbad36abe),
	.w4(32'h3b1fec93),
	.w5(32'h3bb00950),
	.w6(32'h39dd5440),
	.w7(32'h3bde0151),
	.w8(32'h3bd33459),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfda2b),
	.w1(32'h3b443297),
	.w2(32'hbb6ef69c),
	.w3(32'h3bc7fcd8),
	.w4(32'hba669d0c),
	.w5(32'h3a6ad130),
	.w6(32'h3af5b871),
	.w7(32'hbbe74ddc),
	.w8(32'hbaa3eec0),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2da5d),
	.w1(32'hbbd79ae9),
	.w2(32'h39da32d4),
	.w3(32'hbb6b06c7),
	.w4(32'hbabbbc40),
	.w5(32'hba8f7e7b),
	.w6(32'hbb002f09),
	.w7(32'h3ad73929),
	.w8(32'h39b03df7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ba73e),
	.w1(32'hbb7ca5fc),
	.w2(32'hbbca0f01),
	.w3(32'hbba4dbbb),
	.w4(32'hbb9af016),
	.w5(32'hbaf59c7b),
	.w6(32'hbbb3acae),
	.w7(32'hbb641b01),
	.w8(32'hbaed26c6),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa89024),
	.w1(32'h3b8626fd),
	.w2(32'h3b9b9120),
	.w3(32'h3ae2d9b2),
	.w4(32'h3b4a4a87),
	.w5(32'hba99abd0),
	.w6(32'h3bb855ae),
	.w7(32'h3aabd53c),
	.w8(32'hbaaeca02),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81e7f4a),
	.w1(32'h3b0b6fc6),
	.w2(32'h3b204dc2),
	.w3(32'hbb288b3f),
	.w4(32'h3a92a1ac),
	.w5(32'h3a9bce4c),
	.w6(32'hba39f1e5),
	.w7(32'hbb1ac368),
	.w8(32'h3b146324),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402376),
	.w1(32'hbaa76244),
	.w2(32'hb9eb736c),
	.w3(32'hbb735348),
	.w4(32'h3b6a369a),
	.w5(32'h3c0b243c),
	.w6(32'hbb2c2076),
	.w7(32'h3b1a2e7d),
	.w8(32'h3b9c7257),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9339dd),
	.w1(32'h3a3483a4),
	.w2(32'hba616f6d),
	.w3(32'hbb513407),
	.w4(32'hb9a0300c),
	.w5(32'h3bacc131),
	.w6(32'hbc2a4e5c),
	.w7(32'h3a274e06),
	.w8(32'h3b99dee1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d65671),
	.w1(32'h3a22c433),
	.w2(32'h3a91181a),
	.w3(32'h39827f37),
	.w4(32'h3a976b00),
	.w5(32'h3b85e7b2),
	.w6(32'hba170dcd),
	.w7(32'h3b33a2a5),
	.w8(32'h3b8cc66b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9249fe9),
	.w1(32'hba5ca228),
	.w2(32'h3ab70054),
	.w3(32'h3af8e81f),
	.w4(32'h3b1b7496),
	.w5(32'hbb321006),
	.w6(32'h3ae48daf),
	.w7(32'h3ad448c7),
	.w8(32'hbba5bc8a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25693e),
	.w1(32'hbad3d204),
	.w2(32'h3acf7b58),
	.w3(32'hbb089df4),
	.w4(32'h39a41a38),
	.w5(32'h3bc78111),
	.w6(32'hba94baea),
	.w7(32'hba4d2866),
	.w8(32'h3bc90f1c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f7bb1),
	.w1(32'h39b5df4b),
	.w2(32'hbada3cfe),
	.w3(32'h3ad209bc),
	.w4(32'hbaa59554),
	.w5(32'hbaf5c5c4),
	.w6(32'h3b31cd77),
	.w7(32'hba1c3389),
	.w8(32'h39bf51d6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf6a70),
	.w1(32'hbb95dc37),
	.w2(32'hba8ae088),
	.w3(32'hbb48bfff),
	.w4(32'h3adcecdf),
	.w5(32'hba893ed2),
	.w6(32'hbb2fd635),
	.w7(32'h3805a86d),
	.w8(32'hb8519594),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee2b7f),
	.w1(32'hb9b89fd0),
	.w2(32'h3a0358cd),
	.w3(32'hbb493419),
	.w4(32'hba4376c4),
	.w5(32'h3b2dd327),
	.w6(32'hba4313c0),
	.w7(32'h39f80a5d),
	.w8(32'hb96eb03a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fd7d1),
	.w1(32'h3a9bc488),
	.w2(32'hbb7f20b9),
	.w3(32'hbaed02f7),
	.w4(32'h3a8e29de),
	.w5(32'h3a7df3de),
	.w6(32'h38c1e579),
	.w7(32'h3a229e77),
	.w8(32'h3b1d7bd5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992d51c),
	.w1(32'hbb4b4995),
	.w2(32'h39d01205),
	.w3(32'hba807e21),
	.w4(32'hbaa2956a),
	.w5(32'hb9af98da),
	.w6(32'hba2e53ef),
	.w7(32'h39a7ee54),
	.w8(32'hba53c53e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24ad4d),
	.w1(32'h399bf4c9),
	.w2(32'h3a94a511),
	.w3(32'hbb40322f),
	.w4(32'hbb02792e),
	.w5(32'hbb1e354d),
	.w6(32'hba0861ce),
	.w7(32'hb9f1f193),
	.w8(32'hbb4824b5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e42861),
	.w1(32'hbb2cc84d),
	.w2(32'h3a6bc822),
	.w3(32'hbab02dc7),
	.w4(32'hbb04a2da),
	.w5(32'h3bb68f43),
	.w6(32'h3aa99f59),
	.w7(32'hba4d87a5),
	.w8(32'h3bbf9cc1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64e340),
	.w1(32'h3b37e866),
	.w2(32'h39c7a39a),
	.w3(32'h3b4baa2d),
	.w4(32'h3bb9aaf0),
	.w5(32'h3aba63b7),
	.w6(32'h3ac99195),
	.w7(32'h3b0564d6),
	.w8(32'h3b50c60d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99a3fd),
	.w1(32'hbb910903),
	.w2(32'hba19c35e),
	.w3(32'hbb1d8dc5),
	.w4(32'hbb15bc8a),
	.w5(32'h3b6bc581),
	.w6(32'h3adfba62),
	.w7(32'hba190109),
	.w8(32'h3b9dbb98),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85f7ee),
	.w1(32'h3b2fc8a1),
	.w2(32'h3a7e0f11),
	.w3(32'h3b09a4c5),
	.w4(32'h383f1669),
	.w5(32'h3be1d68f),
	.w6(32'h3b9b5aa3),
	.w7(32'h3ab25297),
	.w8(32'h3be94ce7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79aab6),
	.w1(32'h3a6f65e6),
	.w2(32'h39efc9af),
	.w3(32'hbb75fd41),
	.w4(32'h3b57ab43),
	.w5(32'h3b4faf51),
	.w6(32'hbbe28bf7),
	.w7(32'h3baab0af),
	.w8(32'h3b2d3c9b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de6bb),
	.w1(32'h3a454743),
	.w2(32'h3bcc7842),
	.w3(32'h3ae95642),
	.w4(32'h3b8c167f),
	.w5(32'h3b9ad8f0),
	.w6(32'h3b375fa5),
	.w7(32'h3b8a5d82),
	.w8(32'hbadaf143),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4194d),
	.w1(32'hbb3d882d),
	.w2(32'h3b3a13aa),
	.w3(32'hbbb7662a),
	.w4(32'hbbb35646),
	.w5(32'hb9d59ab3),
	.w6(32'hbbd89abc),
	.w7(32'h398fdfd7),
	.w8(32'hb91628f1),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bc9cf),
	.w1(32'hba75fcc2),
	.w2(32'hb7b63626),
	.w3(32'hbac66d55),
	.w4(32'hbaaf0d83),
	.w5(32'hb8df9f54),
	.w6(32'hb9e1b85e),
	.w7(32'h3a9a79e2),
	.w8(32'h393b4e0f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8e80d),
	.w1(32'h39d0bb68),
	.w2(32'h3a329631),
	.w3(32'h3ac24570),
	.w4(32'hb88aaef2),
	.w5(32'h3b25a474),
	.w6(32'h3b996c4a),
	.w7(32'h3a8ec5f9),
	.w8(32'h3b0d6e08),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66dc11),
	.w1(32'h3addadcb),
	.w2(32'h3c0a6093),
	.w3(32'h3b077757),
	.w4(32'hba77889c),
	.w5(32'hba1f800c),
	.w6(32'h3c14bc23),
	.w7(32'h3b8254be),
	.w8(32'hbb42914f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab453c),
	.w1(32'hbb4a8f0e),
	.w2(32'hbaeffc7f),
	.w3(32'hbb40d3ea),
	.w4(32'hbb2d3547),
	.w5(32'h3a9e6bf6),
	.w6(32'hbb9ae993),
	.w7(32'hba3c4480),
	.w8(32'h390564b9),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198acf),
	.w1(32'hbb6fa7e3),
	.w2(32'hbb78d343),
	.w3(32'hbaa9bb20),
	.w4(32'hbb0102bb),
	.w5(32'hbb2adb03),
	.w6(32'hbaa38b93),
	.w7(32'h3a2ceee1),
	.w8(32'hbb213d82),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35720),
	.w1(32'hbb0deb15),
	.w2(32'h3b3f1064),
	.w3(32'hbba23ed1),
	.w4(32'hba8ab168),
	.w5(32'hba69772a),
	.w6(32'hbbb0afe8),
	.w7(32'h3ad7c6b7),
	.w8(32'hba3b4655),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139f65),
	.w1(32'h3a3b7152),
	.w2(32'hba0fe5e8),
	.w3(32'hbacc8ae0),
	.w4(32'hb95f482f),
	.w5(32'h38b94782),
	.w6(32'h3b4fe012),
	.w7(32'hbad25a67),
	.w8(32'hba018dca),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb675054),
	.w1(32'h3a361df2),
	.w2(32'h3ae8e48f),
	.w3(32'hbb62554e),
	.w4(32'hbae5a527),
	.w5(32'h3acfe915),
	.w6(32'hbb32c4b2),
	.w7(32'hbb1bd933),
	.w8(32'h3b8532c3),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabda824),
	.w1(32'hba9ebb60),
	.w2(32'hbaf97469),
	.w3(32'h38c602b4),
	.w4(32'h3a0519f0),
	.w5(32'hbace295a),
	.w6(32'h3ae7049b),
	.w7(32'h3b3710a4),
	.w8(32'hbb32a9ee),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de9bd),
	.w1(32'hbb386e6c),
	.w2(32'hbbe96f79),
	.w3(32'hbb179bc6),
	.w4(32'h3b0d7a02),
	.w5(32'hbb5af200),
	.w6(32'hbb62acc3),
	.w7(32'hba9f83ae),
	.w8(32'hbbb8b8bd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69f65),
	.w1(32'hbb50c6a5),
	.w2(32'h3adecd00),
	.w3(32'hbaf2af35),
	.w4(32'h3b251012),
	.w5(32'hbb3b5610),
	.w6(32'h3ae5d234),
	.w7(32'h3bc0276d),
	.w8(32'h383bbd8c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995e03e),
	.w1(32'h3ab2674d),
	.w2(32'h3b223502),
	.w3(32'hbb18fbc9),
	.w4(32'hbb07cda8),
	.w5(32'hba56d0a8),
	.w6(32'h3a8f6815),
	.w7(32'h3ad70c4d),
	.w8(32'hbb8fe625),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf27855),
	.w1(32'hba7f092e),
	.w2(32'h3ae69e47),
	.w3(32'h3ad81d2f),
	.w4(32'h3a0b4525),
	.w5(32'hbaf41252),
	.w6(32'h3b4e2df9),
	.w7(32'hba55fbe3),
	.w8(32'hbb429bf4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3f5b5),
	.w1(32'h3ab82d00),
	.w2(32'h3b6f7c6d),
	.w3(32'h3af227e3),
	.w4(32'h3b9c2477),
	.w5(32'h3aa4797e),
	.w6(32'h3ab7a78d),
	.w7(32'h3b4b86f4),
	.w8(32'h3a02edef),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9394631),
	.w1(32'h39555ffd),
	.w2(32'hbb21d2de),
	.w3(32'h3a93ca5a),
	.w4(32'h3b44b341),
	.w5(32'h3a89fefb),
	.w6(32'h39948466),
	.w7(32'hb92c830c),
	.w8(32'h3adfa3db),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a774971),
	.w1(32'h392887da),
	.w2(32'hbaa38dc6),
	.w3(32'hb85f1b0b),
	.w4(32'hba90e6db),
	.w5(32'hb6e0789f),
	.w6(32'hbb1afd08),
	.w7(32'hbb158141),
	.w8(32'h37c0d134),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0683),
	.w1(32'h3aacebe8),
	.w2(32'h3a820472),
	.w3(32'h3ada63b9),
	.w4(32'h3b4e1e03),
	.w5(32'hbaa1e407),
	.w6(32'hb8873e7b),
	.w7(32'h3ae9e96c),
	.w8(32'hbb8ac1a4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750343),
	.w1(32'hbace2031),
	.w2(32'h3b62b13d),
	.w3(32'hbb7acdba),
	.w4(32'hbb0c5369),
	.w5(32'h3bc44f99),
	.w6(32'hbb647999),
	.w7(32'h3b9a70bf),
	.w8(32'h3c2b5078),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a6cd0),
	.w1(32'h3aee33c0),
	.w2(32'hbb705aa0),
	.w3(32'h3b77dccf),
	.w4(32'h39dead9d),
	.w5(32'h3ac61adb),
	.w6(32'h3bb2231b),
	.w7(32'hbb824e14),
	.w8(32'h3943f943),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce5a77),
	.w1(32'h3b205539),
	.w2(32'h3b90289e),
	.w3(32'h3b030cb3),
	.w4(32'h3b246822),
	.w5(32'hba741437),
	.w6(32'h3af91a6b),
	.w7(32'h3b528c2c),
	.w8(32'hb9bf6471),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39864bd4),
	.w1(32'h3aa81ecf),
	.w2(32'hba76f4c3),
	.w3(32'h3a17ea84),
	.w4(32'h3b9e9716),
	.w5(32'hbb270397),
	.w6(32'h3b31d67a),
	.w7(32'h3ad344ce),
	.w8(32'hbb6048cc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf1e00),
	.w1(32'hbbf6cb0d),
	.w2(32'hbbaf0c93),
	.w3(32'hbbc0f324),
	.w4(32'hbbced43b),
	.w5(32'h3b26bb30),
	.w6(32'hbb8a5ff6),
	.w7(32'hbadaaf79),
	.w8(32'h3b8161a8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a40fc),
	.w1(32'h3a8a2313),
	.w2(32'h3b112069),
	.w3(32'hba0030b3),
	.w4(32'h3ba44b53),
	.w5(32'h3b645e7b),
	.w6(32'h3b0c23c6),
	.w7(32'h3bf4a22b),
	.w8(32'h3b540374),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b279a50),
	.w1(32'h3ac9dc36),
	.w2(32'h3b97ae2c),
	.w3(32'h3a483f03),
	.w4(32'h3b6361cb),
	.w5(32'hba64f1e1),
	.w6(32'hbb54e676),
	.w7(32'h3b7489c2),
	.w8(32'h3ac916ed),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4665ed),
	.w1(32'hbb05be8d),
	.w2(32'h3a4b997a),
	.w3(32'hbb0227e3),
	.w4(32'h3aad624a),
	.w5(32'h3b9eafd4),
	.w6(32'hba8eacf6),
	.w7(32'hbb5c529b),
	.w8(32'h3b10efdf),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba488523),
	.w1(32'h3a93e349),
	.w2(32'h3b52c05c),
	.w3(32'h3a97cd03),
	.w4(32'h3a302b39),
	.w5(32'h3b0a1f15),
	.w6(32'h3b20ef86),
	.w7(32'h3bacef1b),
	.w8(32'h3aa7f7bb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55d6e8),
	.w1(32'h3b0f803e),
	.w2(32'h3b711687),
	.w3(32'h3a74b01e),
	.w4(32'h389e6e60),
	.w5(32'h3aa73397),
	.w6(32'h3aa5d255),
	.w7(32'h3b7b2aed),
	.w8(32'hb9254604),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d8f14),
	.w1(32'hbb843495),
	.w2(32'h3ad7ce2b),
	.w3(32'hbb21d214),
	.w4(32'hbb86aafd),
	.w5(32'h3b081590),
	.w6(32'h3b91b80b),
	.w7(32'h3b6575ee),
	.w8(32'h3bfc1049),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc7337),
	.w1(32'hbb83d403),
	.w2(32'h3b3e9cfa),
	.w3(32'hbbae52f2),
	.w4(32'hbb6ffb57),
	.w5(32'h3b855a06),
	.w6(32'h3b64114d),
	.w7(32'h3b0495c7),
	.w8(32'h3aaab9f4),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0364f2),
	.w1(32'hbc0f5e2b),
	.w2(32'hbae1f63c),
	.w3(32'hbc1414fa),
	.w4(32'hbbb5620f),
	.w5(32'hbacb5aaf),
	.w6(32'hbc1516ef),
	.w7(32'h3a0a2086),
	.w8(32'h3b495561),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32aa9b),
	.w1(32'hbb321878),
	.w2(32'h39594d94),
	.w3(32'hbb309d49),
	.w4(32'hbb5f7415),
	.w5(32'h3a5a5469),
	.w6(32'hbaaf7e54),
	.w7(32'hbb6c9d40),
	.w8(32'h3956484c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc7fd5),
	.w1(32'h39acdefe),
	.w2(32'hb94c78fb),
	.w3(32'h3ae9d2ae),
	.w4(32'h3ac39919),
	.w5(32'hbb3f47b3),
	.w6(32'h3aa3bbb8),
	.w7(32'hba7524f1),
	.w8(32'hbbc9e376),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd97578),
	.w1(32'h3aeb566e),
	.w2(32'hba525134),
	.w3(32'h3b54e3ae),
	.w4(32'h3b1e7317),
	.w5(32'hbaa27845),
	.w6(32'h3bd5f9b3),
	.w7(32'h3afea17e),
	.w8(32'hbb18ae8c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f7b35),
	.w1(32'h3a1e4447),
	.w2(32'h3a3b904b),
	.w3(32'hbab66971),
	.w4(32'hba9e10b3),
	.w5(32'hba0f39df),
	.w6(32'h3aada82b),
	.w7(32'hbb1707ee),
	.w8(32'h392d8783),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8696e4),
	.w1(32'h3a8032ce),
	.w2(32'h3b5a1f9c),
	.w3(32'hbaaf635c),
	.w4(32'h394da962),
	.w5(32'h3ac48998),
	.w6(32'hbabf9ac3),
	.w7(32'h3af11772),
	.w8(32'h3b0241ea),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa56d4b),
	.w1(32'hbb0fd7b2),
	.w2(32'hbba1dd82),
	.w3(32'hbb1e20cb),
	.w4(32'h393e2c22),
	.w5(32'h3aba8eba),
	.w6(32'hbb156233),
	.w7(32'hbb219ab8),
	.w8(32'hba97523f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3dcf),
	.w1(32'hbb654833),
	.w2(32'hba64261b),
	.w3(32'hbaaca2cf),
	.w4(32'hb8185f69),
	.w5(32'h3a26e6d6),
	.w6(32'hbbc33bfc),
	.w7(32'hbaf1df54),
	.w8(32'h3abe8f10),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79e773c),
	.w1(32'hbad4ef9f),
	.w2(32'h3b3c5365),
	.w3(32'hbaa70eb7),
	.w4(32'h3a2c9e09),
	.w5(32'h3829b0fe),
	.w6(32'hb8afb64f),
	.w7(32'h3b8916ca),
	.w8(32'h3aface9c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aea91),
	.w1(32'hbb57e58e),
	.w2(32'hba2c808a),
	.w3(32'hbaf48b60),
	.w4(32'hbacb78e0),
	.w5(32'hbb47eba5),
	.w6(32'hba86f975),
	.w7(32'hbb4020a2),
	.w8(32'hbb97494e),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c3d7c),
	.w1(32'hbb019b3b),
	.w2(32'hbb587f74),
	.w3(32'hbb91fdbc),
	.w4(32'hbb5f51ca),
	.w5(32'hbadb39b4),
	.w6(32'hbb7b771c),
	.w7(32'hbb8c6996),
	.w8(32'hbb8ca4f5),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ce659),
	.w1(32'hbbcd2bc1),
	.w2(32'hbb7651df),
	.w3(32'hbbcf947c),
	.w4(32'hbbc8e56e),
	.w5(32'h3bb107e9),
	.w6(32'hbb37df3b),
	.w7(32'hba849363),
	.w8(32'h3bfe8b9c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4a505),
	.w1(32'hbacbeae9),
	.w2(32'hbb28170b),
	.w3(32'hbb448234),
	.w4(32'hbb8ab2e0),
	.w5(32'h3a43a178),
	.w6(32'hbaba8dd9),
	.w7(32'hbb0ab878),
	.w8(32'hba3a5f51),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51efc4),
	.w1(32'hbaf1be07),
	.w2(32'hbba2c2c4),
	.w3(32'h3af0dc7f),
	.w4(32'h3b8eaab1),
	.w5(32'h3b22c453),
	.w6(32'hb9e88f5b),
	.w7(32'h3ad7f5f3),
	.w8(32'h3b7f701a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c8f84),
	.w1(32'hbb3e480f),
	.w2(32'h396506a0),
	.w3(32'hbb7b02e0),
	.w4(32'hba053dc0),
	.w5(32'h3bf31262),
	.w6(32'hbb7cc2fb),
	.w7(32'hbb3a6e96),
	.w8(32'h3bbf107e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c1c1d),
	.w1(32'hbb791d68),
	.w2(32'h3aa1893e),
	.w3(32'hba73ca74),
	.w4(32'h39fd4e8d),
	.w5(32'h3b62ce14),
	.w6(32'hbb71c668),
	.w7(32'hba755cde),
	.w8(32'h3aec9884),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b287fa5),
	.w1(32'hba8ac25d),
	.w2(32'h3ba4a513),
	.w3(32'h36461510),
	.w4(32'h3b49d1b0),
	.w5(32'h3b7deb01),
	.w6(32'hbba0d4a0),
	.w7(32'h3a12228f),
	.w8(32'h39389de3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8637ae),
	.w1(32'hbb190370),
	.w2(32'h3b2d855c),
	.w3(32'h3a47be43),
	.w4(32'h3b8305ca),
	.w5(32'h3bd09e60),
	.w6(32'hbb852bb5),
	.w7(32'h3ab9a042),
	.w8(32'h3b12f232),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad78cf),
	.w1(32'h3b8d3803),
	.w2(32'h3b9beed8),
	.w3(32'h3b866e2d),
	.w4(32'h3c0329cb),
	.w5(32'h3a9917a8),
	.w6(32'hbbc7f574),
	.w7(32'h3adc7660),
	.w8(32'h3907c720),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a376ac),
	.w1(32'h39103008),
	.w2(32'hb9584c1d),
	.w3(32'h3b83e572),
	.w4(32'hb9a32deb),
	.w5(32'h3a777887),
	.w6(32'h39a56f49),
	.w7(32'hbb2c7e00),
	.w8(32'hba32f05f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5586f0),
	.w1(32'hbb077d15),
	.w2(32'hbaffc170),
	.w3(32'hbb2ea88b),
	.w4(32'h3a3b5cf4),
	.w5(32'h3c2c7752),
	.w6(32'h39ee0561),
	.w7(32'hba993a1b),
	.w8(32'h3c34c290),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b9e02),
	.w1(32'hba8dc3c5),
	.w2(32'hb9bcde4b),
	.w3(32'h3a1f552f),
	.w4(32'hba5c3a81),
	.w5(32'h3aea689f),
	.w6(32'h3a4dac60),
	.w7(32'h3971207c),
	.w8(32'h3b84d25c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4970b),
	.w1(32'h3a05fd7d),
	.w2(32'h3b6da81a),
	.w3(32'hbb80b772),
	.w4(32'hbafe1af5),
	.w5(32'h3b8a6eb0),
	.w6(32'h378697f2),
	.w7(32'h3a5d9c93),
	.w8(32'h3b20c54b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba152702),
	.w1(32'hbac0c453),
	.w2(32'hba8f9703),
	.w3(32'h3abd4d06),
	.w4(32'hbaef037c),
	.w5(32'h3a7d320f),
	.w6(32'hba0568f5),
	.w7(32'hbac26119),
	.w8(32'hbb052d31),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39928b9a),
	.w1(32'hbb2d6324),
	.w2(32'hbb631fdd),
	.w3(32'hbb062172),
	.w4(32'hbac169ff),
	.w5(32'h3add6dba),
	.w6(32'hb8be2082),
	.w7(32'hbb84c242),
	.w8(32'h3b75a628),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86f718),
	.w1(32'h3b8adcc4),
	.w2(32'hb908178a),
	.w3(32'h3b412a4b),
	.w4(32'h39dda7de),
	.w5(32'hbb9b915f),
	.w6(32'h3bc2f24b),
	.w7(32'hba28b920),
	.w8(32'hbb0029ad),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb677392),
	.w1(32'hbb81c6da),
	.w2(32'hbb78c7f6),
	.w3(32'hbaee9d32),
	.w4(32'hba54224b),
	.w5(32'h3b2dc76b),
	.w6(32'hba6241d6),
	.w7(32'hb8a9e6a6),
	.w8(32'h3a6152bb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01f1fa),
	.w1(32'hbb934f16),
	.w2(32'hb9ba3d4c),
	.w3(32'hbab8f8fc),
	.w4(32'h3b5a9439),
	.w5(32'h3b6c741b),
	.w6(32'hba734213),
	.w7(32'h3b387c66),
	.w8(32'h3b762340),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10e8a5),
	.w1(32'hbb8d7419),
	.w2(32'hba939766),
	.w3(32'hbb1c7ee3),
	.w4(32'hb9ba7ae0),
	.w5(32'hba35fade),
	.w6(32'hbbada541),
	.w7(32'hba01b7fd),
	.w8(32'hbb3b76b7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b728ed),
	.w1(32'hbab3c7dc),
	.w2(32'h3acd6e7c),
	.w3(32'hbab26934),
	.w4(32'h3ba84d18),
	.w5(32'h3c88e417),
	.w6(32'h3a61b0cb),
	.w7(32'h3bac8abd),
	.w8(32'h3c974782),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8de5a7),
	.w1(32'hbb2cff5a),
	.w2(32'hbb29f444),
	.w3(32'hbb8b4700),
	.w4(32'hbb69d236),
	.w5(32'h3c055c4b),
	.w6(32'hba3f2eef),
	.w7(32'hbb5ccfc0),
	.w8(32'h3b0c3748),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26afe8),
	.w1(32'hbbc66c87),
	.w2(32'hbbb3bd4c),
	.w3(32'hb9efdd7c),
	.w4(32'hbb79d9d0),
	.w5(32'h3b4bd8f5),
	.w6(32'hbb7c2707),
	.w7(32'hbb8d7c82),
	.w8(32'h3bc993ba),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc5a2),
	.w1(32'hbb123dc8),
	.w2(32'hb7b042eb),
	.w3(32'hbb02d998),
	.w4(32'h3897583e),
	.w5(32'h3b93b889),
	.w6(32'hbbac6547),
	.w7(32'h3af2c4de),
	.w8(32'h3b3ca5a3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd9345),
	.w1(32'hba006dca),
	.w2(32'hbb281b41),
	.w3(32'h37e7cfcb),
	.w4(32'h391f9092),
	.w5(32'hba7eb782),
	.w6(32'hbabf78d2),
	.w7(32'hbb3ddf03),
	.w8(32'hbb45f139),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bccf9),
	.w1(32'hba55f262),
	.w2(32'h3aab0077),
	.w3(32'hbb0f4a54),
	.w4(32'h3b753ec3),
	.w5(32'h3bde3a3b),
	.w6(32'h39db9913),
	.w7(32'h3b72bbdd),
	.w8(32'h3be7a8fb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab82cd7),
	.w1(32'hba990151),
	.w2(32'hba5cf9c5),
	.w3(32'hbb2ed136),
	.w4(32'hba4b802a),
	.w5(32'h3a352731),
	.w6(32'hbc1c52b8),
	.w7(32'hbba7729b),
	.w8(32'h3aab0ced),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0edae1),
	.w1(32'hb8fcf239),
	.w2(32'h3a8ba0d4),
	.w3(32'hbb41de0b),
	.w4(32'hbb7eacd3),
	.w5(32'h3b893f67),
	.w6(32'h3afbbea3),
	.w7(32'h39d5a0ec),
	.w8(32'h3b0858f0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule