module layer_10_featuremap_233(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb26685),
	.w1(32'h3b34e8d3),
	.w2(32'hbb7515bb),
	.w3(32'h3be43c65),
	.w4(32'h39a22f50),
	.w5(32'h3a30b7f0),
	.w6(32'hbbf1d33f),
	.w7(32'h3af954f6),
	.w8(32'h39c1d0aa),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0eb279),
	.w1(32'hbc91c354),
	.w2(32'hbc1702ef),
	.w3(32'hbbd02c0f),
	.w4(32'hbbb14848),
	.w5(32'hbb44f071),
	.w6(32'h39a03db1),
	.w7(32'hbc33b193),
	.w8(32'hbba6a796),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaefa1),
	.w1(32'h3b2ef6f9),
	.w2(32'hbbaf2394),
	.w3(32'hbaf28317),
	.w4(32'hb9e02626),
	.w5(32'hbb2d2318),
	.w6(32'hbcedbd3b),
	.w7(32'hbb9c3007),
	.w8(32'h3b030318),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb472078),
	.w1(32'h3b12dfa1),
	.w2(32'hbab37bad),
	.w3(32'h3c247a2b),
	.w4(32'hbc6457c7),
	.w5(32'hbba52809),
	.w6(32'hbb52e8bc),
	.w7(32'h3bc4c6f3),
	.w8(32'hbbc53ee3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa573e1),
	.w1(32'hbb6ad95f),
	.w2(32'hb9d6cde7),
	.w3(32'h3a109d60),
	.w4(32'hbaff4692),
	.w5(32'h39d7dc2d),
	.w6(32'h3bace948),
	.w7(32'h3bdd2559),
	.w8(32'h3c06a95f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58bdc4),
	.w1(32'h3b7cba05),
	.w2(32'h3b08bd30),
	.w3(32'h3ab53e7a),
	.w4(32'h3b8aff0c),
	.w5(32'hbb3c1c33),
	.w6(32'h3c88e533),
	.w7(32'h38843985),
	.w8(32'hbba9eb28),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b977abf),
	.w1(32'hbb803271),
	.w2(32'hbc2868ac),
	.w3(32'h3bf8fa24),
	.w4(32'hbc8f0d87),
	.w5(32'h3c1b0503),
	.w6(32'hba957abc),
	.w7(32'h3c6cde66),
	.w8(32'hbc68d5d2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5be502),
	.w1(32'hbc574f32),
	.w2(32'hbc35beaf),
	.w3(32'h3ba24fef),
	.w4(32'hbbe43f11),
	.w5(32'hbb1503bb),
	.w6(32'hbbda06c2),
	.w7(32'hbb8a0c70),
	.w8(32'hbc1a8a7e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e0c8),
	.w1(32'hbbac4a94),
	.w2(32'h3b46f242),
	.w3(32'hba3f4daa),
	.w4(32'hba03bbf5),
	.w5(32'h3b77afd7),
	.w6(32'hba5a0496),
	.w7(32'hbb2aa588),
	.w8(32'h3b2029c7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0598d),
	.w1(32'hba886a49),
	.w2(32'hbac127d8),
	.w3(32'h3b7e5fde),
	.w4(32'hbb98b7a8),
	.w5(32'hbc136456),
	.w6(32'hbbf71c10),
	.w7(32'hbc988ede),
	.w8(32'hbbd78337),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb09b4),
	.w1(32'hbbea576c),
	.w2(32'hbb7d378b),
	.w3(32'hbb3f85b0),
	.w4(32'hbbd561f0),
	.w5(32'h3c8ccf2c),
	.w6(32'h3bed1c3f),
	.w7(32'hbb06837a),
	.w8(32'hb9f9172f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61d2c0),
	.w1(32'h3b15fc68),
	.w2(32'h3c9617e2),
	.w3(32'h3c85aa74),
	.w4(32'h3ca4adae),
	.w5(32'hbb97ddec),
	.w6(32'h3c3aac94),
	.w7(32'h3bb3fc52),
	.w8(32'h37915740),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b296602),
	.w1(32'hbbf07b4f),
	.w2(32'hbc53d3a5),
	.w3(32'h3b77e0a1),
	.w4(32'h3a8d9111),
	.w5(32'hbbd15f10),
	.w6(32'h3ad123ee),
	.w7(32'h3996411c),
	.w8(32'hbc21eee3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c547b27),
	.w1(32'h3bcfb8a8),
	.w2(32'h3ab0004a),
	.w3(32'h3b8fb489),
	.w4(32'hbd12b4ce),
	.w5(32'hbba775e6),
	.w6(32'h3c451ddd),
	.w7(32'hbb955bcf),
	.w8(32'hbb002819),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c2a61),
	.w1(32'hbbdda5b9),
	.w2(32'h395c8448),
	.w3(32'hbc0d16e8),
	.w4(32'h3bc237cb),
	.w5(32'hba9489de),
	.w6(32'hbbd4ceed),
	.w7(32'hbc31999b),
	.w8(32'h3b6ff4f3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc299691),
	.w1(32'hbb16e663),
	.w2(32'hbc4bfce5),
	.w3(32'hbc435e2d),
	.w4(32'hbc2fcddf),
	.w5(32'hbbaec8a9),
	.w6(32'hbc684b49),
	.w7(32'hbc3a9146),
	.w8(32'h3bef4a13),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab23436),
	.w1(32'hbc21a29b),
	.w2(32'hbb9e06e4),
	.w3(32'h3a407cca),
	.w4(32'h389284c6),
	.w5(32'h3a9d1c70),
	.w6(32'hba9bfef2),
	.w7(32'hbb6fac72),
	.w8(32'hbb87cb54),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205410),
	.w1(32'hbcbde834),
	.w2(32'hbc100bb4),
	.w3(32'hb9bf82f0),
	.w4(32'h38bb52b0),
	.w5(32'hbbb43a1b),
	.w6(32'hb985dcf8),
	.w7(32'h3d1a2091),
	.w8(32'hbbf0eced),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01a30),
	.w1(32'h3bd73d97),
	.w2(32'hbaa4ecd9),
	.w3(32'hbaab3e6f),
	.w4(32'hbac33ae4),
	.w5(32'h3b9ea231),
	.w6(32'hbb4d40b9),
	.w7(32'hbac207e0),
	.w8(32'hbb269b23),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae504b0),
	.w1(32'h3b924120),
	.w2(32'hbb86f772),
	.w3(32'hb8d422db),
	.w4(32'hbd1a9d9e),
	.w5(32'h3b4e1d9e),
	.w6(32'h3b5c3f7c),
	.w7(32'h3a973692),
	.w8(32'h3c144619),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ca64d),
	.w1(32'h3ba4867e),
	.w2(32'hbd0d7777),
	.w3(32'hbb97f530),
	.w4(32'hb9aec931),
	.w5(32'h3ae2f578),
	.w6(32'h3b6adb58),
	.w7(32'hbbdf3195),
	.w8(32'h3be53a89),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c8d96),
	.w1(32'h3b0c9393),
	.w2(32'h3b9d8538),
	.w3(32'h39215e74),
	.w4(32'hbb5bf315),
	.w5(32'hbae13eda),
	.w6(32'h3b86e9fc),
	.w7(32'h3a212dff),
	.w8(32'hbb5dd8cb),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0020e),
	.w1(32'h3b201fd3),
	.w2(32'h3c836c5f),
	.w3(32'hbb6fc013),
	.w4(32'hbace0a61),
	.w5(32'h3b6efd1e),
	.w6(32'hbbcef330),
	.w7(32'hbab5fc07),
	.w8(32'h3cd01846),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd64312),
	.w1(32'hbb881dba),
	.w2(32'hbbec534b),
	.w3(32'hbb8e0326),
	.w4(32'h3ad5116d),
	.w5(32'h3a623ebb),
	.w6(32'hbbbfb793),
	.w7(32'hbc9c1de0),
	.w8(32'hbc39edd7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42570e),
	.w1(32'h3a30d440),
	.w2(32'h3c1477a3),
	.w3(32'hbbfb0e50),
	.w4(32'h3cd921ae),
	.w5(32'hbb205d32),
	.w6(32'hbb18097c),
	.w7(32'hbbc510af),
	.w8(32'hbc5628c5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2321c),
	.w1(32'hb9eccd7e),
	.w2(32'h3b979988),
	.w3(32'hbb374962),
	.w4(32'h3c1189b6),
	.w5(32'h3b825048),
	.w6(32'hbc01384e),
	.w7(32'hbb13a8c9),
	.w8(32'h3a8d760d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3cde6),
	.w1(32'hbc221a4b),
	.w2(32'h3c171348),
	.w3(32'hbb6ccf2f),
	.w4(32'hb9bae864),
	.w5(32'hb972e7b5),
	.w6(32'hbac5bd7f),
	.w7(32'h3bb5a7b7),
	.w8(32'h3bedef1b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7f8a3),
	.w1(32'hbb054abb),
	.w2(32'hbc470574),
	.w3(32'hbc5b4275),
	.w4(32'h3cadd9c2),
	.w5(32'hbc4277fd),
	.w6(32'hba3384eb),
	.w7(32'hbbad9cd9),
	.w8(32'hbc1e20da),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0869a),
	.w1(32'hbb844fb0),
	.w2(32'hbb9a6204),
	.w3(32'hbb35fd24),
	.w4(32'hbbe317f8),
	.w5(32'h3b2689b1),
	.w6(32'h3c2fa8fe),
	.w7(32'hb9176060),
	.w8(32'hbb0ea543),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc6c3),
	.w1(32'h3c269fac),
	.w2(32'h3c7461d7),
	.w3(32'h3c182a9b),
	.w4(32'hbc1d6b34),
	.w5(32'hbbc34cab),
	.w6(32'hbba14bea),
	.w7(32'h3b64e7b9),
	.w8(32'hbbc0c8b0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45493e),
	.w1(32'h3bb31d61),
	.w2(32'h3a0524cd),
	.w3(32'h3c02c496),
	.w4(32'h3b8bea9e),
	.w5(32'h3b93c378),
	.w6(32'hbaae23d0),
	.w7(32'h3b6bbf8b),
	.w8(32'h3ca7af6b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9107469),
	.w1(32'hbbbef1a0),
	.w2(32'h3ca0b5b7),
	.w3(32'h3990204e),
	.w4(32'h3cf778da),
	.w5(32'hbaff3883),
	.w6(32'h3c8cfcf8),
	.w7(32'h3bbe51ff),
	.w8(32'hbbc077d3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8b73b),
	.w1(32'hbc108fa3),
	.w2(32'hbcc3a4db),
	.w3(32'h3b678b45),
	.w4(32'h3af132ce),
	.w5(32'hb8e5095e),
	.w6(32'h3bb8b055),
	.w7(32'h3bd0b1a9),
	.w8(32'h3c0999bf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a423c),
	.w1(32'hbb23de75),
	.w2(32'hbc06e072),
	.w3(32'hbc4f2d09),
	.w4(32'h3b2f97d8),
	.w5(32'h3bb30dbb),
	.w6(32'hbbc6e115),
	.w7(32'hbc1524bf),
	.w8(32'hbb9ab2bd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b5091),
	.w1(32'h3bbe7e29),
	.w2(32'h3cc7ad22),
	.w3(32'h3c326edf),
	.w4(32'hbb87c9c2),
	.w5(32'h3d0c5406),
	.w6(32'hbcfe6482),
	.w7(32'hbc8dbbc1),
	.w8(32'hbbabcc21),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf45c5),
	.w1(32'hbc527b58),
	.w2(32'hbcb363a8),
	.w3(32'h3c9811d7),
	.w4(32'h3c50ebfe),
	.w5(32'h3c045567),
	.w6(32'hbc435ce8),
	.w7(32'h3a1548c8),
	.w8(32'hbbadb11d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd138f6e),
	.w1(32'hbcae90ec),
	.w2(32'h3bfd97ee),
	.w3(32'hbc99723e),
	.w4(32'h3b1211f5),
	.w5(32'h3b25101c),
	.w6(32'hbc70f6a0),
	.w7(32'h3c168b72),
	.w8(32'h3c9d7a5f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa0598),
	.w1(32'h3bb9bf14),
	.w2(32'h3bc5323d),
	.w3(32'h3bbb3df4),
	.w4(32'h3bd7d636),
	.w5(32'h3aaac32b),
	.w6(32'h3ad52880),
	.w7(32'hbc1ee5ea),
	.w8(32'hb926ce47),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b584d9f),
	.w1(32'h3cef162c),
	.w2(32'hbc2c0aca),
	.w3(32'h3c8edc9d),
	.w4(32'hbcab3255),
	.w5(32'h3bbbf43c),
	.w6(32'h3ba76d56),
	.w7(32'h3cbdf861),
	.w8(32'h3b6544cd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb90840),
	.w1(32'h3c6f53bb),
	.w2(32'hba76b78e),
	.w3(32'h3bb2f4b8),
	.w4(32'h3b4613d7),
	.w5(32'h3bf60177),
	.w6(32'hbb49a7ee),
	.w7(32'hbc47b8bb),
	.w8(32'h3be5836c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38481f02),
	.w1(32'hbd03062e),
	.w2(32'h3b1623f0),
	.w3(32'h3874aa43),
	.w4(32'h3b490bbc),
	.w5(32'hba9257b9),
	.w6(32'hba0b6212),
	.w7(32'hb996d276),
	.w8(32'h3bacfadc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1208ec),
	.w1(32'hbb06b82c),
	.w2(32'h3c62ceca),
	.w3(32'hbca683a6),
	.w4(32'h3a336d04),
	.w5(32'h3b88c7c0),
	.w6(32'h3a88cc8d),
	.w7(32'hbc11953a),
	.w8(32'h3925b151),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4adfa5),
	.w1(32'h3c194a54),
	.w2(32'hbbe97bcd),
	.w3(32'hbc00f3a1),
	.w4(32'h3bd2d600),
	.w5(32'h3c4520cb),
	.w6(32'h3b5d0c09),
	.w7(32'h3c27b9a2),
	.w8(32'h3b67339a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e64e8),
	.w1(32'h3ba16790),
	.w2(32'hbba9cee9),
	.w3(32'hbbee8b1f),
	.w4(32'hbbe846fa),
	.w5(32'h3be0ca27),
	.w6(32'hbc49614f),
	.w7(32'hbc604481),
	.w8(32'h39d3deef),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc425c5d),
	.w1(32'h3c077e1f),
	.w2(32'h3b9cf912),
	.w3(32'hbbb74581),
	.w4(32'hbc33aee5),
	.w5(32'hbb23de5b),
	.w6(32'hbbb010c9),
	.w7(32'hbc1b8a58),
	.w8(32'hbb14fa06),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74ef26),
	.w1(32'h3a864c29),
	.w2(32'hbc9de473),
	.w3(32'hba874491),
	.w4(32'hbcbdf502),
	.w5(32'h3a699655),
	.w6(32'hbc2dc479),
	.w7(32'hbb88dc76),
	.w8(32'hbc831174),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b88c5),
	.w1(32'h3abea2b4),
	.w2(32'h3b86346b),
	.w3(32'hbb8689d3),
	.w4(32'hbb54f566),
	.w5(32'hb91d9a2d),
	.w6(32'hbb06282b),
	.w7(32'hba570888),
	.w8(32'hbbbba5a6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c0ee),
	.w1(32'h3bf2a705),
	.w2(32'hb7947e54),
	.w3(32'h3c7355cc),
	.w4(32'h3c169d21),
	.w5(32'hbb8220d5),
	.w6(32'h3b4c821b),
	.w7(32'hbba47b22),
	.w8(32'hbb01f8d3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c3322),
	.w1(32'h3b8e3e3e),
	.w2(32'h3b63a476),
	.w3(32'hba8c3a4a),
	.w4(32'hbbd2ad85),
	.w5(32'h39e344f1),
	.w6(32'h3a10ec90),
	.w7(32'h3c4ed6c9),
	.w8(32'h3b95e14b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5995),
	.w1(32'h3bddcae1),
	.w2(32'h3c4b425f),
	.w3(32'hbb9988c9),
	.w4(32'h3bc25574),
	.w5(32'hbbe80063),
	.w6(32'hbc8370e0),
	.w7(32'h3b807811),
	.w8(32'h3bc8f475),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905531b),
	.w1(32'h39f77d63),
	.w2(32'h3a26954c),
	.w3(32'h3b05fee3),
	.w4(32'hbbb16a54),
	.w5(32'hb931fd74),
	.w6(32'hbb3a250a),
	.w7(32'hbb78b1af),
	.w8(32'h3b8d9723),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce00942),
	.w1(32'hbc110599),
	.w2(32'h3c2b810d),
	.w3(32'hbc8d37fa),
	.w4(32'hbbdc842e),
	.w5(32'hbc81f49a),
	.w6(32'hbc1fd197),
	.w7(32'h38dd6d82),
	.w8(32'h3b98606a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0357e2),
	.w1(32'hbb112211),
	.w2(32'h3b8f9f9a),
	.w3(32'hbb5bf21c),
	.w4(32'h3bc5dfb9),
	.w5(32'h3a98ed99),
	.w6(32'hbaf47cd4),
	.w7(32'hbb10fbfc),
	.w8(32'h3b5ec3fc),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91fabb),
	.w1(32'h3a75bc8e),
	.w2(32'h398b2aa6),
	.w3(32'hbb06dc89),
	.w4(32'h3b1c119e),
	.w5(32'hbcabe0d4),
	.w6(32'h3b8b9e9e),
	.w7(32'h3bce1ff8),
	.w8(32'h3ba95f0a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a966955),
	.w1(32'h3c20aeb2),
	.w2(32'h3c2870ba),
	.w3(32'hbbc21718),
	.w4(32'hbcc41b30),
	.w5(32'hbb52e0c0),
	.w6(32'h3b80d0b2),
	.w7(32'hb9f14fb3),
	.w8(32'h3c46be5e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb50a9),
	.w1(32'h39c97a1c),
	.w2(32'hbb400e1a),
	.w3(32'hbb997ac7),
	.w4(32'h3c8d4a85),
	.w5(32'h3bd6a6f9),
	.w6(32'h3900ecca),
	.w7(32'hbc7c70ec),
	.w8(32'hbb7b7e1f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc76f9f),
	.w1(32'h3b43b4d5),
	.w2(32'hbc417e18),
	.w3(32'hbc94dab7),
	.w4(32'hbc00ebb6),
	.w5(32'h3ca08259),
	.w6(32'h3b1ca3f9),
	.w7(32'h3a2f982d),
	.w8(32'hbb92a3c5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11baeb),
	.w1(32'h3c79e8ff),
	.w2(32'hbc8da113),
	.w3(32'hbb35073f),
	.w4(32'h3ac0eb69),
	.w5(32'h3bb153b0),
	.w6(32'hb9f79dae),
	.w7(32'h3cb8940b),
	.w8(32'h3960debc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb877c3f),
	.w1(32'hbc59c4de),
	.w2(32'hb88186ba),
	.w3(32'h3c9e0b06),
	.w4(32'h3c38687f),
	.w5(32'hbc4bdc1d),
	.w6(32'h3c23e96d),
	.w7(32'hbbf2728e),
	.w8(32'h3c4fa26d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab2e67),
	.w1(32'hbbff8ea3),
	.w2(32'h3be1d5c1),
	.w3(32'hbaceb6f5),
	.w4(32'hbb0db1b4),
	.w5(32'hbc455cef),
	.w6(32'hbbf12875),
	.w7(32'h3b525042),
	.w8(32'h3b00c341),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23fd9c),
	.w1(32'hba7bd210),
	.w2(32'hbb5db07f),
	.w3(32'hbbab260b),
	.w4(32'h3c1d4105),
	.w5(32'hbaefa83b),
	.w6(32'hbc836e9c),
	.w7(32'h39c350e8),
	.w8(32'h3bfbea3a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92bdc3),
	.w1(32'h3b24c0d8),
	.w2(32'hba2e3d1d),
	.w3(32'h3a92b621),
	.w4(32'hbbef3ba1),
	.w5(32'hb9aff83b),
	.w6(32'h39967e0d),
	.w7(32'hbc2d2fca),
	.w8(32'h3ba9b208),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc8367),
	.w1(32'h3acfe2d2),
	.w2(32'h3c3d6182),
	.w3(32'h3b84058d),
	.w4(32'hbc070e17),
	.w5(32'hbba32363),
	.w6(32'hbbc339d7),
	.w7(32'hbbe67529),
	.w8(32'hbb29e586),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d38e1),
	.w1(32'hbb516317),
	.w2(32'h3c064bc9),
	.w3(32'hba2106b5),
	.w4(32'h3a842d3f),
	.w5(32'h3bf68d38),
	.w6(32'h3aa33de9),
	.w7(32'hbb01d86e),
	.w8(32'h3c29431e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26143f),
	.w1(32'h3b0db69d),
	.w2(32'h3afd574f),
	.w3(32'h3bc9ebc4),
	.w4(32'h3c4e06c7),
	.w5(32'h3c0482c6),
	.w6(32'h3ccf0cda),
	.w7(32'hba78e731),
	.w8(32'hbc4a3b91),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7d33),
	.w1(32'hbb959498),
	.w2(32'hbbb0e069),
	.w3(32'hbbc0e519),
	.w4(32'hbb384d8b),
	.w5(32'h3a05c8c5),
	.w6(32'h3ba92997),
	.w7(32'h3a2dfac3),
	.w8(32'hbb9787db),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19fba0),
	.w1(32'hbba264f2),
	.w2(32'hbbd16afb),
	.w3(32'h3ab8cbfd),
	.w4(32'hbc20c50c),
	.w5(32'hbb27c9c8),
	.w6(32'h3bbaec0a),
	.w7(32'h3ccf6813),
	.w8(32'hbc9193f2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbee58),
	.w1(32'h3c1eabfe),
	.w2(32'hbbe54f26),
	.w3(32'hbc35587f),
	.w4(32'hbc2919a1),
	.w5(32'hb94a92d2),
	.w6(32'hbbfb8c9d),
	.w7(32'hbc5bb90e),
	.w8(32'hbb49c63f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a895fc2),
	.w1(32'h3bbe3ae4),
	.w2(32'hbbe3560f),
	.w3(32'hbb7d4f3a),
	.w4(32'hbb59f09d),
	.w5(32'h3a321457),
	.w6(32'h3bc9fbe6),
	.w7(32'hbbba086e),
	.w8(32'h3c472ec0),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce6a56),
	.w1(32'hbbb8ed12),
	.w2(32'h3cb18fd0),
	.w3(32'hbc801d39),
	.w4(32'hbc869fd1),
	.w5(32'hbb6ff653),
	.w6(32'hbc2bc396),
	.w7(32'hbce793aa),
	.w8(32'hbb125f74),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f54a5),
	.w1(32'hb9578e69),
	.w2(32'hb9faad2a),
	.w3(32'hbbdeeb08),
	.w4(32'h3b0c2971),
	.w5(32'h3832caaf),
	.w6(32'h3b3341f8),
	.w7(32'h3d1a9cb1),
	.w8(32'hbc0a6a62),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c82c1ac),
	.w1(32'h3a8ca97f),
	.w2(32'h3b8ecede),
	.w3(32'hbb3e6ded),
	.w4(32'hbabbb0eb),
	.w5(32'hbad4824b),
	.w6(32'hbc38e571),
	.w7(32'hbc3af2d9),
	.w8(32'hbc58ff4f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc5f15),
	.w1(32'hbc48ea27),
	.w2(32'h3af828fd),
	.w3(32'hbcae65b6),
	.w4(32'h3af62950),
	.w5(32'h399ce0d3),
	.w6(32'hbc0400b0),
	.w7(32'hbc269570),
	.w8(32'hbc2fd7c9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc22963),
	.w1(32'hb8a0527e),
	.w2(32'h3b878dab),
	.w3(32'hbc1b7888),
	.w4(32'hbadf83da),
	.w5(32'h3c8bec84),
	.w6(32'h3c358ea4),
	.w7(32'h3c92d45e),
	.w8(32'hbacdbf55),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac7cfd),
	.w1(32'hbc817017),
	.w2(32'h35df8a6f),
	.w3(32'h3b3d2786),
	.w4(32'hbb4612d5),
	.w5(32'hbb0b5f73),
	.w6(32'hbba711be),
	.w7(32'hbb419988),
	.w8(32'hba936be4),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d5f4),
	.w1(32'hbc92bfa1),
	.w2(32'h39124ec8),
	.w3(32'hba5f8515),
	.w4(32'h3c22fecc),
	.w5(32'hba046424),
	.w6(32'h3bf6c7e9),
	.w7(32'h3b9f3ceb),
	.w8(32'hbba387ff),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba715f4a),
	.w1(32'hbc33d4dd),
	.w2(32'hbbdaf54c),
	.w3(32'hbbbf05fb),
	.w4(32'hbb597c33),
	.w5(32'h3a71c13d),
	.w6(32'hbba4de08),
	.w7(32'h3c2b6c6f),
	.w8(32'hba558bf6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c836272),
	.w1(32'hbb58ad04),
	.w2(32'h3d080958),
	.w3(32'h3bdf56f5),
	.w4(32'hbaf9d519),
	.w5(32'h3b85a2c9),
	.w6(32'hbc1a03d2),
	.w7(32'hbb355e4a),
	.w8(32'hbb640b16),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9249c9),
	.w1(32'h3a8009a5),
	.w2(32'hbc3ee09c),
	.w3(32'hbc586846),
	.w4(32'hbb380202),
	.w5(32'hbc832aba),
	.w6(32'h3c7bb5b4),
	.w7(32'hbc0cb30d),
	.w8(32'hbc65d4bb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa71c6c),
	.w1(32'hbc115522),
	.w2(32'hbae76fe3),
	.w3(32'h3b7620a1),
	.w4(32'h392b4763),
	.w5(32'h3bb3efc7),
	.w6(32'h3b30b8d3),
	.w7(32'h3b81ed11),
	.w8(32'hbb51087f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba9da5),
	.w1(32'hbbd3315a),
	.w2(32'hba9ff88e),
	.w3(32'hbc7fef75),
	.w4(32'hbc15c496),
	.w5(32'hbc262495),
	.w6(32'hbbb299a3),
	.w7(32'h3c5f1b0d),
	.w8(32'hbc4cd630),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4679),
	.w1(32'hbc43fc25),
	.w2(32'hbc20177a),
	.w3(32'h3cd0944e),
	.w4(32'hbb9fce5e),
	.w5(32'hbc109ca9),
	.w6(32'hb9d19b9a),
	.w7(32'h3ad881fa),
	.w8(32'h3c0e5f17),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14f005),
	.w1(32'hbb5203fa),
	.w2(32'h3c83f665),
	.w3(32'hb980e0e7),
	.w4(32'h3b28aa90),
	.w5(32'hbbb505dd),
	.w6(32'hbbec5469),
	.w7(32'hbbcc6cfc),
	.w8(32'hbcb954d1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6bee3),
	.w1(32'hbba76141),
	.w2(32'hbb1b52ce),
	.w3(32'h3b77513f),
	.w4(32'hbad93852),
	.w5(32'h3b4d0182),
	.w6(32'hbbdbb939),
	.w7(32'hba399dc4),
	.w8(32'h3c0a4153),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eb278),
	.w1(32'h3b961198),
	.w2(32'hbaaeb61e),
	.w3(32'hbb91e3a4),
	.w4(32'h3b0cc514),
	.w5(32'h3c09d8af),
	.w6(32'h3c481ff5),
	.w7(32'hbc9b041f),
	.w8(32'h3beb6483),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8bca),
	.w1(32'h3bba844a),
	.w2(32'hbbd7ce7c),
	.w3(32'hbba8de5e),
	.w4(32'h3b897a6b),
	.w5(32'h3c0896a5),
	.w6(32'hbbe2cf76),
	.w7(32'h3b8745de),
	.w8(32'h3c633d43),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9878e),
	.w1(32'hbc354243),
	.w2(32'hbb91b4fc),
	.w3(32'hbc38081f),
	.w4(32'hbc2e7548),
	.w5(32'h3ba8248d),
	.w6(32'hbb8e2d78),
	.w7(32'h3bd2d9e6),
	.w8(32'hbb842bc1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea89c),
	.w1(32'h3be3f5ed),
	.w2(32'hbabd3702),
	.w3(32'hba2df0b3),
	.w4(32'hba4dbc85),
	.w5(32'h3c58bb46),
	.w6(32'hbba26289),
	.w7(32'hbc25000f),
	.w8(32'hbb9fffe4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c848fe3),
	.w1(32'hbc91608a),
	.w2(32'hbbb3fa60),
	.w3(32'h3bd8c938),
	.w4(32'h3c03e988),
	.w5(32'h393d8ddd),
	.w6(32'hbb03fa58),
	.w7(32'hbc541f0b),
	.w8(32'hbbf9ad6d),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5a53),
	.w1(32'h3b8732c0),
	.w2(32'h3b8f2625),
	.w3(32'h396076d7),
	.w4(32'h3bc63a99),
	.w5(32'hbacc8f85),
	.w6(32'h3d32c1e0),
	.w7(32'hbbd0b6de),
	.w8(32'hba203807),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a4cfb),
	.w1(32'h3c41a667),
	.w2(32'hba369c0f),
	.w3(32'h3b3dad9f),
	.w4(32'h3b93d648),
	.w5(32'h3b1b7f4f),
	.w6(32'h3aaadb52),
	.w7(32'h3c67c748),
	.w8(32'h3c8631dc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad18eb4),
	.w1(32'hbbb024bb),
	.w2(32'hbd4b80dd),
	.w3(32'h3cff1642),
	.w4(32'hbc4785e5),
	.w5(32'hbc031778),
	.w6(32'hb971d1b4),
	.w7(32'h3c50512a),
	.w8(32'h3b0d1563),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7561df),
	.w1(32'h3c69ec68),
	.w2(32'h3c481de8),
	.w3(32'hbbe4db7f),
	.w4(32'hbadc61f5),
	.w5(32'h3aec6ca5),
	.w6(32'h3aedce7f),
	.w7(32'hba86aff1),
	.w8(32'hbc80507a),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad03b),
	.w1(32'hb91a9511),
	.w2(32'hbc5b2629),
	.w3(32'hbc1f21d1),
	.w4(32'hbbedb251),
	.w5(32'hbd1eea47),
	.w6(32'hbc804cf8),
	.w7(32'hbc03fc5e),
	.w8(32'hbc48d5b5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba64c96),
	.w1(32'hbc2ba952),
	.w2(32'hba1f2d52),
	.w3(32'h3b3fc039),
	.w4(32'hbbc2c9c7),
	.w5(32'h3b64c227),
	.w6(32'hbb78525f),
	.w7(32'h3be5ae6b),
	.w8(32'h3bd2da9b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc857d2e),
	.w1(32'hbc016060),
	.w2(32'hbb567772),
	.w3(32'hbc159b1c),
	.w4(32'h3a976a50),
	.w5(32'h3c25a14c),
	.w6(32'h3bcf2294),
	.w7(32'h39a5d6d1),
	.w8(32'h3b45b7ea),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ffc43),
	.w1(32'h3b340e57),
	.w2(32'h3bbf4d00),
	.w3(32'hbc10cb79),
	.w4(32'h3bb66199),
	.w5(32'h3bf90b81),
	.w6(32'hbbe61bd7),
	.w7(32'h3b374aec),
	.w8(32'hb9c70e54),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc100),
	.w1(32'hbc70165c),
	.w2(32'h39a4a3ff),
	.w3(32'hbba62252),
	.w4(32'hba93920f),
	.w5(32'h3a5b9c6c),
	.w6(32'hbc121c55),
	.w7(32'hbbc43c2f),
	.w8(32'hba6893d9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f4889),
	.w1(32'hbbbfaaa9),
	.w2(32'hbb364b29),
	.w3(32'h3ba7f628),
	.w4(32'h3b2f6851),
	.w5(32'h3bfbd751),
	.w6(32'h3c0e4988),
	.w7(32'hbc401553),
	.w8(32'h39fab802),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b666ddc),
	.w1(32'h3b9572a6),
	.w2(32'hbbc35ad2),
	.w3(32'hbbf4ef7d),
	.w4(32'h3bf0dd05),
	.w5(32'hbad7c8e4),
	.w6(32'hb909bcc4),
	.w7(32'h3b1a61de),
	.w8(32'h3b277895),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb962626),
	.w1(32'hba115c8b),
	.w2(32'h3be6145b),
	.w3(32'hbbd023d7),
	.w4(32'hbb6910bf),
	.w5(32'h3bbdcd7f),
	.w6(32'h38a69c74),
	.w7(32'h3bc8cc2c),
	.w8(32'h3c8cb6c0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60920e),
	.w1(32'hb9928db2),
	.w2(32'h3a7936c0),
	.w3(32'hbbb4d8b8),
	.w4(32'hbc26e312),
	.w5(32'h3b1d24d8),
	.w6(32'hbc09caba),
	.w7(32'hbbefaea7),
	.w8(32'hbb372aef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7038ba),
	.w1(32'h3c45e9a3),
	.w2(32'hbc15d165),
	.w3(32'hbb576395),
	.w4(32'hbbbf7968),
	.w5(32'hb9d09245),
	.w6(32'hbc09b1a7),
	.w7(32'hbc4dab08),
	.w8(32'h3bd7f2db),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e6df4),
	.w1(32'hbb0ba97a),
	.w2(32'h3605cc86),
	.w3(32'hb9ff9b04),
	.w4(32'hbbb54881),
	.w5(32'hba103849),
	.w6(32'h39c281fe),
	.w7(32'h3b8a8ac5),
	.w8(32'h3be3927c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29e831),
	.w1(32'hbc9b9a6e),
	.w2(32'hbbcd971f),
	.w3(32'h38c1f517),
	.w4(32'hbc6bfce5),
	.w5(32'h3a50d8b6),
	.w6(32'hbc12bd04),
	.w7(32'hbb52f09c),
	.w8(32'h3b964832),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a766b),
	.w1(32'h3c6b9baf),
	.w2(32'hbbe7ecba),
	.w3(32'h3c01b6c9),
	.w4(32'h3b778c5d),
	.w5(32'h3a0dbfbd),
	.w6(32'h3c408f4f),
	.w7(32'hbb9f2dcf),
	.w8(32'hbb5d5f94),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b887e),
	.w1(32'h3c81ed95),
	.w2(32'h3bb31ee8),
	.w3(32'h3977d2d4),
	.w4(32'hbac82cd3),
	.w5(32'hba2893a0),
	.w6(32'h3c155e9e),
	.w7(32'hbae2a8da),
	.w8(32'hb9c8c10d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbe7a6),
	.w1(32'hba575dca),
	.w2(32'hbb141537),
	.w3(32'h3aaaa703),
	.w4(32'hbbae253e),
	.w5(32'hbb3754da),
	.w6(32'hbbc5d557),
	.w7(32'hbb59b36c),
	.w8(32'hbc1a5e61),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a732580),
	.w1(32'h3c118f4d),
	.w2(32'h3cd1e3fb),
	.w3(32'hbc07563a),
	.w4(32'h3bf50461),
	.w5(32'h3b2d72d7),
	.w6(32'h3bea5bd8),
	.w7(32'h3b3185fe),
	.w8(32'hb95cdc81),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83639),
	.w1(32'h3b55a3ec),
	.w2(32'hbae7cd82),
	.w3(32'h3a8fb5df),
	.w4(32'h3bab4c77),
	.w5(32'h3c81ece1),
	.w6(32'hbc1bf31f),
	.w7(32'h3be6e4de),
	.w8(32'hbc17f300),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985c5c4),
	.w1(32'h3b47dd0a),
	.w2(32'h3c90e5d1),
	.w3(32'hbaa0eb1c),
	.w4(32'hbb4ca7c1),
	.w5(32'hbbdef037),
	.w6(32'hbae904ef),
	.w7(32'h3b8bb15f),
	.w8(32'h3c534c87),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8626db),
	.w1(32'h3d083e02),
	.w2(32'h3bb1d4c8),
	.w3(32'hb9ee0038),
	.w4(32'hbc63dac9),
	.w5(32'h39c10e54),
	.w6(32'hbc058b75),
	.w7(32'h3c54dddc),
	.w8(32'hbc129407),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a11c5),
	.w1(32'hbc8522f7),
	.w2(32'h3c16a958),
	.w3(32'h3b179416),
	.w4(32'h3a56787a),
	.w5(32'hbc322b58),
	.w6(32'hbc21e1cb),
	.w7(32'hbc21a1be),
	.w8(32'hbc4616c4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b032d),
	.w1(32'hbc8c27bf),
	.w2(32'h3cab837b),
	.w3(32'hbbaf39b2),
	.w4(32'hbc5cbe70),
	.w5(32'hbc31ee65),
	.w6(32'hbbd8bd93),
	.w7(32'hbc7bef2d),
	.w8(32'hbc0ea2ed),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace903),
	.w1(32'hbcb49fb3),
	.w2(32'hbb79cfe7),
	.w3(32'hbb56d95a),
	.w4(32'hbb11f637),
	.w5(32'hbc096822),
	.w6(32'h3ccb7fc1),
	.w7(32'hbc0e499f),
	.w8(32'h3c8d6f44),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ad715),
	.w1(32'hbc82465b),
	.w2(32'hbadccc69),
	.w3(32'h3a7a0f02),
	.w4(32'h3bc33ffe),
	.w5(32'hbc45919b),
	.w6(32'h3c8a70d1),
	.w7(32'hbcaebd96),
	.w8(32'hb932d096),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c72e2),
	.w1(32'h3bd37b1a),
	.w2(32'h3bb2f3f3),
	.w3(32'h3aa3bbf3),
	.w4(32'hbcc4cebf),
	.w5(32'hbc89fc3e),
	.w6(32'hba8add9c),
	.w7(32'hbc11133f),
	.w8(32'hbabf48dd),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa1fb4),
	.w1(32'hbbed515c),
	.w2(32'hbcddecdf),
	.w3(32'h3c575d43),
	.w4(32'hbc332470),
	.w5(32'hbcbda243),
	.w6(32'h3cb74c63),
	.w7(32'h3b17c997),
	.w8(32'h3bbac90d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2e438),
	.w1(32'h3ae6eef5),
	.w2(32'h3b8f3f87),
	.w3(32'hbb317fd1),
	.w4(32'hbc264b86),
	.w5(32'hbb893e16),
	.w6(32'hbb86f344),
	.w7(32'h3b52f466),
	.w8(32'hbbe75e76),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c1ec),
	.w1(32'hbc1c09db),
	.w2(32'hbc050e07),
	.w3(32'h3b86889c),
	.w4(32'hbb595016),
	.w5(32'hbb150b21),
	.w6(32'hbb6227fc),
	.w7(32'h3a645368),
	.w8(32'h3c6c0298),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3475cc),
	.w1(32'h3bcf9a5d),
	.w2(32'h3b190349),
	.w3(32'h3a3578c0),
	.w4(32'hbcb4c371),
	.w5(32'hbce3760d),
	.w6(32'h3c01f108),
	.w7(32'hbbaa2c8f),
	.w8(32'h3b44c733),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d7a61),
	.w1(32'h3d0bc2c8),
	.w2(32'hbc4cad4b),
	.w3(32'h3c9de324),
	.w4(32'h3bdee367),
	.w5(32'hbb223e5e),
	.w6(32'h3c5c676f),
	.w7(32'h3bd3009f),
	.w8(32'hbc1ff56a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62bc2d),
	.w1(32'hbc435721),
	.w2(32'hba1c9604),
	.w3(32'hbb560162),
	.w4(32'hbc3c0968),
	.w5(32'h3b30907d),
	.w6(32'hbd260a36),
	.w7(32'hbcb41b3b),
	.w8(32'h3ce57a30),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbe49),
	.w1(32'hbbcc4522),
	.w2(32'hbd5b0e39),
	.w3(32'hb93338a6),
	.w4(32'h3c503eda),
	.w5(32'h3d32d46a),
	.w6(32'h3b0a2851),
	.w7(32'hbb6e3c77),
	.w8(32'hbd2cc723),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd254de),
	.w1(32'hbc39c004),
	.w2(32'hbc579779),
	.w3(32'hbc1a8e46),
	.w4(32'hbc7d8a5f),
	.w5(32'hbb9e6034),
	.w6(32'hbc0a971b),
	.w7(32'hbbc6dece),
	.w8(32'h3d0b2fb0),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc165f),
	.w1(32'h37b04beb),
	.w2(32'h3c870196),
	.w3(32'hbc31c61f),
	.w4(32'hbc82d3cb),
	.w5(32'hbbd62628),
	.w6(32'hbc558e4e),
	.w7(32'h3a314b7d),
	.w8(32'hbb4cfbbc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb91210),
	.w1(32'h3a3e8533),
	.w2(32'hbbe28d61),
	.w3(32'hbc053e03),
	.w4(32'h3c0c1cd8),
	.w5(32'hba9990f5),
	.w6(32'hbc8d416e),
	.w7(32'h3c65e5ec),
	.w8(32'hb83ae396),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39357c3d),
	.w1(32'hbb555635),
	.w2(32'hbada8fca),
	.w3(32'h3c9f21ad),
	.w4(32'hba3f7d2c),
	.w5(32'h3b808496),
	.w6(32'hbc64fb87),
	.w7(32'h3b4f98e2),
	.w8(32'hbc9fdd0d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbc320),
	.w1(32'hbcbb1632),
	.w2(32'hbc1fd017),
	.w3(32'hbc292a73),
	.w4(32'h3b0e2836),
	.w5(32'hbbb35eb9),
	.w6(32'hbc098e7e),
	.w7(32'h3c489e49),
	.w8(32'h3c36ebc1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59988d),
	.w1(32'hbc0fa53a),
	.w2(32'h3b8f98d7),
	.w3(32'hbc434224),
	.w4(32'hba5977bf),
	.w5(32'hbbb3608a),
	.w6(32'hbbf2a57d),
	.w7(32'h3bdde113),
	.w8(32'h3c8414ee),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadafe1e),
	.w1(32'hbbd4191e),
	.w2(32'hbc68138e),
	.w3(32'hbc127490),
	.w4(32'hbcc4b8af),
	.w5(32'hbc19c6b8),
	.w6(32'h3a2f6051),
	.w7(32'hbc34b399),
	.w8(32'hbc5595ee),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14f26a),
	.w1(32'hbc6336ad),
	.w2(32'hbb94d406),
	.w3(32'hbba8aaee),
	.w4(32'hbbcd5ae4),
	.w5(32'h3aeebc51),
	.w6(32'hbb62fcf8),
	.w7(32'h3a460cce),
	.w8(32'h3c19b6dc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c423a),
	.w1(32'h3bbbc4d6),
	.w2(32'hbc6c5636),
	.w3(32'hbb2e8ca0),
	.w4(32'h3a9d717a),
	.w5(32'hbc0148eb),
	.w6(32'hbb20a848),
	.w7(32'h3a77a2ee),
	.w8(32'h3ba1c3db),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc820238),
	.w1(32'hbcbd7193),
	.w2(32'hbb8a576e),
	.w3(32'hbc506a2e),
	.w4(32'h3a61b127),
	.w5(32'h3c095caa),
	.w6(32'hbca2802d),
	.w7(32'hbbdb7b32),
	.w8(32'hbcb774d9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81a9ec),
	.w1(32'hbc1fd20f),
	.w2(32'hbc0a9867),
	.w3(32'hbb27bdf4),
	.w4(32'hba442628),
	.w5(32'hbc3519d9),
	.w6(32'hbc879b62),
	.w7(32'h3c719a7b),
	.w8(32'hbb093fae),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18762d),
	.w1(32'hb9bfa037),
	.w2(32'hbcae250c),
	.w3(32'h3c7216bb),
	.w4(32'hbc03c747),
	.w5(32'hb91f02ae),
	.w6(32'hbc0a9b29),
	.w7(32'hbbdeadbf),
	.w8(32'hbb95ad64),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e324b),
	.w1(32'h3b36f324),
	.w2(32'hbb9511ac),
	.w3(32'hba49ee81),
	.w4(32'hbc221e4e),
	.w5(32'h3af995eb),
	.w6(32'hbc207381),
	.w7(32'h3c7a5c7c),
	.w8(32'hb95ce70f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60d99b),
	.w1(32'h3bc94d40),
	.w2(32'h3ba2656f),
	.w3(32'hbbfdbe15),
	.w4(32'hbc5dc813),
	.w5(32'hbcaca961),
	.w6(32'hbbec4675),
	.w7(32'hbb0a7393),
	.w8(32'hbd0501e3),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc143310),
	.w1(32'hbc868e07),
	.w2(32'h38bc7225),
	.w3(32'h3c48a9c2),
	.w4(32'h3b3a56f0),
	.w5(32'hbb988483),
	.w6(32'h3af14bb2),
	.w7(32'hbc6f23a7),
	.w8(32'h3c0cbcf0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e12ab),
	.w1(32'hbc2ef4ae),
	.w2(32'hbbb3dafb),
	.w3(32'h3cd0fa79),
	.w4(32'h3c0bf7ef),
	.w5(32'h3c8c9d68),
	.w6(32'hbc1582bc),
	.w7(32'h3b4d5db1),
	.w8(32'hbbef0d44),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b8a54),
	.w1(32'h3c86a603),
	.w2(32'hbb53d41b),
	.w3(32'h3a45a741),
	.w4(32'h3bcb0e98),
	.w5(32'hbb3e41a8),
	.w6(32'hbca6670f),
	.w7(32'hbaf60490),
	.w8(32'hba8d7397),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef4250),
	.w1(32'hb9ab1239),
	.w2(32'h3b8f29c7),
	.w3(32'hbbc67145),
	.w4(32'h3b542b49),
	.w5(32'hbb11383b),
	.w6(32'h3be10f85),
	.w7(32'h39804497),
	.w8(32'h3a2f5999),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8efcc),
	.w1(32'h3b57c03e),
	.w2(32'hb9aafe3a),
	.w3(32'h39cf5667),
	.w4(32'h3b363afa),
	.w5(32'h3b9b8417),
	.w6(32'hbbe011dc),
	.w7(32'hbaf70ad4),
	.w8(32'h3b1fddf5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4f97e2),
	.w1(32'h3cc3e2b1),
	.w2(32'hbbae39bb),
	.w3(32'hbac33d20),
	.w4(32'hbb99bd6f),
	.w5(32'h3b0903d9),
	.w6(32'hbc07a33a),
	.w7(32'h3bf4ce98),
	.w8(32'hbc330b12),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba6765),
	.w1(32'hba8b4ce6),
	.w2(32'h3c5d5e64),
	.w3(32'hbbe11338),
	.w4(32'h3afa7e04),
	.w5(32'h3ad76c62),
	.w6(32'h39b12d00),
	.w7(32'hbc6adca7),
	.w8(32'h3cf192cb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ead38),
	.w1(32'hbb77298f),
	.w2(32'hbbf49348),
	.w3(32'hb9a1a468),
	.w4(32'hbae3b1f1),
	.w5(32'hba0a30db),
	.w6(32'h3c67d835),
	.w7(32'h3c02c4e7),
	.w8(32'h3b71e40a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3c42a),
	.w1(32'hba3ba9bc),
	.w2(32'h3b99135f),
	.w3(32'hbbf6bc53),
	.w4(32'hba3d3b24),
	.w5(32'hba0607db),
	.w6(32'h3a927e13),
	.w7(32'h3bf40e48),
	.w8(32'h3abf0c00),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90f1ef),
	.w1(32'hbc0056b6),
	.w2(32'h3a6215d0),
	.w3(32'h3b2fbfc0),
	.w4(32'hbb0e965b),
	.w5(32'h3bbd99be),
	.w6(32'hba28d62c),
	.w7(32'hbb0408b4),
	.w8(32'hbbc4967e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd10cad5),
	.w1(32'h3b348754),
	.w2(32'hbb393d2c),
	.w3(32'hbb7c2304),
	.w4(32'hbc9232dc),
	.w5(32'h3cc849e0),
	.w6(32'h395e6c07),
	.w7(32'h3bbb899b),
	.w8(32'h3ac9c575),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a1eeb),
	.w1(32'hbc1b24af),
	.w2(32'hb9b475da),
	.w3(32'hbc4b4d72),
	.w4(32'h394c1232),
	.w5(32'h3bd8f1d3),
	.w6(32'hbc30a801),
	.w7(32'h3abaabef),
	.w8(32'hb9cb5278),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ac07),
	.w1(32'hbb43d889),
	.w2(32'hbb8af3fb),
	.w3(32'hbb5f44ab),
	.w4(32'h3a96d017),
	.w5(32'hbb1519e3),
	.w6(32'hbc8aa892),
	.w7(32'h3b0937c6),
	.w8(32'hbc154056),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33bc1e),
	.w1(32'hbc2a43d7),
	.w2(32'hbbeb0519),
	.w3(32'h3b24468d),
	.w4(32'hbb40d9f5),
	.w5(32'h3a0c9f93),
	.w6(32'hbb04b9d8),
	.w7(32'h3aa1a78e),
	.w8(32'h3cbe0fbf),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14c86d),
	.w1(32'hbc055ccb),
	.w2(32'h3c365d88),
	.w3(32'hbc451975),
	.w4(32'h3aa7f36b),
	.w5(32'h3b97ba37),
	.w6(32'hbc36b730),
	.w7(32'h3aaab1db),
	.w8(32'hbc478082),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab906d8),
	.w1(32'hb99e60ed),
	.w2(32'hb9843189),
	.w3(32'h3c2badb0),
	.w4(32'hbb9ee9c8),
	.w5(32'hbb15315c),
	.w6(32'h3b79fdc7),
	.w7(32'hbba09ce1),
	.w8(32'hbb9fea72),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dcb86),
	.w1(32'hbafe1dc1),
	.w2(32'h3b9620ae),
	.w3(32'h3c1b7c96),
	.w4(32'hbcb6236b),
	.w5(32'hba3f70b9),
	.w6(32'h3b65ba9b),
	.w7(32'h3b56f785),
	.w8(32'h3ab557bb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a095e),
	.w1(32'h3c10d20c),
	.w2(32'h3bc6af47),
	.w3(32'hbbe1b39d),
	.w4(32'hbbc22f8a),
	.w5(32'hb9a063f5),
	.w6(32'h39bd021b),
	.w7(32'h3c009b3b),
	.w8(32'h3c864b3c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c67b4),
	.w1(32'h3bd66231),
	.w2(32'hbc16ccd4),
	.w3(32'hbb48eb22),
	.w4(32'h3d18cd1d),
	.w5(32'h3c5d6f40),
	.w6(32'hbbdee3f4),
	.w7(32'hbb236346),
	.w8(32'hbc572a03),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48be07),
	.w1(32'hbb99f295),
	.w2(32'hbb5c45af),
	.w3(32'h3a881354),
	.w4(32'hba774ff6),
	.w5(32'h3ab5deec),
	.w6(32'h3b071004),
	.w7(32'hbc0c15a1),
	.w8(32'h3b55081f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44325f),
	.w1(32'hbc177eff),
	.w2(32'hb962ec98),
	.w3(32'hbc0fc72f),
	.w4(32'hbc6ab069),
	.w5(32'h3b54bc40),
	.w6(32'hbb8806e8),
	.w7(32'hba11bf82),
	.w8(32'hbb2aed22),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11e8f1),
	.w1(32'hbbd6a6e7),
	.w2(32'hbbb8e89c),
	.w3(32'h3bf54bd6),
	.w4(32'h3b95d3f3),
	.w5(32'h3b421cc0),
	.w6(32'h3af8cd8e),
	.w7(32'h3b523fd7),
	.w8(32'h3972ba96),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6b380),
	.w1(32'hbb84cca9),
	.w2(32'hbb0ea165),
	.w3(32'h3b105fba),
	.w4(32'h3a1c3a02),
	.w5(32'h3c2f4d86),
	.w6(32'h3a457568),
	.w7(32'hbba8425d),
	.w8(32'hbb6965bf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898bf7),
	.w1(32'h3c23409a),
	.w2(32'h3b89cc4d),
	.w3(32'hbc13044a),
	.w4(32'h3bdf4586),
	.w5(32'h3bbb6258),
	.w6(32'h3b285fb0),
	.w7(32'h3be6154e),
	.w8(32'hbb996c18),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967b87),
	.w1(32'hbb2fbf49),
	.w2(32'h3be6e799),
	.w3(32'hbbee57d7),
	.w4(32'h3bcfcc40),
	.w5(32'h3be728bc),
	.w6(32'h3c4487c9),
	.w7(32'hbbb8c250),
	.w8(32'h3bf0485b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d28a631),
	.w1(32'h3a3f3299),
	.w2(32'hbb3b2435),
	.w3(32'hbb46812c),
	.w4(32'hbc43fc02),
	.w5(32'hba00c094),
	.w6(32'h3b5b0c67),
	.w7(32'h3c3d7aa6),
	.w8(32'hbbf2242b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1f192),
	.w1(32'hbbe6a274),
	.w2(32'hbc21ff54),
	.w3(32'h3a40dc7a),
	.w4(32'hbaca8a37),
	.w5(32'h3b0f07f9),
	.w6(32'hbb9275b1),
	.w7(32'hb879d46e),
	.w8(32'hbc222c8e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04748e),
	.w1(32'hbb7aeb8d),
	.w2(32'hbb61a3fe),
	.w3(32'h3b097541),
	.w4(32'hbb5a4f0f),
	.w5(32'hb9d691d9),
	.w6(32'hbbe5c67f),
	.w7(32'hbbafb82d),
	.w8(32'h3bcbf290),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6973e),
	.w1(32'hbb89ed40),
	.w2(32'hbbe5ad0a),
	.w3(32'hba90b39b),
	.w4(32'h3c11e20d),
	.w5(32'h3bc83588),
	.w6(32'h3c13e412),
	.w7(32'hba88f3e2),
	.w8(32'hbb329b54),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a109b2c),
	.w1(32'hbc627053),
	.w2(32'h3bf71fcf),
	.w3(32'hbc149924),
	.w4(32'hbb986d4f),
	.w5(32'h3b0172e5),
	.w6(32'h3a7c98c8),
	.w7(32'h3b9caeb0),
	.w8(32'h3bb96961),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130537),
	.w1(32'h3b684f03),
	.w2(32'h3be27d2a),
	.w3(32'hbc61d60b),
	.w4(32'hbb3152cc),
	.w5(32'h3c57b512),
	.w6(32'hbbafc8b7),
	.w7(32'hbc4cb1c3),
	.w8(32'hbbb5aad1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214f70),
	.w1(32'h3a0ab0ba),
	.w2(32'hbc17b8e5),
	.w3(32'h3aefa20b),
	.w4(32'hba1a878a),
	.w5(32'hbcd9e800),
	.w6(32'h3b92b8f8),
	.w7(32'h3b3bff6e),
	.w8(32'h3c7acfba),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd45e041),
	.w1(32'hbb7a6de7),
	.w2(32'hbbf71913),
	.w3(32'hbb956795),
	.w4(32'hbb34f48d),
	.w5(32'hba868404),
	.w6(32'hbc319fe5),
	.w7(32'hba7d3905),
	.w8(32'h3ca323cf),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef398e),
	.w1(32'hbb936f66),
	.w2(32'hbd1aae4c),
	.w3(32'h3b7b5d0a),
	.w4(32'h3a8775ee),
	.w5(32'hba81a7e1),
	.w6(32'h39eeff13),
	.w7(32'h3bd248e4),
	.w8(32'h3a9b208c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7052a6),
	.w1(32'hbbb3d8ff),
	.w2(32'h3b450b15),
	.w3(32'h3a6aecf3),
	.w4(32'hba14a0c0),
	.w5(32'hbbb56195),
	.w6(32'hbc0936c4),
	.w7(32'hbaf24d90),
	.w8(32'h3b9ac832),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b388eb5),
	.w1(32'hbb5dcf37),
	.w2(32'hbb40a84b),
	.w3(32'hbc6ec885),
	.w4(32'hbbc27a18),
	.w5(32'hbbad891d),
	.w6(32'hbb73da29),
	.w7(32'hbb123870),
	.w8(32'h3b376a4e),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0891a8),
	.w1(32'hba948472),
	.w2(32'h3b67e8d6),
	.w3(32'hbcbbef09),
	.w4(32'hbc533e82),
	.w5(32'hbc148ed2),
	.w6(32'hbb7e9ac1),
	.w7(32'hbbaf5024),
	.w8(32'hbc661dec),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb57bac),
	.w1(32'hbafdb2e1),
	.w2(32'hba0b7990),
	.w3(32'hbbcbd280),
	.w4(32'h39fb2a00),
	.w5(32'h3a443750),
	.w6(32'hb9d916f0),
	.w7(32'hbaaa0a3a),
	.w8(32'h3a921ebb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03cb76),
	.w1(32'hbac7a5ad),
	.w2(32'h39fb3846),
	.w3(32'hbc10a2ee),
	.w4(32'hbb717858),
	.w5(32'hbc3af877),
	.w6(32'hbbe57eb0),
	.w7(32'hbba88971),
	.w8(32'hbc1cb0fa),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49f1e5),
	.w1(32'hb9d79374),
	.w2(32'hbb703107),
	.w3(32'h3ccb7389),
	.w4(32'h3cb0b142),
	.w5(32'h3b313974),
	.w6(32'h3ad5ae35),
	.w7(32'h3b819973),
	.w8(32'hbb8b050a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf130b0),
	.w1(32'hbb7f3a49),
	.w2(32'hbc450ebc),
	.w3(32'hbbc67f1d),
	.w4(32'hba6d9eca),
	.w5(32'hbab8d549),
	.w6(32'hbb06db01),
	.w7(32'hbbb5e00f),
	.w8(32'hbb00f33b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813c97),
	.w1(32'hbb88f46a),
	.w2(32'hbc7cf43f),
	.w3(32'h3bb7d865),
	.w4(32'h3b4e3a0a),
	.w5(32'h3b538db2),
	.w6(32'h3ba91b5e),
	.w7(32'hbb3298ec),
	.w8(32'h3c5b9bc7),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c6465),
	.w1(32'h3c80da6a),
	.w2(32'hbc90e216),
	.w3(32'h3a0fda36),
	.w4(32'hbc6f596a),
	.w5(32'hbc3eb4fd),
	.w6(32'hbba0536d),
	.w7(32'hbb314b7f),
	.w8(32'hba9ac912),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b4c01),
	.w1(32'h3b9dc903),
	.w2(32'hbb2c6417),
	.w3(32'hbbcac45b),
	.w4(32'hbbbe1a69),
	.w5(32'h3a8ca223),
	.w6(32'hbbe2d6dd),
	.w7(32'hba6c920f),
	.w8(32'h3b109f3e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6e77),
	.w1(32'h3c440c29),
	.w2(32'hbb8c358f),
	.w3(32'h3bb435e3),
	.w4(32'hba432a77),
	.w5(32'hbb2691a2),
	.w6(32'hb821893d),
	.w7(32'h3a7bd09e),
	.w8(32'h3b925042),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67fa80),
	.w1(32'hbbc59128),
	.w2(32'h3d70a07a),
	.w3(32'h3b3d5bbb),
	.w4(32'hbb90a6cb),
	.w5(32'hbad4eebd),
	.w6(32'hbb6694a0),
	.w7(32'hbbad787c),
	.w8(32'h3c792069),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82f10d),
	.w1(32'hb9f22c4d),
	.w2(32'hbabcbcc3),
	.w3(32'h3b9e20fe),
	.w4(32'h3cabd818),
	.w5(32'hbc234eaf),
	.w6(32'hbbeb3f80),
	.w7(32'hbb993e43),
	.w8(32'hbb37bbcd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2fa2e),
	.w1(32'hbb8d2df2),
	.w2(32'hbbd59601),
	.w3(32'h3a8ea83f),
	.w4(32'hbb341d26),
	.w5(32'hbbc5788e),
	.w6(32'hbb7e891f),
	.w7(32'h39628f86),
	.w8(32'hb81e8f67),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c1074),
	.w1(32'hbbb64950),
	.w2(32'hbc13cf27),
	.w3(32'h3bda0c6f),
	.w4(32'hbb882616),
	.w5(32'h3b2958a6),
	.w6(32'hbbb3a3c3),
	.w7(32'h3d167b6f),
	.w8(32'hbbc8c229),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a5d58),
	.w1(32'h3b4fcd03),
	.w2(32'hbc846b6f),
	.w3(32'h3b0f220d),
	.w4(32'hbb21e6c2),
	.w5(32'hbc3a5009),
	.w6(32'hbc33f00b),
	.w7(32'hbc466590),
	.w8(32'hbc7b866d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123996),
	.w1(32'hbcc56225),
	.w2(32'hbb738acb),
	.w3(32'h3b849e2a),
	.w4(32'hba0e8b01),
	.w5(32'h3bbca6d6),
	.w6(32'h3bb80c5d),
	.w7(32'hbae15110),
	.w8(32'h3b6c14d0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc672ca4),
	.w1(32'hbb753c18),
	.w2(32'hbae47346),
	.w3(32'hbbad4763),
	.w4(32'hbc847f04),
	.w5(32'hbb26533d),
	.w6(32'hbbf61c8d),
	.w7(32'h39aef4d0),
	.w8(32'hbbf4243d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dd086),
	.w1(32'hbc28c39f),
	.w2(32'hbbe1f864),
	.w3(32'h3c7f3e9c),
	.w4(32'h3b778cfb),
	.w5(32'hbb1268f3),
	.w6(32'hbbc80722),
	.w7(32'h3c54ffea),
	.w8(32'hbc009474),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dbf47),
	.w1(32'hbc61c747),
	.w2(32'hbc1832af),
	.w3(32'hbb9f4fbe),
	.w4(32'h3a71b8da),
	.w5(32'hba08f1ba),
	.w6(32'hbbf85de3),
	.w7(32'h3bc3a007),
	.w8(32'h3ca71234),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f358),
	.w1(32'h3a4751f7),
	.w2(32'hb9ab0012),
	.w3(32'hbb0388e7),
	.w4(32'hba64ce64),
	.w5(32'hba0aa4a3),
	.w6(32'h38847965),
	.w7(32'hbbed3501),
	.w8(32'h38b5f63d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac330f5),
	.w1(32'h3b547727),
	.w2(32'hbc7bd5b2),
	.w3(32'hbb3e7a3a),
	.w4(32'h3c055e62),
	.w5(32'h3b2eebb3),
	.w6(32'hbbaadcc2),
	.w7(32'h3cd9e023),
	.w8(32'hbb80e79d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc6e97),
	.w1(32'hbb28c953),
	.w2(32'hbb4a0fcc),
	.w3(32'hbaba521a),
	.w4(32'h3bb9bd87),
	.w5(32'hbaa5a798),
	.w6(32'hbcd58d71),
	.w7(32'h3baeb47b),
	.w8(32'hb7ba40e7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1a1c),
	.w1(32'hbb17c54a),
	.w2(32'h3adf1309),
	.w3(32'h3d4ad6a3),
	.w4(32'hbc13b4e5),
	.w5(32'hbb499f04),
	.w6(32'h3ae13879),
	.w7(32'h3c66b38b),
	.w8(32'hbbb399cd),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119649),
	.w1(32'hba7bf7c5),
	.w2(32'hbc22b484),
	.w3(32'hbc86fef7),
	.w4(32'hbc23868f),
	.w5(32'hb9a7912a),
	.w6(32'hbb48b2a5),
	.w7(32'hbb02ad40),
	.w8(32'h3b04c05a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be82605),
	.w1(32'hbc526d63),
	.w2(32'hbc6fd1dc),
	.w3(32'h3b08e1c7),
	.w4(32'hba748950),
	.w5(32'hbba2967b),
	.w6(32'hb9164e33),
	.w7(32'h3c5d69e7),
	.w8(32'h3b39d429),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c259429),
	.w1(32'h3bc8e7ec),
	.w2(32'hba07f82c),
	.w3(32'hbc9c5448),
	.w4(32'h3beb0181),
	.w5(32'hb920820f),
	.w6(32'hbc5d9e71),
	.w7(32'h3bb3254d),
	.w8(32'h3c116e85),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cabb9),
	.w1(32'hbc37fd52),
	.w2(32'hbc44ac07),
	.w3(32'hbc125d83),
	.w4(32'hbcc0be20),
	.w5(32'h3c622bfd),
	.w6(32'hbad18a12),
	.w7(32'h3c0b275e),
	.w8(32'h3c082037),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcf279),
	.w1(32'h3b8251f6),
	.w2(32'h3b6d5e51),
	.w3(32'hbb6832fe),
	.w4(32'h3c2defe2),
	.w5(32'hbc23b2ab),
	.w6(32'hbd8242b3),
	.w7(32'hbd1fa46f),
	.w8(32'h3b9b16d7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ba3e5),
	.w1(32'h3c84c660),
	.w2(32'hbc6c403d),
	.w3(32'h3cd3ec0b),
	.w4(32'h3c24f6b2),
	.w5(32'h3cf63ec4),
	.w6(32'hbbc2b980),
	.w7(32'hbb24d7c6),
	.w8(32'hba0dd207),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25d73c),
	.w1(32'hbc25cd1a),
	.w2(32'hbc2014c7),
	.w3(32'hbc1235f3),
	.w4(32'hbc48f550),
	.w5(32'h3a646846),
	.w6(32'hbbcc01c7),
	.w7(32'h3cb841a9),
	.w8(32'hbaa6734a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e8119),
	.w1(32'hbbb8b8a2),
	.w2(32'h3c2211c6),
	.w3(32'h3bb694f4),
	.w4(32'h3c90fae2),
	.w5(32'h3b03a389),
	.w6(32'h3bef9495),
	.w7(32'hbc3d8974),
	.w8(32'hbac3e184),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc425e2e),
	.w1(32'h3c04dbeb),
	.w2(32'h3989c22d),
	.w3(32'h3b402993),
	.w4(32'hbc790f10),
	.w5(32'hbcaf722e),
	.w6(32'hbc834c2d),
	.w7(32'hbb045013),
	.w8(32'h3d97f3f2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ff09),
	.w1(32'h3a44f809),
	.w2(32'hbcf19136),
	.w3(32'hbae2e2c4),
	.w4(32'hbcab376d),
	.w5(32'hbcac4c81),
	.w6(32'hbc159215),
	.w7(32'hbc15a713),
	.w8(32'hbaf3f9e7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd26aca),
	.w1(32'h3c817854),
	.w2(32'hbb905bfb),
	.w3(32'hbd014f9f),
	.w4(32'h3c4cd17a),
	.w5(32'hbc01df43),
	.w6(32'h3bc99a6e),
	.w7(32'h3c28085a),
	.w8(32'hbc40d07d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d080f95),
	.w1(32'h3aff8d4a),
	.w2(32'hbbec19d3),
	.w3(32'h3aa46627),
	.w4(32'hbc34fc1a),
	.w5(32'h3b304b6f),
	.w6(32'h3cc69dbe),
	.w7(32'h3bcc79ef),
	.w8(32'hbb88d50c),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48975f),
	.w1(32'h3cb83d70),
	.w2(32'hbc6b8083),
	.w3(32'hbafb9fe3),
	.w4(32'hbae679c3),
	.w5(32'h35bf1148),
	.w6(32'h3b9147ea),
	.w7(32'hbb060978),
	.w8(32'hbcd4737d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eadf9),
	.w1(32'hbb5ec61c),
	.w2(32'hbc347a88),
	.w3(32'h3a38463d),
	.w4(32'hbb889de6),
	.w5(32'hbc52f4fb),
	.w6(32'hbce12013),
	.w7(32'h3b869b92),
	.w8(32'h3b53042d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ba515),
	.w1(32'h3bf65f8d),
	.w2(32'h38cce504),
	.w3(32'hbba4a233),
	.w4(32'hba48eb53),
	.w5(32'h3b1626f1),
	.w6(32'hbb5c680c),
	.w7(32'h3c59c93f),
	.w8(32'h3ae8dc9f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9696fb),
	.w1(32'h3af065b2),
	.w2(32'h3cfa319d),
	.w3(32'h3c91d3aa),
	.w4(32'h3c0a409e),
	.w5(32'h3c6ce588),
	.w6(32'h3b85e547),
	.w7(32'hbc0443f4),
	.w8(32'h3c12afb4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0fce9),
	.w1(32'h3b9ded04),
	.w2(32'h3b5b3ccb),
	.w3(32'hbc8f7af7),
	.w4(32'hbb443b81),
	.w5(32'h3c386ad6),
	.w6(32'h3afc0a38),
	.w7(32'hbc48d680),
	.w8(32'hbc014580),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2ff9b),
	.w1(32'hbcc189d5),
	.w2(32'hbc1c5bcd),
	.w3(32'hbc1b5d12),
	.w4(32'hbceffc13),
	.w5(32'h3c595cd7),
	.w6(32'hbb9157f3),
	.w7(32'hbb3a392a),
	.w8(32'hbc215d38),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b39e6),
	.w1(32'hbc5756a1),
	.w2(32'h3c773de9),
	.w3(32'h3c2e944e),
	.w4(32'hbb97c42e),
	.w5(32'hbcc4b3a6),
	.w6(32'h3cac9937),
	.w7(32'h3a6a7fd6),
	.w8(32'h3bfa3e30),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04cc89),
	.w1(32'h3b8d3e11),
	.w2(32'hbac48b72),
	.w3(32'h3b73a7ac),
	.w4(32'hbaad354f),
	.w5(32'h3c7402f8),
	.w6(32'hbccf6aa9),
	.w7(32'hb9c2727d),
	.w8(32'h398957b4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d5cb3),
	.w1(32'hbc6b9fee),
	.w2(32'hbb8c0feb),
	.w3(32'h3bc0cc60),
	.w4(32'hbc2ba3d3),
	.w5(32'hbcc4b8e2),
	.w6(32'h3b61cf0a),
	.w7(32'hbbcde844),
	.w8(32'h3b894dc3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf462b5),
	.w1(32'h3d1d0664),
	.w2(32'h3b50a734),
	.w3(32'h3c6fdb4d),
	.w4(32'h3b456f89),
	.w5(32'hbc2d723b),
	.w6(32'h3c3ad2a9),
	.w7(32'h3a7753bc),
	.w8(32'hbb4e99b6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9939b4),
	.w1(32'h3a09c91b),
	.w2(32'hbcc69a60),
	.w3(32'h3bd78c01),
	.w4(32'h3a9f3dc1),
	.w5(32'h3b9d344b),
	.w6(32'hba199a68),
	.w7(32'h3c91e50f),
	.w8(32'h3b5eb9ce),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa363f),
	.w1(32'hbc850f34),
	.w2(32'h3c2b87ff),
	.w3(32'hbbb7bf9f),
	.w4(32'h3ae3723d),
	.w5(32'h3b56e065),
	.w6(32'h3cb77655),
	.w7(32'hb9e4d895),
	.w8(32'h3b012da3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd0280),
	.w1(32'hbae4812f),
	.w2(32'h3af50a84),
	.w3(32'hbce23b86),
	.w4(32'hbba7a545),
	.w5(32'h3b60c42b),
	.w6(32'hbab34e40),
	.w7(32'h3a03edbf),
	.w8(32'hbbd7b3a4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20ccd2),
	.w1(32'h3a0ee97e),
	.w2(32'h3b09d6cf),
	.w3(32'h3cdca197),
	.w4(32'hbbda2ee8),
	.w5(32'h3c5ed122),
	.w6(32'h3bccb699),
	.w7(32'hbc3c3d24),
	.w8(32'h3cb018ad),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced287b),
	.w1(32'hbcaf733d),
	.w2(32'h3ad2f2dc),
	.w3(32'hbb5587ba),
	.w4(32'hbc13e4ad),
	.w5(32'h3c37f1d8),
	.w6(32'hbc589417),
	.w7(32'hbcb25ca6),
	.w8(32'h3b45f410),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d050b57),
	.w1(32'h3c9d6b60),
	.w2(32'h3c0e153e),
	.w3(32'hbc16ba56),
	.w4(32'h3a7da75f),
	.w5(32'h3c01e0e9),
	.w6(32'hbca9792a),
	.w7(32'h3bd29de5),
	.w8(32'hba2e1792),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d6784d),
	.w1(32'hbbc30678),
	.w2(32'h3c24afd4),
	.w3(32'h3cd6259f),
	.w4(32'h3a8e008b),
	.w5(32'hbc928738),
	.w6(32'h3c32882b),
	.w7(32'hbe10ea92),
	.w8(32'h3cc332fa),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91866c),
	.w1(32'hbb9974c6),
	.w2(32'hbcad2424),
	.w3(32'h3a04f9e1),
	.w4(32'hbc3c62a0),
	.w5(32'hbb43d2d6),
	.w6(32'h3c6b62df),
	.w7(32'h3c7f52ac),
	.w8(32'hb996a3c5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554636),
	.w1(32'hbb25819a),
	.w2(32'hbc9da8fe),
	.w3(32'h3ab16551),
	.w4(32'hbac9fe81),
	.w5(32'hbb0bc64f),
	.w6(32'hbb1903ef),
	.w7(32'h3c0b4d9c),
	.w8(32'hbc14901a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e5240),
	.w1(32'h39a44c57),
	.w2(32'hbb82e71b),
	.w3(32'hbbaeed74),
	.w4(32'hbc30df4e),
	.w5(32'h3bc7dd88),
	.w6(32'hbb477c83),
	.w7(32'hbbfa6b0e),
	.w8(32'hbbbfe1c8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b69eb),
	.w1(32'hbb2b53d2),
	.w2(32'h3ba5dde1),
	.w3(32'hbbe2d36b),
	.w4(32'hbb86a57f),
	.w5(32'hbb253971),
	.w6(32'hbb42ac18),
	.w7(32'hbd8107f8),
	.w8(32'hbbe0c4f6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04561c),
	.w1(32'hb9aa937f),
	.w2(32'hb80ee0a8),
	.w3(32'hbbf63f20),
	.w4(32'h3b8d1f6b),
	.w5(32'h3c9670d9),
	.w6(32'h3c3de573),
	.w7(32'hbbb60395),
	.w8(32'hbbdcad74),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc519e80),
	.w1(32'hbb8842c2),
	.w2(32'hbb8965d7),
	.w3(32'h3c026a2e),
	.w4(32'hbae84fb0),
	.w5(32'h3bb62661),
	.w6(32'hbb83d272),
	.w7(32'h383c876c),
	.w8(32'hbc35d4a2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28fdb9),
	.w1(32'h3ab20014),
	.w2(32'hbb72e701),
	.w3(32'h3bc5b020),
	.w4(32'hba5b3901),
	.w5(32'hbb21adb4),
	.w6(32'hbac01527),
	.w7(32'hbb79ce91),
	.w8(32'h3beed708),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8abfb5),
	.w1(32'h397e1e03),
	.w2(32'h3c05b316),
	.w3(32'h39534660),
	.w4(32'hbc30f69f),
	.w5(32'hbbb9ec3f),
	.w6(32'h3af068f9),
	.w7(32'h3b8ba18e),
	.w8(32'hbc0d4efb),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d58b39),
	.w1(32'hbbb4fbeb),
	.w2(32'hba5d0bd3),
	.w3(32'hb9d35072),
	.w4(32'h3bb9dce3),
	.w5(32'hbb092e9f),
	.w6(32'hbae3b0bc),
	.w7(32'hba9d44ae),
	.w8(32'h3b4a5849),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292bc9),
	.w1(32'h3cad3bcc),
	.w2(32'h3bc3e21e),
	.w3(32'hbb63519b),
	.w4(32'h3b8963a5),
	.w5(32'hbc15bc72),
	.w6(32'hba6bd1ae),
	.w7(32'hb6c5378d),
	.w8(32'hbbb30b80),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841536f),
	.w1(32'h3a8d5417),
	.w2(32'hbba18341),
	.w3(32'h3a0dbb78),
	.w4(32'hba4d3a21),
	.w5(32'hbc0c9452),
	.w6(32'hbb7198a8),
	.w7(32'hbc5020fe),
	.w8(32'h3c895b05),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fce09),
	.w1(32'hb974b43f),
	.w2(32'h3a3e6563),
	.w3(32'h399ef0d0),
	.w4(32'h3a0dfc50),
	.w5(32'hbc86c173),
	.w6(32'h3bd444b8),
	.w7(32'hbc6dab06),
	.w8(32'h392a1593),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3be3),
	.w1(32'h3a351a31),
	.w2(32'hbc1f0fe6),
	.w3(32'hbc0a0660),
	.w4(32'hbc0f4cd8),
	.w5(32'hba45ab60),
	.w6(32'h3a75a55a),
	.w7(32'hbaaa150a),
	.w8(32'hbb0d3534),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80abe7),
	.w1(32'hbaef1dce),
	.w2(32'h3b2b4577),
	.w3(32'h3a2256f0),
	.w4(32'h3a8a07bb),
	.w5(32'h3b0470ce),
	.w6(32'h3b737995),
	.w7(32'hbbf76e10),
	.w8(32'h3b87ffa7),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabeb124),
	.w1(32'hbb33fdc9),
	.w2(32'hbbdc4139),
	.w3(32'hbb4de630),
	.w4(32'hba86973f),
	.w5(32'hbac52e7f),
	.w6(32'hbc9e7017),
	.w7(32'hbbeaa6ab),
	.w8(32'hbb576432),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe86792),
	.w1(32'hbc01af25),
	.w2(32'hbc97c2e6),
	.w3(32'hbc12108d),
	.w4(32'hbb7cef03),
	.w5(32'hbb37de61),
	.w6(32'h3ab238af),
	.w7(32'h3d28a4f9),
	.w8(32'hbc038345),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bb8c8),
	.w1(32'h3adcf489),
	.w2(32'h39a0526f),
	.w3(32'hbbb3f222),
	.w4(32'h3be52b85),
	.w5(32'h3b1c6569),
	.w6(32'h3ba96f9d),
	.w7(32'hbbee5aa3),
	.w8(32'hb9c567a3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90553b),
	.w1(32'h3b9eb476),
	.w2(32'h3a97c37c),
	.w3(32'hbbcd39a9),
	.w4(32'h3ab6adc0),
	.w5(32'h3bb5d617),
	.w6(32'h3a149b8c),
	.w7(32'hb8e1ae68),
	.w8(32'h3b52015d),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57f346),
	.w1(32'hbb4fa7cf),
	.w2(32'h3ac4ed93),
	.w3(32'hbadc4bda),
	.w4(32'h3cb7449c),
	.w5(32'h3aed19f3),
	.w6(32'h3c0344f1),
	.w7(32'hb9c72299),
	.w8(32'h3ba6182e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1bd9e),
	.w1(32'h39ad2cd1),
	.w2(32'h3a3b3407),
	.w3(32'hbb87e82d),
	.w4(32'h3b030840),
	.w5(32'hbc394145),
	.w6(32'h3b2ebea5),
	.w7(32'hbb57014f),
	.w8(32'hbcf79409),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc690e),
	.w1(32'h386cdf73),
	.w2(32'h3b7a59fc),
	.w3(32'hbbafc411),
	.w4(32'h3a8863f6),
	.w5(32'h3b929b60),
	.w6(32'hbca88258),
	.w7(32'hba8dcb01),
	.w8(32'hbc32e0b7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba688d0),
	.w1(32'hbb48df04),
	.w2(32'hbc26d688),
	.w3(32'hbb0ba0e2),
	.w4(32'hbbf41a9c),
	.w5(32'hba4e60b6),
	.w6(32'h3abd9060),
	.w7(32'h3b46e69f),
	.w8(32'hbac42847),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c808690),
	.w1(32'h3bddd0d4),
	.w2(32'h39806dcc),
	.w3(32'hbb55a0c6),
	.w4(32'h3be13eba),
	.w5(32'hbb993b39),
	.w6(32'hbbda5caa),
	.w7(32'hbc28d166),
	.w8(32'hbb40a772),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3c620),
	.w1(32'h3a86f14e),
	.w2(32'hba8a73d6),
	.w3(32'hba30682d),
	.w4(32'h3b8ea181),
	.w5(32'hbc0dc7a7),
	.w6(32'hbb8f3b0a),
	.w7(32'hbc6c8ba6),
	.w8(32'hba0674bd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9642ef),
	.w1(32'hbaab4a91),
	.w2(32'hbb682651),
	.w3(32'h36d9f5ea),
	.w4(32'h3a0e90bc),
	.w5(32'hbab1b122),
	.w6(32'h3b520c29),
	.w7(32'hb8833227),
	.w8(32'hbab11a26),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b014e64),
	.w1(32'hba5c44d7),
	.w2(32'h3bda4ecd),
	.w3(32'hbb8f69fd),
	.w4(32'hbb09481a),
	.w5(32'hbb33a787),
	.w6(32'h3c0cc5a4),
	.w7(32'hbb4f3e53),
	.w8(32'hbbd9f3b7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bc0c9),
	.w1(32'h3bbb59e5),
	.w2(32'hbb501a68),
	.w3(32'hbc68052d),
	.w4(32'h3b95d4a7),
	.w5(32'hbb6d8219),
	.w6(32'h3aa27cd3),
	.w7(32'h38a7d799),
	.w8(32'h3beab17a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5fdba),
	.w1(32'hbb6f5ab1),
	.w2(32'hbbb4f2f3),
	.w3(32'hbb3d5363),
	.w4(32'hbcda67b4),
	.w5(32'hbab545e8),
	.w6(32'h3ad0b640),
	.w7(32'hbb8c08b0),
	.w8(32'hbc10124b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe890c1),
	.w1(32'hbc2b563a),
	.w2(32'hbb743d71),
	.w3(32'hba47f267),
	.w4(32'hbba0d8d5),
	.w5(32'hbbf2d96f),
	.w6(32'h3c0f222f),
	.w7(32'hbb472fba),
	.w8(32'h3bd13912),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4466eb),
	.w1(32'hbb0243c1),
	.w2(32'h3b6e8b9b),
	.w3(32'hbae970e8),
	.w4(32'h3c2ea531),
	.w5(32'hbbd3cfc4),
	.w6(32'h3bc72a00),
	.w7(32'h3aac16f8),
	.w8(32'h3c303578),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38e4fa),
	.w1(32'hb89dc0e8),
	.w2(32'h3c006217),
	.w3(32'hbb1a7393),
	.w4(32'h3c51d4e2),
	.w5(32'hbbfc21de),
	.w6(32'hbb82a712),
	.w7(32'h3beb8f3d),
	.w8(32'h3c5e82e1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule