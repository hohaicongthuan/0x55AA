module layer_8_featuremap_144(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803f6c),
	.w1(32'hbc197104),
	.w2(32'hbbe9c6b2),
	.w3(32'h3be8f0ea),
	.w4(32'hbc0b705e),
	.w5(32'hbbe28494),
	.w6(32'hbc1a6983),
	.w7(32'h3a49708a),
	.w8(32'h3b104be3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b980a1f),
	.w1(32'h3864bed4),
	.w2(32'hbb87e958),
	.w3(32'hb8cdcb39),
	.w4(32'hbb50a79e),
	.w5(32'hbbc24d73),
	.w6(32'hbb8aa43f),
	.w7(32'h3bd52b02),
	.w8(32'h3c5f033f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f618c),
	.w1(32'hbb4cd9ba),
	.w2(32'hbcbbc16b),
	.w3(32'h3b719a97),
	.w4(32'hbbd4cd95),
	.w5(32'hbbbf691c),
	.w6(32'hbbf1dcd9),
	.w7(32'hbad90839),
	.w8(32'h3c3fdd16),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99ec10),
	.w1(32'hbc3d2da7),
	.w2(32'h3c8389da),
	.w3(32'h3ca761ab),
	.w4(32'h3c14a0e7),
	.w5(32'hbc88580f),
	.w6(32'hbc9926b0),
	.w7(32'h3c9cfff7),
	.w8(32'h3c3a638c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1877ba),
	.w1(32'h3ba69cac),
	.w2(32'h3c5dd1a1),
	.w3(32'hbcbbad30),
	.w4(32'hbb33fe45),
	.w5(32'h3ca2913c),
	.w6(32'hbcf632c0),
	.w7(32'hbc3ef993),
	.w8(32'hbc9ded87),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd2e7),
	.w1(32'h3b4c148e),
	.w2(32'h3bd7fa85),
	.w3(32'h3cbf0dd7),
	.w4(32'h3bbc7dbf),
	.w5(32'hbc975d56),
	.w6(32'h3cefaa7d),
	.w7(32'h3ccfc0d8),
	.w8(32'h3c271907),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087310),
	.w1(32'h3c529957),
	.w2(32'hbc22d0e3),
	.w3(32'hbc865478),
	.w4(32'h39c3366d),
	.w5(32'hbb913f56),
	.w6(32'hbc522ae7),
	.w7(32'h3c3ccf7f),
	.w8(32'h3c23c851),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95e98e),
	.w1(32'hbc30aa6a),
	.w2(32'h3b658434),
	.w3(32'hbc1c8c6e),
	.w4(32'h3abe0fff),
	.w5(32'hbbdca193),
	.w6(32'hbbf5dede),
	.w7(32'h3b3c59e4),
	.w8(32'hbbaae63c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b774022),
	.w1(32'hbb8fe91d),
	.w2(32'h3b98f3f4),
	.w3(32'hbaabec02),
	.w4(32'hbc568078),
	.w5(32'hbc8809c5),
	.w6(32'hbc65c8f5),
	.w7(32'hbbd53f4d),
	.w8(32'hbae76522),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a4cfd),
	.w1(32'h3c32e222),
	.w2(32'hbc02aea6),
	.w3(32'hbb66c749),
	.w4(32'hbb455ac9),
	.w5(32'hbbe92c4f),
	.w6(32'hbafa9609),
	.w7(32'hbbe1c4d5),
	.w8(32'h3c0eef5e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d4ecc),
	.w1(32'h3c6c7e9b),
	.w2(32'hbc8d9594),
	.w3(32'h3c40b25b),
	.w4(32'hbc8f102e),
	.w5(32'h3b9a5187),
	.w6(32'hbc897621),
	.w7(32'hbd021de9),
	.w8(32'hbc655625),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd126e6d),
	.w1(32'hbcaff5a1),
	.w2(32'h3c378c1f),
	.w3(32'h3c9629b2),
	.w4(32'hba87d333),
	.w5(32'hbc6f0413),
	.w6(32'h3c8e45ae),
	.w7(32'h3c36112c),
	.w8(32'hbc7ef28b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4484),
	.w1(32'hbc6b418b),
	.w2(32'h3b65a7f9),
	.w3(32'h3baf186d),
	.w4(32'h3b13595f),
	.w5(32'hbb82fc07),
	.w6(32'h3ba5fe0d),
	.w7(32'h3ab67b3d),
	.w8(32'hbaf0bad4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0f5a),
	.w1(32'h3b871fd4),
	.w2(32'h3b03f955),
	.w3(32'hbb17c2e8),
	.w4(32'h3ad9c54f),
	.w5(32'hbbd5c288),
	.w6(32'hb83bb711),
	.w7(32'h3b15d978),
	.w8(32'hbba1df33),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168afc),
	.w1(32'hba205f50),
	.w2(32'h3b890af3),
	.w3(32'hbc212172),
	.w4(32'h3b0a7831),
	.w5(32'hbbfb0741),
	.w6(32'hbbaf433a),
	.w7(32'h3b65eda3),
	.w8(32'hbbc3a72c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbd6df),
	.w1(32'h39be8e23),
	.w2(32'hbbee85f2),
	.w3(32'hbc0fcaee),
	.w4(32'h3c14f82f),
	.w5(32'h3c66e88a),
	.w6(32'hbbe4a3fc),
	.w7(32'hbbabd30d),
	.w8(32'hbb96bef0),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae5dbb),
	.w1(32'hbb4f444b),
	.w2(32'hbc05a038),
	.w3(32'hbc317275),
	.w4(32'hbb82f13e),
	.w5(32'h3bd4e2e4),
	.w6(32'h3cda8e6d),
	.w7(32'h3bba492f),
	.w8(32'h3c67c9e8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58b5d7),
	.w1(32'hbafa95bf),
	.w2(32'hbc25750f),
	.w3(32'h3c14dde5),
	.w4(32'hbbce1277),
	.w5(32'h3c65a842),
	.w6(32'h3bd39b6a),
	.w7(32'hbc6253f2),
	.w8(32'hbc9d7d87),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdcc752),
	.w1(32'hbc00a1c4),
	.w2(32'h3c60b385),
	.w3(32'h3ba6a294),
	.w4(32'hbc1712f8),
	.w5(32'h3c045dc9),
	.w6(32'h3bfe0432),
	.w7(32'h395624f5),
	.w8(32'hbc46f1cc),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3252ab),
	.w1(32'hbcb33b8e),
	.w2(32'h3c295244),
	.w3(32'h3c350d11),
	.w4(32'hbcb538f0),
	.w5(32'hb9db926f),
	.w6(32'h3be9f5a7),
	.w7(32'hbc0ad992),
	.w8(32'hbc185d70),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b480b49),
	.w1(32'hbbe945ab),
	.w2(32'hbb1b3a6c),
	.w3(32'h3cb57d95),
	.w4(32'hbbd27d5c),
	.w5(32'h3a665800),
	.w6(32'h3c1915b6),
	.w7(32'hbc0e00b3),
	.w8(32'hba8ad578),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266d38),
	.w1(32'h3c496ba9),
	.w2(32'hbd07e38a),
	.w3(32'hbc00e630),
	.w4(32'h3bef3bec),
	.w5(32'hbb971288),
	.w6(32'h3c0e04c1),
	.w7(32'hbb6edc40),
	.w8(32'h3c95dcd4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b746329),
	.w1(32'h3aff7cca),
	.w2(32'h3bace7db),
	.w3(32'hbbfc2241),
	.w4(32'hbc68357d),
	.w5(32'hbb3f7a99),
	.w6(32'hbc3344e1),
	.w7(32'hbc1c5acd),
	.w8(32'hbbc14a0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38b4b6),
	.w1(32'h3ad7af3e),
	.w2(32'h3bccfbe7),
	.w3(32'hba24d949),
	.w4(32'h3c3db881),
	.w5(32'hbbcc1d64),
	.w6(32'h3c0c2d78),
	.w7(32'h3c19fa43),
	.w8(32'hbc3ffb76),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fe3a0),
	.w1(32'hbc77e0a6),
	.w2(32'hbbc275ec),
	.w3(32'hbbc8277a),
	.w4(32'h3a929c5b),
	.w5(32'h3c4fe7e4),
	.w6(32'hbc46b673),
	.w7(32'hbbf68731),
	.w8(32'hbb6a5e52),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f1322),
	.w1(32'hbaa9965a),
	.w2(32'h3cb888e2),
	.w3(32'h3c1b406d),
	.w4(32'h3b539af5),
	.w5(32'hbccbe38a),
	.w6(32'h3bf272f3),
	.w7(32'h3ce27c0b),
	.w8(32'h3c1261f8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a7756),
	.w1(32'hbc26eb71),
	.w2(32'hbbbc5a56),
	.w3(32'hbcbb60b8),
	.w4(32'hbbcdb24c),
	.w5(32'h3c37d042),
	.w6(32'hbcb7b999),
	.w7(32'hbc92a8cc),
	.w8(32'hbc12be87),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe80615),
	.w1(32'h3a1fc958),
	.w2(32'hbc80dc56),
	.w3(32'h3c98ab1b),
	.w4(32'hbb0f3800),
	.w5(32'h3aa1a1fa),
	.w6(32'h3cb74e93),
	.w7(32'hbc0e0020),
	.w8(32'h3c6ae772),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac864ff),
	.w1(32'h3ba9c1fa),
	.w2(32'h3c95d33e),
	.w3(32'hbbb06ecf),
	.w4(32'h3b0fa258),
	.w5(32'hbcbeb667),
	.w6(32'h3c120159),
	.w7(32'h3cfc37c8),
	.w8(32'hbacacc2e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08a651),
	.w1(32'hb9d2f4a4),
	.w2(32'hbc0150aa),
	.w3(32'h3a8ff0e5),
	.w4(32'h3bc68ba8),
	.w5(32'h3bc8f3eb),
	.w6(32'hbd0c9774),
	.w7(32'hbb2279ff),
	.w8(32'hbb0d030f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28d30a),
	.w1(32'h3c1dc98b),
	.w2(32'h3c029875),
	.w3(32'h3a55a32d),
	.w4(32'hbadc6f65),
	.w5(32'hbb3524e0),
	.w6(32'h3cb12764),
	.w7(32'h3b4a1d19),
	.w8(32'h3aee541f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02302e),
	.w1(32'h3b34b6da),
	.w2(32'hbd256364),
	.w3(32'hbbda9d87),
	.w4(32'h3bc9cd99),
	.w5(32'h3c7ad2ca),
	.w6(32'hbb975d98),
	.w7(32'hbcc8311d),
	.w8(32'hbb516ec5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20f300),
	.w1(32'h3c602125),
	.w2(32'h3c94c6d7),
	.w3(32'h3ca54ea1),
	.w4(32'h3bc8a929),
	.w5(32'h3ba83bb2),
	.w6(32'h3d04b8b1),
	.w7(32'h3c804fc9),
	.w8(32'h3c3fe1f1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d067535),
	.w1(32'hbbbe68d6),
	.w2(32'hbb9dfbfb),
	.w3(32'hbb5907dd),
	.w4(32'h3b525159),
	.w5(32'h3bf7e0d8),
	.w6(32'hbcc6d5f3),
	.w7(32'hbae1775b),
	.w8(32'hbbe3ab27),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e1d25),
	.w1(32'hbc6db9ca),
	.w2(32'h3c8872d1),
	.w3(32'h3c978ee4),
	.w4(32'h3beb31ec),
	.w5(32'hbbd1ef2a),
	.w6(32'hbb5b620e),
	.w7(32'h3c84a2f5),
	.w8(32'h3b773955),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb34585),
	.w1(32'h3b9f2a04),
	.w2(32'h3ad2499f),
	.w3(32'hbc99bb17),
	.w4(32'hb99e9a11),
	.w5(32'hbc6e670d),
	.w6(32'hbc44d261),
	.w7(32'h3b8835fd),
	.w8(32'h3b4a109f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd2451e),
	.w1(32'h3cf12e7d),
	.w2(32'hbb35f98e),
	.w3(32'hbcc4f54b),
	.w4(32'h3be5ddd5),
	.w5(32'h3c6eb889),
	.w6(32'hbca2bbd2),
	.w7(32'h3c2746f1),
	.w8(32'h3bb69113),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03973),
	.w1(32'h3ac14475),
	.w2(32'hba7babad),
	.w3(32'h3c28aa94),
	.w4(32'hbb736901),
	.w5(32'h3cb85fab),
	.w6(32'h3be083f1),
	.w7(32'h3c28587d),
	.w8(32'h3c72e646),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ee8ed),
	.w1(32'hbc957e54),
	.w2(32'hbcbbe687),
	.w3(32'h3c3dfd18),
	.w4(32'hbbd6a2b9),
	.w5(32'h3c19b089),
	.w6(32'hb9f252ce),
	.w7(32'hbc76a9bc),
	.w8(32'h3b595876),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc473cc3),
	.w1(32'hbc2c4771),
	.w2(32'h3c16c392),
	.w3(32'h3c4c2738),
	.w4(32'hbc625d4f),
	.w5(32'hbb7fa8bb),
	.w6(32'h3ba858ed),
	.w7(32'h3c1948e0),
	.w8(32'h3b04a637),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d8248),
	.w1(32'hbb860427),
	.w2(32'hbcc00f49),
	.w3(32'h3b1efad4),
	.w4(32'hbbfbea67),
	.w5(32'h3c12e128),
	.w6(32'h3c2a9a5f),
	.w7(32'hbca84d1f),
	.w8(32'hbc9e1128),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfcc422),
	.w1(32'hbc113537),
	.w2(32'h3b1d9bce),
	.w3(32'h3c08cb4a),
	.w4(32'hbc9acd11),
	.w5(32'h3a010c53),
	.w6(32'h3c08d765),
	.w7(32'hbc6f7fc1),
	.w8(32'hbbe13e82),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cc6b),
	.w1(32'h3c801c28),
	.w2(32'h3b8b06da),
	.w3(32'h3c1fcac6),
	.w4(32'h3bab621a),
	.w5(32'hbbefb3ea),
	.w6(32'h3cf7e62f),
	.w7(32'h3c853a3c),
	.w8(32'hbb71c0e1),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7da90b),
	.w1(32'h38a2f5f9),
	.w2(32'h3b71ec0e),
	.w3(32'hbc8ec93a),
	.w4(32'h3a4b00f0),
	.w5(32'hbbc7809d),
	.w6(32'hbb906af0),
	.w7(32'h3a626683),
	.w8(32'hbb2c8862),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45d3a1),
	.w1(32'h3aeffcb0),
	.w2(32'hbc59e348),
	.w3(32'hbbb82a1d),
	.w4(32'h3bcbc599),
	.w5(32'hbc8ed941),
	.w6(32'hbb53049c),
	.w7(32'h3c616d79),
	.w8(32'h3c53c0f1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68cdbb),
	.w1(32'h3c382d6b),
	.w2(32'hbb53c895),
	.w3(32'hbbb76058),
	.w4(32'h3b34a74b),
	.w5(32'hbb809336),
	.w6(32'hbc3a14fe),
	.w7(32'h3b2d538d),
	.w8(32'h3b848cd7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8e87),
	.w1(32'h3a737caf),
	.w2(32'h3cbc361e),
	.w3(32'hbc626c59),
	.w4(32'h3ad7db9f),
	.w5(32'hbceb953f),
	.w6(32'hbc08493a),
	.w7(32'h3cee01e5),
	.w8(32'h39a4bb40),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01d79f),
	.w1(32'h3c194753),
	.w2(32'hba3ef23d),
	.w3(32'hbc3a05f1),
	.w4(32'h3c7174b8),
	.w5(32'hbc81e89c),
	.w6(32'hbcbb81e7),
	.w7(32'h3c9c07c9),
	.w8(32'h3ac21501),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf23e1b),
	.w1(32'h3c14520a),
	.w2(32'hbd2f7240),
	.w3(32'hbc46b021),
	.w4(32'hbbd3fe03),
	.w5(32'h3c975184),
	.w6(32'hbd06d0ed),
	.w7(32'hbd2fe80e),
	.w8(32'h3b3d1919),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1c2bf7),
	.w1(32'h3afb5988),
	.w2(32'hbd8fe98c),
	.w3(32'h3c81a6fc),
	.w4(32'hbbd563c1),
	.w5(32'h3d16b964),
	.w6(32'h3d02b87f),
	.w7(32'hbd36cbe9),
	.w8(32'h3b10c74c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8ae584),
	.w1(32'hbcae40c1),
	.w2(32'h3bf6ad3f),
	.w3(32'h3d68ea20),
	.w4(32'hbb0ee350),
	.w5(32'h3d002128),
	.w6(32'h3d3c5b12),
	.w7(32'hba690d4c),
	.w8(32'hbc14f517),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cd34a),
	.w1(32'hbc1f50d2),
	.w2(32'h3ba7e599),
	.w3(32'h3c92bd5b),
	.w4(32'h3ba2fabb),
	.w5(32'hbc9af4e2),
	.w6(32'h3bc47e64),
	.w7(32'h3c8da7ad),
	.w8(32'h3b863e17),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1614e4),
	.w1(32'h3cea933f),
	.w2(32'hbc364bef),
	.w3(32'hbc67258e),
	.w4(32'hbc2f171f),
	.w5(32'h3c77c5ff),
	.w6(32'h3b3d8190),
	.w7(32'hbc19f5f4),
	.w8(32'hbabe2485),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc007e9),
	.w1(32'h3b311677),
	.w2(32'h3915e200),
	.w3(32'hb99acbce),
	.w4(32'h3a834d08),
	.w5(32'hbb80ea04),
	.w6(32'hbb2beaa4),
	.w7(32'hb88ffe68),
	.w8(32'hba1a2862),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbb0b4),
	.w1(32'h3aab80d4),
	.w2(32'hbb8e4e7d),
	.w3(32'hbb97cf46),
	.w4(32'hb93acc5d),
	.w5(32'hbb39dfa9),
	.w6(32'hbb3c1be8),
	.w7(32'h3c76f3fc),
	.w8(32'hba943ce8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab43f2),
	.w1(32'hbb7b0f65),
	.w2(32'hbceb3853),
	.w3(32'h3bc3e986),
	.w4(32'hbaef2944),
	.w5(32'h3c583c5b),
	.w6(32'hbc651c66),
	.w7(32'hbc921f22),
	.w8(32'h3bc8c934),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd62385),
	.w1(32'hbc11fa9b),
	.w2(32'hbbbbbddf),
	.w3(32'h3c660c3b),
	.w4(32'hbbaec836),
	.w5(32'hbbd00335),
	.w6(32'h3b26065b),
	.w7(32'hbbcc43cc),
	.w8(32'hbb8b41e1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90973b),
	.w1(32'hba75536f),
	.w2(32'h3c477bdb),
	.w3(32'h3b881bcb),
	.w4(32'h3c44e96a),
	.w5(32'h3c944882),
	.w6(32'h3bc41caa),
	.w7(32'h3c8cc3eb),
	.w8(32'h3b7c8e5d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d0605),
	.w1(32'hbca68fd5),
	.w2(32'h3b008298),
	.w3(32'hba144bff),
	.w4(32'h3a14e74b),
	.w5(32'hbb7d9536),
	.w6(32'hbc6ab1f7),
	.w7(32'h394c8cb3),
	.w8(32'hbad8f6d8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdf95e),
	.w1(32'h3a6c4400),
	.w2(32'h3b19712d),
	.w3(32'hbb8d1adf),
	.w4(32'h3b3d2cfe),
	.w5(32'h3af4dade),
	.w6(32'hbb5bf606),
	.w7(32'hbb4f1dbf),
	.w8(32'hbbc4c770),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97b148),
	.w1(32'h3b1e1a54),
	.w2(32'hbc96ab9c),
	.w3(32'h3c2d65a8),
	.w4(32'h3bba28b6),
	.w5(32'h3c92c96e),
	.w6(32'hba0de74c),
	.w7(32'hbc4b1708),
	.w8(32'h3b926906),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07e07),
	.w1(32'h3c50bcc5),
	.w2(32'hbbb63af1),
	.w3(32'h3c8cb87f),
	.w4(32'hbba44a3a),
	.w5(32'hbc262f96),
	.w6(32'h3c5aff11),
	.w7(32'hbbcf5593),
	.w8(32'hbcb5ba2a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ebe8d),
	.w1(32'hbc940499),
	.w2(32'h3b3d582d),
	.w3(32'h3b471017),
	.w4(32'h3bd3f953),
	.w5(32'h3b7eaa26),
	.w6(32'hbc3fbc91),
	.w7(32'h3be0b5bd),
	.w8(32'h3b5542a3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43437),
	.w1(32'hbbeb604a),
	.w2(32'hbb8fdf8c),
	.w3(32'hbbf04acb),
	.w4(32'hbbba08cc),
	.w5(32'hbb3aa684),
	.w6(32'hbc2f2510),
	.w7(32'h3abb1411),
	.w8(32'h3c9edd8b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bb949),
	.w1(32'hbb5d35f3),
	.w2(32'h3cda4caa),
	.w3(32'hbbcdf302),
	.w4(32'hbbaa8394),
	.w5(32'hbc664455),
	.w6(32'h3ae60478),
	.w7(32'h3ca653f0),
	.w8(32'hbaa54509),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf4223),
	.w1(32'h3bbe6658),
	.w2(32'h3c86d999),
	.w3(32'hbc8b4161),
	.w4(32'h3c3287ca),
	.w5(32'h3c820bf7),
	.w6(32'hbbc850e8),
	.w7(32'h3c9fb9b3),
	.w8(32'h3bacf561),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2bf80),
	.w1(32'hbcad5251),
	.w2(32'h3c6739ac),
	.w3(32'h3b896edf),
	.w4(32'hbbd01c84),
	.w5(32'h3baf0264),
	.w6(32'hbc1f0a2f),
	.w7(32'hbaf1c3a9),
	.w8(32'h39e3ac23),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5fced),
	.w1(32'hbccc2f7e),
	.w2(32'hbbb23913),
	.w3(32'h3cae5df4),
	.w4(32'hbc114676),
	.w5(32'h3c3613cb),
	.w6(32'hbc5c4fed),
	.w7(32'hbc9b100e),
	.w8(32'h3b255065),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa94cbc),
	.w1(32'h3c1e41b5),
	.w2(32'hbcdcb1f2),
	.w3(32'h3c258fa0),
	.w4(32'hbb66768e),
	.w5(32'h3c1d5a14),
	.w6(32'h3cacfd59),
	.w7(32'hbcbf4f04),
	.w8(32'h3b2cfa6d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcac307d),
	.w1(32'h3baa648c),
	.w2(32'hbc719c87),
	.w3(32'h3a100971),
	.w4(32'h3c5974c3),
	.w5(32'h3ce1720f),
	.w6(32'h3c9d4a4f),
	.w7(32'hbbbb658a),
	.w8(32'h398311da),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce83976),
	.w1(32'hbb910cc2),
	.w2(32'hbca10575),
	.w3(32'h3cd9cbef),
	.w4(32'h3bed361f),
	.w5(32'h3caff8b7),
	.w6(32'h3c2db3f0),
	.w7(32'hbc7a5a4c),
	.w8(32'h3a81b990),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07a918),
	.w1(32'h3cc3cba2),
	.w2(32'hbcd661b3),
	.w3(32'h3d32226b),
	.w4(32'h3c2d6b01),
	.w5(32'h3c299f1d),
	.w6(32'h3d1eb3a5),
	.w7(32'hbbb2ad2e),
	.w8(32'h3c8930fe),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc7750d),
	.w1(32'hbbac4956),
	.w2(32'hbc531ed3),
	.w3(32'hbc1c8923),
	.w4(32'hbc030ba2),
	.w5(32'hbb4fee82),
	.w6(32'h3b656c58),
	.w7(32'hbc8e05c2),
	.w8(32'hbc057600),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2dbae),
	.w1(32'hbbce9b0f),
	.w2(32'h3a3a9775),
	.w3(32'h3bc40159),
	.w4(32'hbbb87fb2),
	.w5(32'h3c29c0fb),
	.w6(32'h3bda1173),
	.w7(32'hbbcd98c3),
	.w8(32'hbbfb819d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff801a),
	.w1(32'h3b447931),
	.w2(32'h3ba6c138),
	.w3(32'h3c5112fa),
	.w4(32'h3b92a0c9),
	.w5(32'h3c8f196e),
	.w6(32'h3cdc11e6),
	.w7(32'hbb753123),
	.w8(32'hbc8b5e7c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf54c72),
	.w1(32'hba4c3b32),
	.w2(32'hbcb14e47),
	.w3(32'h3ce1fbf6),
	.w4(32'h3c4e3563),
	.w5(32'h3c0a6914),
	.w6(32'h3c3ce4be),
	.w7(32'hbc31da4a),
	.w8(32'h3b8e206e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca64b2c),
	.w1(32'h3c05cd20),
	.w2(32'hbb41df85),
	.w3(32'hbb906f15),
	.w4(32'h3a86d3e4),
	.w5(32'h3b7c3d76),
	.w6(32'h3b1a71cf),
	.w7(32'h3ad6e5ab),
	.w8(32'h3b5517fa),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46fbb3),
	.w1(32'hbb55d506),
	.w2(32'h3c13605f),
	.w3(32'h39c6f7ac),
	.w4(32'h3ade97ea),
	.w5(32'h3c161068),
	.w6(32'h3ad49795),
	.w7(32'h3beaaa00),
	.w8(32'h3c61dfcf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c266c58),
	.w1(32'h3c135c8e),
	.w2(32'h3c0d0a3a),
	.w3(32'h3be3b703),
	.w4(32'h3b209855),
	.w5(32'h3bf52704),
	.w6(32'h3c803c08),
	.w7(32'h3bda617d),
	.w8(32'h3c29183c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b847),
	.w1(32'h3b8745f6),
	.w2(32'h3b07d644),
	.w3(32'h3ad89a50),
	.w4(32'hbc18d2fc),
	.w5(32'hbc7509e3),
	.w6(32'h3b8bfd22),
	.w7(32'hbbb0fbd9),
	.w8(32'hbb9e9cb4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f1919),
	.w1(32'h3c4e7f07),
	.w2(32'hbbc071cf),
	.w3(32'hbab5e4f9),
	.w4(32'hbbf98460),
	.w5(32'hbc248b78),
	.w6(32'h3b9fc650),
	.w7(32'hbba0b699),
	.w8(32'hbc7cd07c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e8ebc),
	.w1(32'hbc4bba48),
	.w2(32'h3ba0a135),
	.w3(32'hbb99976f),
	.w4(32'h3bb6d854),
	.w5(32'h3c8639c7),
	.w6(32'hbbf5de81),
	.w7(32'h3c0f9b88),
	.w8(32'h3c875c0c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7553b8),
	.w1(32'hbc13de2f),
	.w2(32'h3c829342),
	.w3(32'hbb3a94b5),
	.w4(32'h3cb65816),
	.w5(32'h3bece94d),
	.w6(32'h3acdff9d),
	.w7(32'h3cefb1c2),
	.w8(32'h3b83858b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3c620),
	.w1(32'h3cbfa45c),
	.w2(32'h3c19e5af),
	.w3(32'h3c4374d5),
	.w4(32'h3af3320a),
	.w5(32'h3c032813),
	.w6(32'h3cecac4a),
	.w7(32'h3c1dd948),
	.w8(32'h39c58eb5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3816df),
	.w1(32'h3cd5474f),
	.w2(32'hbc432cc4),
	.w3(32'h3c7b25d7),
	.w4(32'hbbe30551),
	.w5(32'h3bb39626),
	.w6(32'hbb574593),
	.w7(32'hbc037ba5),
	.w8(32'h3d33ce0e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574494),
	.w1(32'hbc867d3f),
	.w2(32'h3cb38d4e),
	.w3(32'hbbe90000),
	.w4(32'hbc00e21c),
	.w5(32'h3c524962),
	.w6(32'h3c64d93c),
	.w7(32'h3b9b5730),
	.w8(32'h3d5288df),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1de040),
	.w1(32'hba304acb),
	.w2(32'hbba98813),
	.w3(32'hbab8b097),
	.w4(32'hbbcc48f4),
	.w5(32'h3bf7459f),
	.w6(32'h3d1692cc),
	.w7(32'h39a6c10d),
	.w8(32'h3d69d565),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c983aeb),
	.w1(32'hbc1ca385),
	.w2(32'h3b5ee5fc),
	.w3(32'hbaa8ed68),
	.w4(32'h3c56004a),
	.w5(32'hbaf94e0c),
	.w6(32'h3c86b5d4),
	.w7(32'h3c61a6b0),
	.w8(32'h3b81b06b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0377f7),
	.w1(32'h3be96ef6),
	.w2(32'h3c01ad89),
	.w3(32'hbae8aa0b),
	.w4(32'hbbbafa6b),
	.w5(32'hbbaa0acb),
	.w6(32'h3b142154),
	.w7(32'h3be45b8b),
	.w8(32'h3c2ec91c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b335c),
	.w1(32'hbca2451f),
	.w2(32'hbc60644c),
	.w3(32'hbc802abd),
	.w4(32'h3a728635),
	.w5(32'hbadb6c82),
	.w6(32'hbc21f11e),
	.w7(32'hbbb6c839),
	.w8(32'h3c568c44),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9fbbc),
	.w1(32'hbca224eb),
	.w2(32'h3c70f6e4),
	.w3(32'hbc559e0f),
	.w4(32'h3b990dc2),
	.w5(32'hbbdd5044),
	.w6(32'hbb94c2d8),
	.w7(32'h3c192a53),
	.w8(32'hbcad5e5d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9c865),
	.w1(32'h3c9df014),
	.w2(32'hbbad4bd3),
	.w3(32'h3ba4ddf3),
	.w4(32'hbc0cc894),
	.w5(32'h3b344f2e),
	.w6(32'hbc6ed35a),
	.w7(32'hbb0d2834),
	.w8(32'h3c8b8e3c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331f46),
	.w1(32'hbc86f527),
	.w2(32'hbc5a04b1),
	.w3(32'hb9dcbe98),
	.w4(32'hbb2a72d3),
	.w5(32'h3bedffee),
	.w6(32'h3bf487aa),
	.w7(32'hbbfe60f5),
	.w8(32'hbb844def),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdf9c4b),
	.w1(32'hbbfb1662),
	.w2(32'hbc68fed6),
	.w3(32'hbc9a2123),
	.w4(32'hbb64cab3),
	.w5(32'hb98ca3d6),
	.w6(32'hbb0d0266),
	.w7(32'hbbe5b8b1),
	.w8(32'hbba55ff5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93fa81),
	.w1(32'hbc60c130),
	.w2(32'h3a8432a2),
	.w3(32'h3967d61f),
	.w4(32'h3a00b5b1),
	.w5(32'h3b134a2e),
	.w6(32'hbc18135b),
	.w7(32'h39a6c65a),
	.w8(32'h3b34de37),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817084),
	.w1(32'h3b0fbdb5),
	.w2(32'hbbc178a8),
	.w3(32'h3ab1fa3f),
	.w4(32'hb9e097fe),
	.w5(32'h3a57922a),
	.w6(32'h3aa432f0),
	.w7(32'hbc8a5ca0),
	.w8(32'hbc84757c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a7312),
	.w1(32'hbc22226f),
	.w2(32'hbc26fbe7),
	.w3(32'hbb1fca68),
	.w4(32'h3b9c5f1a),
	.w5(32'hbc3fd668),
	.w6(32'hbc6e789c),
	.w7(32'hbaacae18),
	.w8(32'h3c1358a2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb73027),
	.w1(32'hbbeae938),
	.w2(32'h39b275a2),
	.w3(32'hbb2e0cc4),
	.w4(32'h3aa1fad7),
	.w5(32'hbc485450),
	.w6(32'h3b5fdc7e),
	.w7(32'h3af1632d),
	.w8(32'hbc47cdd1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8118eb),
	.w1(32'h3a47b841),
	.w2(32'hbb8f8d75),
	.w3(32'hbb94b7e1),
	.w4(32'h39b92823),
	.w5(32'h3aa90869),
	.w6(32'hbc118c88),
	.w7(32'hbac99523),
	.w8(32'h3c4a7d8c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76e40b),
	.w1(32'h3b8478af),
	.w2(32'hbb0f3d9d),
	.w3(32'h3b894864),
	.w4(32'hbb971006),
	.w5(32'h3bbd7d8c),
	.w6(32'h3baa7d58),
	.w7(32'hbc2a1fbc),
	.w8(32'h3cba1938),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5a289),
	.w1(32'hbacfd149),
	.w2(32'hbc063860),
	.w3(32'hbb8dd21a),
	.w4(32'hbb0494df),
	.w5(32'hbbfd9c47),
	.w6(32'h3c03b640),
	.w7(32'hbbc11f63),
	.w8(32'h3aa4f2dc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c637a7e),
	.w1(32'hbbbb040e),
	.w2(32'hbba4441d),
	.w3(32'hbc878b77),
	.w4(32'hbbc3546e),
	.w5(32'hbc3b8125),
	.w6(32'hbc092e46),
	.w7(32'hbb6b7165),
	.w8(32'hbc1c332a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc67b8fc),
	.w1(32'hbbbd99b2),
	.w2(32'h3bafc95c),
	.w3(32'hbc456dd7),
	.w4(32'h3b9ceb63),
	.w5(32'hbbd0a261),
	.w6(32'hbae2e14c),
	.w7(32'h3ae7a9c7),
	.w8(32'hbceec103),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ae777),
	.w1(32'h3b0e628e),
	.w2(32'hbb6f8885),
	.w3(32'h3b98a0ed),
	.w4(32'h3b017c3d),
	.w5(32'hbba3a93d),
	.w6(32'hbac10658),
	.w7(32'h3bb9597a),
	.w8(32'h3bf34406),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3325f),
	.w1(32'h3b53aea1),
	.w2(32'h3c3f1fa5),
	.w3(32'hbbf00cbf),
	.w4(32'hbbe010a5),
	.w5(32'h3ae88a76),
	.w6(32'h3a7eab1a),
	.w7(32'h39525b2b),
	.w8(32'hbc8a911e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2a66d),
	.w1(32'h3c95dd74),
	.w2(32'hbbdef720),
	.w3(32'h3c81ec50),
	.w4(32'hbb2fb582),
	.w5(32'h398c821a),
	.w6(32'h3bbf97b0),
	.w7(32'hbbce423f),
	.w8(32'h3c9a8d87),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe13e7),
	.w1(32'hbbeb2d99),
	.w2(32'hbc147997),
	.w3(32'hbaa9e5d6),
	.w4(32'hba11bcf7),
	.w5(32'h3b78ad5f),
	.w6(32'hbc9c3940),
	.w7(32'hbc091b18),
	.w8(32'h3aed9d5e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc548558),
	.w1(32'hbc7a1a8d),
	.w2(32'hbb161caa),
	.w3(32'hbc36337f),
	.w4(32'h3aefd768),
	.w5(32'h3ae7f766),
	.w6(32'hbb01e5b9),
	.w7(32'h3b56e99d),
	.w8(32'h3af1b310),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cd5d7),
	.w1(32'hbb04e06a),
	.w2(32'hbbc7cb90),
	.w3(32'hb9e9d977),
	.w4(32'hbc9bbfda),
	.w5(32'h3c4cb88f),
	.w6(32'h3ab9af2b),
	.w7(32'hbbefb9e4),
	.w8(32'hbb98e323),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3500),
	.w1(32'hbc21ff2a),
	.w2(32'hbc227c0b),
	.w3(32'hbbe4d0ba),
	.w4(32'hbae9c6b5),
	.w5(32'hbc8779b4),
	.w6(32'h3b95bf69),
	.w7(32'h3a33841f),
	.w8(32'h3b920c59),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bbcfd),
	.w1(32'hbc9c9e8e),
	.w2(32'hbc0a3720),
	.w3(32'hbc35d16c),
	.w4(32'hbbb85c7a),
	.w5(32'hb914ca59),
	.w6(32'hbc49ea9e),
	.w7(32'hbbc5c3ff),
	.w8(32'h3bda91ad),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2dac),
	.w1(32'hbb3cec14),
	.w2(32'h3c08cdfb),
	.w3(32'hbc2a0715),
	.w4(32'hbb56f3af),
	.w5(32'h3c6a38aa),
	.w6(32'hbbcddf8b),
	.w7(32'h3c3244ec),
	.w8(32'h3c8d744e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54e633),
	.w1(32'hbc53f988),
	.w2(32'h3c5d30bd),
	.w3(32'hbc3eb9e8),
	.w4(32'h3c11e44e),
	.w5(32'h3c1c44ef),
	.w6(32'hba1c394c),
	.w7(32'hba606e5b),
	.w8(32'h3ab88580),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb04d7),
	.w1(32'h3b910c75),
	.w2(32'h3c5d7f16),
	.w3(32'h3b2056bd),
	.w4(32'hbacf7dc9),
	.w5(32'h3ba831fc),
	.w6(32'hbaf4e82c),
	.w7(32'h3bb326a2),
	.w8(32'hbc731813),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cc1f3),
	.w1(32'h3ad4ce21),
	.w2(32'hbc5af5c9),
	.w3(32'hbbcd577c),
	.w4(32'hbb2ea6bd),
	.w5(32'hbc1d46ca),
	.w6(32'hbb0f12d9),
	.w7(32'hbb28486a),
	.w8(32'h3a4cc42d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f3d72),
	.w1(32'h3b6b6f39),
	.w2(32'hbbd9d54c),
	.w3(32'h3b1c9866),
	.w4(32'hba2aeb5d),
	.w5(32'hbb01fdf0),
	.w6(32'hbb927dc2),
	.w7(32'hbb87f492),
	.w8(32'h3cc9d46e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7a99),
	.w1(32'hbc22a01f),
	.w2(32'h3cc7b0f6),
	.w3(32'hbb80b80c),
	.w4(32'h3c6387e2),
	.w5(32'h3bd81d49),
	.w6(32'h3b0c9544),
	.w7(32'h3c933e7d),
	.w8(32'h3b761d76),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaf52c),
	.w1(32'h3a91e6f5),
	.w2(32'hbaf567bf),
	.w3(32'hbb3c99ac),
	.w4(32'hb9b67fa0),
	.w5(32'h3a84f9f2),
	.w6(32'hbb01bf99),
	.w7(32'h3a1fc509),
	.w8(32'h3a4f6272),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b117a2),
	.w1(32'hba34d276),
	.w2(32'hbc248fb1),
	.w3(32'hb9a27305),
	.w4(32'h3b7c2c1f),
	.w5(32'h3c0e5d22),
	.w6(32'h3aef371e),
	.w7(32'h3c151603),
	.w8(32'h3bf24d29),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3178a),
	.w1(32'h3b51c459),
	.w2(32'h3c3cfe50),
	.w3(32'hbb96b9bf),
	.w4(32'h3c2dc427),
	.w5(32'hbbb25f65),
	.w6(32'h3c1822d7),
	.w7(32'h3c3911c8),
	.w8(32'hbcb39caa),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a9ec5),
	.w1(32'hb8efdc22),
	.w2(32'hba2cf785),
	.w3(32'h3a022b02),
	.w4(32'hbc1f9539),
	.w5(32'hba12a385),
	.w6(32'h3a237cca),
	.w7(32'h3b00cea8),
	.w8(32'h3c0f9ef2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c333e1),
	.w1(32'hbb1ceb71),
	.w2(32'hbb6367d6),
	.w3(32'h3b1558e0),
	.w4(32'h3bd51ce7),
	.w5(32'h3a77bd27),
	.w6(32'h3b7067b9),
	.w7(32'h3ab6a3d7),
	.w8(32'h3c12ec30),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6172c3),
	.w1(32'hbc580309),
	.w2(32'hbb311fc1),
	.w3(32'hbb225920),
	.w4(32'h3adf12be),
	.w5(32'h39ccb390),
	.w6(32'h3a649df2),
	.w7(32'h3afc7c25),
	.w8(32'hba8ac297),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4837aa),
	.w1(32'hba887259),
	.w2(32'hbc08c16f),
	.w3(32'hba43e4f3),
	.w4(32'hbb755be6),
	.w5(32'hbc3070aa),
	.w6(32'h38d0c4bd),
	.w7(32'hbb8a9e25),
	.w8(32'hbbdb1663),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a3ab2),
	.w1(32'hbbd7ed13),
	.w2(32'h3a8d5986),
	.w3(32'hb911e46b),
	.w4(32'hbb2e474a),
	.w5(32'h3c476202),
	.w6(32'hbc710579),
	.w7(32'hbbee0e12),
	.w8(32'h38b1c7ac),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40a732),
	.w1(32'h3c2560fc),
	.w2(32'hbc00936f),
	.w3(32'h3b9a0dbd),
	.w4(32'h3babaf00),
	.w5(32'h3bc03be2),
	.w6(32'h38dc31d1),
	.w7(32'h3c006b7c),
	.w8(32'h3c95f1d0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910b05),
	.w1(32'h3c3f6c6f),
	.w2(32'h3c34b7e8),
	.w3(32'h399c9bae),
	.w4(32'h3b79f448),
	.w5(32'h3ccf27d8),
	.w6(32'h3c3d5015),
	.w7(32'h3cb45032),
	.w8(32'h3cde9b80),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ff1c8),
	.w1(32'h3c7f9836),
	.w2(32'h3a6cf691),
	.w3(32'hbb6248ef),
	.w4(32'h3c4acde4),
	.w5(32'h3b377800),
	.w6(32'h3cd0ec4d),
	.w7(32'h3c0237ef),
	.w8(32'hbaf3d3c5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule