module layer_8_featuremap_34(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00e00),
	.w1(32'h3a9dd83a),
	.w2(32'h3a210dd3),
	.w3(32'h39ade552),
	.w4(32'h3934de01),
	.w5(32'h39283495),
	.w6(32'h3a824b21),
	.w7(32'hb897f589),
	.w8(32'hba06d288),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83ca83f),
	.w1(32'h38ae1e78),
	.w2(32'h3944dbb2),
	.w3(32'hb910b021),
	.w4(32'h38646efd),
	.w5(32'h3919a0d4),
	.w6(32'hb896109d),
	.w7(32'h38d45b23),
	.w8(32'h3950c7e7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996d6c5),
	.w1(32'hb900d8a1),
	.w2(32'h38f6f19e),
	.w3(32'hb97ef317),
	.w4(32'hb92b4a04),
	.w5(32'h385115be),
	.w6(32'hb95837e3),
	.w7(32'h382d712a),
	.w8(32'h38c6b24f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881c2d),
	.w1(32'h3a6851f8),
	.w2(32'h39fadffd),
	.w3(32'h3a25b838),
	.w4(32'h3a8bcb3f),
	.w5(32'hb91999ca),
	.w6(32'hb8c7adc9),
	.w7(32'hb8ff58d0),
	.w8(32'h39570a03),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9618cf6),
	.w1(32'hb9715be8),
	.w2(32'hb87195d8),
	.w3(32'hb98af7d5),
	.w4(32'hb9bb20b4),
	.w5(32'hb93ae056),
	.w6(32'h36ce5b26),
	.w7(32'h38b528f8),
	.w8(32'h39566013),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46661e),
	.w1(32'hb8cf1e16),
	.w2(32'h3a285e37),
	.w3(32'hb8ce0ab4),
	.w4(32'h3970f1aa),
	.w5(32'h3a2cbbc7),
	.w6(32'hb95f83f5),
	.w7(32'h3a2ebe2f),
	.w8(32'h3b0b8f22),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f351aa),
	.w1(32'h36da766f),
	.w2(32'h368b22d3),
	.w3(32'hb5a073ea),
	.w4(32'h367a8f3c),
	.w5(32'hb455032c),
	.w6(32'hb7041b94),
	.w7(32'hb6d170bc),
	.w8(32'hb712303a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6272b5),
	.w1(32'h3a57ad52),
	.w2(32'h39ff24c4),
	.w3(32'h39a052ab),
	.w4(32'h3a82be77),
	.w5(32'h39ed4bac),
	.w6(32'h3953068d),
	.w7(32'h39f79f72),
	.w8(32'h385e6f05),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4b3dc),
	.w1(32'hb8e6d9fc),
	.w2(32'h38e2e4d1),
	.w3(32'hb96d36f6),
	.w4(32'hb966fd18),
	.w5(32'hb9588fc4),
	.w6(32'hb9db3212),
	.w7(32'hb96b02f3),
	.w8(32'h37438e97),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b30b2),
	.w1(32'h3abf87f2),
	.w2(32'h3a570a72),
	.w3(32'h39b96ba9),
	.w4(32'h3a33df2f),
	.w5(32'h3a346f92),
	.w6(32'h3a8b2386),
	.w7(32'h3a5dfac9),
	.w8(32'h39d1987a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9708c3),
	.w1(32'h3a33444d),
	.w2(32'h395c6559),
	.w3(32'h39d50264),
	.w4(32'h3a3fce34),
	.w5(32'h391c5067),
	.w6(32'h3985b132),
	.w7(32'hb9fbd76b),
	.w8(32'hb9b52ef4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad38ed),
	.w1(32'h3a894fb9),
	.w2(32'h3a2b7751),
	.w3(32'h3a206734),
	.w4(32'h3a282809),
	.w5(32'h395b744c),
	.w6(32'h3a720fd2),
	.w7(32'hb9afa5ed),
	.w8(32'hb9664716),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cca37a),
	.w1(32'h3905139c),
	.w2(32'h39a5371e),
	.w3(32'h38418bdc),
	.w4(32'h37939abc),
	.w5(32'h38cf5625),
	.w6(32'h39fe06e1),
	.w7(32'h3a25d029),
	.w8(32'h3a3127d3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5134fce),
	.w1(32'h36410b1c),
	.w2(32'h361fbe69),
	.w3(32'hb6411ffc),
	.w4(32'h35baeaa4),
	.w5(32'hb55350f0),
	.w6(32'hb736885d),
	.w7(32'hb6d40865),
	.w8(32'hb6ed8400),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f2ffc7),
	.w1(32'h359e0db9),
	.w2(32'h361fae07),
	.w3(32'hb60ac491),
	.w4(32'h359442d5),
	.w5(32'h35913eb5),
	.w6(32'hb70ae3b7),
	.w7(32'hb6a496e9),
	.w8(32'hb69939c0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377a5921),
	.w1(32'hb578fb15),
	.w2(32'h379e031a),
	.w3(32'hb6bbe0e2),
	.w4(32'h34e2cfe4),
	.w5(32'h36b82b86),
	.w6(32'hb717a24c),
	.w7(32'hb6206d75),
	.w8(32'h36bcb1b6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7da31),
	.w1(32'h39cd4d5e),
	.w2(32'h39edc0b7),
	.w3(32'hb84d72dc),
	.w4(32'h38c59381),
	.w5(32'h3a168cec),
	.w6(32'h3838fc66),
	.w7(32'h396dbdb2),
	.w8(32'h399ef654),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2070a0),
	.w1(32'h3a81e8ef),
	.w2(32'h3a0111f0),
	.w3(32'h39f4a009),
	.w4(32'h39e7696c),
	.w5(32'h3a4d463d),
	.w6(32'h3a5bc0fc),
	.w7(32'h3a42e0e9),
	.w8(32'h3a1ace56),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943278),
	.w1(32'h3b556638),
	.w2(32'h3acca08d),
	.w3(32'h39137397),
	.w4(32'h3b460dcd),
	.w5(32'h3a8a83ad),
	.w6(32'h3aeaa473),
	.w7(32'hba6c5b8e),
	.w8(32'hbad95518),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94daee5),
	.w1(32'hb9fc78d5),
	.w2(32'hb9eb839a),
	.w3(32'h39841b75),
	.w4(32'hba823c23),
	.w5(32'hba951b12),
	.w6(32'h3af94933),
	.w7(32'h3a8d45cc),
	.w8(32'h39c010b5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d40d30),
	.w1(32'h39ed9c67),
	.w2(32'h3a885b09),
	.w3(32'hb9f138f9),
	.w4(32'hba2ffce4),
	.w5(32'h39c11715),
	.w6(32'h39fabc58),
	.w7(32'hb72a8c22),
	.w8(32'h3a327d03),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abf6fa),
	.w1(32'hb8f4c0ba),
	.w2(32'h399a37e2),
	.w3(32'hb92fa733),
	.w4(32'hb6bb25cc),
	.w5(32'h391a3a03),
	.w6(32'h38123c5c),
	.w7(32'h39c8845d),
	.w8(32'h3a042f46),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ea950),
	.w1(32'h3b2a4121),
	.w2(32'h3ad0f6ec),
	.w3(32'h3964fddd),
	.w4(32'h3af061ad),
	.w5(32'h39dd8012),
	.w6(32'h3aef8b00),
	.w7(32'hb98461bd),
	.w8(32'hba8c7c0c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38879b06),
	.w1(32'hb7795da6),
	.w2(32'h38a492cb),
	.w3(32'h3984562f),
	.w4(32'hb9814033),
	.w5(32'hb95bd226),
	.w6(32'h39c9c7f0),
	.w7(32'h3918a1b3),
	.w8(32'h39cf2fab),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d7efab),
	.w1(32'h36f65f5b),
	.w2(32'h36f40ebf),
	.w3(32'h3720cab8),
	.w4(32'h37426606),
	.w5(32'h37a3f791),
	.w6(32'hb6c14941),
	.w7(32'h374ab48d),
	.w8(32'h3782fa7f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa97840),
	.w1(32'h3a4373cc),
	.w2(32'h399fe6b0),
	.w3(32'h3a4f7467),
	.w4(32'h38e45bc8),
	.w5(32'h390d46e2),
	.w6(32'h3a8d4296),
	.w7(32'hb9236aaa),
	.w8(32'hb96c5e8d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b44b37),
	.w1(32'h36af7d82),
	.w2(32'h368a7aff),
	.w3(32'hb627b1dc),
	.w4(32'h36315a38),
	.w5(32'hb57c7d6c),
	.w6(32'hb6fcd341),
	.w7(32'hb50cd992),
	.w8(32'hb600032f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c275782),
	.w1(32'h3c041d6d),
	.w2(32'h3bb794fa),
	.w3(32'h3b0b9e46),
	.w4(32'h3bdafda0),
	.w5(32'h3c042111),
	.w6(32'h3bbb5f2d),
	.w7(32'h39b1633d),
	.w8(32'h3b0c427c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5785ec),
	.w1(32'h3a3dc69a),
	.w2(32'h39d7617a),
	.w3(32'h39bf00c4),
	.w4(32'h395c35a5),
	.w5(32'hb916e080),
	.w6(32'h3a062437),
	.w7(32'h384970b3),
	.w8(32'hb9272c6d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84dc20f),
	.w1(32'h37602246),
	.w2(32'h38e9204f),
	.w3(32'hb89f23aa),
	.w4(32'h37c4a178),
	.w5(32'h38632adf),
	.w6(32'h36491582),
	.w7(32'h3931e42e),
	.w8(32'h39700276),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84ccd52),
	.w1(32'h394bf4af),
	.w2(32'h37bf0d35),
	.w3(32'hb5cde35f),
	.w4(32'h39a81eec),
	.w5(32'h385c4255),
	.w6(32'h38cb2504),
	.w7(32'h399b39c6),
	.w8(32'h38eb99a5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3897d61b),
	.w1(32'h389070a2),
	.w2(32'h3982766a),
	.w3(32'hb8e755b7),
	.w4(32'hb9bda237),
	.w5(32'hb817269a),
	.w6(32'h3888dcb3),
	.w7(32'h3837767c),
	.w8(32'h39ae6f06),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37212dcc),
	.w1(32'h375f2f65),
	.w2(32'h37199681),
	.w3(32'hb77bd0eb),
	.w4(32'hb6dd424f),
	.w5(32'hb7139a5b),
	.w6(32'hb7702311),
	.w7(32'hb7513539),
	.w8(32'hb7792566),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b81c2e),
	.w1(32'h3660b111),
	.w2(32'hb39d0130),
	.w3(32'hb54e53bd),
	.w4(32'hb5b1580c),
	.w5(32'hb68ae620),
	.w6(32'hb6ac9b78),
	.w7(32'hb6fa55d5),
	.w8(32'hb7982fae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcfeba),
	.w1(32'hb793be30),
	.w2(32'hb92ab2ed),
	.w3(32'hb95c2812),
	.w4(32'hb8f4f57f),
	.w5(32'hb90ff1f3),
	.w6(32'h3a4a7395),
	.w7(32'h3a89580b),
	.w8(32'h3a37f56e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91d583),
	.w1(32'h3a8c45cc),
	.w2(32'h3a53cac8),
	.w3(32'h38a42ce0),
	.w4(32'h3a28d5ed),
	.w5(32'h39e926a4),
	.w6(32'h3a600514),
	.w7(32'h383e8a5b),
	.w8(32'hb9171ecd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37012a64),
	.w1(32'h3730a1ab),
	.w2(32'hb25cea62),
	.w3(32'hb64eff9f),
	.w4(32'h36a073c4),
	.w5(32'h361a0081),
	.w6(32'hb62de682),
	.w7(32'h36e6cf85),
	.w8(32'hb6e3328a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97502eb),
	.w1(32'h378c9d75),
	.w2(32'h38da66c6),
	.w3(32'hb91ed8c3),
	.w4(32'h38f1116e),
	.w5(32'h38d55e8b),
	.w6(32'hb9b2520f),
	.w7(32'hb80cc139),
	.w8(32'h3924a613),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f77a26),
	.w1(32'hb69fc973),
	.w2(32'hb59f693b),
	.w3(32'hb6b8da2a),
	.w4(32'hb686593f),
	.w5(32'hb6616043),
	.w6(32'hb771ec82),
	.w7(32'hb6f822f7),
	.w8(32'hb6f34a08),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3555e756),
	.w1(32'hb74b1b62),
	.w2(32'hb6cbd1a9),
	.w3(32'h37321c86),
	.w4(32'h37d01b8b),
	.w5(32'h371b5993),
	.w6(32'hb6a967c0),
	.w7(32'hb726db3d),
	.w8(32'hb722902b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9416b1),
	.w1(32'h3b733609),
	.w2(32'h3a82c3cb),
	.w3(32'h3b53a463),
	.w4(32'h3b0ead42),
	.w5(32'h39a31a4a),
	.w6(32'h3b68f707),
	.w7(32'h3a33120d),
	.w8(32'hbb85f58e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ec5e9),
	.w1(32'h3acaff2c),
	.w2(32'h3a1977b8),
	.w3(32'hbc063746),
	.w4(32'h3b1285a9),
	.w5(32'hbbad560d),
	.w6(32'hbc0550b9),
	.w7(32'hbb7c04c5),
	.w8(32'h3c10dd21),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f75d2),
	.w1(32'hbb40b53c),
	.w2(32'h3cb5e83e),
	.w3(32'hbbffcd22),
	.w4(32'hbca7160c),
	.w5(32'h3ceca54f),
	.w6(32'h3d191427),
	.w7(32'hbbb0b7b6),
	.w8(32'hbbe6440e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eddb25),
	.w1(32'h3a3c3f59),
	.w2(32'hb9a1a80c),
	.w3(32'h3b5fc50e),
	.w4(32'h3c806039),
	.w5(32'h3b3562d1),
	.w6(32'hbc763215),
	.w7(32'hbbbb74e6),
	.w8(32'hbbfc2832),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdadbd4),
	.w1(32'h3b4036c1),
	.w2(32'h3b813f51),
	.w3(32'h3c3752a6),
	.w4(32'h3cab2526),
	.w5(32'h3c2bad43),
	.w6(32'hbc9d22c7),
	.w7(32'hbc2792a4),
	.w8(32'h39033169),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ea287),
	.w1(32'hbc0319dd),
	.w2(32'hbc097ee4),
	.w3(32'hbb8856b3),
	.w4(32'h3b8f21bd),
	.w5(32'h3b0b959c),
	.w6(32'hbc639c37),
	.w7(32'hbc5659a0),
	.w8(32'hbc3e0209),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11c4d7),
	.w1(32'hb9a7ac67),
	.w2(32'hbc9479cd),
	.w3(32'hbc8f231e),
	.w4(32'h3c3232c4),
	.w5(32'h3a7e7c0a),
	.w6(32'h3c05360a),
	.w7(32'h39e42387),
	.w8(32'hbc8d2d22),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e2e9e),
	.w1(32'hbb8f8201),
	.w2(32'h3ab2b8ff),
	.w3(32'hbc526edd),
	.w4(32'h3c53a03e),
	.w5(32'h3bcb7996),
	.w6(32'hbcd1afd4),
	.w7(32'hbbf2d8bc),
	.w8(32'h3cd18bc0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6b291),
	.w1(32'h3b32899c),
	.w2(32'hbc110ac0),
	.w3(32'hbca48a68),
	.w4(32'hbd2857eb),
	.w5(32'hbd03c926),
	.w6(32'h3d4f2dd3),
	.w7(32'h3cc3cebb),
	.w8(32'hbbe42e84),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d782),
	.w1(32'hbb3ef7fb),
	.w2(32'hbab294b4),
	.w3(32'h3c0225ee),
	.w4(32'h3cabf333),
	.w5(32'h3c2a098b),
	.w6(32'hbcb0dece),
	.w7(32'hbc59154d),
	.w8(32'hbba59dfe),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1fa82),
	.w1(32'hbab4e868),
	.w2(32'h3aad3697),
	.w3(32'h3b7c38da),
	.w4(32'h3be099f0),
	.w5(32'h3b881dfb),
	.w6(32'hbc20edee),
	.w7(32'hbb84231d),
	.w8(32'hbc2d979c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3081dc),
	.w1(32'h3aeb6d99),
	.w2(32'h3b31ec4e),
	.w3(32'h3bb328a2),
	.w4(32'h3c99e97e),
	.w5(32'h3bb3d75d),
	.w6(32'hbcbc599d),
	.w7(32'hbc148cd8),
	.w8(32'hbc27461e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb12b0),
	.w1(32'hbc951861),
	.w2(32'hb99def5e),
	.w3(32'h3bfa2f7a),
	.w4(32'hbc1d02d5),
	.w5(32'hbca6575d),
	.w6(32'h3aed6bfc),
	.w7(32'h3c2b05a1),
	.w8(32'h3b027024),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df10c),
	.w1(32'h3ae6a304),
	.w2(32'hbac6a010),
	.w3(32'h3af3b10a),
	.w4(32'hbc2da951),
	.w5(32'hbb89aa47),
	.w6(32'h3c286c3a),
	.w7(32'h399760d3),
	.w8(32'h3ccdbede),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9b60d),
	.w1(32'hbbfbb32f),
	.w2(32'hbbb2c80e),
	.w3(32'hbbcf4bd3),
	.w4(32'h3c7bf9c9),
	.w5(32'h3cc3a9b0),
	.w6(32'h3c0d510c),
	.w7(32'hbc43349f),
	.w8(32'h3b1bf026),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2b3d0),
	.w1(32'h3b272ff0),
	.w2(32'h3bb9f604),
	.w3(32'h3beff1fd),
	.w4(32'h3b711eab),
	.w5(32'hbbc70c66),
	.w6(32'hbc29400c),
	.w7(32'h3c3365d2),
	.w8(32'hb8a8245d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5fa72c),
	.w1(32'h3bbe8c99),
	.w2(32'hbb84c4a1),
	.w3(32'h3bb89c6b),
	.w4(32'h3bca708e),
	.w5(32'hbb8e1f1f),
	.w6(32'hbb4ec10e),
	.w7(32'h3a59384c),
	.w8(32'h3af06218),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc6870),
	.w1(32'hbbd20a68),
	.w2(32'h3bf32ce2),
	.w3(32'hbb087e97),
	.w4(32'hbbc63c82),
	.w5(32'h3c530079),
	.w6(32'hbc8e413f),
	.w7(32'h3b24d589),
	.w8(32'h3b961ecb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01681),
	.w1(32'h3b411f4e),
	.w2(32'hbba31b8f),
	.w3(32'hb721f121),
	.w4(32'h3c42e5df),
	.w5(32'hbb506c07),
	.w6(32'h3c141502),
	.w7(32'h3b79e865),
	.w8(32'hbbfd5c06),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c5c6b),
	.w1(32'hbb2623ad),
	.w2(32'hb9bdcd0a),
	.w3(32'h3b843a8c),
	.w4(32'hbbd078a9),
	.w5(32'h3c231ced),
	.w6(32'hbb010b63),
	.w7(32'hbbf9a2ab),
	.w8(32'hbba8bfc5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb30a8),
	.w1(32'h3b878301),
	.w2(32'hbc47688e),
	.w3(32'hbb9dfb38),
	.w4(32'hbb858eb2),
	.w5(32'h3c5865c8),
	.w6(32'h3c822992),
	.w7(32'hbc481403),
	.w8(32'hbc0501cf),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ecec5),
	.w1(32'hbc3c2ee7),
	.w2(32'hbc957c55),
	.w3(32'hbc5a6beb),
	.w4(32'h3b45b571),
	.w5(32'hbbbb9d4a),
	.w6(32'hbca086ef),
	.w7(32'hbc3e8a96),
	.w8(32'hbc06670a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ddb72),
	.w1(32'h3b0f34a5),
	.w2(32'h3721023c),
	.w3(32'h3caa2c8c),
	.w4(32'h3cceeb21),
	.w5(32'h3c82b76e),
	.w6(32'hbc7eecfc),
	.w7(32'hbc559085),
	.w8(32'h3b638ee4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23eb4e),
	.w1(32'h3b255833),
	.w2(32'hbb624a45),
	.w3(32'hbc1fe9a2),
	.w4(32'hbc2ce267),
	.w5(32'hbc76861a),
	.w6(32'hbc8b705f),
	.w7(32'hbce09669),
	.w8(32'hbb73ba3e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafc01d),
	.w1(32'h38ac6faa),
	.w2(32'hb939b361),
	.w3(32'h3bb8dbff),
	.w4(32'h3c3eeb7b),
	.w5(32'h3a866992),
	.w6(32'hbc39d74d),
	.w7(32'hbb8f41b2),
	.w8(32'hbb4d79ea),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b065cc7),
	.w1(32'h3b2004d6),
	.w2(32'h3b0e1759),
	.w3(32'h3b1cacce),
	.w4(32'h3c10d0f5),
	.w5(32'h3ae5e73c),
	.w6(32'hbbe7ef96),
	.w7(32'hbb1f4fdd),
	.w8(32'hbb8690b7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38753391),
	.w1(32'hb9034e53),
	.w2(32'h3ac3aafc),
	.w3(32'h3b1272d7),
	.w4(32'h3b7c0a2c),
	.w5(32'h3ad33a4e),
	.w6(32'hbbfa11a4),
	.w7(32'hbb6eb115),
	.w8(32'h3b984296),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf499d8),
	.w1(32'h3a08551d),
	.w2(32'hbbd01a72),
	.w3(32'hbcae1c9f),
	.w4(32'h3b7c6fee),
	.w5(32'hbc21c348),
	.w6(32'hbb759d9a),
	.w7(32'hbbe22be8),
	.w8(32'hbbaf07df),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b4882),
	.w1(32'hbb26a640),
	.w2(32'h3983b6fe),
	.w3(32'h3bd61160),
	.w4(32'h3c5bffb9),
	.w5(32'h3c07e2a9),
	.w6(32'hbc8ddd00),
	.w7(32'hbc34e0f7),
	.w8(32'hbcc11049),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a2fc9),
	.w1(32'h3a8cac66),
	.w2(32'h3a721b38),
	.w3(32'h3cb193ea),
	.w4(32'h3d85cc13),
	.w5(32'h3d069198),
	.w6(32'hbd23c346),
	.w7(32'hbca047b5),
	.w8(32'hbb3954a4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11aef7),
	.w1(32'h3b019e32),
	.w2(32'h3abe74ce),
	.w3(32'hba260ed6),
	.w4(32'h3bc25897),
	.w5(32'hba9559cf),
	.w6(32'hbbfd5c0a),
	.w7(32'hbb82c78a),
	.w8(32'hbbb2bec5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3af4c4),
	.w1(32'hbb968795),
	.w2(32'hb9bb2316),
	.w3(32'h3bc54172),
	.w4(32'h3c881ff0),
	.w5(32'h3c311690),
	.w6(32'hbc9ea229),
	.w7(32'hbc46679f),
	.w8(32'hbb58d4e3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952630),
	.w1(32'h3b3a5e88),
	.w2(32'h3b3d5c0d),
	.w3(32'h3b32ccee),
	.w4(32'h3c1e319c),
	.w5(32'h3af65123),
	.w6(32'hbc4e8796),
	.w7(32'hbbc6b2e0),
	.w8(32'hbad0de40),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc94043),
	.w1(32'hbb18f2f4),
	.w2(32'hbc5c3dc7),
	.w3(32'hbc3e377e),
	.w4(32'h3b535873),
	.w5(32'hbc49a04f),
	.w6(32'hbace56bc),
	.w7(32'hbc4077b6),
	.w8(32'hbc0f14dc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77e546),
	.w1(32'hbb8a22a2),
	.w2(32'hbb7a4991),
	.w3(32'hbb22c84f),
	.w4(32'h3abb4c59),
	.w5(32'hbb193de1),
	.w6(32'hbcaa02c7),
	.w7(32'hbc8c7279),
	.w8(32'hbb8a5f6b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f16c53),
	.w1(32'hba5361da),
	.w2(32'h38f701f2),
	.w3(32'h3ac72895),
	.w4(32'h3c026aff),
	.w5(32'h3a7f716c),
	.w6(32'hbc2ec199),
	.w7(32'hbb92bf3f),
	.w8(32'hbbc4193f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5f86),
	.w1(32'hbb05ab81),
	.w2(32'hbb4299be),
	.w3(32'hbbd585e0),
	.w4(32'h3b214a46),
	.w5(32'hbbb26f9e),
	.w6(32'hbc4afde2),
	.w7(32'hbbfd25d4),
	.w8(32'hbccae0cf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f0102),
	.w1(32'h3a5c5ad6),
	.w2(32'hba7c3324),
	.w3(32'h3cbcdc36),
	.w4(32'h3d90f824),
	.w5(32'h3d03f9bf),
	.w6(32'hbd2cb1d3),
	.w7(32'hbcad7fc8),
	.w8(32'hbc8a8bbc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7aa2),
	.w1(32'hbb09750c),
	.w2(32'hb97a60b0),
	.w3(32'h3c64b4c8),
	.w4(32'h3d2d5504),
	.w5(32'h3cbf2cbd),
	.w6(32'hbd086e19),
	.w7(32'hbc73deed),
	.w8(32'hbbadfdf3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ef9a3),
	.w1(32'h3b8586a6),
	.w2(32'h3a5cf6c5),
	.w3(32'h3b6fc1f1),
	.w4(32'h3c2b184c),
	.w5(32'hbb0b038b),
	.w6(32'hbc156048),
	.w7(32'hba411118),
	.w8(32'hbc33ece7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf8d43),
	.w1(32'hb958ff74),
	.w2(32'hbc633730),
	.w3(32'h3b800a11),
	.w4(32'hbbea7ba2),
	.w5(32'hbb9fd25a),
	.w6(32'hbbe039c9),
	.w7(32'hbcb19f64),
	.w8(32'hbbfb51c2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb4713),
	.w1(32'hbbe2052b),
	.w2(32'hbbd99711),
	.w3(32'hbbdc128e),
	.w4(32'hbaaabed0),
	.w5(32'hbb74da4b),
	.w6(32'hbc6725e9),
	.w7(32'hbc0cb58a),
	.w8(32'hbb9a0dce),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab79b7a),
	.w1(32'h3a794ccd),
	.w2(32'hba277940),
	.w3(32'h3c145fd9),
	.w4(32'h3cd31652),
	.w5(32'h3bc1b1df),
	.w6(32'hbcc9b728),
	.w7(32'hbc431eb9),
	.w8(32'hbc7d13e7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf2c5),
	.w1(32'h3b79c9a4),
	.w2(32'h3b0c74ea),
	.w3(32'hbbc8c09a),
	.w4(32'hbc97b6e8),
	.w5(32'hbc933065),
	.w6(32'hbc77bddf),
	.w7(32'h3c643b70),
	.w8(32'hbbed0573),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aeee50),
	.w1(32'hba3c3abd),
	.w2(32'hb91b378a),
	.w3(32'h3b560ab7),
	.w4(32'hbb33c445),
	.w5(32'h3b4198f8),
	.w6(32'hbb3b3717),
	.w7(32'hbb87e421),
	.w8(32'hbc2f7482),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93900d),
	.w1(32'hb7b7cbaa),
	.w2(32'h38bf07fb),
	.w3(32'h3c1b2b52),
	.w4(32'h3c9a9846),
	.w5(32'h3c27fecb),
	.w6(32'hbcb6c189),
	.w7(32'hbc69214d),
	.w8(32'h3d0ee06a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176ff8),
	.w1(32'h3b6cda53),
	.w2(32'hbc4237a8),
	.w3(32'hbcd9361a),
	.w4(32'hbd5e5f4d),
	.w5(32'hbd2eb384),
	.w6(32'h3d88ad4e),
	.w7(32'h3d0142b3),
	.w8(32'hba7e5313),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b8f54),
	.w1(32'hbb335858),
	.w2(32'h3a775ba3),
	.w3(32'h3bb196f2),
	.w4(32'h3ca41455),
	.w5(32'h3c0e9d73),
	.w6(32'hbc89c632),
	.w7(32'hbbc143df),
	.w8(32'hbc84ef9a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0736d1),
	.w1(32'h3a37cd23),
	.w2(32'hbbcd9b8d),
	.w3(32'h3b45815d),
	.w4(32'hba1f5e1e),
	.w5(32'h3b83f72e),
	.w6(32'hbc05cf4e),
	.w7(32'hbca2b730),
	.w8(32'h3d056712),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160e14),
	.w1(32'h3b5f9289),
	.w2(32'hbc3457d7),
	.w3(32'hbccae1d2),
	.w4(32'hbd5040d8),
	.w5(32'hbd237e67),
	.w6(32'h3d8006ec),
	.w7(32'h3cf1e829),
	.w8(32'h3ce4b08b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2aa95a),
	.w1(32'h3b618dd5),
	.w2(32'hbc1521f9),
	.w3(32'hbcaabb0d),
	.w4(32'hbd31898e),
	.w5(32'hbd0af9a5),
	.w6(32'h3d5c79a9),
	.w7(32'h3ccff72a),
	.w8(32'hbbf74e07),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e9b1a),
	.w1(32'hbb5bdc3b),
	.w2(32'hbb5232da),
	.w3(32'h39899be2),
	.w4(32'hbc0f825e),
	.w5(32'hb90acc02),
	.w6(32'hbb172bb2),
	.w7(32'hbbd64ac9),
	.w8(32'hbb2735e6),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eda07),
	.w1(32'hbc03c0ba),
	.w2(32'h3c397484),
	.w3(32'h3c48eafb),
	.w4(32'h3caa0d3c),
	.w5(32'hbca27076),
	.w6(32'hbc76b8ad),
	.w7(32'h3d0b3c51),
	.w8(32'hbb515d2d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9680505),
	.w1(32'hb8e870d2),
	.w2(32'h3a42ff5d),
	.w3(32'h3ad57911),
	.w4(32'h3ba6a59f),
	.w5(32'h3aeda340),
	.w6(32'hbbf49bcc),
	.w7(32'hbb66f4da),
	.w8(32'hbbf7a294),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd402e7),
	.w1(32'h3c4a1a51),
	.w2(32'hbcb2e571),
	.w3(32'hbca3bec8),
	.w4(32'hbc3394e2),
	.w5(32'hbc8c313e),
	.w6(32'hbb6298c2),
	.w7(32'hbb2a9da7),
	.w8(32'hbcfcfc05),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1acd07),
	.w1(32'hbb8073df),
	.w2(32'hbbe745c7),
	.w3(32'h3b5227fe),
	.w4(32'hbc01f215),
	.w5(32'h3ba7721c),
	.w6(32'hbca19c7f),
	.w7(32'hbce7901e),
	.w8(32'hb691e414),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba1ed7),
	.w1(32'hbc05974e),
	.w2(32'hbcb78187),
	.w3(32'hbd01d13c),
	.w4(32'h3b57519b),
	.w5(32'hbb9e93fc),
	.w6(32'hbaeb1883),
	.w7(32'hbb81bbdf),
	.w8(32'hbb86abb7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11f144),
	.w1(32'h3ba8ca9d),
	.w2(32'h3aefa1b9),
	.w3(32'hbb3424f8),
	.w4(32'hbb9779c6),
	.w5(32'hbbf392d1),
	.w6(32'h3bc5d969),
	.w7(32'hbbc8196b),
	.w8(32'hbcb28d9d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52a55e),
	.w1(32'hb9bb5e7a),
	.w2(32'hba9af90b),
	.w3(32'h3ca3b153),
	.w4(32'h3d7ccf03),
	.w5(32'h3ce75efa),
	.w6(32'hbd1bf181),
	.w7(32'hbc961876),
	.w8(32'hba621337),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf89d0),
	.w1(32'h3b0fa834),
	.w2(32'h3a63d0ae),
	.w3(32'h3b2da887),
	.w4(32'h3c8b69de),
	.w5(32'h3b97ef52),
	.w6(32'hbc7a4752),
	.w7(32'hbbb311b3),
	.w8(32'hbbf6408d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22d9e4),
	.w1(32'hbb9afe3e),
	.w2(32'hbbc71c67),
	.w3(32'h3ba86d56),
	.w4(32'hbc179f99),
	.w5(32'h3be65f27),
	.w6(32'hbb8c3312),
	.w7(32'hbc896b66),
	.w8(32'hbbcdaea7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdfbb0),
	.w1(32'hbb23aad7),
	.w2(32'h3af1a790),
	.w3(32'h3b5e1ecc),
	.w4(32'h3bc9a8a4),
	.w5(32'h3b9682c9),
	.w6(32'hbc49ee7b),
	.w7(32'hbbb718e7),
	.w8(32'hbcec95cd),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6fd261),
	.w1(32'hbc3e72c4),
	.w2(32'hbb8ac04b),
	.w3(32'h3cc06cdf),
	.w4(32'h3d9c7a2b),
	.w5(32'h3d3883a2),
	.w6(32'hbd8cea45),
	.w7(32'hbcfea5d7),
	.w8(32'hbc2afbcb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5336d),
	.w1(32'hba8a50eb),
	.w2(32'hbb385dd9),
	.w3(32'hb992fffd),
	.w4(32'hbbd0b208),
	.w5(32'h3b203720),
	.w6(32'hbb6b37d7),
	.w7(32'hbc329510),
	.w8(32'h3c6224b9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89ba5c),
	.w1(32'h3aa5ac45),
	.w2(32'hbb8b2d4d),
	.w3(32'hbc27d07c),
	.w4(32'hbcafd2fe),
	.w5(32'hbc84cb02),
	.w6(32'h3ccf0e1f),
	.w7(32'h3c46565b),
	.w8(32'h3908839c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac58cd3),
	.w1(32'h3adcb08d),
	.w2(32'h3aba4a77),
	.w3(32'hba0c7bb8),
	.w4(32'h39adabc5),
	.w5(32'h3a658dee),
	.w6(32'h39d0a734),
	.w7(32'hb828f9cf),
	.w8(32'hba33972d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8d9f6),
	.w1(32'hba718a5e),
	.w2(32'h3af3422e),
	.w3(32'h39d27481),
	.w4(32'h3b3369e2),
	.w5(32'hb993c2bd),
	.w6(32'hbab6ed26),
	.w7(32'h38718c77),
	.w8(32'hb99dc483),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02456d),
	.w1(32'hba123087),
	.w2(32'hb95b6653),
	.w3(32'hba28dd03),
	.w4(32'hbaa9bf74),
	.w5(32'hba11215b),
	.w6(32'h38ef02dc),
	.w7(32'hb90bd220),
	.w8(32'h3a0d12da),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396be486),
	.w1(32'h39fba596),
	.w2(32'h3a9aad99),
	.w3(32'h394bfb0d),
	.w4(32'h39f7a5ca),
	.w5(32'h3aa41fc6),
	.w6(32'hb9332a1a),
	.w7(32'h39e2085c),
	.w8(32'h39ae1e95),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fc705),
	.w1(32'h3b14eb21),
	.w2(32'h3addee8e),
	.w3(32'hbaa47d69),
	.w4(32'hbaa01494),
	.w5(32'hb804aba7),
	.w6(32'h3a0fd374),
	.w7(32'h3a0d5681),
	.w8(32'h3b3e63d8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c9be0),
	.w1(32'hbb2d4a88),
	.w2(32'hbbcf0d17),
	.w3(32'hb9f61574),
	.w4(32'hbb987cc4),
	.w5(32'hbb4aebd8),
	.w6(32'h3b68da45),
	.w7(32'h39ef10fc),
	.w8(32'hb98e88c1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b8d33),
	.w1(32'h39412a2e),
	.w2(32'h3b8295d0),
	.w3(32'hbb20d10b),
	.w4(32'hbb16c9cd),
	.w5(32'h3a4a1a64),
	.w6(32'h3a21f302),
	.w7(32'h3b09350b),
	.w8(32'h399ae16d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2efb0c),
	.w1(32'hb9a934bd),
	.w2(32'hb81b8f2e),
	.w3(32'hb9ed80dc),
	.w4(32'h392fdb82),
	.w5(32'hb98145f0),
	.w6(32'hb9665def),
	.w7(32'h3a27e722),
	.w8(32'h39c21ac3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a36743d),
	.w1(32'h3a70c702),
	.w2(32'h3a8fa6f4),
	.w3(32'hb9dc48a1),
	.w4(32'hb9addfa5),
	.w5(32'h3a2f6378),
	.w6(32'h3943922d),
	.w7(32'h380ec2bd),
	.w8(32'hba0b808f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30759a),
	.w1(32'hb9e4fa55),
	.w2(32'hb8c3a346),
	.w3(32'hba7fee9a),
	.w4(32'hba33b205),
	.w5(32'hba00cce6),
	.w6(32'hb95bbb8a),
	.w7(32'hb9157e2c),
	.w8(32'hba38dc9c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84a6c4),
	.w1(32'hba8c6180),
	.w2(32'hba507ae3),
	.w3(32'hbad982fa),
	.w4(32'hbb0b0c35),
	.w5(32'hbacf131c),
	.w6(32'hba4c2b04),
	.w7(32'hba42163d),
	.w8(32'hbb0d4b8c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa741b7),
	.w1(32'h3bc7a896),
	.w2(32'hbb0bf2cc),
	.w3(32'hba627eb0),
	.w4(32'h3c0270ec),
	.w5(32'h3a1fa6a3),
	.w6(32'h3b6c9964),
	.w7(32'hba367eb6),
	.w8(32'h39d78908),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95d69),
	.w1(32'h3a796d60),
	.w2(32'h39498fdd),
	.w3(32'hb91a27c2),
	.w4(32'hb9e9b4a0),
	.w5(32'hb9f0b22b),
	.w6(32'h391ab18e),
	.w7(32'hb9951983),
	.w8(32'hbaa3c090),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ce42d),
	.w1(32'hbb83bde3),
	.w2(32'hbb8c9ff7),
	.w3(32'hba6cf98b),
	.w4(32'hbb0acad1),
	.w5(32'hbb69260e),
	.w6(32'hbb23ce91),
	.w7(32'h398255fe),
	.w8(32'h3b3422f8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9a70d),
	.w1(32'h3c09d71f),
	.w2(32'h3bac29d5),
	.w3(32'hbb5f7052),
	.w4(32'hbbcfc005),
	.w5(32'h3ac26c25),
	.w6(32'h3ba1bd6f),
	.w7(32'h3a7c00b0),
	.w8(32'h39954595),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a18239),
	.w1(32'h3a2ec711),
	.w2(32'hba6902b5),
	.w3(32'h39c18717),
	.w4(32'hbab4982b),
	.w5(32'hba41c86c),
	.w6(32'h3b008716),
	.w7(32'h38e7720b),
	.w8(32'h3a2f44a2),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28dc2b),
	.w1(32'h3a564d11),
	.w2(32'h3c0186a5),
	.w3(32'h3961f8af),
	.w4(32'hba9e3313),
	.w5(32'h3b1bb6ac),
	.w6(32'h3b17effb),
	.w7(32'h3bcbf0d3),
	.w8(32'h39b72c64),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a79c2d),
	.w1(32'hba14dfe0),
	.w2(32'hb8e0d6b9),
	.w3(32'hb7294420),
	.w4(32'hb91f9117),
	.w5(32'h3734bc26),
	.w6(32'h388cce5f),
	.w7(32'h38efb59a),
	.w8(32'hbb809ab3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d29f),
	.w1(32'hba674fbe),
	.w2(32'hbb2f241d),
	.w3(32'hb99e6659),
	.w4(32'h3b2a7a6f),
	.w5(32'hba3bae6c),
	.w6(32'hbb6693d1),
	.w7(32'hbb30971f),
	.w8(32'hba56c4b1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adee51b),
	.w1(32'h3b022616),
	.w2(32'hbad5f513),
	.w3(32'h3ac7cb22),
	.w4(32'hbbd5149f),
	.w5(32'hbbea3400),
	.w6(32'h3b71c36a),
	.w7(32'h39747187),
	.w8(32'h3a922022),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea42a7),
	.w1(32'h3b196552),
	.w2(32'h3b26462b),
	.w3(32'hbac8b279),
	.w4(32'hbb1b1184),
	.w5(32'hba67f8d3),
	.w6(32'h3adb5373),
	.w7(32'h3ad0f938),
	.w8(32'h38fb2301),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dffb37),
	.w1(32'hbac811ce),
	.w2(32'hba23da82),
	.w3(32'hba9ed9ba),
	.w4(32'hbb3fad42),
	.w5(32'hbad147e3),
	.w6(32'hb7e15e8a),
	.w7(32'hb9cc7f6b),
	.w8(32'h3ac09669),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4821dd),
	.w1(32'hbb9827db),
	.w2(32'h3ae2356f),
	.w3(32'h3875e0f7),
	.w4(32'h3ae4d766),
	.w5(32'h3b7ecc36),
	.w6(32'h3aa9f4cc),
	.w7(32'h3b24417a),
	.w8(32'h37b56b5a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule