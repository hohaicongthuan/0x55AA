module layer_8_featuremap_42(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7995a2),
	.w1(32'h385218d9),
	.w2(32'h3b32065e),
	.w3(32'hbbb212e9),
	.w4(32'hbad1171e),
	.w5(32'h3b12aefe),
	.w6(32'hbb6f9fd6),
	.w7(32'hba33e666),
	.w8(32'h3b53d360),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037e40),
	.w1(32'h3bd25a43),
	.w2(32'h3b958ead),
	.w3(32'h3bd0f44f),
	.w4(32'h3ba5b39f),
	.w5(32'h3b844fcf),
	.w6(32'h3bc3ad78),
	.w7(32'h3ba812b1),
	.w8(32'h3b9ca60f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3afb0c),
	.w1(32'h3c098268),
	.w2(32'h3c01530c),
	.w3(32'h3c2e62ef),
	.w4(32'h3c0966fe),
	.w5(32'h3bee0dd1),
	.w6(32'h3c426de6),
	.w7(32'h3c22e728),
	.w8(32'h3c1976a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b22d25),
	.w1(32'h3818b803),
	.w2(32'hb92b8f12),
	.w3(32'h38af0a5b),
	.w4(32'h38689cd8),
	.w5(32'hb906f657),
	.w6(32'hb5f54e88),
	.w7(32'hb76cbb91),
	.w8(32'hb937675a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6e659),
	.w1(32'h3ba96fb6),
	.w2(32'h3bb04120),
	.w3(32'h3b7cc050),
	.w4(32'h3b663518),
	.w5(32'h3b96b2a0),
	.w6(32'h3b570951),
	.w7(32'h3b7c3279),
	.w8(32'h3bc62b18),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b030410),
	.w1(32'h398e8001),
	.w2(32'h3ba340cd),
	.w3(32'h3aee777b),
	.w4(32'hb66ada28),
	.w5(32'h3b718761),
	.w6(32'h3b0e5b88),
	.w7(32'h3aa2f85f),
	.w8(32'h3bafd961),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7c6f3),
	.w1(32'h3897e0a9),
	.w2(32'hb91b7a01),
	.w3(32'h39048f18),
	.w4(32'h387014c0),
	.w5(32'hb915d016),
	.w6(32'h381fb986),
	.w7(32'h36c49ea4),
	.w8(32'hb956758d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c309967),
	.w1(32'h3bf3b218),
	.w2(32'h3c0e4036),
	.w3(32'h3be792dc),
	.w4(32'h3ba36f5f),
	.w5(32'h3bde7257),
	.w6(32'h3c0cdda8),
	.w7(32'h3c19f873),
	.w8(32'h3c388ada),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22136b),
	.w1(32'h3c0b50bf),
	.w2(32'h3ba271ee),
	.w3(32'h3c1450d6),
	.w4(32'h3be6d5de),
	.w5(32'h3b63b347),
	.w6(32'h3c23b756),
	.w7(32'h3c1f4468),
	.w8(32'h3c1be9f3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be18c3c),
	.w1(32'h3bd8d306),
	.w2(32'h3bd495d8),
	.w3(32'h3b8632f0),
	.w4(32'h3b76d67a),
	.w5(32'h3bab8d0b),
	.w6(32'h3bbd7c7e),
	.w7(32'h3bae6805),
	.w8(32'h3bef2a58),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad45d1),
	.w1(32'hbb2593f4),
	.w2(32'h3b18e54a),
	.w3(32'hbbd430c2),
	.w4(32'hbb3fb04b),
	.w5(32'h3b283d06),
	.w6(32'hbbc554ce),
	.w7(32'hbb521d1e),
	.w8(32'h3b04482a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ea71a),
	.w1(32'h3aeaec8f),
	.w2(32'h3b296fcb),
	.w3(32'h3a9512ca),
	.w4(32'h3a8bfd63),
	.w5(32'h3af274ac),
	.w6(32'h3a982e3d),
	.w7(32'h3ab441c2),
	.w8(32'h3b312823),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b84c1),
	.w1(32'h3be078ff),
	.w2(32'h3b7b7422),
	.w3(32'h3c1690fe),
	.w4(32'h3bc8be72),
	.w5(32'h3b203b2d),
	.w6(32'h3c27acf1),
	.w7(32'h3bff2764),
	.w8(32'h3bc87cd0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f962d6),
	.w1(32'hb8ccc465),
	.w2(32'hb90091e4),
	.w3(32'h38748c14),
	.w4(32'hb90f6236),
	.w5(32'hb906694d),
	.w6(32'h37513310),
	.w7(32'hb95c85af),
	.w8(32'hb9040c70),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ec649),
	.w1(32'hb798b277),
	.w2(32'hb90b8993),
	.w3(32'h37e7ac12),
	.w4(32'hb6d6ee65),
	.w5(32'hb901c78d),
	.w6(32'hb7927d21),
	.w7(32'hb80db6aa),
	.w8(32'hb914b1b1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890ddb3),
	.w1(32'h39da4c0d),
	.w2(32'h3947c85b),
	.w3(32'hb65282f2),
	.w4(32'h394d0bd9),
	.w5(32'h38b15c22),
	.w6(32'hb7456efe),
	.w7(32'h39b6d266),
	.w8(32'h39974d99),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9006a2),
	.w1(32'h3a4e9c4c),
	.w2(32'h3a8d7db1),
	.w3(32'h3a451cbe),
	.w4(32'h3a0184f2),
	.w5(32'h3a2f85e8),
	.w6(32'h3a64703d),
	.w7(32'h3a5fc37d),
	.w8(32'h3a986a2b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf4ba4),
	.w1(32'h3ba286aa),
	.w2(32'h3bc78e93),
	.w3(32'h3b86a652),
	.w4(32'h3b7f2bda),
	.w5(32'h3ba72c3c),
	.w6(32'h3bab3410),
	.w7(32'h3b87fd94),
	.w8(32'h3bd0efe7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b75c9),
	.w1(32'hbbbd3532),
	.w2(32'h3be075d3),
	.w3(32'hbc8785e0),
	.w4(32'hbbe8e8fa),
	.w5(32'h3bac9d02),
	.w6(32'hbc73965c),
	.w7(32'hbc05381b),
	.w8(32'h3bb3746c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f690),
	.w1(32'hbc044641),
	.w2(32'h3ba2385c),
	.w3(32'hbc7431c2),
	.w4(32'hbc1dca32),
	.w5(32'h3af82498),
	.w6(32'hbc4eb24d),
	.w7(32'hbc34b876),
	.w8(32'h3b50b6f3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a5c59),
	.w1(32'hbb1628d9),
	.w2(32'h3ab884c3),
	.w3(32'hbb2367fb),
	.w4(32'hbb128604),
	.w5(32'h3aa000a8),
	.w6(32'hbadb712a),
	.w7(32'hbb0f0c78),
	.w8(32'h3a8d40d0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57f4bf),
	.w1(32'h3c28072c),
	.w2(32'h3c02b37f),
	.w3(32'h3c3e5c14),
	.w4(32'h3bec7f02),
	.w5(32'h3bc73e08),
	.w6(32'h3c403ba2),
	.w7(32'h3bf369d6),
	.w8(32'h3bd93c97),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33e30a),
	.w1(32'h3c6a0bd6),
	.w2(32'h3c72bd02),
	.w3(32'h3bdc23fa),
	.w4(32'h3c2b5c89),
	.w5(32'h3c6442fd),
	.w6(32'h3bc529f7),
	.w7(32'h3c39e16b),
	.w8(32'h3c7a09f0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d4442),
	.w1(32'hb90308d1),
	.w2(32'h3b18cc78),
	.w3(32'hbb44fe41),
	.w4(32'hbb068c27),
	.w5(32'h3ad3fd02),
	.w6(32'hbb6c80d0),
	.w7(32'hba0b974b),
	.w8(32'h3b58a57e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04e248),
	.w1(32'hb9a3f2b5),
	.w2(32'h3975f8c7),
	.w3(32'hb9c88dd4),
	.w4(32'hba29219c),
	.w5(32'h394814a2),
	.w6(32'hb925c82e),
	.w7(32'hb9c9c5a8),
	.w8(32'h39a9e210),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac518f5),
	.w1(32'h3b821f2e),
	.w2(32'h3bcb638b),
	.w3(32'hbb1d496b),
	.w4(32'h3b1e49aa),
	.w5(32'h3bd24839),
	.w6(32'hbb3f6d26),
	.w7(32'h398a27a2),
	.w8(32'h3bc1d9dc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f95898),
	.w1(32'hb7ae6ee3),
	.w2(32'h385050dd),
	.w3(32'hb7ff2668),
	.w4(32'hb8839b23),
	.w5(32'h37ad2be8),
	.w6(32'hb770b23e),
	.w7(32'hb7203452),
	.w8(32'hb7bcbea3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb4a9f),
	.w1(32'hbc76aabd),
	.w2(32'h3ba6a483),
	.w3(32'hbcadeb54),
	.w4(32'hbce3cae9),
	.w5(32'hba5fb48c),
	.w6(32'hbb3034af),
	.w7(32'hbcb408cf),
	.w8(32'h3b9740e8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6104d0),
	.w1(32'h3ac97c16),
	.w2(32'h3b7aabb2),
	.w3(32'hbb015f5b),
	.w4(32'hba2a3671),
	.w5(32'h3b2ca865),
	.w6(32'hba656eb7),
	.w7(32'h39318d7c),
	.w8(32'h3b62d28c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b305284),
	.w1(32'h3acc8bd7),
	.w2(32'h3abc7496),
	.w3(32'h3b188b1a),
	.w4(32'h3aa10842),
	.w5(32'h3a73000c),
	.w6(32'h3b2a3826),
	.w7(32'h3b034299),
	.w8(32'h3b008d21),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07c10c),
	.w1(32'h3ab3428e),
	.w2(32'h3b89039a),
	.w3(32'h3ad63841),
	.w4(32'h3a0696a4),
	.w5(32'h3b50dcb2),
	.w6(32'h3b5b1493),
	.w7(32'h3b14a17c),
	.w8(32'h3b8da7c6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227c9f),
	.w1(32'h3b0a8ce2),
	.w2(32'h3b306e83),
	.w3(32'h39af78cf),
	.w4(32'h3a889eee),
	.w5(32'h3b1919be),
	.w6(32'h3adaabd9),
	.w7(32'h3b0779fc),
	.w8(32'h3b59299f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d380ab),
	.w1(32'hb7e5980f),
	.w2(32'hb96ea82e),
	.w3(32'h382ac334),
	.w4(32'h36ec229c),
	.w5(32'hb954816b),
	.w6(32'hb8883328),
	.w7(32'hb8934997),
	.w8(32'hb9967e82),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38059d24),
	.w1(32'hb6f5bba1),
	.w2(32'hb9666561),
	.w3(32'h387f166e),
	.w4(32'h37b9ee75),
	.w5(32'hb9461245),
	.w6(32'hb7938511),
	.w7(32'hb860b348),
	.w8(32'hb98482f7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392ab50c),
	.w1(32'hbb86e2a4),
	.w2(32'h398cfc72),
	.w3(32'h3a4027eb),
	.w4(32'hbb515c94),
	.w5(32'h3984e60e),
	.w6(32'h3b0d60df),
	.w7(32'hbb022155),
	.w8(32'h3a88ef38),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cfdcf),
	.w1(32'hbab3e728),
	.w2(32'h3aa918e6),
	.w3(32'hbba2aca3),
	.w4(32'hbb348ffe),
	.w5(32'h3a05b402),
	.w6(32'hbb9f21ad),
	.w7(32'hbb1a8459),
	.w8(32'h3a837c45),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2f070),
	.w1(32'hb89356ca),
	.w2(32'hb926ae17),
	.w3(32'hb7d7a851),
	.w4(32'hb894ea27),
	.w5(32'hb92fd629),
	.w6(32'hb876e86d),
	.w7(32'hb7a1c24c),
	.w8(32'hb9459b37),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190a5c),
	.w1(32'h3c0104d8),
	.w2(32'h3b96a152),
	.w3(32'h3bde4756),
	.w4(32'h3bb71dec),
	.w5(32'h3b8638df),
	.w6(32'h3be1f66e),
	.w7(32'h3bb7b1b5),
	.w8(32'h3b8b437a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86bc2c7),
	.w1(32'hb8b6dc13),
	.w2(32'hb98b58d0),
	.w3(32'h386e022c),
	.w4(32'hb7e450bb),
	.w5(32'hb94b1a1d),
	.w6(32'h3872b0a0),
	.w7(32'hb8bc8c52),
	.w8(32'hb99ff05d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa41df),
	.w1(32'hb9346255),
	.w2(32'hb980a121),
	.w3(32'hb8c7d922),
	.w4(32'hb96c6288),
	.w5(32'hb995b35e),
	.w6(32'hb91ab3e4),
	.w7(32'hb98570c0),
	.w8(32'hb9a798e0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6fd58),
	.w1(32'h3b910c24),
	.w2(32'h3bb7402f),
	.w3(32'h3b9c1fde),
	.w4(32'h3bbbe401),
	.w5(32'h3be6c946),
	.w6(32'h3bc1e0b2),
	.w7(32'h3bbe95bc),
	.w8(32'h3bcfd71b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d140e0),
	.w1(32'hba032aa2),
	.w2(32'h3a57ff94),
	.w3(32'hb98e0f04),
	.w4(32'hba475765),
	.w5(32'h3a1b7be8),
	.w6(32'hb88a42ac),
	.w7(32'hb99d4a49),
	.w8(32'hbaa544e7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aad90),
	.w1(32'hbb3396cc),
	.w2(32'hbabbbfee),
	.w3(32'hbb321219),
	.w4(32'hbb3f6d01),
	.w5(32'hbaeebee5),
	.w6(32'hbb69c5fc),
	.w7(32'hbb11f733),
	.w8(32'hb9c3963a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb634f0b),
	.w1(32'hbadc6144),
	.w2(32'h3ad224f7),
	.w3(32'hbb7f7195),
	.w4(32'hbb05a77e),
	.w5(32'h3aa794f8),
	.w6(32'hbb33e409),
	.w7(32'hba97eaad),
	.w8(32'h3b26460c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0977),
	.w1(32'hb9c21699),
	.w2(32'h3b59ca21),
	.w3(32'hbbd3a364),
	.w4(32'hbb5cb71d),
	.w5(32'h39e58db0),
	.w6(32'hbbbe1dde),
	.w7(32'hbb564fb5),
	.w8(32'h3b77e244),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9cb50),
	.w1(32'h3ac22e7d),
	.w2(32'h3a2cb93a),
	.w3(32'h3ae64bff),
	.w4(32'h3ab30f7f),
	.w5(32'h39ed4622),
	.w6(32'h3aa34c2d),
	.w7(32'h3a63742a),
	.w8(32'hbac5d744),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a375f7b),
	.w1(32'h3a1cffa7),
	.w2(32'h3a998f85),
	.w3(32'h38f0968d),
	.w4(32'h3a89da25),
	.w5(32'h390f79f0),
	.w6(32'hba640390),
	.w7(32'h385b2f61),
	.w8(32'h3a9056c5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a1bc0),
	.w1(32'h39c698f1),
	.w2(32'h3b2e9f48),
	.w3(32'hbbbd7dd7),
	.w4(32'hbb07e328),
	.w5(32'h3ad5c2c4),
	.w6(32'hbb946daf),
	.w7(32'hbb366aea),
	.w8(32'h3b0d6435),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b747a54),
	.w1(32'h3b47d0cf),
	.w2(32'h3be8f231),
	.w3(32'h3b39e292),
	.w4(32'h3b048f32),
	.w5(32'h3bd3c5b4),
	.w6(32'h3b3c808f),
	.w7(32'h3b53921c),
	.w8(32'h3bde96bf),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d323),
	.w1(32'h39de8eef),
	.w2(32'h3a9373c9),
	.w3(32'hb89f2d5d),
	.w4(32'hb966a5c5),
	.w5(32'h3a3abdf3),
	.w6(32'h38d46fab),
	.w7(32'h387a8bd7),
	.w8(32'h3b033855),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c859ed0),
	.w1(32'h3c5a9c22),
	.w2(32'h3bac7ddb),
	.w3(32'h3c49ac85),
	.w4(32'h3c24fac7),
	.w5(32'h3b898526),
	.w6(32'h3c3c219e),
	.w7(32'h3c16e734),
	.w8(32'h3b97e862),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5080),
	.w1(32'hbad3991f),
	.w2(32'h3c60ee9b),
	.w3(32'hbc0cad7e),
	.w4(32'hbb882eda),
	.w5(32'h3c073a55),
	.w6(32'hbbd88209),
	.w7(32'hbb145818),
	.w8(32'h3c5d6f52),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7e54),
	.w1(32'hbb186a91),
	.w2(32'h3b883e37),
	.w3(32'hbc00db47),
	.w4(32'hbb679edd),
	.w5(32'h3b4f45d1),
	.w6(32'hbbffed7d),
	.w7(32'hbb04356d),
	.w8(32'h3aa18545),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8fe54),
	.w1(32'hba53c29f),
	.w2(32'h3a20f27e),
	.w3(32'hbb5f5cf6),
	.w4(32'hbb10a062),
	.w5(32'hb9c64633),
	.w6(32'hbb4d8b5c),
	.w7(32'hbadf7c63),
	.w8(32'h3afe89b0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ee4320),
	.w1(32'h39fabec9),
	.w2(32'h3a2d807d),
	.w3(32'hb9275f97),
	.w4(32'h37fff586),
	.w5(32'hb9d53396),
	.w6(32'hb9e0d163),
	.w7(32'hb8aab008),
	.w8(32'hbaf6fdf4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7704ed),
	.w1(32'h3bdc60b5),
	.w2(32'h3b8bb573),
	.w3(32'hb92097b5),
	.w4(32'h3b277373),
	.w5(32'h3b26bc8d),
	.w6(32'h3a35abf2),
	.w7(32'h3aa40d41),
	.w8(32'h3b99468b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9b71b),
	.w1(32'h3901009b),
	.w2(32'h3b45193d),
	.w3(32'hb9393fe1),
	.w4(32'hbad8f871),
	.w5(32'h3a9438c2),
	.w6(32'h3a9d5430),
	.w7(32'h3901e18d),
	.w8(32'h3b53f964),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00b745),
	.w1(32'h3bf9b363),
	.w2(32'h3c374223),
	.w3(32'h3bc1d171),
	.w4(32'h3be437da),
	.w5(32'h3c15af88),
	.w6(32'h3bdd7af5),
	.w7(32'h3bfe6aea),
	.w8(32'h3c51bc63),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac304c7),
	.w1(32'h3b03d62c),
	.w2(32'h3b9f0ee0),
	.w3(32'h3a93fae9),
	.w4(32'h3af4d00c),
	.w5(32'h3b995822),
	.w6(32'h3abf7feb),
	.w7(32'h3b65e1da),
	.w8(32'h3b35b890),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cfb7b),
	.w1(32'hbbaa092e),
	.w2(32'hbb6f2101),
	.w3(32'hbaf0ef87),
	.w4(32'hbb6a2252),
	.w5(32'hbb63c62a),
	.w6(32'hbb760af0),
	.w7(32'hbb39c269),
	.w8(32'hba218ad3),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49d42b),
	.w1(32'h3b046685),
	.w2(32'h3a8af1ee),
	.w3(32'h39af61dd),
	.w4(32'h393f22e2),
	.w5(32'hb9f97030),
	.w6(32'hb92c2f21),
	.w7(32'hb8cc1589),
	.w8(32'h3a7cb625),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1758a),
	.w1(32'h3af24ab5),
	.w2(32'h3a679787),
	.w3(32'h3aaed56d),
	.w4(32'h3aaa50e7),
	.w5(32'h3a771cbe),
	.w6(32'h3aea69cd),
	.w7(32'h3a9b6432),
	.w8(32'hba87583d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32cbbe),
	.w1(32'h3a442fa2),
	.w2(32'h3c0501d6),
	.w3(32'hbbc24236),
	.w4(32'hbb3cce97),
	.w5(32'h3ba552d6),
	.w6(32'hbb283831),
	.w7(32'hba784bd6),
	.w8(32'h3c0349d1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b334e2e),
	.w1(32'h3ab0f638),
	.w2(32'h3ab1ea0d),
	.w3(32'h3b43527a),
	.w4(32'h3abfe12d),
	.w5(32'hb743e035),
	.w6(32'h3b1b6bbc),
	.w7(32'h397de088),
	.w8(32'h3b02171b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dc7a7),
	.w1(32'hbb252dad),
	.w2(32'hbac00ead),
	.w3(32'hbb366d22),
	.w4(32'hbb581d0c),
	.w5(32'hbb22fe43),
	.w6(32'hbb19f94b),
	.w7(32'hbb3fb155),
	.w8(32'hba642d3d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed6c4),
	.w1(32'h3babf21c),
	.w2(32'h3b9391d0),
	.w3(32'h3bbdd5cd),
	.w4(32'h3bb607f1),
	.w5(32'h3b8f79df),
	.w6(32'h3bcc30bb),
	.w7(32'h3bebab3e),
	.w8(32'h3bdd48fd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2114e),
	.w1(32'h3bab5305),
	.w2(32'h3bd96241),
	.w3(32'h3bbf8b1a),
	.w4(32'h3b8f99f6),
	.w5(32'h3bafc503),
	.w6(32'h3bf8cc77),
	.w7(32'h3be5c0c4),
	.w8(32'h3c0ffba1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99fc0c3),
	.w1(32'h39587bc3),
	.w2(32'h3ae00194),
	.w3(32'hbaf13097),
	.w4(32'hba704a9b),
	.w5(32'h3a46ddbd),
	.w6(32'h3905d018),
	.w7(32'h3a2f2dc5),
	.w8(32'h3ab19e2b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a0b9f2),
	.w1(32'hba119930),
	.w2(32'hba489921),
	.w3(32'hba09e38e),
	.w4(32'hba2194b8),
	.w5(32'hba3d9cd6),
	.w6(32'hba35a282),
	.w7(32'hba202679),
	.w8(32'h3a079236),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61c787),
	.w1(32'hbc2dcd6b),
	.w2(32'h3a960383),
	.w3(32'hbc794c9b),
	.w4(32'hbc2b9150),
	.w5(32'h3b2911c0),
	.w6(32'hbc68a0da),
	.w7(32'hbc24f4c5),
	.w8(32'h3b41440b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41647c),
	.w1(32'hba971eaa),
	.w2(32'hba7abc3a),
	.w3(32'hba20fd2f),
	.w4(32'hba739b10),
	.w5(32'hba477bb5),
	.w6(32'hba53c34a),
	.w7(32'hba62b7d6),
	.w8(32'h380af607),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999dba8),
	.w1(32'h3a6cbcf4),
	.w2(32'h3b981d70),
	.w3(32'hbae1e191),
	.w4(32'hb90d7f0b),
	.w5(32'h3b8b8f80),
	.w6(32'hb908f9e7),
	.w7(32'h3a674ce6),
	.w8(32'h3bbef9b6),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba185eed),
	.w1(32'hbab7557b),
	.w2(32'hbac1abde),
	.w3(32'hb9eb4fc4),
	.w4(32'hba90edc9),
	.w5(32'hbaaafdee),
	.w6(32'hba473184),
	.w7(32'hba6b25bc),
	.w8(32'hba742d19),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c135676),
	.w1(32'h3bdb5aa4),
	.w2(32'h3b298a0b),
	.w3(32'h3ba73473),
	.w4(32'h3ba0fd55),
	.w5(32'h3b448435),
	.w6(32'h3ba04475),
	.w7(32'h3b4bbd1b),
	.w8(32'h3ba0e867),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87f954),
	.w1(32'h3a1b9b29),
	.w2(32'h3945b301),
	.w3(32'h3a7763fc),
	.w4(32'h3a536847),
	.w5(32'h393a1121),
	.w6(32'h3a62df61),
	.w7(32'h39e09338),
	.w8(32'hb991fb83),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8daf85),
	.w1(32'h3b9f0772),
	.w2(32'h3c0c22f0),
	.w3(32'h3b09161c),
	.w4(32'h3b4e1b41),
	.w5(32'h3bfaa287),
	.w6(32'h3b81c477),
	.w7(32'h3b9a91c8),
	.w8(32'h3c20a8e5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36988fb0),
	.w1(32'hb9b7e7b0),
	.w2(32'hba0a6c04),
	.w3(32'h382be03b),
	.w4(32'hb958a8bc),
	.w5(32'hb9dd36d9),
	.w6(32'hb807118c),
	.w7(32'hb99aacf5),
	.w8(32'h3a519b13),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd0aae),
	.w1(32'hbb386896),
	.w2(32'h3ae64af4),
	.w3(32'hbc0d9d3b),
	.w4(32'hbb9a8938),
	.w5(32'h3a9ac506),
	.w6(32'hbbc3afd7),
	.w7(32'hbb299af4),
	.w8(32'h3b05fea9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a4313),
	.w1(32'h3b11aff0),
	.w2(32'h391a393f),
	.w3(32'h3b02a70d),
	.w4(32'h3a22a063),
	.w5(32'hb99dc92b),
	.w6(32'h3b0aeb17),
	.w7(32'h3ab61336),
	.w8(32'hb9942d31),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88719f4),
	.w1(32'hba32f6a1),
	.w2(32'hb9a6f4b3),
	.w3(32'hb9d05057),
	.w4(32'hba2720d8),
	.w5(32'hb9ae54a2),
	.w6(32'hb99eca36),
	.w7(32'hba07b360),
	.w8(32'h3b0a6ede),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab322a0),
	.w1(32'h3ad93543),
	.w2(32'h3aa8ff79),
	.w3(32'h3aa20445),
	.w4(32'h3aa5e092),
	.w5(32'h3a86ddae),
	.w6(32'h3ad02a27),
	.w7(32'h3ae4b1a9),
	.w8(32'h3a6018ef),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22554e),
	.w1(32'h3ae4af16),
	.w2(32'h3b3b8130),
	.w3(32'h3b0b01d8),
	.w4(32'h3a9e6d64),
	.w5(32'h3b17b9c5),
	.w6(32'h3b3a7746),
	.w7(32'h3b037fbb),
	.w8(32'h3b8a284c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda2bfa),
	.w1(32'hbb7c347b),
	.w2(32'hb99f2b69),
	.w3(32'hbc04f3f6),
	.w4(32'hbb8901f5),
	.w5(32'hba322d2d),
	.w6(32'hbbf0c24f),
	.w7(32'hbba08a66),
	.w8(32'h3b72d5a1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f4a5),
	.w1(32'h3b0d7d45),
	.w2(32'h3c332668),
	.w3(32'h3ad375e3),
	.w4(32'h3af6935f),
	.w5(32'h3c16484d),
	.w6(32'h3b7cde73),
	.w7(32'h3b6d3a96),
	.w8(32'h3bfdafc4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc133041),
	.w1(32'hbb5631d0),
	.w2(32'h3b6922f1),
	.w3(32'hbc641cb3),
	.w4(32'hbbd63f9f),
	.w5(32'h3b4e9105),
	.w6(32'hbc40e2aa),
	.w7(32'hbbb6a1cd),
	.w8(32'h3be0f3b2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009f24),
	.w1(32'hbb2272fa),
	.w2(32'h3b048dac),
	.w3(32'hbc2616a3),
	.w4(32'hbb85ee84),
	.w5(32'h3a95a5c3),
	.w6(32'hbbf916d3),
	.w7(32'hbb64bf23),
	.w8(32'h3b623fc5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab22fb9),
	.w1(32'h39e6eda9),
	.w2(32'hb8805bff),
	.w3(32'h3b00aab0),
	.w4(32'h3a8ed435),
	.w5(32'h3a08d271),
	.w6(32'h38cb7223),
	.w7(32'h39efb2c8),
	.w8(32'hba7b3d24),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c091fc),
	.w1(32'hb9a6f03b),
	.w2(32'hbab1d77d),
	.w3(32'h39af72a3),
	.w4(32'hb91a5379),
	.w5(32'hba96eb3b),
	.w6(32'hb9e9dd3c),
	.w7(32'hba70aaa6),
	.w8(32'hbb633fb4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb436411),
	.w1(32'hbbb02861),
	.w2(32'hbb963b41),
	.w3(32'hbb313a4e),
	.w4(32'hbb86374f),
	.w5(32'hbb8b6fe2),
	.w6(32'hbb83aa86),
	.w7(32'hbb799fe5),
	.w8(32'h3a0469a8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42ec75),
	.w1(32'hba2765dc),
	.w2(32'h3a647c4d),
	.w3(32'hbb6b0653),
	.w4(32'hbac4294d),
	.w5(32'h3ab9febf),
	.w6(32'hbb8e2e41),
	.w7(32'hba9305b7),
	.w8(32'h3a98b60c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9d17c),
	.w1(32'h3a6f3b9c),
	.w2(32'h3acfe9e6),
	.w3(32'h3ae8a074),
	.w4(32'h3a9bd6c4),
	.w5(32'h3af0e0d0),
	.w6(32'h3a88c187),
	.w7(32'h3abd0027),
	.w8(32'hbae731cd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f3799),
	.w1(32'hbb791c65),
	.w2(32'hbb10f059),
	.w3(32'hbb401ca3),
	.w4(32'hbb409305),
	.w5(32'hbac45d93),
	.w6(32'hbb3d0850),
	.w7(32'hbb382cef),
	.w8(32'h3a3de041),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f18b0e),
	.w1(32'hbb37e860),
	.w2(32'hba2ee10f),
	.w3(32'hbab34dbd),
	.w4(32'hbb3218f9),
	.w5(32'hb9b88062),
	.w6(32'hbacc3569),
	.w7(32'hbb39608c),
	.w8(32'h3b3fe30e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d6cba),
	.w1(32'h3ace201b),
	.w2(32'h3ba98fe1),
	.w3(32'hbb097803),
	.w4(32'hba820ccb),
	.w5(32'h3b72d9bb),
	.w6(32'h386235a6),
	.w7(32'h39c057d0),
	.w8(32'h3ba393fa),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b593a73),
	.w1(32'h3b3c5d24),
	.w2(32'h3a48da9b),
	.w3(32'h3b3588c7),
	.w4(32'h3b14b125),
	.w5(32'hb8869e4c),
	.w6(32'h3b5342ef),
	.w7(32'h3a92b7d4),
	.w8(32'hbbbd54ce),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc044cbf),
	.w1(32'hbc167e49),
	.w2(32'hbb99dcb2),
	.w3(32'hbc2325cb),
	.w4(32'hbc1c3dc3),
	.w5(32'hbbae0c77),
	.w6(32'hbc20ac05),
	.w7(32'hbc128fad),
	.w8(32'h3ab2bdf1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44674a),
	.w1(32'h3b5885b4),
	.w2(32'h3b8f5015),
	.w3(32'hbb795551),
	.w4(32'hb9886344),
	.w5(32'h3b4d5650),
	.w6(32'hbaece07a),
	.w7(32'h3aa55364),
	.w8(32'h3ba48468),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139af3),
	.w1(32'hbad8d589),
	.w2(32'hbb08ffe6),
	.w3(32'hbaa8e8ba),
	.w4(32'hba8b07df),
	.w5(32'hbb0450d4),
	.w6(32'hbab608e6),
	.w7(32'hbaab66eb),
	.w8(32'h3a16b417),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba003405),
	.w1(32'hba22a1c9),
	.w2(32'hbab03e31),
	.w3(32'hb9cc39f9),
	.w4(32'hba6dfe3b),
	.w5(32'hba80ca89),
	.w6(32'h3989ddeb),
	.w7(32'h38af1038),
	.w8(32'hba958c03),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f615c0),
	.w1(32'hba9dc246),
	.w2(32'hbb05b94c),
	.w3(32'hb9aeb607),
	.w4(32'hba85875f),
	.w5(32'hbaed98a3),
	.w6(32'hba6c71ad),
	.w7(32'hbab76aab),
	.w8(32'hbb107544),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd7092),
	.w1(32'hbb4043f0),
	.w2(32'hbb0845ca),
	.w3(32'hba9438e9),
	.w4(32'hbadaa8e4),
	.w5(32'hbb060c56),
	.w6(32'hbb2075a7),
	.w7(32'hbb091195),
	.w8(32'h3a7827e5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b950b79),
	.w1(32'h3b88a4b2),
	.w2(32'h3b035033),
	.w3(32'h3b62ae85),
	.w4(32'h3b65bf92),
	.w5(32'h3b006190),
	.w6(32'h3b77dcac),
	.w7(32'h3b5777fa),
	.w8(32'h3aa9faf7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f4b5),
	.w1(32'hba4f9611),
	.w2(32'hb92666f9),
	.w3(32'hbafec26a),
	.w4(32'hbb060de9),
	.w5(32'hba6047ac),
	.w6(32'hba7dd093),
	.w7(32'hba75d0c4),
	.w8(32'hbb864e02),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35a6fc),
	.w1(32'hbb86aff0),
	.w2(32'hbb1e3270),
	.w3(32'hbb10b5ea),
	.w4(32'hbb916898),
	.w5(32'hbb706af7),
	.w6(32'hbb0d920e),
	.w7(32'hbb309d77),
	.w8(32'h3b6d2636),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a650e8e),
	.w1(32'h39ef50b7),
	.w2(32'h3b01c68f),
	.w3(32'h3a2c7c74),
	.w4(32'h390fc362),
	.w5(32'h3af54df7),
	.w6(32'h3a660fd4),
	.w7(32'h3a3d9195),
	.w8(32'hbb66bb2e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb72273),
	.w1(32'hbb3cfeb0),
	.w2(32'h3cd6236f),
	.w3(32'hbc992ab7),
	.w4(32'hba560b6d),
	.w5(32'h3c8b9337),
	.w6(32'hbbf5300e),
	.w7(32'h3c139b9f),
	.w8(32'hbbdf0d96),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc641651),
	.w1(32'h3c87bf0f),
	.w2(32'h3c58ec7b),
	.w3(32'hbc9b1f5b),
	.w4(32'h3b6aec2e),
	.w5(32'h3b96ae99),
	.w6(32'h3be6c8bf),
	.w7(32'h3bb397f0),
	.w8(32'hbb7121b4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc878a11),
	.w1(32'hbb3d4a5a),
	.w2(32'h3ccf8ff4),
	.w3(32'hbc21f87c),
	.w4(32'hbb0ea53b),
	.w5(32'h3c45b864),
	.w6(32'h3a7e4aa2),
	.w7(32'h3c6f78f4),
	.w8(32'hbbf376b6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1b4ab),
	.w1(32'h3b92ec96),
	.w2(32'h3d14153d),
	.w3(32'hbc9f5ed8),
	.w4(32'h3a6f23f1),
	.w5(32'h3cca98b7),
	.w6(32'h3c0983b7),
	.w7(32'h3cb5bf70),
	.w8(32'hbc2188bb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca87ed5),
	.w1(32'h3b41fdf1),
	.w2(32'h3cd03d77),
	.w3(32'hbc9b006e),
	.w4(32'hba0baf14),
	.w5(32'h3c970fae),
	.w6(32'h3b46e54f),
	.w7(32'h3c49d847),
	.w8(32'h3c5a3785),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c829b),
	.w1(32'h3c9348e2),
	.w2(32'h3c8daee5),
	.w3(32'hba139f0f),
	.w4(32'hbb711c21),
	.w5(32'h3c470f41),
	.w6(32'h3cb8585a),
	.w7(32'hbc5338ed),
	.w8(32'h3abeb334),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a337cb7),
	.w1(32'hbbe8d9db),
	.w2(32'h3c291be2),
	.w3(32'hbb0ccfa4),
	.w4(32'hba609f09),
	.w5(32'h3bd08f3f),
	.w6(32'hbc819de1),
	.w7(32'hbbd889ed),
	.w8(32'h3d2b3038),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7ba9e0),
	.w1(32'h3ac9108f),
	.w2(32'hbd295e65),
	.w3(32'h3d2914ff),
	.w4(32'hbb360890),
	.w5(32'hbca9232a),
	.w6(32'hbc046d51),
	.w7(32'hbd0703e6),
	.w8(32'hbbfe0bb8),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc6138f),
	.w1(32'h3a22a9ed),
	.w2(32'h3d0b026f),
	.w3(32'hbcb554b2),
	.w4(32'h393a3ff4),
	.w5(32'h3cb906cd),
	.w6(32'h3aa8c9c8),
	.w7(32'h3cb36468),
	.w8(32'hbc245e0a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860269),
	.w1(32'h3910911d),
	.w2(32'h3c56317f),
	.w3(32'hbc33d708),
	.w4(32'h3a8d765c),
	.w5(32'h3beaaf69),
	.w6(32'h3b3ca72e),
	.w7(32'h3c14f9da),
	.w8(32'hbc990a29),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd068ce7),
	.w1(32'h3ae2f0b6),
	.w2(32'h3d0bb326),
	.w3(32'hbcc689b8),
	.w4(32'h3b172d1f),
	.w5(32'h3c86e1f4),
	.w6(32'h3c1a59ef),
	.w7(32'h3cc0a2a4),
	.w8(32'hbb0c11e9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0988f),
	.w1(32'hbccbce86),
	.w2(32'h3c597c17),
	.w3(32'hbcc848c1),
	.w4(32'hbce6df76),
	.w5(32'h3b56681c),
	.w6(32'hbc47e6d9),
	.w7(32'hbaa5e235),
	.w8(32'h3bfe074c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ead87),
	.w1(32'h3bd24235),
	.w2(32'h3bf8220d),
	.w3(32'hbbc3cab8),
	.w4(32'h396fcd0c),
	.w5(32'h3c5ae8c0),
	.w6(32'h3b96bd67),
	.w7(32'h3c35637c),
	.w8(32'h3c07cbe9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26f490),
	.w1(32'h3c594c8d),
	.w2(32'h3b4960c7),
	.w3(32'h3a3bbae0),
	.w4(32'hbbac6cea),
	.w5(32'hbb87a137),
	.w6(32'h3bb549b4),
	.w7(32'hbb631836),
	.w8(32'h3b9d339d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3469a1),
	.w1(32'hbc894438),
	.w2(32'h3b218299),
	.w3(32'h3bca9fa2),
	.w4(32'hbc640e19),
	.w5(32'hbc79cdc8),
	.w6(32'hbc9edf5b),
	.w7(32'hbc36fad0),
	.w8(32'h3bf1875d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b98b),
	.w1(32'hbc19d838),
	.w2(32'hbc2101bf),
	.w3(32'hbb589357),
	.w4(32'hbc768ffb),
	.w5(32'hbc636cda),
	.w6(32'h3aafb971),
	.w7(32'h3c41fa57),
	.w8(32'h38c13a45),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad509b),
	.w1(32'h3c2f6319),
	.w2(32'h3c8b24d3),
	.w3(32'hbb199037),
	.w4(32'h3bbbe676),
	.w5(32'hbb226c39),
	.w6(32'hbc29f740),
	.w7(32'h3c2589da),
	.w8(32'h3be65d28),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6da674),
	.w1(32'hba0d4855),
	.w2(32'h3c9b0355),
	.w3(32'h3b97fb16),
	.w4(32'hbc21c93d),
	.w5(32'h3bb2f03a),
	.w6(32'hbc2f8602),
	.w7(32'h3bb4dd3c),
	.w8(32'hbc222c1f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9b861),
	.w1(32'h3ab5e2d7),
	.w2(32'h3cdfc029),
	.w3(32'hbc869825),
	.w4(32'hbba3a99f),
	.w5(32'h3cbff5fc),
	.w6(32'h3c06b816),
	.w7(32'h3cdcb096),
	.w8(32'h3c5020c9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d19e4),
	.w1(32'h3c2a23e5),
	.w2(32'h3c49275d),
	.w3(32'h3b8dd110),
	.w4(32'h3bb9c1e6),
	.w5(32'h3c350c22),
	.w6(32'h3c210e35),
	.w7(32'hbc35bfaa),
	.w8(32'hbc80ca05),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce4d7fe),
	.w1(32'hba8b8f0a),
	.w2(32'h3cd16095),
	.w3(32'hbca070f0),
	.w4(32'hbc0bfd44),
	.w5(32'h3bffd8d4),
	.w6(32'hbb53d354),
	.w7(32'h3c5e0008),
	.w8(32'hba90bee0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed77df),
	.w1(32'h3ca85470),
	.w2(32'h3d6148d5),
	.w3(32'hbbf617b6),
	.w4(32'h3cb47895),
	.w5(32'h3d3286a7),
	.w6(32'h3cccfca5),
	.w7(32'h3d41ceea),
	.w8(32'hbbe27959),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09620e),
	.w1(32'h3c65ce36),
	.w2(32'h3bd678a0),
	.w3(32'hbb8066fd),
	.w4(32'h3be62005),
	.w5(32'hbbf4a111),
	.w6(32'h3b43915a),
	.w7(32'h3c9c5316),
	.w8(32'h3b342ef5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule