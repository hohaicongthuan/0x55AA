module layer_10_featuremap_433(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h352fd80d),
	.w1(32'h3ae480ea),
	.w2(32'hba8af842),
	.w3(32'h39591190),
	.w4(32'hbaa3e0b2),
	.w5(32'hbafc591a),
	.w6(32'hbba08295),
	.w7(32'hba8ba573),
	.w8(32'h3aad0f22),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269bc4),
	.w1(32'hba82f1d1),
	.w2(32'hbb07ccc6),
	.w3(32'hbc176ff2),
	.w4(32'hbaee97ce),
	.w5(32'hba8590e1),
	.w6(32'hbb6806ef),
	.w7(32'h3a48f6ca),
	.w8(32'h3a07d32e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a3cb),
	.w1(32'hbbc78a4c),
	.w2(32'hb8cbab2d),
	.w3(32'hbbb05d44),
	.w4(32'hbb32fdaf),
	.w5(32'hbb6edc9c),
	.w6(32'hbb09aa69),
	.w7(32'hbbda1b91),
	.w8(32'hbba36840),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa2919),
	.w1(32'h3b1cfa9b),
	.w2(32'h3b22f34b),
	.w3(32'h3a5e0cc1),
	.w4(32'h3bfb9ba6),
	.w5(32'h3b6befde),
	.w6(32'hbbdd3ad6),
	.w7(32'h3b1d80c0),
	.w8(32'h3bb17b79),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb712747),
	.w1(32'h3b9ae8d0),
	.w2(32'h3a8628f7),
	.w3(32'hbacc1802),
	.w4(32'h3b2551ac),
	.w5(32'h3bf32ac5),
	.w6(32'hbb7a863a),
	.w7(32'h3b3bc010),
	.w8(32'h3ba2153b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27d8a8),
	.w1(32'hbb17a4af),
	.w2(32'h3a365694),
	.w3(32'h3ac14e81),
	.w4(32'h3a384c6a),
	.w5(32'hbb952622),
	.w6(32'h39878534),
	.w7(32'h3b3626a5),
	.w8(32'hb98d700e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc08789),
	.w1(32'hbb322d81),
	.w2(32'hb984b663),
	.w3(32'hbbd4693a),
	.w4(32'hbae54fce),
	.w5(32'h3ac1a212),
	.w6(32'hbba8cd6c),
	.w7(32'h3a278393),
	.w8(32'h3bb86da8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad1201),
	.w1(32'hbada2eb8),
	.w2(32'h3abd074b),
	.w3(32'h3c8460dc),
	.w4(32'h3be5c72f),
	.w5(32'hbb17f81b),
	.w6(32'h3a3e6dcf),
	.w7(32'hb95c328d),
	.w8(32'hbbb33109),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9647f6),
	.w1(32'hbb17b192),
	.w2(32'h3bb2465f),
	.w3(32'hbb8f76ab),
	.w4(32'hba75abd8),
	.w5(32'h3bbb9121),
	.w6(32'hbbe666cb),
	.w7(32'hba747352),
	.w8(32'h3bd36be2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fd91e),
	.w1(32'hbb53acba),
	.w2(32'hbc098741),
	.w3(32'hbb22aea3),
	.w4(32'h3b55b87a),
	.w5(32'hbb8b0785),
	.w6(32'h3906566a),
	.w7(32'h3b9b4700),
	.w8(32'h3bd4e9c8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e02dc),
	.w1(32'h3b05774c),
	.w2(32'hba8f45af),
	.w3(32'h3b72aa3e),
	.w4(32'hba679018),
	.w5(32'hbb57589a),
	.w6(32'h3ac57cac),
	.w7(32'hbb1bf10c),
	.w8(32'hbb1c835e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa50fa1),
	.w1(32'hbb8615b1),
	.w2(32'h3b575763),
	.w3(32'hbb84c4be),
	.w4(32'hbbab35e6),
	.w5(32'hbbab0e03),
	.w6(32'hbb538f0b),
	.w7(32'hba491a0c),
	.w8(32'h3a0261c3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004135),
	.w1(32'h3aa7ae60),
	.w2(32'hbba33db1),
	.w3(32'h3b4c9a1b),
	.w4(32'h3b42dda0),
	.w5(32'hbba06ff5),
	.w6(32'h3a142f32),
	.w7(32'h3b9d82f5),
	.w8(32'hba4b010d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf7cf5),
	.w1(32'h3ba960f9),
	.w2(32'h3a2d331f),
	.w3(32'hbaeac557),
	.w4(32'h3bb92fdd),
	.w5(32'h3c1f9225),
	.w6(32'h3912dcf3),
	.w7(32'h3ace0d5e),
	.w8(32'h3aefb180),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc109d25),
	.w1(32'hbbb237d6),
	.w2(32'h3a7f0948),
	.w3(32'hbb2b5dbb),
	.w4(32'hbb873c2c),
	.w5(32'hbb8973e5),
	.w6(32'hbadeaa51),
	.w7(32'h3b4ece69),
	.w8(32'hbabfebf6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f114),
	.w1(32'h3ab307b2),
	.w2(32'h3a92a9ef),
	.w3(32'h3c56e266),
	.w4(32'h3b1462a3),
	.w5(32'hbaa57636),
	.w6(32'h3c6464a5),
	.w7(32'h3bd03d01),
	.w8(32'hb86ce0b7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8596e0),
	.w1(32'hbb37cbb2),
	.w2(32'hbb998cf3),
	.w3(32'h3b10dde5),
	.w4(32'hbb002af7),
	.w5(32'hbbba5786),
	.w6(32'h3ab6b21a),
	.w7(32'hba19164f),
	.w8(32'hbb9b27d3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01a58d),
	.w1(32'h3c19f0be),
	.w2(32'h3be382d1),
	.w3(32'h3c1f1695),
	.w4(32'h3c112deb),
	.w5(32'h3aea17b5),
	.w6(32'h3b86f10b),
	.w7(32'h3a84e928),
	.w8(32'h3a4a70f2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ece50),
	.w1(32'h39abbc72),
	.w2(32'hbb01a191),
	.w3(32'h3b8842ed),
	.w4(32'h3ae892bb),
	.w5(32'hbb0d30c1),
	.w6(32'hbbac83eb),
	.w7(32'hb9bda814),
	.w8(32'hbafcd77d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8231dc),
	.w1(32'h3b001801),
	.w2(32'hbc04673f),
	.w3(32'hbb03fe90),
	.w4(32'h3c3251ea),
	.w5(32'hbbd599e8),
	.w6(32'h39e104d0),
	.w7(32'hba21c238),
	.w8(32'h3b232a12),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9399f1),
	.w1(32'hbaa9294e),
	.w2(32'h3ac66868),
	.w3(32'hbc087af9),
	.w4(32'hba971374),
	.w5(32'hbb1fd3f7),
	.w6(32'hb92867a4),
	.w7(32'hbb47ceff),
	.w8(32'hbb62bba9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fa465),
	.w1(32'h3b5825cd),
	.w2(32'hbc440c6d),
	.w3(32'hbaa9276c),
	.w4(32'h3c106213),
	.w5(32'hbc379278),
	.w6(32'hbb6b2379),
	.w7(32'h3bd4eb80),
	.w8(32'hbafc6c1f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e099f),
	.w1(32'h3c3fc163),
	.w2(32'hb99ac238),
	.w3(32'h3c5fb941),
	.w4(32'h3b216408),
	.w5(32'hbbb50b04),
	.w6(32'h3c71d984),
	.w7(32'h3c114a91),
	.w8(32'h3b1c2a57),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9ccc3),
	.w1(32'hbbb87715),
	.w2(32'hbbde49f1),
	.w3(32'hbc323edd),
	.w4(32'h39032b70),
	.w5(32'hba85e008),
	.w6(32'hbae0beee),
	.w7(32'h3b1c72f4),
	.w8(32'h3b200124),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca788),
	.w1(32'hbb9fe994),
	.w2(32'hbc2b16f5),
	.w3(32'hbc3ddfda),
	.w4(32'hbc3e6d4d),
	.w5(32'hbc3c40da),
	.w6(32'hbad44a27),
	.w7(32'hb8697fe8),
	.w8(32'h3a9aea18),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb938642),
	.w1(32'hbc13369e),
	.w2(32'hbbc0348a),
	.w3(32'hbbdb2343),
	.w4(32'hbab64631),
	.w5(32'hba8366a6),
	.w6(32'h3a8c9d9e),
	.w7(32'hba055f9b),
	.w8(32'hbb7c7b25),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba14aa8),
	.w1(32'hbb83262f),
	.w2(32'hbb81a669),
	.w3(32'hbb98d37f),
	.w4(32'hbb3866e1),
	.w5(32'h3b2223a8),
	.w6(32'hbb3e0dd9),
	.w7(32'hbb894dec),
	.w8(32'hbb88fa56),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49afd4),
	.w1(32'hbbc98174),
	.w2(32'hbb51962f),
	.w3(32'hbc284a1d),
	.w4(32'hbc68b03f),
	.w5(32'hbb451773),
	.w6(32'hbc2b6a6e),
	.w7(32'hbb9a75fe),
	.w8(32'hbb759bee),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a67f8),
	.w1(32'hbb956d5c),
	.w2(32'hbbd6f09d),
	.w3(32'hb9be8b6e),
	.w4(32'hbc33c17d),
	.w5(32'hbc30fc30),
	.w6(32'hbb086b97),
	.w7(32'hbb99c003),
	.w8(32'hb942701f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232bab),
	.w1(32'hbba9fd16),
	.w2(32'h3ac46de4),
	.w3(32'hbc0231c0),
	.w4(32'hbbc529be),
	.w5(32'hbab2cc17),
	.w6(32'hbba46cfd),
	.w7(32'h3b643077),
	.w8(32'h3b930a2f),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d2ced),
	.w1(32'hbba96553),
	.w2(32'hbb22d5e1),
	.w3(32'h3bb91930),
	.w4(32'h3a832456),
	.w5(32'hbbd3d62b),
	.w6(32'h3bf6281d),
	.w7(32'h3b668917),
	.w8(32'h3a87aa69),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a79a),
	.w1(32'hb97ece60),
	.w2(32'hb9dced48),
	.w3(32'hbab41e90),
	.w4(32'h3a0cde98),
	.w5(32'hba8deaa2),
	.w6(32'hbb074b43),
	.w7(32'h3b4a8468),
	.w8(32'h3a82e46c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3abeb6),
	.w1(32'hba8457ff),
	.w2(32'hbb6a0ecd),
	.w3(32'hbb4db503),
	.w4(32'hbaaf2409),
	.w5(32'h3b6725cb),
	.w6(32'hb9da9a3b),
	.w7(32'hbbf10453),
	.w8(32'hbb1784b4),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a19b),
	.w1(32'hbbad352e),
	.w2(32'hbc067ad6),
	.w3(32'hbb9e967b),
	.w4(32'hbb0c6a7d),
	.w5(32'hbb316ec2),
	.w6(32'hbb398be9),
	.w7(32'h3ab68ac8),
	.w8(32'h3b46704e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0dcdc),
	.w1(32'hbb8fc149),
	.w2(32'hbbdff665),
	.w3(32'h39839cf5),
	.w4(32'hbb31f5a9),
	.w5(32'h3b9c3850),
	.w6(32'hbb99b694),
	.w7(32'hbc0156f1),
	.w8(32'hbb4c016c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd32d),
	.w1(32'hbabb02f3),
	.w2(32'h3ae940bc),
	.w3(32'hb9bbd626),
	.w4(32'hb8289b54),
	.w5(32'hbab1fcf8),
	.w6(32'h3a4ee97e),
	.w7(32'h3b252c0e),
	.w8(32'h3b509822),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0491ae),
	.w1(32'h3c15b341),
	.w2(32'h3be40b3b),
	.w3(32'hbb2f9940),
	.w4(32'h3a8188d5),
	.w5(32'hbbca0c6c),
	.w6(32'h3a27a97f),
	.w7(32'hba643761),
	.w8(32'h3c1295ee),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bfe80),
	.w1(32'hbb606673),
	.w2(32'h3ac6304c),
	.w3(32'hbbf4d0a7),
	.w4(32'hb9eba630),
	.w5(32'h3bee6b10),
	.w6(32'h3b7bcd36),
	.w7(32'h3bfa5b8e),
	.w8(32'h3bce0442),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe69565),
	.w1(32'hbc569a7c),
	.w2(32'h3a719ea9),
	.w3(32'hbc8b3e99),
	.w4(32'hbc7403ca),
	.w5(32'h3bafda7a),
	.w6(32'hbc3d5fd8),
	.w7(32'hbc251bbe),
	.w8(32'h3bcb67f2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad559e7),
	.w1(32'hb9ec8193),
	.w2(32'h3b228e17),
	.w3(32'h3bc381d1),
	.w4(32'hbacca26f),
	.w5(32'h3a616a9b),
	.w6(32'h3b16af94),
	.w7(32'hbb58e120),
	.w8(32'hbace4b2c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac12ca),
	.w1(32'hba64cdac),
	.w2(32'hbbd16dab),
	.w3(32'hbb598f7e),
	.w4(32'hbb4d4eea),
	.w5(32'hbbad18ed),
	.w6(32'hba974ab8),
	.w7(32'hba66c76e),
	.w8(32'hbc0b4f19),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb554342),
	.w1(32'hbb797f26),
	.w2(32'hba237072),
	.w3(32'hbb9e468f),
	.w4(32'hbb8aff45),
	.w5(32'hbb3e3698),
	.w6(32'hbbcc976d),
	.w7(32'hba903090),
	.w8(32'hba714d53),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81286a),
	.w1(32'h3a031162),
	.w2(32'hba91ecd6),
	.w3(32'h3b184f96),
	.w4(32'h3a8305fe),
	.w5(32'hbae56503),
	.w6(32'h3aa46b52),
	.w7(32'h3b184fff),
	.w8(32'h3b00765a),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eda36e),
	.w1(32'h3abab33f),
	.w2(32'h38f98ba1),
	.w3(32'h3aa8d6a3),
	.w4(32'hb9829a67),
	.w5(32'h3c723e7f),
	.w6(32'h3b014cb7),
	.w7(32'hbba2bc51),
	.w8(32'h3c252a61),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b88817),
	.w1(32'hbbbf78a3),
	.w2(32'h3a11f9b7),
	.w3(32'hbbe897bf),
	.w4(32'hbb892059),
	.w5(32'h3af95318),
	.w6(32'hbb057606),
	.w7(32'hba40fb66),
	.w8(32'hbb099c1f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50d45c),
	.w1(32'hba35ec92),
	.w2(32'hbbb0c0ac),
	.w3(32'hba6d9d17),
	.w4(32'hbbaaeefa),
	.w5(32'hbc151ec2),
	.w6(32'hba77297b),
	.w7(32'hbb3ca2ee),
	.w8(32'hba0b5c70),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7232d3a),
	.w1(32'h3b61c06d),
	.w2(32'hbb056c20),
	.w3(32'h3bb0c903),
	.w4(32'hbb349f24),
	.w5(32'hbb9e439b),
	.w6(32'h3bb1fbb5),
	.w7(32'hbacd9b3a),
	.w8(32'hbbef8abd),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c386fe9),
	.w1(32'h3c583dea),
	.w2(32'h3bc22ed3),
	.w3(32'h3c8e4170),
	.w4(32'h3c6d6158),
	.w5(32'h393021ba),
	.w6(32'h3bd4a4a4),
	.w7(32'h3bef2c00),
	.w8(32'h39a48f70),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac23e22),
	.w1(32'hbb0585fc),
	.w2(32'h3a5ec63e),
	.w3(32'h39cdd547),
	.w4(32'hbb824f8a),
	.w5(32'h3bea4fd2),
	.w6(32'hba0be2c2),
	.w7(32'hbb419179),
	.w8(32'h3b87220b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ed246),
	.w1(32'hb8615402),
	.w2(32'h3ba8981e),
	.w3(32'hbb48a69f),
	.w4(32'hb9b40f38),
	.w5(32'hb9b964e5),
	.w6(32'hbaf6f201),
	.w7(32'h3b97b983),
	.w8(32'h3a6514f7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1911b5),
	.w1(32'hbb00eda4),
	.w2(32'h3a925499),
	.w3(32'hbbe4e10b),
	.w4(32'hba524913),
	.w5(32'hb9a853cf),
	.w6(32'hbba9a0ea),
	.w7(32'hbb6d6c5b),
	.w8(32'hba955372),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae115f8),
	.w1(32'h3b0db816),
	.w2(32'hba676acc),
	.w3(32'hbb45d10e),
	.w4(32'hb981fdbf),
	.w5(32'h3bd4a5a8),
	.w6(32'hbb2230b2),
	.w7(32'hbbb628d0),
	.w8(32'h3b1fbded),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4c2a),
	.w1(32'hb9011467),
	.w2(32'h39bc7055),
	.w3(32'hb975318d),
	.w4(32'h3b1a6321),
	.w5(32'hba9926f1),
	.w6(32'h3ba2cd88),
	.w7(32'h3ac73d4d),
	.w8(32'hbac0e18e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12918e),
	.w1(32'h3c7b1506),
	.w2(32'h3b809560),
	.w3(32'h3c5dd7d0),
	.w4(32'h3c4e5ae6),
	.w5(32'h3c318d67),
	.w6(32'h3b75a5aa),
	.w7(32'h3bd25cba),
	.w8(32'h3bdf1b10),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cca73),
	.w1(32'h3b8c0d49),
	.w2(32'h3b8b84f7),
	.w3(32'hbb0fc9c7),
	.w4(32'h3a666c24),
	.w5(32'h3a936d59),
	.w6(32'hbb81a767),
	.w7(32'hbae9f1ab),
	.w8(32'hbb62e6f4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b989e33),
	.w1(32'h3b855e2d),
	.w2(32'h3b64d7cd),
	.w3(32'h3aee1048),
	.w4(32'h3ae4d252),
	.w5(32'h3c26e429),
	.w6(32'h3b000ca3),
	.w7(32'hbb047528),
	.w8(32'h3b8638ad),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3995d),
	.w1(32'h39f303b0),
	.w2(32'hbb407601),
	.w3(32'hbba9d349),
	.w4(32'hbb7d29fa),
	.w5(32'hbbc35f90),
	.w6(32'hbb5868f1),
	.w7(32'hbac64e53),
	.w8(32'hbbb090af),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb445eae),
	.w1(32'hbb7bfe5c),
	.w2(32'h3bfc316c),
	.w3(32'hbb7071e9),
	.w4(32'hbab0e097),
	.w5(32'hbb98b211),
	.w6(32'hbba24b10),
	.w7(32'h3ac96668),
	.w8(32'h3a346cbd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b487dce),
	.w1(32'hba9fdff5),
	.w2(32'hbb9c444a),
	.w3(32'h395da023),
	.w4(32'h3a6c1091),
	.w5(32'hbbbe0386),
	.w6(32'h3ba21472),
	.w7(32'hbacea25e),
	.w8(32'hbb9caf87),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf73ddc),
	.w1(32'hbb1d3d80),
	.w2(32'hbba98b97),
	.w3(32'hbc74602a),
	.w4(32'h3a40497a),
	.w5(32'hbbe9273b),
	.w6(32'hbc160a6f),
	.w7(32'h3adbaf4d),
	.w8(32'hbb24d6d7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004a8e),
	.w1(32'h3b410737),
	.w2(32'h3b0cab5e),
	.w3(32'h3b316624),
	.w4(32'h3bce383f),
	.w5(32'hbb98589a),
	.w6(32'h3b1555af),
	.w7(32'hbb5d6c4e),
	.w8(32'hbc26e171),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace0ad),
	.w1(32'h3a566776),
	.w2(32'h3b0e42bf),
	.w3(32'h3bb862e6),
	.w4(32'hbb851553),
	.w5(32'h3c1c5a95),
	.w6(32'hbba199a1),
	.w7(32'h3a81d01a),
	.w8(32'hba867862),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c67d),
	.w1(32'hbb275b9e),
	.w2(32'hbbab5ce1),
	.w3(32'h3aa1ee23),
	.w4(32'hba88d619),
	.w5(32'hbc14c58e),
	.w6(32'hbb2a68fd),
	.w7(32'hbb5f7624),
	.w8(32'hbb0f119d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb86da),
	.w1(32'hb947276a),
	.w2(32'h38938f57),
	.w3(32'hbbf5c7c1),
	.w4(32'hbacb0e22),
	.w5(32'hbb9b3697),
	.w6(32'hbb8a24df),
	.w7(32'hba7bb2a8),
	.w8(32'hbb1550b7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cab08),
	.w1(32'h3b013526),
	.w2(32'hb9744ffa),
	.w3(32'hba6d3dd8),
	.w4(32'h3b5be2fb),
	.w5(32'h3be8b5ec),
	.w6(32'hbb1d965a),
	.w7(32'h3b148313),
	.w8(32'hb9999f49),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf5ad7),
	.w1(32'h393f42d1),
	.w2(32'h3bed0ec9),
	.w3(32'hbba414c7),
	.w4(32'hbb475dc5),
	.w5(32'h3bb41803),
	.w6(32'hbb8d29b3),
	.w7(32'hbb0db117),
	.w8(32'h3b908c5c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6448b),
	.w1(32'h3c104f9e),
	.w2(32'h3ab7a2c8),
	.w3(32'h3be4c9a1),
	.w4(32'hba269e04),
	.w5(32'hbba1ba6f),
	.w6(32'h3b8af94a),
	.w7(32'h3c0511d0),
	.w8(32'hbaf6de5f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8285a56),
	.w1(32'hbba73158),
	.w2(32'hbb61496c),
	.w3(32'hbbf8112b),
	.w4(32'h3b7b32da),
	.w5(32'h39ce9180),
	.w6(32'hbbb599a8),
	.w7(32'hbb326e54),
	.w8(32'h38d5f4aa),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15c774),
	.w1(32'hb8bda07f),
	.w2(32'h3b17c009),
	.w3(32'hbb46a746),
	.w4(32'hbbf65d94),
	.w5(32'h3b9b47f9),
	.w6(32'hba938b89),
	.w7(32'hbc0d63d0),
	.w8(32'h3afe1c28),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbf4f8),
	.w1(32'hbc0591a3),
	.w2(32'hba4f84bd),
	.w3(32'hbbd1b2fd),
	.w4(32'hbc1b5b77),
	.w5(32'hba8fad62),
	.w6(32'h39aa3a89),
	.w7(32'h3b0c7415),
	.w8(32'h3bb3b75f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd370f),
	.w1(32'h3b953eeb),
	.w2(32'h3c020728),
	.w3(32'hbb953e38),
	.w4(32'hbbc72e16),
	.w5(32'h3a7e8976),
	.w6(32'hbba86cb5),
	.w7(32'hbb7bda86),
	.w8(32'hbbb1f3ba),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2216b0),
	.w1(32'h3b74adc9),
	.w2(32'h3af23ef1),
	.w3(32'h3b8d13d4),
	.w4(32'h3b927df7),
	.w5(32'hbb6f4c0d),
	.w6(32'h3981c6e5),
	.w7(32'h3a9699f3),
	.w8(32'hbb490472),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35cf01),
	.w1(32'hbaf5d62f),
	.w2(32'h3c0050f5),
	.w3(32'hbb489e71),
	.w4(32'hbb82e9d5),
	.w5(32'h3c41192e),
	.w6(32'h3b1e2a37),
	.w7(32'hbb12a19b),
	.w8(32'hbb4a6fb6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d97e1),
	.w1(32'h3a8dea0c),
	.w2(32'hba70b409),
	.w3(32'h3b89926c),
	.w4(32'h3aafe049),
	.w5(32'hba695bc2),
	.w6(32'h3ba7f9e1),
	.w7(32'hbb00580c),
	.w8(32'hb9702b09),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca78c5),
	.w1(32'hbc42f49a),
	.w2(32'hbb99d8cf),
	.w3(32'hbb1b36a7),
	.w4(32'hbba7eb8a),
	.w5(32'hbbcf9571),
	.w6(32'h3b301537),
	.w7(32'hba12f05a),
	.w8(32'hbb80a74e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5db632),
	.w1(32'h3c1e3b58),
	.w2(32'h39a1485b),
	.w3(32'h3c4e8523),
	.w4(32'h3b8e746f),
	.w5(32'h3bd4f5a3),
	.w6(32'hbaf7abe5),
	.w7(32'hbbf70014),
	.w8(32'h3b02ea0d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35507f),
	.w1(32'h3b95634d),
	.w2(32'h3bf0dd5b),
	.w3(32'h3b011c7f),
	.w4(32'h3c1df3ca),
	.w5(32'hbbca312a),
	.w6(32'h3c62aa8e),
	.w7(32'h3b5f83ed),
	.w8(32'h3af68e72),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a51b9),
	.w1(32'hbc4ad032),
	.w2(32'hbbc3cfc9),
	.w3(32'hbc21874a),
	.w4(32'hbc05128f),
	.w5(32'h3b8ff643),
	.w6(32'hbb277d63),
	.w7(32'hbb2a1495),
	.w8(32'hbb329493),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86d879),
	.w1(32'hbc165cc5),
	.w2(32'hbc01519f),
	.w3(32'h3c2078fb),
	.w4(32'hbc00eea0),
	.w5(32'hbc7112d4),
	.w6(32'hbb3265f2),
	.w7(32'hbb217310),
	.w8(32'hbc3e952b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58b092),
	.w1(32'h3b649195),
	.w2(32'hbbdd5300),
	.w3(32'hbb92c0d7),
	.w4(32'hbbc10cfb),
	.w5(32'hbbd9cd50),
	.w6(32'hbbd5c9e1),
	.w7(32'h3c2e81c4),
	.w8(32'h3aef403a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b206e),
	.w1(32'h3bab9dfc),
	.w2(32'hb9e506a3),
	.w3(32'hbb58f729),
	.w4(32'h3c332ec2),
	.w5(32'h3919853b),
	.w6(32'h3c292dc6),
	.w7(32'h3c5292be),
	.w8(32'h3c7e8490),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb95bd),
	.w1(32'h3b8e3876),
	.w2(32'h3b41d304),
	.w3(32'h3b771707),
	.w4(32'h3ba82e37),
	.w5(32'h3ba3a6ef),
	.w6(32'h3c0fef65),
	.w7(32'h3b1a79e5),
	.w8(32'h3bcf3211),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8eca9),
	.w1(32'hb7b140e9),
	.w2(32'hbb88e1d0),
	.w3(32'h3b1a927b),
	.w4(32'hba19e956),
	.w5(32'hbc1f0c64),
	.w6(32'h3a7cea2c),
	.w7(32'h39e73cdb),
	.w8(32'hb6603a6e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3528eb),
	.w1(32'hba180fd4),
	.w2(32'hba2b56e1),
	.w3(32'hbbdcd9c8),
	.w4(32'hbb98da3f),
	.w5(32'hbc1c628e),
	.w6(32'h3a985630),
	.w7(32'hbbbc4104),
	.w8(32'hba4ee756),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa891a9),
	.w1(32'h383fa9a8),
	.w2(32'h3b9eca78),
	.w3(32'h39ae4852),
	.w4(32'h3b632f76),
	.w5(32'h3c50f066),
	.w6(32'hbb4c8f9a),
	.w7(32'h3b9296d1),
	.w8(32'h3c20a0be),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6e36),
	.w1(32'h3aa51086),
	.w2(32'h3b83edeb),
	.w3(32'h3b6d7b01),
	.w4(32'h3a8b7efc),
	.w5(32'h3b96bcb0),
	.w6(32'h3bc2aa4f),
	.w7(32'hbad484ae),
	.w8(32'h3c28a9c2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0abb),
	.w1(32'h390190ec),
	.w2(32'hbbb4d233),
	.w3(32'hbc16b4fe),
	.w4(32'h3b4d96b3),
	.w5(32'hba45cd9a),
	.w6(32'hb8a5ebc2),
	.w7(32'h3c23e5c3),
	.w8(32'h3b324b20),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75f2e8),
	.w1(32'h3b517c40),
	.w2(32'hbb667baa),
	.w3(32'hbb8e1a5d),
	.w4(32'h3b90cfc6),
	.w5(32'hbb948b51),
	.w6(32'hbb02f7a2),
	.w7(32'h3bd4d16f),
	.w8(32'hbb05e6ab),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed3db1),
	.w1(32'hba27e3bc),
	.w2(32'h3b28ec13),
	.w3(32'hbbb124fe),
	.w4(32'hbbd0a3b7),
	.w5(32'hbbe22be3),
	.w6(32'hbb304e41),
	.w7(32'hbb7a2997),
	.w8(32'hbb7fde6c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44cc60),
	.w1(32'h3b918a5b),
	.w2(32'hbb1e3497),
	.w3(32'h3c85c7c1),
	.w4(32'h3bb01569),
	.w5(32'hbbc38f9d),
	.w6(32'h3c4903e0),
	.w7(32'h3c188312),
	.w8(32'hba5ef629),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedc295),
	.w1(32'hba379a8b),
	.w2(32'h3b710c30),
	.w3(32'hbb2d7461),
	.w4(32'hbb08b1c3),
	.w5(32'h39eaeaa3),
	.w6(32'hba145afc),
	.w7(32'hbb435f13),
	.w8(32'h3a0d3ad6),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ebd61),
	.w1(32'h3bbcf9dd),
	.w2(32'h3b81d4f0),
	.w3(32'h3b491181),
	.w4(32'hbc0ffe55),
	.w5(32'hbb71e952),
	.w6(32'h3b17c52e),
	.w7(32'h3a001fc5),
	.w8(32'hbb22bea9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5448fc),
	.w1(32'hb7c0bd5e),
	.w2(32'h3baa0cda),
	.w3(32'h3b57dec6),
	.w4(32'h3ac35ad1),
	.w5(32'h3bd0dae3),
	.w6(32'hbba912b9),
	.w7(32'hba83ad94),
	.w8(32'h3b46780f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5667d4),
	.w1(32'h3c3b8458),
	.w2(32'h3c32895e),
	.w3(32'h3c11fd8c),
	.w4(32'h3b171bf6),
	.w5(32'h3ba0d4fa),
	.w6(32'h3b5a228a),
	.w7(32'hbb463a97),
	.w8(32'h3bbdd400),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a3c66),
	.w1(32'h3b427246),
	.w2(32'h3aa5a5ad),
	.w3(32'h3b521add),
	.w4(32'hbb768e6c),
	.w5(32'h395b1624),
	.w6(32'h3beff65d),
	.w7(32'h3b913023),
	.w8(32'hbb32a5a4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be42d2d),
	.w1(32'hbbb51aad),
	.w2(32'h3c324afe),
	.w3(32'hbb8ee8ca),
	.w4(32'hbc8f4c22),
	.w5(32'h3bd6a9ec),
	.w6(32'h3aa81241),
	.w7(32'hbc487327),
	.w8(32'hbc086012),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07d2aa),
	.w1(32'h3ae0006e),
	.w2(32'hb9c101c6),
	.w3(32'h3c8773a7),
	.w4(32'hbb016942),
	.w5(32'hbbd41e39),
	.w6(32'h3ab62704),
	.w7(32'hbb1d3be8),
	.w8(32'hbb11fe3c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9b129),
	.w1(32'h39d78779),
	.w2(32'h3bd2c17e),
	.w3(32'h3b80881a),
	.w4(32'h3a304ef0),
	.w5(32'h3b0b6b84),
	.w6(32'h3ac3f495),
	.w7(32'hba527a26),
	.w8(32'h3ada9765),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad15f09),
	.w1(32'h3a9e7bcf),
	.w2(32'h3bb5c0c9),
	.w3(32'hbb1e722e),
	.w4(32'hbca3fad2),
	.w5(32'hbc1c869e),
	.w6(32'h3c1b4098),
	.w7(32'hbb854f9c),
	.w8(32'hbc25482b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bd463),
	.w1(32'h3bc9d377),
	.w2(32'hbb373519),
	.w3(32'h3c8a8097),
	.w4(32'h3c5dbe4f),
	.w5(32'hbb7c131e),
	.w6(32'h3c8d676c),
	.w7(32'hba71f6c9),
	.w8(32'hbb5161aa),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba43efe),
	.w1(32'h3b043215),
	.w2(32'h3b72341f),
	.w3(32'hbc84d401),
	.w4(32'hbbc4391b),
	.w5(32'h3a8fff10),
	.w6(32'h3a889c84),
	.w7(32'hbbe5fcbb),
	.w8(32'h3ae82845),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24fd34),
	.w1(32'hbb93e0e2),
	.w2(32'h3bc50863),
	.w3(32'hbba8d1b1),
	.w4(32'h3ae1729b),
	.w5(32'h3cbc9b6e),
	.w6(32'h3b16e3ca),
	.w7(32'h3b9d3b70),
	.w8(32'h3c775c4b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7651),
	.w1(32'h3b0f2dfc),
	.w2(32'h3c1336e7),
	.w3(32'h3b8a616f),
	.w4(32'hbc578d9c),
	.w5(32'hbc77dfa1),
	.w6(32'h3bde60b9),
	.w7(32'hbc321231),
	.w8(32'hbc04378a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca76684),
	.w1(32'hbbb4daae),
	.w2(32'hbaca6037),
	.w3(32'h3c5cf648),
	.w4(32'hbbd97037),
	.w5(32'h3a0aa09e),
	.w6(32'h3b6dedd6),
	.w7(32'hba733749),
	.w8(32'hbc0dfdf0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae2719),
	.w1(32'h3ccb5970),
	.w2(32'h3cca2599),
	.w3(32'h3ca8c7be),
	.w4(32'h3c8b454f),
	.w5(32'h3c65663b),
	.w6(32'h3c2da9cd),
	.w7(32'h3bb9d2b9),
	.w8(32'h3c38926e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5d039),
	.w1(32'hbb7d18f7),
	.w2(32'h3b850fe5),
	.w3(32'h3b5950ac),
	.w4(32'hbc1bd844),
	.w5(32'h3b44cf5c),
	.w6(32'h3c054a5c),
	.w7(32'hbbd53271),
	.w8(32'h3b9361ea),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1861),
	.w1(32'h3a1cda7f),
	.w2(32'hbc24e3c8),
	.w3(32'h3aeac595),
	.w4(32'h3ba28b58),
	.w5(32'hbb20a75c),
	.w6(32'h39938214),
	.w7(32'h39af5a83),
	.w8(32'hba08aaf6),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf1d9a),
	.w1(32'hba065179),
	.w2(32'h3816f863),
	.w3(32'hbba0da70),
	.w4(32'hb7d2e9ec),
	.w5(32'h39f30a72),
	.w6(32'hb9cf1f69),
	.w7(32'h3bece458),
	.w8(32'h3a201cb8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8432e2),
	.w1(32'hbbf58b56),
	.w2(32'h3b08db4f),
	.w3(32'h3b6719a6),
	.w4(32'hbb8f7506),
	.w5(32'h3c2d6dff),
	.w6(32'hbafddbbb),
	.w7(32'h3b2894a2),
	.w8(32'h3a4beee2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e09f1),
	.w1(32'hbb8da402),
	.w2(32'h3c3ec350),
	.w3(32'hbb80012d),
	.w4(32'hbb9cf419),
	.w5(32'h3d0cfcd7),
	.w6(32'hbae7fc28),
	.w7(32'hbc5773f7),
	.w8(32'hbb199b48),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39244cb1),
	.w1(32'h3ad9547a),
	.w2(32'h3b45d0b2),
	.w3(32'h3c82aad4),
	.w4(32'hbc1b979d),
	.w5(32'hbb5b2b65),
	.w6(32'h3bfe3640),
	.w7(32'hbb50f01e),
	.w8(32'h3a93d615),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73e5d7),
	.w1(32'hbb4dcd79),
	.w2(32'hbaf9089e),
	.w3(32'h3b677917),
	.w4(32'hba82510b),
	.w5(32'h3bbde0dd),
	.w6(32'h3a59d81a),
	.w7(32'hb988beaf),
	.w8(32'h3aaddaa6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1cce7),
	.w1(32'hbb858e99),
	.w2(32'hba1a3a14),
	.w3(32'h399e4370),
	.w4(32'h385453b1),
	.w5(32'hb95fb117),
	.w6(32'h3bc228d4),
	.w7(32'hbb7fb84c),
	.w8(32'hb999907c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8760e),
	.w1(32'hb932ab02),
	.w2(32'hbc4f4744),
	.w3(32'h3c13e248),
	.w4(32'h3c901b5a),
	.w5(32'h3aec9a05),
	.w6(32'h3c6330df),
	.w7(32'h3b138942),
	.w8(32'h3c076d48),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2952bf),
	.w1(32'hbbf4df3c),
	.w2(32'hbb09dbc8),
	.w3(32'hbc8b3514),
	.w4(32'h3ac1417f),
	.w5(32'hbc1f5837),
	.w6(32'h3bdb3520),
	.w7(32'h3be61dbc),
	.w8(32'hbb52e2e6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34a1cf),
	.w1(32'h391aa87f),
	.w2(32'h3bed32b0),
	.w3(32'hbc06e21f),
	.w4(32'hbb2722bd),
	.w5(32'h3b8647bf),
	.w6(32'hbb6eb5a5),
	.w7(32'hbb62caa7),
	.w8(32'h3a0590ed),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b948917),
	.w1(32'hbae34290),
	.w2(32'h3c1ae4eb),
	.w3(32'h3c07960b),
	.w4(32'h3b7011cc),
	.w5(32'h3c9606f0),
	.w6(32'h3b3fdf3f),
	.w7(32'hbb65a661),
	.w8(32'h3b127b68),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc03050),
	.w1(32'h3c0bf664),
	.w2(32'h3b228a5e),
	.w3(32'h3a16d805),
	.w4(32'h3c113395),
	.w5(32'h3bd36c0c),
	.w6(32'h3b039efb),
	.w7(32'h3b72cba1),
	.w8(32'h3c50083a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0effd1),
	.w1(32'hba4be4e2),
	.w2(32'hba909022),
	.w3(32'h3b37ef49),
	.w4(32'hbbf6787a),
	.w5(32'hbb6edba7),
	.w6(32'h3c312e6b),
	.w7(32'hbbb55ffd),
	.w8(32'hbbfabc7b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e0d76),
	.w1(32'h3bd5ff43),
	.w2(32'h3c3af9de),
	.w3(32'h3b44ad67),
	.w4(32'hbbeddf04),
	.w5(32'h3ce0f7b3),
	.w6(32'hba9637e9),
	.w7(32'hbc77b6df),
	.w8(32'hbbc6b900),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb27fdc1),
	.w1(32'h384f3e1d),
	.w2(32'h3a07308d),
	.w3(32'h3c92884c),
	.w4(32'hb9bc861c),
	.w5(32'hbb77af23),
	.w6(32'h3bda6cb9),
	.w7(32'hba6f118a),
	.w8(32'hbb8986bb),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdb5fc),
	.w1(32'h3b2d95e3),
	.w2(32'hbb52d126),
	.w3(32'h3bf5a8d0),
	.w4(32'hba2b1971),
	.w5(32'hbb884679),
	.w6(32'h3b8437b1),
	.w7(32'h3bc60c00),
	.w8(32'h3aded42d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa343e8),
	.w1(32'hbaa0b860),
	.w2(32'h3973d406),
	.w3(32'hbbb6812e),
	.w4(32'hbb9ea475),
	.w5(32'hbbc35d74),
	.w6(32'hbb50cce3),
	.w7(32'h3b783d96),
	.w8(32'h3b9fd2c0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafef513),
	.w1(32'hbb21f2f0),
	.w2(32'hbb019116),
	.w3(32'hbb807379),
	.w4(32'h3bb28a49),
	.w5(32'h3c4c7efc),
	.w6(32'hbb4ba744),
	.w7(32'h3b80ec28),
	.w8(32'h3b8b0407),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8f857),
	.w1(32'hbbba39ca),
	.w2(32'hbbb812cc),
	.w3(32'h3b45e8ef),
	.w4(32'h3b027528),
	.w5(32'h3c8db78d),
	.w6(32'h3a672a79),
	.w7(32'h3bff3e8e),
	.w8(32'h3bd502e2),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ef64c),
	.w1(32'h3a42a1c5),
	.w2(32'hbb514fca),
	.w3(32'hbc354fa4),
	.w4(32'h3b02e2b4),
	.w5(32'hbb81ffd3),
	.w6(32'h3a409252),
	.w7(32'hbc19372d),
	.w8(32'hbbed2712),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa775ac),
	.w1(32'hbb7afaea),
	.w2(32'h3ba0af71),
	.w3(32'h3b7c2e3c),
	.w4(32'hbc273daa),
	.w5(32'hbb227739),
	.w6(32'h3b538c8f),
	.w7(32'hbbf7f002),
	.w8(32'hbba8a68b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab49133),
	.w1(32'h3aac72ea),
	.w2(32'h3c2e1d4e),
	.w3(32'h3ba63347),
	.w4(32'hbb958ec9),
	.w5(32'h3b4314db),
	.w6(32'h3b855551),
	.w7(32'hbb3ec8d6),
	.w8(32'h39c12211),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c785355),
	.w1(32'h39cdc464),
	.w2(32'hba86fe15),
	.w3(32'h3be1ecb1),
	.w4(32'hbb0d87aa),
	.w5(32'hbbb9e453),
	.w6(32'h3b0a0587),
	.w7(32'hba133231),
	.w8(32'hbb43c8c3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb88c5),
	.w1(32'hbb07ba68),
	.w2(32'hbbb41980),
	.w3(32'h3b597a2b),
	.w4(32'hbab9ef1c),
	.w5(32'hbb1a7fca),
	.w6(32'h3b7f89f5),
	.w7(32'hbb555d40),
	.w8(32'hbb4a4a1c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beaeb22),
	.w1(32'h3a7c3e13),
	.w2(32'h3babd179),
	.w3(32'h3b6aa7e3),
	.w4(32'hbc093201),
	.w5(32'h3ceae701),
	.w6(32'h3ba075a1),
	.w7(32'hbca7c45c),
	.w8(32'hb9ce856b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d4963),
	.w1(32'h3ad3244a),
	.w2(32'h3a2dd9d1),
	.w3(32'hba813b0b),
	.w4(32'h3bd7bd2b),
	.w5(32'hbbb31b48),
	.w6(32'h3be39bfd),
	.w7(32'h3ba624e2),
	.w8(32'h3b803096),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a48039),
	.w1(32'hbb9eab21),
	.w2(32'hbb8252c0),
	.w3(32'hbbcb82f5),
	.w4(32'hbaeb63bb),
	.w5(32'h3bb2c0ab),
	.w6(32'h3b6d5d95),
	.w7(32'hbb105fea),
	.w8(32'hbb9a3e89),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebbd8b),
	.w1(32'hba600a1e),
	.w2(32'h3ae80e7d),
	.w3(32'h3ae4b274),
	.w4(32'h3a8527b4),
	.w5(32'hbb8578a3),
	.w6(32'h3b201111),
	.w7(32'h3c173262),
	.w8(32'hb7e787f8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e8976),
	.w1(32'h3bc79886),
	.w2(32'h3bcc595e),
	.w3(32'h3bb3ba21),
	.w4(32'hbbaa5a55),
	.w5(32'hbbb6452b),
	.w6(32'h3bbb712e),
	.w7(32'hba00283c),
	.w8(32'hbb22f1ca),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169a19),
	.w1(32'h3b843646),
	.w2(32'h3b9e6498),
	.w3(32'h3bdc0cbd),
	.w4(32'hba593caf),
	.w5(32'h3ad23227),
	.w6(32'h3b851877),
	.w7(32'hba3b3a80),
	.w8(32'h3ade6278),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a2d0f),
	.w1(32'hba56b416),
	.w2(32'hbbc440fa),
	.w3(32'h3afcad8c),
	.w4(32'h3acc791f),
	.w5(32'hbbd650fe),
	.w6(32'h3bce0c42),
	.w7(32'hba9d0d63),
	.w8(32'hbc3305f5),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea62ba),
	.w1(32'h3bc0d512),
	.w2(32'h3b96495b),
	.w3(32'h3bd09adb),
	.w4(32'h3aaef8ec),
	.w5(32'hbbbf64da),
	.w6(32'hba374b18),
	.w7(32'h3b6e6f1c),
	.w8(32'hbbefb590),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1846e8),
	.w1(32'hbc138c4c),
	.w2(32'hba986758),
	.w3(32'hbb279232),
	.w4(32'hbc06eb95),
	.w5(32'hbb4a54c9),
	.w6(32'h3a958d17),
	.w7(32'hbae11df1),
	.w8(32'hbbd1c434),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a9c55),
	.w1(32'hbaa8c13f),
	.w2(32'h3b107497),
	.w3(32'h3bd48029),
	.w4(32'hbb42b45c),
	.w5(32'h3b9978d4),
	.w6(32'h3aac695e),
	.w7(32'hbb5d7926),
	.w8(32'h3ac8fd83),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb51e79),
	.w1(32'hba760b76),
	.w2(32'hba23efa1),
	.w3(32'h3a603647),
	.w4(32'hbbe9b87a),
	.w5(32'hbbf9f1a0),
	.w6(32'h3b495988),
	.w7(32'hbc153f6e),
	.w8(32'hbc11cce7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a318893),
	.w1(32'hba018261),
	.w2(32'h3be350b0),
	.w3(32'h3aee252a),
	.w4(32'hbbfa6d29),
	.w5(32'h3bf33385),
	.w6(32'hba03f06b),
	.w7(32'h3b6a5f8b),
	.w8(32'h3c460af3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6320b0),
	.w1(32'hba870ebc),
	.w2(32'h3a2ad7ae),
	.w3(32'h380c0b04),
	.w4(32'h3af2925d),
	.w5(32'h3cc2c166),
	.w6(32'h3a911123),
	.w7(32'hbac81af3),
	.w8(32'h3ada73c8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c1874),
	.w1(32'hb9ad1699),
	.w2(32'h3b16478c),
	.w3(32'hbbabfe89),
	.w4(32'hba984d90),
	.w5(32'h3b8cb32c),
	.w6(32'hb7c70a32),
	.w7(32'hbbc840e8),
	.w8(32'h3b4c0550),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dcf41),
	.w1(32'hbb6ad6c5),
	.w2(32'hbacad138),
	.w3(32'h3b08b286),
	.w4(32'hb9900e13),
	.w5(32'h3bb23342),
	.w6(32'h3b4f7afe),
	.w7(32'h3baf11dd),
	.w8(32'h3b412051),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0867f),
	.w1(32'h3b2e38b5),
	.w2(32'h3ab1f3e5),
	.w3(32'h3b746a49),
	.w4(32'hbac82030),
	.w5(32'hbb91833b),
	.w6(32'hbad6222b),
	.w7(32'h39a534ce),
	.w8(32'hb909aea0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3984af2d),
	.w1(32'hbb690d50),
	.w2(32'hbb7482fb),
	.w3(32'hbb0c45ea),
	.w4(32'hb97b7bc0),
	.w5(32'hbabf251c),
	.w6(32'h3b61801b),
	.w7(32'h3b6d156a),
	.w8(32'hbab863a7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cdecf),
	.w1(32'h3ad9e788),
	.w2(32'h3badbbbc),
	.w3(32'hbaedca87),
	.w4(32'hbb2cadf1),
	.w5(32'h3bc0fd14),
	.w6(32'hbb677d18),
	.w7(32'h3ac2332a),
	.w8(32'hbb663450),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91c04e),
	.w1(32'h3b9a6f1b),
	.w2(32'h3a94a9a2),
	.w3(32'h3bcb1724),
	.w4(32'h3b8742ef),
	.w5(32'hba460b6d),
	.w6(32'h3b598eaf),
	.w7(32'h3bd5a267),
	.w8(32'h3b80bcea),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fdc7),
	.w1(32'hbb51820f),
	.w2(32'hbb27263b),
	.w3(32'h3a9c0cc6),
	.w4(32'h3a6ae505),
	.w5(32'hbbf6df87),
	.w6(32'h3bdd6e2f),
	.w7(32'h3b9f419e),
	.w8(32'h3ae6bb0e),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f6c13),
	.w1(32'hbc071f9a),
	.w2(32'hbb2c1947),
	.w3(32'hbb925ac4),
	.w4(32'hbb26e1ca),
	.w5(32'hbb547028),
	.w6(32'hbaeb04cc),
	.w7(32'hba5e4c41),
	.w8(32'h39016bf8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02a787),
	.w1(32'h3bd6bf4d),
	.w2(32'h3b2bd51f),
	.w3(32'hbb174dd9),
	.w4(32'h3b19a911),
	.w5(32'h3b01b0ff),
	.w6(32'hbb76f391),
	.w7(32'h3bcf5019),
	.w8(32'h3b26905a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4aa5e6),
	.w1(32'hbbb9e400),
	.w2(32'hbae4a3b5),
	.w3(32'h3b1dc46c),
	.w4(32'hbc2c880a),
	.w5(32'h3ac22fde),
	.w6(32'hbb9f0f6a),
	.w7(32'h3b2a87b3),
	.w8(32'h3a7867dd),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e905a),
	.w1(32'h3af06c5f),
	.w2(32'hbb98235a),
	.w3(32'h3aceba23),
	.w4(32'hbba6fee5),
	.w5(32'hbc72d491),
	.w6(32'h39a9c1e0),
	.w7(32'h3b3080f4),
	.w8(32'hbb7b7568),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fb397),
	.w1(32'hbace4cdc),
	.w2(32'hbbae3007),
	.w3(32'hbc10083e),
	.w4(32'hbb00eff3),
	.w5(32'hbc4e03da),
	.w6(32'hbc0b074a),
	.w7(32'hbb82c03b),
	.w8(32'hbb9ffd4a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6f6e),
	.w1(32'h3a11c81e),
	.w2(32'h3ae9c919),
	.w3(32'hbb988c5e),
	.w4(32'hbad52aa0),
	.w5(32'hbb1f4c3d),
	.w6(32'hbb48abdb),
	.w7(32'h3b726c89),
	.w8(32'hb9afe1c4),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdc48a),
	.w1(32'hbbf75fae),
	.w2(32'h3b1f9178),
	.w3(32'h3a580f98),
	.w4(32'hbbf8dc7b),
	.w5(32'hbbadc147),
	.w6(32'hba862d61),
	.w7(32'h3a3b94c7),
	.w8(32'h3ba60436),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999a644),
	.w1(32'hb9c97837),
	.w2(32'h3aa517a7),
	.w3(32'h3af4d4b3),
	.w4(32'hba058dd2),
	.w5(32'hbb299f32),
	.w6(32'h39a0b841),
	.w7(32'h3b0a7193),
	.w8(32'h3af93518),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93a737),
	.w1(32'h3bbfb51c),
	.w2(32'h3be0687d),
	.w3(32'h3bdbf160),
	.w4(32'hbaeb4c8b),
	.w5(32'hbb8e8670),
	.w6(32'h3b01d0bb),
	.w7(32'hbafb127b),
	.w8(32'hbacf6976),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb056f),
	.w1(32'h3bbcb4e3),
	.w2(32'h3c02a9df),
	.w3(32'hb9c37559),
	.w4(32'h3bad4c9b),
	.w5(32'h3d0dd4ca),
	.w6(32'hbb13ed5c),
	.w7(32'hbb8dc4ec),
	.w8(32'h3c04cfa0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd215),
	.w1(32'h3bc0f888),
	.w2(32'h3b2d0b6b),
	.w3(32'h3c108074),
	.w4(32'h39f57d22),
	.w5(32'hba8d3ac4),
	.w6(32'h3beb7eaf),
	.w7(32'h3c0feb0e),
	.w8(32'hbab2a8cf),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb199f),
	.w1(32'hbbaa3ddf),
	.w2(32'h3910725a),
	.w3(32'h3a90a91e),
	.w4(32'hbbd5dec2),
	.w5(32'hbc19c70b),
	.w6(32'h3b5d351d),
	.w7(32'h3a3219f7),
	.w8(32'hbbaa8de3),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3739ec),
	.w1(32'hbbd6b934),
	.w2(32'hbb8104a5),
	.w3(32'h3bf6fa90),
	.w4(32'hbc52ee03),
	.w5(32'hbc9e07dd),
	.w6(32'h3a2f5c45),
	.w7(32'h3b3fea98),
	.w8(32'hbbaad423),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32ab04),
	.w1(32'hba0b1c1e),
	.w2(32'hbbc97cf6),
	.w3(32'hbc3e1718),
	.w4(32'h3a8fc424),
	.w5(32'hbc64f1ac),
	.w6(32'hbbc3bba2),
	.w7(32'h3bc243a0),
	.w8(32'hbad1e4b1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d17a2),
	.w1(32'hbbd4b843),
	.w2(32'hbb905947),
	.w3(32'hbc70f261),
	.w4(32'hba8a0f7b),
	.w5(32'hbb8817ee),
	.w6(32'hbb5bd835),
	.w7(32'h3c2a2df5),
	.w8(32'hbb7569a6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49e0b0),
	.w1(32'hba696ad9),
	.w2(32'hbb13356f),
	.w3(32'hbc15ceaf),
	.w4(32'h3b52f154),
	.w5(32'h3c526569),
	.w6(32'hbbae1a4b),
	.w7(32'hb94c5665),
	.w8(32'h3b4c8a1d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e9305),
	.w1(32'h3a4be188),
	.w2(32'h3c27ed7b),
	.w3(32'h3b7635be),
	.w4(32'hbbd9ce41),
	.w5(32'h3c8780f3),
	.w6(32'h3b9e9d09),
	.w7(32'hbc2ff40c),
	.w8(32'hbc002bb8),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf173b),
	.w1(32'h3b336639),
	.w2(32'h3b841e10),
	.w3(32'h3c81cd17),
	.w4(32'h3b8c7a40),
	.w5(32'hbba67a62),
	.w6(32'h3bf6199d),
	.w7(32'h3bdcb57b),
	.w8(32'h3b2bc0ab),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cd3d1),
	.w1(32'hbbacd9a6),
	.w2(32'h3bfdc4e7),
	.w3(32'h3bab8a03),
	.w4(32'hbc5f06aa),
	.w5(32'hbb996c7c),
	.w6(32'h3bee201e),
	.w7(32'hbc4b4307),
	.w8(32'hbbff6199),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c057866),
	.w1(32'h3b20f3a8),
	.w2(32'h3bcb3c70),
	.w3(32'h3c2bbb36),
	.w4(32'h3b8186cb),
	.w5(32'h3c04a413),
	.w6(32'hbbadc85b),
	.w7(32'h3ae3130a),
	.w8(32'h3b18f255),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5464a4),
	.w1(32'hbb583eeb),
	.w2(32'hbb1ef8e8),
	.w3(32'h3a4c5a1a),
	.w4(32'hbba726ac),
	.w5(32'hbb8c8555),
	.w6(32'hbaefa605),
	.w7(32'hbba5b931),
	.w8(32'hbb9fd77e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb217d88),
	.w1(32'h3b5ad66c),
	.w2(32'h3b63d0e7),
	.w3(32'hbb814c5a),
	.w4(32'h3aaae276),
	.w5(32'h38b464ef),
	.w6(32'hbb3ccabe),
	.w7(32'h3b6fab96),
	.w8(32'h3a6fabcb),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c798794),
	.w1(32'h3bb5b2a1),
	.w2(32'h3be6abb0),
	.w3(32'h3c6ddc7a),
	.w4(32'h3781a29e),
	.w5(32'h3bb57a96),
	.w6(32'h3beec6c2),
	.w7(32'h3b876753),
	.w8(32'h3a871067),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc4c0d),
	.w1(32'h3bba482a),
	.w2(32'h3c20765d),
	.w3(32'h3beeae10),
	.w4(32'hbab5ed67),
	.w5(32'h3c263ef9),
	.w6(32'hb7d01e7b),
	.w7(32'hbbe60bee),
	.w8(32'h3b0b3146),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2330e8),
	.w1(32'h3afc9e88),
	.w2(32'h3b892630),
	.w3(32'h3c8d6311),
	.w4(32'hbb1e4709),
	.w5(32'hbb53b376),
	.w6(32'h3c44e8b8),
	.w7(32'hbb316062),
	.w8(32'hba12f4ab),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa119cc),
	.w1(32'h3b535549),
	.w2(32'h3c0436e1),
	.w3(32'h3afa148c),
	.w4(32'hbb9bc8d1),
	.w5(32'h3be8e259),
	.w6(32'hb99b475a),
	.w7(32'hbbc90fa5),
	.w8(32'hbac8dbac),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7c47c),
	.w1(32'hbc5ac1fa),
	.w2(32'hbc3e1d36),
	.w3(32'h3c3bc916),
	.w4(32'hbb1445cd),
	.w5(32'hbc8fee61),
	.w6(32'h3c3cef64),
	.w7(32'hb9514c61),
	.w8(32'hbbb65a00),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698f4f),
	.w1(32'h3c34e20c),
	.w2(32'h3c2f442b),
	.w3(32'hbc22a16b),
	.w4(32'h3c1438c1),
	.w5(32'h3ca0bcdc),
	.w6(32'hbbd0e8d5),
	.w7(32'hbadbe7b8),
	.w8(32'h3b9be332),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4840e8),
	.w1(32'hbbdfe4e8),
	.w2(32'hbb8a4bd8),
	.w3(32'h3c1a7eab),
	.w4(32'hbc00598d),
	.w5(32'hbb7f7444),
	.w6(32'h3c08291d),
	.w7(32'hbbdcd700),
	.w8(32'hbb59628d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba6abe),
	.w1(32'hb931027e),
	.w2(32'hbb511c87),
	.w3(32'hba6fe487),
	.w4(32'h3b02d458),
	.w5(32'hbb858cf0),
	.w6(32'hbad097e7),
	.w7(32'h3b063723),
	.w8(32'hbb7d6213),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2860b0),
	.w1(32'h3aefd877),
	.w2(32'h3b96955b),
	.w3(32'h3be6e6fb),
	.w4(32'h3b93af5a),
	.w5(32'hbac86d70),
	.w6(32'h3c067781),
	.w7(32'h3c14a647),
	.w8(32'h3a90f010),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a543332),
	.w1(32'hbb2a19e5),
	.w2(32'hbbd80cbd),
	.w3(32'h3b882870),
	.w4(32'hbb621a8b),
	.w5(32'hbc8c2995),
	.w6(32'h3abb7ad1),
	.w7(32'h3c0ea2f4),
	.w8(32'hbb9964c5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32c92),
	.w1(32'h3a8254f4),
	.w2(32'h3bcf614d),
	.w3(32'hbc26fb08),
	.w4(32'hbb09fb93),
	.w5(32'hb8f56667),
	.w6(32'hbc0c6791),
	.w7(32'hbba0d5f9),
	.w8(32'hbbc9f32e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e1fd5),
	.w1(32'hbc334faf),
	.w2(32'hbc1e21f7),
	.w3(32'h3c0e872f),
	.w4(32'hbc304ba7),
	.w5(32'hbaf1ce5e),
	.w6(32'h3b8e799b),
	.w7(32'hbaa46ddd),
	.w8(32'hbc35363e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b559c1b),
	.w1(32'h3afb1bbf),
	.w2(32'hbc024502),
	.w3(32'hbbbe62f7),
	.w4(32'hbb836ed6),
	.w5(32'hbb1bc1b4),
	.w6(32'hbbc2dcc5),
	.w7(32'h3bfa6150),
	.w8(32'h3b5f4405),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7bf96),
	.w1(32'h3aec5d97),
	.w2(32'h3bd4ca67),
	.w3(32'h3aecee81),
	.w4(32'h3b0803fb),
	.w5(32'h3ba2eef4),
	.w6(32'h3b1a2603),
	.w7(32'hbb4dae38),
	.w8(32'h3bc7c3b5),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16af4a),
	.w1(32'hba26fbab),
	.w2(32'hbbd65fc3),
	.w3(32'hbc4c30d6),
	.w4(32'hbbba2ebc),
	.w5(32'hbc37cf1b),
	.w6(32'hbb17171e),
	.w7(32'hbb2ac12a),
	.w8(32'hbc54fe48),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c128594),
	.w1(32'h3c0817e6),
	.w2(32'hba969237),
	.w3(32'h3aba9965),
	.w4(32'h3a91d717),
	.w5(32'h3b103bb1),
	.w6(32'hbb663f83),
	.w7(32'h3c066343),
	.w8(32'hbb6f1b83),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4a30),
	.w1(32'hbbba88ed),
	.w2(32'hbb85e4de),
	.w3(32'h3bff7f61),
	.w4(32'hbca98bf9),
	.w5(32'hbc577ae8),
	.w6(32'h3c44c507),
	.w7(32'h3bab6fd2),
	.w8(32'hbb67d71e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad81993),
	.w1(32'hbbbde4ee),
	.w2(32'h3b5239f5),
	.w3(32'h3c380879),
	.w4(32'hbba9baaa),
	.w5(32'h3c80a9c9),
	.w6(32'h3b126548),
	.w7(32'hbbc484c4),
	.w8(32'hbb1cb80e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0312a1),
	.w1(32'h3b7d5b98),
	.w2(32'hbb5a7d03),
	.w3(32'h3c05ab2d),
	.w4(32'h3b33976b),
	.w5(32'hbba382d5),
	.w6(32'h3b64450f),
	.w7(32'hb989b873),
	.w8(32'hbba46fff),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9fddb),
	.w1(32'hb98d5d83),
	.w2(32'h38b47e96),
	.w3(32'hbae45492),
	.w4(32'hbc06ecda),
	.w5(32'hb919ba60),
	.w6(32'hbb825b7f),
	.w7(32'hbba7d02b),
	.w8(32'hbba930b3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ec95b),
	.w1(32'h3ba54daf),
	.w2(32'hbbd1d58c),
	.w3(32'h3b1b0512),
	.w4(32'h3c7170cc),
	.w5(32'hb970b4ca),
	.w6(32'hbaccb98f),
	.w7(32'h3c5b0449),
	.w8(32'h3c0b2015),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb365762),
	.w1(32'h3a17edb7),
	.w2(32'h3c61f91e),
	.w3(32'hbab0357e),
	.w4(32'hba46ffe7),
	.w5(32'h3c828be7),
	.w6(32'h3ad17037),
	.w7(32'hbba03698),
	.w8(32'h3b36059b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46001a),
	.w1(32'hbb5f9b54),
	.w2(32'hba6c6807),
	.w3(32'h3c35f564),
	.w4(32'hbb887330),
	.w5(32'hbb4a7e3e),
	.w6(32'h3b3d7976),
	.w7(32'hbbdb17d2),
	.w8(32'h393348fd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc224125),
	.w1(32'hbb0e9b84),
	.w2(32'h3b99e9a0),
	.w3(32'hbacf08cd),
	.w4(32'hbb9772c8),
	.w5(32'hbba43282),
	.w6(32'hbab3a2e6),
	.w7(32'h3b8b79ba),
	.w8(32'h3aebaf6b),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd55a68),
	.w1(32'hbb84a5bc),
	.w2(32'hbb8845c7),
	.w3(32'h3c3baa5c),
	.w4(32'hbc2b7b7c),
	.w5(32'hbbbd6d03),
	.w6(32'h3bb1edcf),
	.w7(32'hbb993082),
	.w8(32'hbbe01284),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec2730),
	.w1(32'hbc112a67),
	.w2(32'h3b327fcf),
	.w3(32'h3afa13dc),
	.w4(32'hbc195fb3),
	.w5(32'h3b7c338d),
	.w6(32'h3c0007b7),
	.w7(32'hbb46b0b9),
	.w8(32'h3c11ae7b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b7a34),
	.w1(32'h3c72b277),
	.w2(32'h3c26e7fa),
	.w3(32'hbb4d25e8),
	.w4(32'h3c1f6587),
	.w5(32'h39a88bf8),
	.w6(32'h39ee99d4),
	.w7(32'hb95bc732),
	.w8(32'hbb987553),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3dfd7),
	.w1(32'h3c4b1e6a),
	.w2(32'h3b576b44),
	.w3(32'hbb14682f),
	.w4(32'h3c8467d3),
	.w5(32'h3c4fa7cf),
	.w6(32'hbb0979b6),
	.w7(32'h3c5a4daa),
	.w8(32'h3b914d9f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9c81),
	.w1(32'h3c18389f),
	.w2(32'h3b5cffc2),
	.w3(32'h3c2929b0),
	.w4(32'h3b6111d8),
	.w5(32'h3bf31dd3),
	.w6(32'h3b8b1b79),
	.w7(32'h3b3b2e0c),
	.w8(32'h3b831679),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8082),
	.w1(32'hbbd0a09a),
	.w2(32'hbb8e2b32),
	.w3(32'hbb462e25),
	.w4(32'hbb782fe2),
	.w5(32'hbb15cda1),
	.w6(32'hbb4a76df),
	.w7(32'hbb5fe152),
	.w8(32'hbbbc20a5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59964),
	.w1(32'h3a543e52),
	.w2(32'h3c27fb36),
	.w3(32'hb924ab34),
	.w4(32'hb9797a55),
	.w5(32'h3bff0a7c),
	.w6(32'hbbf31ab8),
	.w7(32'hbb041dfc),
	.w8(32'hbad062bf),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042467),
	.w1(32'hbbac06d8),
	.w2(32'hba95e8f0),
	.w3(32'hbb9ec1f0),
	.w4(32'hbb86d9e2),
	.w5(32'h387fa64f),
	.w6(32'hbb113f12),
	.w7(32'h3bd1a957),
	.w8(32'h3ae06e9e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9149c),
	.w1(32'h3bb76526),
	.w2(32'h3bca50d6),
	.w3(32'hbb9d5780),
	.w4(32'h3b2715a3),
	.w5(32'h3c2ebe8a),
	.w6(32'hbb1ba19d),
	.w7(32'h399cb958),
	.w8(32'h3bd44460),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ae267),
	.w1(32'hbc0d7afd),
	.w2(32'hbcad8248),
	.w3(32'h3b3d1966),
	.w4(32'hbbfd58c4),
	.w5(32'hbcaf09bb),
	.w6(32'h3b214bb5),
	.w7(32'hbbbf658a),
	.w8(32'hbbeae414),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb6248),
	.w1(32'hbb788c8f),
	.w2(32'h39d684fb),
	.w3(32'hbcb8bbd9),
	.w4(32'hbbd66e24),
	.w5(32'h3a3c2bb7),
	.w6(32'hbc9046bb),
	.w7(32'hbbde79fa),
	.w8(32'hbb68ca3b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3fcc9),
	.w1(32'hb918985a),
	.w2(32'h3ab7e33b),
	.w3(32'h3bfb5f3b),
	.w4(32'hbb846427),
	.w5(32'h39aff09a),
	.w6(32'h3b877d24),
	.w7(32'h3b42c392),
	.w8(32'hbb853e3f),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc14f3f),
	.w1(32'hbb37a877),
	.w2(32'h3b2e2e89),
	.w3(32'h3adef24c),
	.w4(32'h3ad7e4ff),
	.w5(32'h3c28b9e0),
	.w6(32'hbb007197),
	.w7(32'hbb18bf17),
	.w8(32'h3c25568e),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace9736),
	.w1(32'h3b9a85fe),
	.w2(32'h3b60114b),
	.w3(32'h3c145add),
	.w4(32'h3bd83dac),
	.w5(32'h3b9d59ee),
	.w6(32'h3c053b5d),
	.w7(32'h3be38652),
	.w8(32'h3b6e57c7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a659dc7),
	.w1(32'hbad3957f),
	.w2(32'hbbb3f13a),
	.w3(32'h39ccb22d),
	.w4(32'hbb537874),
	.w5(32'hbbc835f9),
	.w6(32'hb7b8ce61),
	.w7(32'hbbf596b2),
	.w8(32'hbc3581aa),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb868b31),
	.w1(32'hbb64d9f5),
	.w2(32'hbbd1138f),
	.w3(32'hbc1dcacf),
	.w4(32'h3b8582cb),
	.w5(32'hba639f92),
	.w6(32'hbc69efad),
	.w7(32'h3b550d59),
	.w8(32'h3b3add99),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb88daa),
	.w1(32'h3c28ae4a),
	.w2(32'h3ba18edd),
	.w3(32'h3bffb920),
	.w4(32'h3c317980),
	.w5(32'h3c267dde),
	.w6(32'h3c6363ca),
	.w7(32'h3c46c14f),
	.w8(32'h3c5814e4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dce34),
	.w1(32'h3be161f5),
	.w2(32'hba76c029),
	.w3(32'hba1ac118),
	.w4(32'h3bf03ece),
	.w5(32'h3ba0aa2c),
	.w6(32'h3bb54822),
	.w7(32'h39e0476c),
	.w8(32'h3b02ec50),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01f357),
	.w1(32'h3ba55ecd),
	.w2(32'hbb634ca4),
	.w3(32'hbb283b0c),
	.w4(32'h3ba3df40),
	.w5(32'h3b800a22),
	.w6(32'hb9e7ca7c),
	.w7(32'h3c92376e),
	.w8(32'h3c03b459),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92ac39),
	.w1(32'h3c3d5f46),
	.w2(32'h3b723b4d),
	.w3(32'h3b25137d),
	.w4(32'h3c87ab1e),
	.w5(32'h3caa8cc6),
	.w6(32'h3b8035ff),
	.w7(32'h3c99c573),
	.w8(32'h3c38c4f9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24913a),
	.w1(32'h3b198c4d),
	.w2(32'h3b1ff0e9),
	.w3(32'h3ba43214),
	.w4(32'hbacc8dfc),
	.w5(32'hbad0e69b),
	.w6(32'h3982c3ff),
	.w7(32'hbb2bff3f),
	.w8(32'hbae4418f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b1863),
	.w1(32'hbbeac1e3),
	.w2(32'h39c88a71),
	.w3(32'hbc285362),
	.w4(32'h3a6df599),
	.w5(32'h3b255a4e),
	.w6(32'h3ad11569),
	.w7(32'h39cf0766),
	.w8(32'h3b666b5f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b062816),
	.w1(32'h3baf8a0b),
	.w2(32'h3b9899ba),
	.w3(32'h3bb00e74),
	.w4(32'h3befbfe8),
	.w5(32'h3c114d05),
	.w6(32'h398d70fa),
	.w7(32'h3c54d196),
	.w8(32'h3c12b817),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e37a1),
	.w1(32'h3b7f720c),
	.w2(32'h3bba9985),
	.w3(32'h3bdf7e98),
	.w4(32'h3bd8f938),
	.w5(32'h3a912c39),
	.w6(32'h3c039136),
	.w7(32'h3b3feb4a),
	.w8(32'h3b1575bf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4b1f),
	.w1(32'hbc135780),
	.w2(32'hbabd533c),
	.w3(32'hba32785f),
	.w4(32'hbb2e73aa),
	.w5(32'h3bc7e663),
	.w6(32'hb9900213),
	.w7(32'hbb9ed061),
	.w8(32'h3ad1b291),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1608a),
	.w1(32'hbae1fd31),
	.w2(32'h3aa40f28),
	.w3(32'h3b75f3b5),
	.w4(32'hbb5cb2c3),
	.w5(32'h385e913f),
	.w6(32'h3b5203d9),
	.w7(32'h3b9bb915),
	.w8(32'h3a262974),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c94f),
	.w1(32'h3ba7122b),
	.w2(32'h3b824d42),
	.w3(32'hba8555e5),
	.w4(32'hbb8bceea),
	.w5(32'hbabcb673),
	.w6(32'hbb492c63),
	.w7(32'h3b337041),
	.w8(32'hbb4b87dc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25047d),
	.w1(32'hbccf3d23),
	.w2(32'hbc858925),
	.w3(32'hbb965f95),
	.w4(32'hbcb2dc39),
	.w5(32'hbc1e77a3),
	.w6(32'h3b21b72e),
	.w7(32'hbca0d6f6),
	.w8(32'hbc280267),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc66177b),
	.w1(32'hb9495f72),
	.w2(32'h3a5b0a02),
	.w3(32'hbb478794),
	.w4(32'hbaf0b756),
	.w5(32'h3c1332e4),
	.w6(32'hbc2fa7d6),
	.w7(32'h3b59fd3f),
	.w8(32'h3b61cc6a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4ef07),
	.w1(32'hbb2b8099),
	.w2(32'h3b4ab8d2),
	.w3(32'h3b9d8e95),
	.w4(32'hbad96921),
	.w5(32'h3b3478e9),
	.w6(32'h3afb48a6),
	.w7(32'hb9c2bd72),
	.w8(32'h3912d6c5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf37c71),
	.w1(32'h3bac57c1),
	.w2(32'h3c5e37cf),
	.w3(32'h3b8e09a4),
	.w4(32'hbba7001f),
	.w5(32'hb910a00b),
	.w6(32'h3b933c6f),
	.w7(32'h3b62a754),
	.w8(32'h3b8a7a38),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d706c),
	.w1(32'hbb8155bd),
	.w2(32'hbaf1835b),
	.w3(32'h3c19868f),
	.w4(32'h3a0a3039),
	.w5(32'hbb01794b),
	.w6(32'h3b9c86d4),
	.w7(32'hbb029225),
	.w8(32'h3b34ede2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b63b9),
	.w1(32'h3bc44a15),
	.w2(32'h3c0e1a18),
	.w3(32'hbb7848bb),
	.w4(32'h3bdc6a06),
	.w5(32'h3c437e2d),
	.w6(32'hbba43a71),
	.w7(32'h3b949285),
	.w8(32'h3ba7e547),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20bc64),
	.w1(32'hbb4cb9a4),
	.w2(32'h3bb80a1e),
	.w3(32'h3c1ea676),
	.w4(32'h39bef20e),
	.w5(32'h3c868180),
	.w6(32'h3bd441b5),
	.w7(32'hbb96c0f5),
	.w8(32'h3c0e9673),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5183c),
	.w1(32'h3c4ae5c6),
	.w2(32'h3bd1637b),
	.w3(32'h3c92299d),
	.w4(32'h3bb30a6c),
	.w5(32'h3b12d4ec),
	.w6(32'h3c633af1),
	.w7(32'h3bffcd5e),
	.w8(32'h3c6d7dff),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9c010),
	.w1(32'h3c3786d2),
	.w2(32'h3a4f8cf7),
	.w3(32'h3b8df914),
	.w4(32'h3c9cbbb5),
	.w5(32'h3bd11bc8),
	.w6(32'h3baed8b8),
	.w7(32'h3c04a798),
	.w8(32'h3c1b0071),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd8420),
	.w1(32'h3a76066d),
	.w2(32'hb9b63086),
	.w3(32'hbc0b1763),
	.w4(32'hbc06a074),
	.w5(32'hbc326cf5),
	.w6(32'hbadd950a),
	.w7(32'hbc6c7c78),
	.w8(32'hbc95872a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a4701),
	.w1(32'h3be934ba),
	.w2(32'h3bf64348),
	.w3(32'hbbcc2ba9),
	.w4(32'h3b2a4721),
	.w5(32'h3be6ba95),
	.w6(32'hbc202532),
	.w7(32'h3b49eb8d),
	.w8(32'h3b4716b9),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f7a0),
	.w1(32'hbbb39271),
	.w2(32'hbc3bcd9d),
	.w3(32'hbb1dde35),
	.w4(32'hbc0f308b),
	.w5(32'hbc8ef44c),
	.w6(32'hbb513c2d),
	.w7(32'hbc15a36e),
	.w8(32'hbc6d4cd6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b3064),
	.w1(32'hbc2b836c),
	.w2(32'h3b8b0af6),
	.w3(32'hbb4c66b9),
	.w4(32'hbc2a0e22),
	.w5(32'h3b228677),
	.w6(32'hbba2961b),
	.w7(32'hbc3b1d00),
	.w8(32'h38485a14),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f40e0),
	.w1(32'h3b1491aa),
	.w2(32'h37e513a4),
	.w3(32'h3ba4af7e),
	.w4(32'h3baae050),
	.w5(32'h3bb6cf8e),
	.w6(32'hbaae6b11),
	.w7(32'h3b6deda5),
	.w8(32'h3b92b8ef),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093f88),
	.w1(32'hbb82f2d6),
	.w2(32'h3bac24f2),
	.w3(32'h3b023c86),
	.w4(32'hbbb5f1b1),
	.w5(32'h3bec8a31),
	.w6(32'h3b8415ed),
	.w7(32'hbc67cca2),
	.w8(32'hbc392809),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b8444),
	.w1(32'hba430c5c),
	.w2(32'h3b8cb021),
	.w3(32'hbb5144f3),
	.w4(32'hbb91b5b3),
	.w5(32'hbadea2ca),
	.w6(32'hbc521c92),
	.w7(32'hbb22f1f2),
	.w8(32'hba7e7f17),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf22186),
	.w1(32'hbb5b093e),
	.w2(32'h3b236c71),
	.w3(32'h3aaed229),
	.w4(32'hbbaa7a31),
	.w5(32'h3bcb1d4f),
	.w6(32'h3a7985a9),
	.w7(32'h3b3001e0),
	.w8(32'h3c307a80),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e598f),
	.w1(32'h3b552e93),
	.w2(32'h3b90bb22),
	.w3(32'h3b86cdec),
	.w4(32'h3b9a296a),
	.w5(32'h3c51c025),
	.w6(32'h3afb9c8a),
	.w7(32'h3beb828e),
	.w8(32'h3c2a4139),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a339c),
	.w1(32'hbbc75789),
	.w2(32'hbb7bdc5a),
	.w3(32'h3c411c13),
	.w4(32'h3afbc0a0),
	.w5(32'hb7fdd787),
	.w6(32'h3bb5dec7),
	.w7(32'h3b9b95e0),
	.w8(32'hbb8756fa),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c4f12),
	.w1(32'hbc0a0a27),
	.w2(32'hbbc7beb3),
	.w3(32'h3979b8f1),
	.w4(32'hbc19760b),
	.w5(32'hbc005825),
	.w6(32'h393131a2),
	.w7(32'hbba4c4d3),
	.w8(32'hbc22f5d5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d3550),
	.w1(32'h3c9882c2),
	.w2(32'h3c0a4876),
	.w3(32'hba11afd2),
	.w4(32'h3cd58f08),
	.w5(32'h3c963404),
	.w6(32'h3b763d18),
	.w7(32'h3cb09eb0),
	.w8(32'h3c5377fe),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ac123),
	.w1(32'h3b7dcb8e),
	.w2(32'h3b73ec46),
	.w3(32'hbafca4ef),
	.w4(32'h3a79bee8),
	.w5(32'h3c3ed3f9),
	.w6(32'hbaf25b2f),
	.w7(32'h3b9f5da7),
	.w8(32'h3bfb23c4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be8de5),
	.w1(32'h38100855),
	.w2(32'hb99e0b3f),
	.w3(32'h3b4e30a4),
	.w4(32'h3a932ad5),
	.w5(32'hbba3e27d),
	.w6(32'h3b7e050e),
	.w7(32'h3a524373),
	.w8(32'hbb8cbe34),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f8f12),
	.w1(32'hbc16cbb9),
	.w2(32'hbc0fc968),
	.w3(32'h3b0dd253),
	.w4(32'hbc22c60f),
	.w5(32'hbc374ed8),
	.w6(32'hbb8f1d07),
	.w7(32'hbb8d6f45),
	.w8(32'hbb39be50),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc386ae8),
	.w1(32'h396b6d85),
	.w2(32'h3a4d5302),
	.w3(32'hbc1b5e15),
	.w4(32'hbbca4e29),
	.w5(32'h3b2b6376),
	.w6(32'hbc356a19),
	.w7(32'h3b878c6c),
	.w8(32'h3ad8d2d9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2ab9d),
	.w1(32'hbb6f0df9),
	.w2(32'hbb69cef0),
	.w3(32'h3ad951e9),
	.w4(32'hbb12203f),
	.w5(32'h3a9bc1b0),
	.w6(32'hba485bd4),
	.w7(32'hbb39f14c),
	.w8(32'h3a9bab97),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926dc1),
	.w1(32'hbc670602),
	.w2(32'hbb8d77be),
	.w3(32'hb94f7558),
	.w4(32'hbb35b0cb),
	.w5(32'h3b22a2cd),
	.w6(32'hba3dac87),
	.w7(32'hbaab9bf0),
	.w8(32'h3c20696d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13cb05),
	.w1(32'h3bfe373d),
	.w2(32'h3addb48b),
	.w3(32'h3b3af83f),
	.w4(32'h3bdc9bd9),
	.w5(32'h3c2af851),
	.w6(32'h3b77138f),
	.w7(32'h3ade7ac4),
	.w8(32'h38150c6f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3a153),
	.w1(32'hb9ff8163),
	.w2(32'h3bd2e8fc),
	.w3(32'h3b77e531),
	.w4(32'h3bb673e2),
	.w5(32'h3c9aa2e4),
	.w6(32'hbb193457),
	.w7(32'h3b04a024),
	.w8(32'h3c715137),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c30b7),
	.w1(32'h3c32c55d),
	.w2(32'h3c25abd1),
	.w3(32'h3c320467),
	.w4(32'h3c9a55a4),
	.w5(32'h3c9a1d59),
	.w6(32'h3c08a07d),
	.w7(32'h3c7b45d0),
	.w8(32'h3c7e40f1),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd11d23),
	.w1(32'hbbe10653),
	.w2(32'h3a958b81),
	.w3(32'h3c5dd1fc),
	.w4(32'hba6d6a33),
	.w5(32'h3c2fa777),
	.w6(32'h3c51c18b),
	.w7(32'h3bcc19cd),
	.w8(32'h3b421642),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c7701),
	.w1(32'h3c129dcc),
	.w2(32'hbac81c0b),
	.w3(32'h3c1a01ea),
	.w4(32'h3bef3e7d),
	.w5(32'hbc022c12),
	.w6(32'h3bbe3952),
	.w7(32'h3a5967da),
	.w8(32'hbc3eb04a),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0355a1),
	.w1(32'h3c85d0d0),
	.w2(32'h3c3585bd),
	.w3(32'hbc10b750),
	.w4(32'h3b52204e),
	.w5(32'hbbcb1fc0),
	.w6(32'hbbbe98d9),
	.w7(32'hbb1a5ffe),
	.w8(32'hbbc5a4a3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule