module layer_10_featuremap_8(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa06d8),
	.w1(32'h3b5c9dc9),
	.w2(32'h3b2ce810),
	.w3(32'h3b2fceaa),
	.w4(32'h3b4eb6a7),
	.w5(32'h3834314e),
	.w6(32'hbb724183),
	.w7(32'hba201699),
	.w8(32'h3ba23357),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebf8ab),
	.w1(32'h3bcec5d2),
	.w2(32'h3c276961),
	.w3(32'hbc22c902),
	.w4(32'hba2bb869),
	.w5(32'hbb364cf7),
	.w6(32'h3b3b571d),
	.w7(32'hbb4b6fed),
	.w8(32'hbbcd608a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a7006),
	.w1(32'h3adae164),
	.w2(32'h3a98d803),
	.w3(32'hbbaf3c2c),
	.w4(32'hbbc8bd68),
	.w5(32'hb89c1072),
	.w6(32'hbc34f51d),
	.w7(32'hbb705b22),
	.w8(32'h39321faf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef4200),
	.w1(32'hbbb0a8f6),
	.w2(32'h3bad224e),
	.w3(32'hbbdc97c2),
	.w4(32'hbc064554),
	.w5(32'hbb187383),
	.w6(32'hbbf0a9cd),
	.w7(32'hbba0d7bb),
	.w8(32'hbbcbe974),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09c6f1),
	.w1(32'hbb5b84a3),
	.w2(32'h391d8b39),
	.w3(32'hbc0442de),
	.w4(32'hbb796592),
	.w5(32'h3b811bff),
	.w6(32'hbbb7469d),
	.w7(32'hbb0ddf20),
	.w8(32'h3b12a56a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46a493),
	.w1(32'h3b6a52da),
	.w2(32'h3b7a81ed),
	.w3(32'h3bb9a5de),
	.w4(32'h3c04c86b),
	.w5(32'h3c13ea82),
	.w6(32'h3b7d6951),
	.w7(32'h3bb116c3),
	.w8(32'h3b9dc1ce),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c261d37),
	.w1(32'h3bcdb4f4),
	.w2(32'hbbb67f12),
	.w3(32'h3b982315),
	.w4(32'h3c558e7e),
	.w5(32'h3b0c209b),
	.w6(32'h3b95135b),
	.w7(32'h3c4257a5),
	.w8(32'h382c1e42),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb76dc),
	.w1(32'h3d46c48e),
	.w2(32'h3bc3c7b9),
	.w3(32'h3c79f624),
	.w4(32'h3cb04a25),
	.w5(32'hbaf05f4b),
	.w6(32'h3bd63455),
	.w7(32'h3c3c46e2),
	.w8(32'hba9a8653),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb755e08),
	.w1(32'hbb13bfdb),
	.w2(32'h39f32151),
	.w3(32'hbbb6e49f),
	.w4(32'hbb8978c1),
	.w5(32'hba9d9b15),
	.w6(32'h3b990c81),
	.w7(32'h3831200e),
	.w8(32'hba76f920),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0308a4),
	.w1(32'hba2553b3),
	.w2(32'hbc721859),
	.w3(32'hbc02a627),
	.w4(32'hbb4d3788),
	.w5(32'hbca2ec61),
	.w6(32'hba7bf9ba),
	.w7(32'h3b683967),
	.w8(32'hbc81aa4a),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62304b),
	.w1(32'hbc1461d0),
	.w2(32'h38f19794),
	.w3(32'hbcce5689),
	.w4(32'hbc96c2b8),
	.w5(32'h3acf7cbb),
	.w6(32'hbcb4e0a3),
	.w7(32'hbc913945),
	.w8(32'hbb4613de),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb39771),
	.w1(32'h3bb175f5),
	.w2(32'hbb0f5556),
	.w3(32'hbbbc2d41),
	.w4(32'h3a0f45e6),
	.w5(32'h3c96d068),
	.w6(32'hba45cb19),
	.w7(32'h3bb9a15b),
	.w8(32'h3c9ff427),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62798b),
	.w1(32'h3bffcfb5),
	.w2(32'hbb97f1ec),
	.w3(32'h3cc243c2),
	.w4(32'h3cbefc84),
	.w5(32'h3a9f24db),
	.w6(32'h3cad32a3),
	.w7(32'h3cc4c694),
	.w8(32'hbba98820),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c26c),
	.w1(32'h3c4e29ce),
	.w2(32'h3ba0ff2a),
	.w3(32'h3baa39fa),
	.w4(32'h3bfef6df),
	.w5(32'h3ba35630),
	.w6(32'hba816f32),
	.w7(32'h3bc556f8),
	.w8(32'hbbbd151e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0afa70),
	.w1(32'hbada5e14),
	.w2(32'h3bb391fd),
	.w3(32'hbb83ce5e),
	.w4(32'hbb0bca3b),
	.w5(32'h3a6237ba),
	.w6(32'hbb6b7ac8),
	.w7(32'hbb07ddc9),
	.w8(32'hbabcd2b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa6126),
	.w1(32'h3c477a6e),
	.w2(32'hbc217f6f),
	.w3(32'h3b6ee306),
	.w4(32'h3c6c550f),
	.w5(32'hbcd38c0d),
	.w6(32'hbb5d70b3),
	.w7(32'h3c0afdcf),
	.w8(32'hbcdcaba4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab3ec0),
	.w1(32'hbc786610),
	.w2(32'h3aee4c62),
	.w3(32'hbd187536),
	.w4(32'hbced1942),
	.w5(32'h3b0ab1a1),
	.w6(32'hbd1122d5),
	.w7(32'hbce23cdb),
	.w8(32'hbaa94c45),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8b12),
	.w1(32'hbb0bf95e),
	.w2(32'hbc39daeb),
	.w3(32'h3ab5ec34),
	.w4(32'h3c42eba5),
	.w5(32'hbc41e14c),
	.w6(32'h3bcc9f39),
	.w7(32'h3c5a2b20),
	.w8(32'hbc08a6d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade7f24),
	.w1(32'h3a999b6a),
	.w2(32'hbc097d0c),
	.w3(32'h3ad21eee),
	.w4(32'h3bad9f26),
	.w5(32'hbc1d57bc),
	.w6(32'h3ba620bc),
	.w7(32'h3c1a5a59),
	.w8(32'hbbdc8c86),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f4e5),
	.w1(32'hbb9b89c4),
	.w2(32'hba2474ef),
	.w3(32'hbb6bc378),
	.w4(32'hbc1f52c0),
	.w5(32'hbb27658f),
	.w6(32'hbb9f9c85),
	.w7(32'hbb487b85),
	.w8(32'hbb10cae8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774fa4),
	.w1(32'hbb24e325),
	.w2(32'h3b92e3fd),
	.w3(32'hbb6809d8),
	.w4(32'h3ac76093),
	.w5(32'h3b193ccb),
	.w6(32'hba977017),
	.w7(32'h3ac551d3),
	.w8(32'hba08f007),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07779e),
	.w1(32'h39c7ae09),
	.w2(32'hba0fe636),
	.w3(32'hb967380f),
	.w4(32'h3b160e55),
	.w5(32'h38c09d18),
	.w6(32'h3b15065f),
	.w7(32'h39bd786a),
	.w8(32'h39059a64),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68bf00),
	.w1(32'h3b8c9e61),
	.w2(32'hbbe54c03),
	.w3(32'hbc7d009c),
	.w4(32'h3be1217b),
	.w5(32'hba61f90d),
	.w6(32'hbbbdb559),
	.w7(32'h3c47d915),
	.w8(32'hbae67402),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2fea),
	.w1(32'hb9c58003),
	.w2(32'h3aa2add7),
	.w3(32'h3b7fadff),
	.w4(32'h3b4b7870),
	.w5(32'hbb5a6cd4),
	.w6(32'h3b9b51f4),
	.w7(32'h3babdc34),
	.w8(32'h3bc0929d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ec93a),
	.w1(32'hbb7d7017),
	.w2(32'h3bf71de2),
	.w3(32'hbc4aa399),
	.w4(32'hb95713a8),
	.w5(32'h3b6cd158),
	.w6(32'hbbf033ab),
	.w7(32'hbb36873d),
	.w8(32'h3a3840ef),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ea299),
	.w1(32'hbbab2342),
	.w2(32'hbb154abe),
	.w3(32'hbbeff3a2),
	.w4(32'hbbef5296),
	.w5(32'hbb617af9),
	.w6(32'h39c62772),
	.w7(32'hbb230481),
	.w8(32'hbb920f78),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5dd82e),
	.w1(32'hbadc3f29),
	.w2(32'h3a2f811c),
	.w3(32'hbb95b71e),
	.w4(32'h38447036),
	.w5(32'h3ab2b9d9),
	.w6(32'hbb7cdf63),
	.w7(32'hbacb3adf),
	.w8(32'h3a1a3cd7),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37ffe2),
	.w1(32'hbbacb618),
	.w2(32'hbb8a99d5),
	.w3(32'h3b40cd79),
	.w4(32'h3be107d7),
	.w5(32'h3c4afd98),
	.w6(32'h3c2165ad),
	.w7(32'h3bc87526),
	.w8(32'hbab3a910),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a519dbb),
	.w1(32'h3aa7fed6),
	.w2(32'h3c12fda0),
	.w3(32'h3be6ebf1),
	.w4(32'h3c014147),
	.w5(32'hbc9697b6),
	.w6(32'h3b76fa93),
	.w7(32'h3ba6707e),
	.w8(32'hbca269c4),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca68bd),
	.w1(32'h3cbb4454),
	.w2(32'hbbd60042),
	.w3(32'hbcf2ccdc),
	.w4(32'h3c0817d8),
	.w5(32'hbbd7fb79),
	.w6(32'hbcaba49c),
	.w7(32'hbc55e38b),
	.w8(32'hbc08b5a5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315039),
	.w1(32'hb933adb5),
	.w2(32'hbb92d5d2),
	.w3(32'h3b1a1358),
	.w4(32'h3b9f7396),
	.w5(32'hbc794f09),
	.w6(32'h39bb3707),
	.w7(32'h3b4376bb),
	.w8(32'hbbf68aa6),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f9bc),
	.w1(32'hb9445c9b),
	.w2(32'h3932ea65),
	.w3(32'hbcb80fe6),
	.w4(32'hbbc7337f),
	.w5(32'hbcaf033a),
	.w6(32'hbc09ac09),
	.w7(32'h3b08dc0b),
	.w8(32'hbc9c22dd),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c150795),
	.w1(32'h3c4d4aac),
	.w2(32'hbbd26c74),
	.w3(32'hbccd7d91),
	.w4(32'h3afc7417),
	.w5(32'hbba7b989),
	.w6(32'hbc900573),
	.w7(32'hbc02f48d),
	.w8(32'hbb259deb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba832cc9),
	.w1(32'h3b940c1d),
	.w2(32'h3b8c2723),
	.w3(32'hba974b3b),
	.w4(32'h3b6a467a),
	.w5(32'hbac94dc1),
	.w6(32'hbb5b7ecd),
	.w7(32'hba04eb81),
	.w8(32'hbbf06d18),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf07bae),
	.w1(32'hbbef3580),
	.w2(32'hbb6ba776),
	.w3(32'hbbbfbfd5),
	.w4(32'h3a2180be),
	.w5(32'hbabdca9b),
	.w6(32'h3ae8e601),
	.w7(32'h3c12fe6f),
	.w8(32'h3ab10be9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8288fe),
	.w1(32'hb9cba8da),
	.w2(32'h3cd44191),
	.w3(32'hbba82f43),
	.w4(32'h3a9edf95),
	.w5(32'h3c8609d2),
	.w6(32'hbb80ec3c),
	.w7(32'h3a8b95fe),
	.w8(32'h3c6f2190),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb918ee1),
	.w1(32'h3d603efe),
	.w2(32'h3cd1a655),
	.w3(32'hbca81842),
	.w4(32'h3bd89f90),
	.w5(32'h3d42f285),
	.w6(32'hbc92ab3e),
	.w7(32'h3c232800),
	.w8(32'h3d4343b7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb487bd),
	.w1(32'hbb423b9f),
	.w2(32'hbb6f3a71),
	.w3(32'hbc304980),
	.w4(32'h3b9d8834),
	.w5(32'hbc5fa369),
	.w6(32'hbbbdb2fb),
	.w7(32'h3b64ff9a),
	.w8(32'hbb10ceb8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c64f4),
	.w1(32'hbbb94c0b),
	.w2(32'hbc5b84c3),
	.w3(32'hb9fae64e),
	.w4(32'hbae54040),
	.w5(32'hbbbb0f73),
	.w6(32'h3c9a1c9b),
	.w7(32'h3b4387c6),
	.w8(32'hbc004ab6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5f54),
	.w1(32'h3bdd35a1),
	.w2(32'h3b6da559),
	.w3(32'h3aba84d3),
	.w4(32'h3aa5b26e),
	.w5(32'hba8faa68),
	.w6(32'hbbdbbb0c),
	.w7(32'hbbc83f05),
	.w8(32'hba2105bc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2aef3),
	.w1(32'hbaedd211),
	.w2(32'hbbc8a8b0),
	.w3(32'hbb850ae0),
	.w4(32'hbc0ac783),
	.w5(32'hbc1320f1),
	.w6(32'hbc2f07e4),
	.w7(32'hbc2b482c),
	.w8(32'hbbdab289),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d093a),
	.w1(32'hbac02893),
	.w2(32'hbc12aca7),
	.w3(32'hbb9aa4eb),
	.w4(32'h3a8e6cfb),
	.w5(32'hbbe74079),
	.w6(32'hbab8ef1b),
	.w7(32'h3ba3e9ed),
	.w8(32'h3bab299d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a149636),
	.w1(32'h3b66e614),
	.w2(32'hb9eccabb),
	.w3(32'hbc06bca6),
	.w4(32'h3ad912df),
	.w5(32'h3baa4f27),
	.w6(32'hbb01a06a),
	.w7(32'hbb581555),
	.w8(32'h3b7ccf31),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd22303),
	.w1(32'hbc5203ca),
	.w2(32'hbcb3ea59),
	.w3(32'hba3cf88d),
	.w4(32'h3c1025b5),
	.w5(32'hbc994520),
	.w6(32'h3896c019),
	.w7(32'h3c4974c1),
	.w8(32'hbcb894a0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13db1a),
	.w1(32'hbb338631),
	.w2(32'h3c39c498),
	.w3(32'hbc107b59),
	.w4(32'hbba0f075),
	.w5(32'hba9a28e6),
	.w6(32'h3b89ae1d),
	.w7(32'hbb4810c9),
	.w8(32'hbb9b4321),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64ee10),
	.w1(32'h3c2475cd),
	.w2(32'h3b1ab32c),
	.w3(32'hbbf373ab),
	.w4(32'hbb5bb060),
	.w5(32'hbc2429ec),
	.w6(32'hbc97e383),
	.w7(32'hbb94b25d),
	.w8(32'hbc855bdf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3622c),
	.w1(32'hbb926744),
	.w2(32'hbc42994f),
	.w3(32'hbcc916b3),
	.w4(32'hbbc96410),
	.w5(32'hbc6a2627),
	.w6(32'hbc26ca3b),
	.w7(32'h3c086e8f),
	.w8(32'hbc12a1c7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13688f),
	.w1(32'h39a0c04a),
	.w2(32'hbc8160a4),
	.w3(32'hbc8507bb),
	.w4(32'h3bab3f68),
	.w5(32'hbbc36cad),
	.w6(32'hbb87752d),
	.w7(32'h3ca00223),
	.w8(32'hbb23479a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a2c5),
	.w1(32'h36e12bc7),
	.w2(32'hbb99cc03),
	.w3(32'hbaca39a9),
	.w4(32'h3a6027cd),
	.w5(32'hbc5ee8ee),
	.w6(32'h3a354462),
	.w7(32'h3b0bc10f),
	.w8(32'hbb966ea7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1dbc9),
	.w1(32'h3bbdd315),
	.w2(32'hbbfb4da6),
	.w3(32'hbbc83aef),
	.w4(32'hbb95ccc7),
	.w5(32'hbb61a0e7),
	.w6(32'h386f9e22),
	.w7(32'hbaa4233f),
	.w8(32'h3b150cf4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ee71b),
	.w1(32'h3b8abb0e),
	.w2(32'hbbd71e64),
	.w3(32'h38b1c1ef),
	.w4(32'h3c3300a6),
	.w5(32'hbbc394ad),
	.w6(32'h3c38435e),
	.w7(32'h3bef8c35),
	.w8(32'h3a3cb62e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48cda3),
	.w1(32'hbbdb6376),
	.w2(32'hbb558863),
	.w3(32'h3b4234b0),
	.w4(32'h3c28b64d),
	.w5(32'hbb23e8f4),
	.w6(32'h3c85f0e2),
	.w7(32'h3b68b6c1),
	.w8(32'hbbb192c8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b918e9b),
	.w1(32'h3ae4bd10),
	.w2(32'h3a6a6a81),
	.w3(32'h3bead6d4),
	.w4(32'h3b7ed6ef),
	.w5(32'hbc397c74),
	.w6(32'h3babcd77),
	.w7(32'hbb878a7b),
	.w8(32'hbb5a767f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb825),
	.w1(32'h3c216319),
	.w2(32'hbc5e2952),
	.w3(32'hbbd4b4b4),
	.w4(32'h3bce5edb),
	.w5(32'hbcaf484b),
	.w6(32'h3c2a45ad),
	.w7(32'h3c7650a5),
	.w8(32'hbbe36d3f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0de3b9),
	.w1(32'h3c2ecc04),
	.w2(32'h3b64ff6f),
	.w3(32'hbbb7326d),
	.w4(32'h3c432241),
	.w5(32'hbcb03e42),
	.w6(32'h3a6db3f9),
	.w7(32'hba149735),
	.w8(32'hbcae597c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9551d8),
	.w1(32'h3b94d91b),
	.w2(32'hbc1b5933),
	.w3(32'hbccc42eb),
	.w4(32'hbc355324),
	.w5(32'hbcd55ee8),
	.w6(32'hbc9f1bcf),
	.w7(32'hbc544425),
	.w8(32'hbc1b4e6c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe38ac7),
	.w1(32'h3c43abdd),
	.w2(32'hbb6c4703),
	.w3(32'hbcc5a054),
	.w4(32'hba87727c),
	.w5(32'h3b0c1563),
	.w6(32'hbc993587),
	.w7(32'h3a88f62d),
	.w8(32'hbabac2ce),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39c950),
	.w1(32'hbbc51116),
	.w2(32'h3a9abd76),
	.w3(32'hbbadd90f),
	.w4(32'hbb3b05eb),
	.w5(32'h3b2d861c),
	.w6(32'hbbc6634c),
	.w7(32'hbbb38698),
	.w8(32'hbae6de07),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85006e),
	.w1(32'hb9f5ddac),
	.w2(32'h3ab9220a),
	.w3(32'h3ac85286),
	.w4(32'h3b124458),
	.w5(32'hb8bc8bbc),
	.w6(32'hbbc5bbc9),
	.w7(32'hbbf36013),
	.w8(32'h3b90fcc2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba852a7e),
	.w1(32'h39b474b5),
	.w2(32'hbbdc3821),
	.w3(32'h3b1c4351),
	.w4(32'h3af7efb4),
	.w5(32'h3c1637e3),
	.w6(32'hb8af1cbe),
	.w7(32'h3a993ffb),
	.w8(32'h3bddda50),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a994969),
	.w1(32'hbc1f99a0),
	.w2(32'hbbf94236),
	.w3(32'h3c94f455),
	.w4(32'h3c866454),
	.w5(32'hbc438f64),
	.w6(32'h3c8f09c7),
	.w7(32'h3ca645ea),
	.w8(32'hbbda818b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac77a8a),
	.w1(32'hbb8cbb05),
	.w2(32'h3a84c023),
	.w3(32'hbc891064),
	.w4(32'hbaa8cbb5),
	.w5(32'hbaa07f17),
	.w6(32'hbb5b4081),
	.w7(32'h3c4d74c7),
	.w8(32'hbc1e1d99),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891259c),
	.w1(32'h3b7bec3d),
	.w2(32'h3c145e20),
	.w3(32'h39d454aa),
	.w4(32'h3c03fedd),
	.w5(32'h3cb63026),
	.w6(32'hbbb42521),
	.w7(32'h3b0f9995),
	.w8(32'h3c70c4fa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5d2f2e),
	.w1(32'h3bbfda5b),
	.w2(32'h3b86791c),
	.w3(32'h3ce0ab6c),
	.w4(32'h3cb08606),
	.w5(32'h3c5d7b87),
	.w6(32'h3c9c8339),
	.w7(32'h3c08e980),
	.w8(32'h3bb5b253),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9c710),
	.w1(32'hbae3dfa8),
	.w2(32'h3b8f823e),
	.w3(32'h3c143336),
	.w4(32'h3a48fcfc),
	.w5(32'hb8f65b80),
	.w6(32'h3bd2a040),
	.w7(32'h3b147507),
	.w8(32'hbb43ef31),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8dacf),
	.w1(32'h3b6ab0c6),
	.w2(32'hbab7ae22),
	.w3(32'h3a97accc),
	.w4(32'h3b0c89e4),
	.w5(32'h3b78ab48),
	.w6(32'hbb8e520f),
	.w7(32'hbb4955b0),
	.w8(32'h3afcb95f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7e03),
	.w1(32'hbbc028a2),
	.w2(32'hbc514089),
	.w3(32'hbb9f4f8a),
	.w4(32'hbb47036a),
	.w5(32'hbc119c7b),
	.w6(32'h3c29007b),
	.w7(32'h3c78deee),
	.w8(32'hbbf89d26),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bd832),
	.w1(32'h3c871752),
	.w2(32'h3c022089),
	.w3(32'h3c53515f),
	.w4(32'h3c078196),
	.w5(32'hbbec39d8),
	.w6(32'h3bf9e648),
	.w7(32'hbbb6ebaf),
	.w8(32'hbc9f2409),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11b5ac),
	.w1(32'hbc0eea45),
	.w2(32'h3a93db92),
	.w3(32'hbc39d25d),
	.w4(32'hbb4035a4),
	.w5(32'h3827b97e),
	.w6(32'hbbd766f7),
	.w7(32'hbc396a44),
	.w8(32'hbc0a259b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe05d69),
	.w1(32'hb9545d50),
	.w2(32'h3ba79bb9),
	.w3(32'hbc4c146b),
	.w4(32'hbb5179b7),
	.w5(32'h3b99d1da),
	.w6(32'hbbebfdf9),
	.w7(32'hbba42918),
	.w8(32'h3c1b1f56),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908574),
	.w1(32'hbb9114b7),
	.w2(32'h3b131387),
	.w3(32'h3bf1f1f8),
	.w4(32'hb9ed1627),
	.w5(32'hba8a23bd),
	.w6(32'h3c1a9cef),
	.w7(32'hba8ea945),
	.w8(32'hba8da36b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97d312),
	.w1(32'h3b34db38),
	.w2(32'hbbe7c3a7),
	.w3(32'hba095f5d),
	.w4(32'hbb96a36d),
	.w5(32'hbc2e227f),
	.w6(32'hbae87eee),
	.w7(32'hbc1b0e9b),
	.w8(32'h36c20eea),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc349e15),
	.w1(32'hbbe4158f),
	.w2(32'hbb42d94b),
	.w3(32'hbc51b32e),
	.w4(32'hbbd0587f),
	.w5(32'h3c5b44f7),
	.w6(32'h3af13660),
	.w7(32'h3c82daea),
	.w8(32'h3b24ccc4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf39c87),
	.w1(32'h3b9a458f),
	.w2(32'hbb2842af),
	.w3(32'h3c5c5592),
	.w4(32'h3c64f2c3),
	.w5(32'h3af49f58),
	.w6(32'h3c1e7e68),
	.w7(32'h3c5ec0a9),
	.w8(32'hbb3e65fc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ccdc83),
	.w1(32'h3b74d559),
	.w2(32'hbbffd10d),
	.w3(32'h3b7ac864),
	.w4(32'h3ba8ec65),
	.w5(32'hbb330d0a),
	.w6(32'h3b459da0),
	.w7(32'h3bda12ea),
	.w8(32'h3c15aeff),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a840),
	.w1(32'hbb852971),
	.w2(32'hbc07d837),
	.w3(32'hbb5567a2),
	.w4(32'hbbe13749),
	.w5(32'hbc08790b),
	.w6(32'h3be0e8ce),
	.w7(32'h3c353e18),
	.w8(32'hbbccbdce),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79f063),
	.w1(32'h3a3ec603),
	.w2(32'hbbda95c1),
	.w3(32'hbbd248df),
	.w4(32'h3b41a576),
	.w5(32'hbc4207a3),
	.w6(32'hbc9c8a58),
	.w7(32'h3c0db3fc),
	.w8(32'hbb2b0f91),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2ba1bd),
	.w1(32'hbcde8ad8),
	.w2(32'hbb1416c5),
	.w3(32'hbce000ef),
	.w4(32'hbc7028d7),
	.w5(32'hbc1c32aa),
	.w6(32'hbbcade37),
	.w7(32'h3bc7e575),
	.w8(32'hbc3680ca),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafcf5d),
	.w1(32'h3ba6cb81),
	.w2(32'hba449225),
	.w3(32'hbbf25cdd),
	.w4(32'hba475db2),
	.w5(32'h3ad0a5e7),
	.w6(32'hb8617e6c),
	.w7(32'h3bdd5426),
	.w8(32'hbabb0cca),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc97f8),
	.w1(32'h3be8932b),
	.w2(32'hbae26d7b),
	.w3(32'hbc2a8106),
	.w4(32'hbb313b16),
	.w5(32'hbbbbe661),
	.w6(32'hbbacc321),
	.w7(32'h3b842ab2),
	.w8(32'hbb38e15d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b772c00),
	.w1(32'hbb260152),
	.w2(32'hbb402e8b),
	.w3(32'hb93353f7),
	.w4(32'h39ff513a),
	.w5(32'hbb358509),
	.w6(32'h3afe780a),
	.w7(32'h3a27b0ef),
	.w8(32'hbbcee855),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2e08d),
	.w1(32'h3999f1fb),
	.w2(32'hb8c79a96),
	.w3(32'h3b36826a),
	.w4(32'h3bbd3030),
	.w5(32'h3c328c7f),
	.w6(32'hba9ccec5),
	.w7(32'h3b23ae76),
	.w8(32'h3c13b911),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17485d),
	.w1(32'hbc0be84d),
	.w2(32'h3abba006),
	.w3(32'h3ac50b7a),
	.w4(32'hbad8ca59),
	.w5(32'hbb80de9a),
	.w6(32'h3b74bbab),
	.w7(32'h3ba7b309),
	.w8(32'hbbba80e1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbda577),
	.w1(32'hbbb8012c),
	.w2(32'hbb9bfbd7),
	.w3(32'hbca26d18),
	.w4(32'hbc80da7e),
	.w5(32'hbaaeaaed),
	.w6(32'hbc5716c9),
	.w7(32'hbc6a3c64),
	.w8(32'hbb10df89),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc331166),
	.w1(32'h3ae86494),
	.w2(32'h3bcb5227),
	.w3(32'hbc4f88b7),
	.w4(32'h3b8d103c),
	.w5(32'h3c03a0a9),
	.w6(32'h3a857267),
	.w7(32'h3c1d4807),
	.w8(32'h3bd3c071),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e0b99),
	.w1(32'hbbd58a9e),
	.w2(32'hbb2c6bd3),
	.w3(32'h3aee4dec),
	.w4(32'hbbb9ea76),
	.w5(32'hb988f6d4),
	.w6(32'h3ba26813),
	.w7(32'hbb51d3e6),
	.w8(32'hb9eb884b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c9bb),
	.w1(32'h39982f99),
	.w2(32'h3c5f6196),
	.w3(32'hbb05adbd),
	.w4(32'hbb46fe01),
	.w5(32'h3c3f366c),
	.w6(32'hbb619e05),
	.w7(32'hbb8e5520),
	.w8(32'h3bf1a9a6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c2fe1),
	.w1(32'h3aaeba5c),
	.w2(32'hbc2eccce),
	.w3(32'h3b7b7bcb),
	.w4(32'h3b0a18c9),
	.w5(32'hbb2dd8b1),
	.w6(32'h3b4e1aa9),
	.w7(32'h3aa25a90),
	.w8(32'h3b3911a5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc289),
	.w1(32'h3b6b471e),
	.w2(32'h3c5282a7),
	.w3(32'h3a211548),
	.w4(32'h3b4ac654),
	.w5(32'hbbb6b904),
	.w6(32'h3be5b127),
	.w7(32'hbc3a2465),
	.w8(32'hbc401eac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb74e18),
	.w1(32'h3c0a133d),
	.w2(32'h3b6d669f),
	.w3(32'hbc7a689a),
	.w4(32'hbb9d18be),
	.w5(32'h3bada7e5),
	.w6(32'hbc2de8c1),
	.w7(32'hbb1238f0),
	.w8(32'h3be2408d),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf6182),
	.w1(32'h3b049cc1),
	.w2(32'hb9899eb0),
	.w3(32'hbba5ac53),
	.w4(32'h3b6e1b08),
	.w5(32'h3c8ccdb9),
	.w6(32'h3b90deb7),
	.w7(32'h3bfd4183),
	.w8(32'h3b7ef119),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e1860),
	.w1(32'h3c372111),
	.w2(32'hbc2bca2b),
	.w3(32'h3b81d128),
	.w4(32'h3c823812),
	.w5(32'hbb8ea551),
	.w6(32'hb9114740),
	.w7(32'h3bd7d004),
	.w8(32'h3b6ed58d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc75773),
	.w1(32'h39c49d23),
	.w2(32'hbb76220e),
	.w3(32'hbbbd0cc8),
	.w4(32'hbb907fb9),
	.w5(32'h39d8cc0a),
	.w6(32'h3b579018),
	.w7(32'h3adb0e23),
	.w8(32'h3b15d691),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92e9f9),
	.w1(32'hbb85e25e),
	.w2(32'hbb567b60),
	.w3(32'h3bed55c7),
	.w4(32'h3bcba15c),
	.w5(32'hbc008f42),
	.w6(32'h3b921687),
	.w7(32'h3be0a8a9),
	.w8(32'hbc9ff0eb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215518),
	.w1(32'hbc128537),
	.w2(32'hbc9ff23d),
	.w3(32'hbc94b3de),
	.w4(32'hbc14a223),
	.w5(32'hbca6d21a),
	.w6(32'hbc86fef7),
	.w7(32'hbc1b7884),
	.w8(32'hbc3666e6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a71e8),
	.w1(32'hbcb24211),
	.w2(32'h3988dc3c),
	.w3(32'hbd0acef9),
	.w4(32'hbd03ac1a),
	.w5(32'hbaa59ce5),
	.w6(32'hbccdf7cd),
	.w7(32'hbc8c7adb),
	.w8(32'h3b0b9d8d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13d144),
	.w1(32'h3a70884f),
	.w2(32'hbc40476b),
	.w3(32'hbb8e3bc0),
	.w4(32'hbbb3877c),
	.w5(32'hbbcae13a),
	.w6(32'h3b440b61),
	.w7(32'h3b6e9f46),
	.w8(32'hba2104bb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd094),
	.w1(32'h3c4048f1),
	.w2(32'hbcbfc990),
	.w3(32'hbbd72616),
	.w4(32'h3c0a6f85),
	.w5(32'hbd113733),
	.w6(32'hbb1aa398),
	.w7(32'h3ca06f7f),
	.w8(32'hbbcfe856),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf3766b),
	.w1(32'hbc7751ce),
	.w2(32'hbc8bf456),
	.w3(32'hbcb108f4),
	.w4(32'hbc1e047a),
	.w5(32'hbbc6f9a5),
	.w6(32'hbbe36655),
	.w7(32'h3c7e34b2),
	.w8(32'hbbbb2dff),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41221f),
	.w1(32'h3cd46305),
	.w2(32'h3d5135cf),
	.w3(32'h3ba18926),
	.w4(32'h3ca3f1ca),
	.w5(32'h3d5de888),
	.w6(32'hbb4ec6a7),
	.w7(32'h3c4fc802),
	.w8(32'h3d07ee7c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5c68),
	.w1(32'h3b8295f9),
	.w2(32'h3c28678b),
	.w3(32'h3bd5fc5d),
	.w4(32'h3b6cb042),
	.w5(32'h3c1d9d26),
	.w6(32'h3aeaf4df),
	.w7(32'h3b2dab8d),
	.w8(32'h3bc95b9d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2915f8),
	.w1(32'hbbc2241c),
	.w2(32'h3bdbeb48),
	.w3(32'hbc88d743),
	.w4(32'hba948ab2),
	.w5(32'hbb84022e),
	.w6(32'hbc02d3cd),
	.w7(32'hbb8270fd),
	.w8(32'hbb8d36d7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991324),
	.w1(32'h3c67c5dc),
	.w2(32'hbb0bd9de),
	.w3(32'hbc4db608),
	.w4(32'hba82dbb8),
	.w5(32'h3b80ec47),
	.w6(32'hbc2eb521),
	.w7(32'h3bc54837),
	.w8(32'h3c5ed2ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986e326),
	.w1(32'hbb4dac0a),
	.w2(32'hbb596294),
	.w3(32'hbaafe1b2),
	.w4(32'hbbaf473c),
	.w5(32'hbad54c13),
	.w6(32'h3b03fbb5),
	.w7(32'h39083aa3),
	.w8(32'h3bf93692),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66328c),
	.w1(32'h3d05c10d),
	.w2(32'h3cae2c07),
	.w3(32'h3c21cf0e),
	.w4(32'h3c068afe),
	.w5(32'h3d17c155),
	.w6(32'h3997741c),
	.w7(32'h3cd57b12),
	.w8(32'h3cf35224),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f5fc4),
	.w1(32'hb9c971d4),
	.w2(32'h3b2b8eb2),
	.w3(32'h3bb431a4),
	.w4(32'hbb6dd7c3),
	.w5(32'h3c1c0661),
	.w6(32'h3b7c6130),
	.w7(32'hbba63d78),
	.w8(32'h3c6d0b8f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac44880),
	.w1(32'h3bbe0281),
	.w2(32'h3b0428e2),
	.w3(32'h3bbfa607),
	.w4(32'h3baab885),
	.w5(32'hbc574a9e),
	.w6(32'h3bf740bc),
	.w7(32'h3ba02b29),
	.w8(32'hbb7a23b2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd20e09),
	.w1(32'h3c795037),
	.w2(32'hbbd6a24e),
	.w3(32'hbc3f2397),
	.w4(32'hbb8cf96e),
	.w5(32'hbc26d7d7),
	.w6(32'hbb8ac970),
	.w7(32'hb85c0b41),
	.w8(32'hbc1fd3c3),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba963c52),
	.w1(32'h3c1abcdd),
	.w2(32'hbc377482),
	.w3(32'hbb97d848),
	.w4(32'h3be7cfd7),
	.w5(32'hbc872c71),
	.w6(32'hbb08e8a2),
	.w7(32'h3bbd1f75),
	.w8(32'hbc42ed60),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d108a),
	.w1(32'hbbe94665),
	.w2(32'h3bd32dc4),
	.w3(32'hbcc1c525),
	.w4(32'hbc884d5c),
	.w5(32'h3c03be0f),
	.w6(32'hbbc8e5da),
	.w7(32'hbb893424),
	.w8(32'h3b0870c9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf759c8),
	.w1(32'h3c04ecbe),
	.w2(32'hbba2ddd8),
	.w3(32'h3c7a65fa),
	.w4(32'h3bd74cbd),
	.w5(32'hbaf590d8),
	.w6(32'h3c0726b9),
	.w7(32'h3bd7cefd),
	.w8(32'hbbc447ed),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17c2b9),
	.w1(32'hbb62f433),
	.w2(32'h3c823fac),
	.w3(32'h3baa6b07),
	.w4(32'hbb67bacb),
	.w5(32'h3be8ed2c),
	.w6(32'h3c0425a1),
	.w7(32'h3c40c1e0),
	.w8(32'h3b78955d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78b333),
	.w1(32'hbc6d009d),
	.w2(32'hbbad2cac),
	.w3(32'hbc5dac24),
	.w4(32'hba8b0cdd),
	.w5(32'hbc9b0655),
	.w6(32'hbc407d10),
	.w7(32'hbc058362),
	.w8(32'hbcadd0f0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01f4d9),
	.w1(32'h3c63522e),
	.w2(32'hbbfff55f),
	.w3(32'hbcb8ebf3),
	.w4(32'h3ba86934),
	.w5(32'hbbd7ded3),
	.w6(32'hbc4d38cd),
	.w7(32'hbb1fdefa),
	.w8(32'hbc19a880),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96861a),
	.w1(32'hba97bd03),
	.w2(32'h3b33f877),
	.w3(32'hbc85aafa),
	.w4(32'hbbc9223e),
	.w5(32'h39ac4129),
	.w6(32'hbbceeef3),
	.w7(32'h3b5a4c89),
	.w8(32'h3bdaa2e7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70c6d6),
	.w1(32'h3bcefee5),
	.w2(32'h3a8a705e),
	.w3(32'h3ba51a9d),
	.w4(32'h3bb8d7a6),
	.w5(32'hbb558546),
	.w6(32'h3c162ac0),
	.w7(32'h3bc09c80),
	.w8(32'hbbc34489),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f57bd),
	.w1(32'h3b299bd7),
	.w2(32'h3bbf8c37),
	.w3(32'hbbf8f9b0),
	.w4(32'hbb31b2d4),
	.w5(32'hbb250fe6),
	.w6(32'hbc141652),
	.w7(32'hbc182434),
	.w8(32'h3a008035),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b747770),
	.w1(32'h3b56f498),
	.w2(32'hbc043836),
	.w3(32'hb90818af),
	.w4(32'h3b9a3b52),
	.w5(32'hbc96f565),
	.w6(32'hb9b744b3),
	.w7(32'h3ae3410c),
	.w8(32'hbbcb2163),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc928dfb),
	.w1(32'hbc42f5d4),
	.w2(32'h3b8b2a22),
	.w3(32'hbc4f811b),
	.w4(32'hbb7868a8),
	.w5(32'h3c1cee81),
	.w6(32'hbb47df73),
	.w7(32'hbb7ef37f),
	.w8(32'h3ba870c4),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b492249),
	.w1(32'h3b134560),
	.w2(32'h3adebd98),
	.w3(32'h3bc8a16e),
	.w4(32'h3a89051f),
	.w5(32'h3b8dc76d),
	.w6(32'h3bb79037),
	.w7(32'h3bcd6248),
	.w8(32'hbb91a82c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b907f4f),
	.w1(32'h3c0a64e9),
	.w2(32'hbb4deee5),
	.w3(32'h3c180078),
	.w4(32'h3b8f93c3),
	.w5(32'hbb2e412f),
	.w6(32'h3a57f6f7),
	.w7(32'h3b1c6043),
	.w8(32'hbb4ddbe1),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ec03),
	.w1(32'h3b1554fa),
	.w2(32'hbbf36d6d),
	.w3(32'h3a119bc8),
	.w4(32'h3a4ba655),
	.w5(32'hbb97a87b),
	.w6(32'hb9a0dc16),
	.w7(32'h39cec2d6),
	.w8(32'hbb07f8b1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc819978),
	.w1(32'hbc459271),
	.w2(32'h3bd5f918),
	.w3(32'hbc41d6e9),
	.w4(32'hbc281ab3),
	.w5(32'h3c7bae3a),
	.w6(32'hbbcd8e6f),
	.w7(32'hbc0dd585),
	.w8(32'h3baa0ae0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52923b),
	.w1(32'h3b5623b5),
	.w2(32'h3b1b3212),
	.w3(32'h3ce319ae),
	.w4(32'h3bf7ba8b),
	.w5(32'h3b5ec3b3),
	.w6(32'h3c9f40a1),
	.w7(32'h3bbe23a9),
	.w8(32'h38ff5784),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2e85),
	.w1(32'h3ba0a215),
	.w2(32'h3b20129e),
	.w3(32'h3b1d3d55),
	.w4(32'h3b8b46cb),
	.w5(32'h3c1d3e7b),
	.w6(32'hbb391329),
	.w7(32'h39621b93),
	.w8(32'h3c7bdc77),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60b03),
	.w1(32'h398fd045),
	.w2(32'h3b8d6174),
	.w3(32'h3c475830),
	.w4(32'h3b8ed749),
	.w5(32'hbbc1e5cb),
	.w6(32'h3c979355),
	.w7(32'h3aeba57f),
	.w8(32'h3c0105af),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf36367),
	.w1(32'hbc0661f1),
	.w2(32'h3bee2aa9),
	.w3(32'h3bf74703),
	.w4(32'h3b4775b0),
	.w5(32'h3b1c6ce3),
	.w6(32'h3c35eed3),
	.w7(32'h3c1db160),
	.w8(32'h3b8ca76a),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c937a),
	.w1(32'h3c5e901f),
	.w2(32'hbc4c9e00),
	.w3(32'hbc2a85a8),
	.w4(32'h3c59a8e7),
	.w5(32'hbbe01aa7),
	.w6(32'hba23ef7f),
	.w7(32'hba48bdc7),
	.w8(32'hbcaa1dfd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfaffe4),
	.w1(32'h3bea480e),
	.w2(32'hbd2685a0),
	.w3(32'hbcd500e0),
	.w4(32'hbae46443),
	.w5(32'hbcecc75d),
	.w6(32'hbc5d49d3),
	.w7(32'hbb2e86fe),
	.w8(32'hbc884957),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf6541b),
	.w1(32'hbc262531),
	.w2(32'h394da9d1),
	.w3(32'hbcc2f260),
	.w4(32'hbcc13126),
	.w5(32'h3b0b4254),
	.w6(32'hbc98acea),
	.w7(32'hbc7183d4),
	.w8(32'hbb4b161c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba134b15),
	.w1(32'h3bbe3d12),
	.w2(32'h3c2acbfc),
	.w3(32'hbbb43699),
	.w4(32'h3b23757a),
	.w5(32'h3c847c2b),
	.w6(32'hbca9d71f),
	.w7(32'hbbb1303c),
	.w8(32'h3bea2b96),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd27b),
	.w1(32'h3c41f2fe),
	.w2(32'hbb1a2105),
	.w3(32'h3c7da143),
	.w4(32'h3bbb2510),
	.w5(32'hbc3c334b),
	.w6(32'h3c3361e4),
	.w7(32'h3b99212f),
	.w8(32'hbbf19cff),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4e73),
	.w1(32'hbc4cbf02),
	.w2(32'h3b7c0f9b),
	.w3(32'hbc32c377),
	.w4(32'hbc1ee726),
	.w5(32'hbbcc3293),
	.w6(32'hbbdfc91c),
	.w7(32'hbc23ca05),
	.w8(32'hbb568cbe),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39546511),
	.w1(32'hbb9f9833),
	.w2(32'hbac09e50),
	.w3(32'hbc0f76e9),
	.w4(32'h3a772641),
	.w5(32'h3b1d291c),
	.w6(32'hb9de19ad),
	.w7(32'hbbf01751),
	.w8(32'hbb717209),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb165e09),
	.w1(32'hba3350a8),
	.w2(32'hbc8edf2a),
	.w3(32'hbb4a696e),
	.w4(32'h3c08c341),
	.w5(32'hbc9a19a6),
	.w6(32'h3b94a420),
	.w7(32'h3c3e19be),
	.w8(32'hbbf09172),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4333),
	.w1(32'h3b8401d2),
	.w2(32'hba2cebd7),
	.w3(32'hbbf090e7),
	.w4(32'h39b1da1c),
	.w5(32'hbc189974),
	.w6(32'hbb69f9f2),
	.w7(32'h3b66d05d),
	.w8(32'h3b8e412e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9460be),
	.w1(32'h3c30950d),
	.w2(32'h3b8f0411),
	.w3(32'hbc6745a8),
	.w4(32'hbb00e969),
	.w5(32'h3c242d91),
	.w6(32'hbbb78104),
	.w7(32'h3aff88c9),
	.w8(32'h3a272bd3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7aab6),
	.w1(32'h3b2429da),
	.w2(32'hbc09ae61),
	.w3(32'h386e086f),
	.w4(32'hbaf4a543),
	.w5(32'h3b078157),
	.w6(32'hbb808fc1),
	.w7(32'hbbe32ea6),
	.w8(32'h3b30b022),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb66bf9),
	.w1(32'h39ebf452),
	.w2(32'h3c8ede50),
	.w3(32'hba862815),
	.w4(32'h3b67fb64),
	.w5(32'h3c28188f),
	.w6(32'hbaca8303),
	.w7(32'hb6bb3f26),
	.w8(32'h3bc39020),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58afea),
	.w1(32'h3cbf1d3d),
	.w2(32'hbbd407ae),
	.w3(32'h3bf9ebc3),
	.w4(32'h3ac3dc92),
	.w5(32'hbbf918bc),
	.w6(32'h3c7802d6),
	.w7(32'hba75736f),
	.w8(32'hbb138d76),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb602578),
	.w1(32'hbb7a34aa),
	.w2(32'h3ba8d932),
	.w3(32'hbae080e3),
	.w4(32'hbb527345),
	.w5(32'hbb3abe9b),
	.w6(32'hb9453d3f),
	.w7(32'hb8aafd96),
	.w8(32'hbbeec290),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932166),
	.w1(32'h3c396079),
	.w2(32'hbc51584d),
	.w3(32'h3c0a3a7c),
	.w4(32'h3bce7a07),
	.w5(32'hbc815ef0),
	.w6(32'h3a649b3f),
	.w7(32'h3906f272),
	.w8(32'h3a91ca1d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58927c),
	.w1(32'hbbf043bb),
	.w2(32'h3bfb113c),
	.w3(32'hbc771de6),
	.w4(32'hbb17c4b1),
	.w5(32'hbbcdffbf),
	.w6(32'h3a872781),
	.w7(32'h3bd174d6),
	.w8(32'hbac64d67),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a414a),
	.w1(32'h3c1deeb6),
	.w2(32'hbb32d141),
	.w3(32'h39e42cd0),
	.w4(32'h3bb2c2ba),
	.w5(32'h39cbb39f),
	.w6(32'hbb3daa6e),
	.w7(32'hbad342b9),
	.w8(32'hb73d0b99),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66ec10),
	.w1(32'hbb1a0c06),
	.w2(32'h3ba44271),
	.w3(32'h3b029733),
	.w4(32'h3aefb247),
	.w5(32'h3b63384c),
	.w6(32'h3b03a002),
	.w7(32'h3a84622d),
	.w8(32'h3a6e2597),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baefcae),
	.w1(32'h3c0d92e2),
	.w2(32'h3a865e9b),
	.w3(32'h3ac9b870),
	.w4(32'h3c1e35bf),
	.w5(32'h3b4f8220),
	.w6(32'h3adad6e2),
	.w7(32'h3c2829cb),
	.w8(32'h3b4569f1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f159b),
	.w1(32'h3b82d270),
	.w2(32'hbbc71ff0),
	.w3(32'hbc01c03d),
	.w4(32'h3b5d54b9),
	.w5(32'hbc41fef0),
	.w6(32'hbbbf8141),
	.w7(32'hb9eadc55),
	.w8(32'hbb171991),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64bdb8),
	.w1(32'hbb57bc8d),
	.w2(32'hb9346309),
	.w3(32'hbc9c3285),
	.w4(32'hbbf4330c),
	.w5(32'hba3b2e6e),
	.w6(32'hbc3347cf),
	.w7(32'h3bd5fc6f),
	.w8(32'h3a8329ce),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d2f08),
	.w1(32'hbaa40e9e),
	.w2(32'hba8169d6),
	.w3(32'hba193b73),
	.w4(32'hba48ccfd),
	.w5(32'h3b5c99ae),
	.w6(32'h3a6fd79c),
	.w7(32'hb88a9a1f),
	.w8(32'h3ae4093d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ae6f6),
	.w1(32'h3c930a80),
	.w2(32'hbc6692c9),
	.w3(32'h3ba5208d),
	.w4(32'h3c8fd227),
	.w5(32'hbc5294ad),
	.w6(32'h3c03c56e),
	.w7(32'h3ca379c7),
	.w8(32'hbc09f766),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22b763),
	.w1(32'hbbdcf497),
	.w2(32'hbb98b28f),
	.w3(32'hbc1f44d5),
	.w4(32'hbbb8a2ee),
	.w5(32'hbb43bc5e),
	.w6(32'hbbe25c3a),
	.w7(32'hbbdc2667),
	.w8(32'hbbaddd51),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0342aa),
	.w1(32'h3bba8844),
	.w2(32'hbb92caf7),
	.w3(32'hbb6cde11),
	.w4(32'h3ba895fc),
	.w5(32'hb9404014),
	.w6(32'hba3ca9c4),
	.w7(32'h3bb9b12e),
	.w8(32'h396e3ec6),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b644696),
	.w1(32'hbc4da136),
	.w2(32'hbcd42a25),
	.w3(32'hbb068fce),
	.w4(32'hbb866b82),
	.w5(32'hbca42e40),
	.w6(32'hbbaa00d7),
	.w7(32'h39b455da),
	.w8(32'hbc2f1078),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9acf0e),
	.w1(32'hbc923c45),
	.w2(32'h39864a20),
	.w3(32'hbcd4e486),
	.w4(32'hbc960b7c),
	.w5(32'hbc8a3f7d),
	.w6(32'hbc17e519),
	.w7(32'h3b6b2b98),
	.w8(32'hbbf4e896),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91c943),
	.w1(32'hbc0b099b),
	.w2(32'h3ab4565f),
	.w3(32'hbc5b49f0),
	.w4(32'h3b23b837),
	.w5(32'hbb9b5a4d),
	.w6(32'hbc4ba100),
	.w7(32'hbad4e5be),
	.w8(32'h3a607c8c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb302e52),
	.w1(32'hba3bf922),
	.w2(32'hba2e8a75),
	.w3(32'hbc37e06c),
	.w4(32'hbc160028),
	.w5(32'hbbe429dd),
	.w6(32'hbba6020e),
	.w7(32'hbb5d3ad9),
	.w8(32'h3a53e738),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeb086),
	.w1(32'hbbabcc50),
	.w2(32'h3b2ac0dc),
	.w3(32'hbbffaeb0),
	.w4(32'hbc14a2c4),
	.w5(32'h3d0280c2),
	.w6(32'h39f18121),
	.w7(32'h3be6c5fa),
	.w8(32'hbc7fab8d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc780ccf),
	.w1(32'hbc907b87),
	.w2(32'h3b41d64f),
	.w3(32'h3d03e57d),
	.w4(32'h3c61ef89),
	.w5(32'h3b0cbce5),
	.w6(32'hbcdda142),
	.w7(32'hbc0392b8),
	.w8(32'h3a88445f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86073a),
	.w1(32'h3a621b11),
	.w2(32'h3a110c1e),
	.w3(32'hb9da7d02),
	.w4(32'h3ad39565),
	.w5(32'h3c749eec),
	.w6(32'hbaa8f14e),
	.w7(32'h392dd8b9),
	.w8(32'hbca4669f),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1867ab),
	.w1(32'h3be0ab49),
	.w2(32'hbbca6e25),
	.w3(32'h3c6287cf),
	.w4(32'h3c10329a),
	.w5(32'h3c3de429),
	.w6(32'hbc81f001),
	.w7(32'hbc5b93e6),
	.w8(32'h3a6fa0c6),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebaba8),
	.w1(32'hbc42d602),
	.w2(32'hbaf1703b),
	.w3(32'h3b366fc2),
	.w4(32'h3b923570),
	.w5(32'hba8ff255),
	.w6(32'hb92ba759),
	.w7(32'h3c82949f),
	.w8(32'hbb9d2771),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032b81),
	.w1(32'h3ae338de),
	.w2(32'hb9cc6102),
	.w3(32'hb9d6ed0c),
	.w4(32'h3b8cb1f3),
	.w5(32'hbc256456),
	.w6(32'hbc03bf21),
	.w7(32'hbb74a45f),
	.w8(32'hbbacd135),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932cb07),
	.w1(32'hbb8e58f0),
	.w2(32'hbb0e23e7),
	.w3(32'hbc992b17),
	.w4(32'hbc50b004),
	.w5(32'hbb39ec85),
	.w6(32'h3bc0b4bb),
	.w7(32'h3bae8b86),
	.w8(32'hbb595ccd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42d0a7),
	.w1(32'hbb88a78a),
	.w2(32'hbc86fb68),
	.w3(32'hbaed82c6),
	.w4(32'hba8f9bf2),
	.w5(32'h3c8fda8c),
	.w6(32'hbaa5c232),
	.w7(32'hb9a68666),
	.w8(32'h3bdeb01a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd14074),
	.w1(32'hbcffbbd1),
	.w2(32'hbbfb19ca),
	.w3(32'h3c9629be),
	.w4(32'h3cef4c77),
	.w5(32'hbad3ea52),
	.w6(32'hbc194014),
	.w7(32'hbc034b7a),
	.w8(32'hbba281c1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaeba2),
	.w1(32'hbbc6f176),
	.w2(32'h3c44d288),
	.w3(32'hba91f84d),
	.w4(32'h3b55e80f),
	.w5(32'h3aec2cd5),
	.w6(32'hbbf5f44d),
	.w7(32'hbb397afe),
	.w8(32'h3c145df5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf2604),
	.w1(32'hbb57c0eb),
	.w2(32'hb97cb929),
	.w3(32'hbbd65e15),
	.w4(32'hbc1c7d8d),
	.w5(32'hba7f70e5),
	.w6(32'h3c8526ee),
	.w7(32'h3c486f0c),
	.w8(32'hbb0e8752),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53564a),
	.w1(32'h3b212758),
	.w2(32'h3b5e5468),
	.w3(32'h3ae13d32),
	.w4(32'h3adcfaf3),
	.w5(32'h3acd2bfe),
	.w6(32'hbbaa8309),
	.w7(32'hba24d8a7),
	.w8(32'hbac3794b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0808ec),
	.w1(32'h3c38a07c),
	.w2(32'h3b40f683),
	.w3(32'hbc08518b),
	.w4(32'h3bc859c9),
	.w5(32'h3c2a4ea7),
	.w6(32'hbc594a2b),
	.w7(32'h3a967d07),
	.w8(32'h39b073cd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a187),
	.w1(32'hbbbc6176),
	.w2(32'h3be972b5),
	.w3(32'h3b21c98e),
	.w4(32'hba614c92),
	.w5(32'hba1bb8c5),
	.w6(32'h3b8dc3b2),
	.w7(32'h3bcc284a),
	.w8(32'hbca71338),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc3776),
	.w1(32'hbc809d7e),
	.w2(32'hbbf33fc1),
	.w3(32'hbb86c532),
	.w4(32'hbb8ef4f7),
	.w5(32'hbb98f3a6),
	.w6(32'hbcda0c6d),
	.w7(32'hbca5197a),
	.w8(32'hbb1e5c3d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663fb8),
	.w1(32'hbc140f7b),
	.w2(32'hb9e835de),
	.w3(32'h3ab2bff0),
	.w4(32'hbae14b14),
	.w5(32'h3b9d9232),
	.w6(32'h3c0b9fe5),
	.w7(32'h3bacd46b),
	.w8(32'hbc66a2e4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadb416),
	.w1(32'hbc83da02),
	.w2(32'hbc64b84c),
	.w3(32'h3c399f83),
	.w4(32'h3c14ea75),
	.w5(32'h3b36c18e),
	.w6(32'hbc0f318d),
	.w7(32'h3ab23d12),
	.w8(32'hbc565cc6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe82569),
	.w1(32'h3bc8f1e0),
	.w2(32'hbc04b1f3),
	.w3(32'h3c4384bd),
	.w4(32'hba4bb519),
	.w5(32'hbb080e33),
	.w6(32'hbbc48b6c),
	.w7(32'h3ba57c44),
	.w8(32'h3c0e3bfe),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0746),
	.w1(32'h3b9a8140),
	.w2(32'hba96dd00),
	.w3(32'hbba52e94),
	.w4(32'h3bff667d),
	.w5(32'hbc146aed),
	.w6(32'h3bb2e70d),
	.w7(32'h3c3ac723),
	.w8(32'hbbf2b47d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32bb0e),
	.w1(32'hba2702b1),
	.w2(32'hbb2dc39b),
	.w3(32'hbc4f3dc4),
	.w4(32'hbb829af2),
	.w5(32'hba7d1c0d),
	.w6(32'h3b460fb5),
	.w7(32'h3b38e0e9),
	.w8(32'hbba2276f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a952e08),
	.w1(32'hbb3c08ea),
	.w2(32'h3bb624f9),
	.w3(32'hbba78bcd),
	.w4(32'hbb8c59a1),
	.w5(32'hbc1a1541),
	.w6(32'hbaa4b2a2),
	.w7(32'h3a5926e8),
	.w8(32'hbc55b056),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487592),
	.w1(32'h3c355b37),
	.w2(32'h3b6ee27f),
	.w3(32'hbc661e69),
	.w4(32'hbc252e76),
	.w5(32'hbbb3d072),
	.w6(32'hbc3c8ad9),
	.w7(32'hbbe4e1e8),
	.w8(32'h3c4e1d2a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60eb3a),
	.w1(32'hbb84de71),
	.w2(32'hbb4a5273),
	.w3(32'hbbad5c10),
	.w4(32'hbb4ab268),
	.w5(32'hba325e06),
	.w6(32'h3c77cae8),
	.w7(32'h3c737c38),
	.w8(32'h3b33524f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe08dea),
	.w1(32'h3b17d415),
	.w2(32'h3b951a23),
	.w3(32'h3a8dbdc2),
	.w4(32'h39ed3f0a),
	.w5(32'hbbfbe303),
	.w6(32'hbac724d6),
	.w7(32'hbc18a71f),
	.w8(32'h3c94e402),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb8073),
	.w1(32'hbbf4b0ff),
	.w2(32'hb9e32c2a),
	.w3(32'hbb8323d5),
	.w4(32'h3b02e854),
	.w5(32'h39e3d03b),
	.w6(32'h3cb23bd3),
	.w7(32'h3caff949),
	.w8(32'hbcbc2ed9),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8e7aa),
	.w1(32'h3b567b8a),
	.w2(32'hbbb4677f),
	.w3(32'h3bcaf407),
	.w4(32'h3b96b008),
	.w5(32'h3c5f1010),
	.w6(32'hbc964800),
	.w7(32'hbc8b5016),
	.w8(32'hbc707321),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc187b15),
	.w1(32'hbc320487),
	.w2(32'hbc276287),
	.w3(32'h3cca5e05),
	.w4(32'h3c442b69),
	.w5(32'h3be33c4f),
	.w6(32'hbc500ef0),
	.w7(32'hbbec9566),
	.w8(32'h3c8c3ded),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f3a99),
	.w1(32'hbc699c1c),
	.w2(32'h3b8a3b18),
	.w3(32'h3b20c34b),
	.w4(32'h3c11c632),
	.w5(32'h3b8ee78e),
	.w6(32'h3c5ca383),
	.w7(32'h3c4b2651),
	.w8(32'hb944f0b6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e1a24),
	.w1(32'h3b597be6),
	.w2(32'hbbeefc54),
	.w3(32'h3a3e40ce),
	.w4(32'hb9f0372b),
	.w5(32'h3b651f18),
	.w6(32'hbb247e82),
	.w7(32'hbb4f1783),
	.w8(32'h3c0977d5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0bca5),
	.w1(32'h3be2dd9c),
	.w2(32'h3c7a8b2f),
	.w3(32'h3b47ba7d),
	.w4(32'hbaa660a8),
	.w5(32'h3c580f00),
	.w6(32'h3b516aa0),
	.w7(32'h3c14bdb8),
	.w8(32'h3c617a24),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e78b3e),
	.w1(32'h3bd81894),
	.w2(32'hbb78d674),
	.w3(32'hbab3e508),
	.w4(32'h3c252b79),
	.w5(32'h3a9a1a66),
	.w6(32'hbc0040d1),
	.w7(32'h3ac5c4df),
	.w8(32'hbb4c196a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab39d5b),
	.w1(32'hbbe3fd24),
	.w2(32'hbc783204),
	.w3(32'h3b2417c4),
	.w4(32'h3bee8fa3),
	.w5(32'hbc2e9a4f),
	.w6(32'hbb8ffa05),
	.w7(32'h3b0e6149),
	.w8(32'hbc1817eb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7047d),
	.w1(32'hbbf27316),
	.w2(32'hbbd760b2),
	.w3(32'h3c0ed9b7),
	.w4(32'hbbaf79c3),
	.w5(32'hbb814896),
	.w6(32'h3c941218),
	.w7(32'h3bf9d450),
	.w8(32'hbbbff798),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacbbce),
	.w1(32'h3be40f81),
	.w2(32'h3c127bc8),
	.w3(32'hbc30cc4e),
	.w4(32'hbb9f1c35),
	.w5(32'hbc35eab5),
	.w6(32'hbafafdb8),
	.w7(32'h3b678158),
	.w8(32'h3c35d64e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3924d3),
	.w1(32'h3bf47bab),
	.w2(32'h3b9a8955),
	.w3(32'hbc91dcec),
	.w4(32'hbc41908b),
	.w5(32'hbc1272b3),
	.w6(32'h3bf30745),
	.w7(32'h3c843d84),
	.w8(32'hbb0f1e40),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636a23),
	.w1(32'hb9279fc3),
	.w2(32'hbb145a26),
	.w3(32'hbb925a32),
	.w4(32'hbb889bf8),
	.w5(32'h3b475214),
	.w6(32'hbb29a068),
	.w7(32'hbb21aec1),
	.w8(32'h3c4fd01d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba899399),
	.w1(32'h3abbf5f8),
	.w2(32'hbb5b02d8),
	.w3(32'h3c825a8c),
	.w4(32'h3cd55a10),
	.w5(32'hbb28a985),
	.w6(32'h3b4c63d9),
	.w7(32'hbc22157a),
	.w8(32'h3afe3f99),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a56f),
	.w1(32'h3b87e943),
	.w2(32'hbb2f06e8),
	.w3(32'hbb8ece8d),
	.w4(32'h3b902001),
	.w5(32'h3bc4bca1),
	.w6(32'hb998667c),
	.w7(32'h3c0218ae),
	.w8(32'h3c35c100),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02189b),
	.w1(32'hbb973afb),
	.w2(32'hbb02d057),
	.w3(32'h3b04c61b),
	.w4(32'h3b9d62a4),
	.w5(32'hb92a68bb),
	.w6(32'h3b264899),
	.w7(32'h3b3e9b27),
	.w8(32'hb9e02d31),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc300295),
	.w1(32'hbb84bc8e),
	.w2(32'h3c66afbe),
	.w3(32'hbac3a893),
	.w4(32'h3a163fc3),
	.w5(32'hbb45f638),
	.w6(32'h3a9f2474),
	.w7(32'hbb1cc679),
	.w8(32'h3c99721a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb243d2b),
	.w1(32'h3b0bf91e),
	.w2(32'hbb5581c7),
	.w3(32'hbc9124ea),
	.w4(32'hbc954d2f),
	.w5(32'hbc1b69f2),
	.w6(32'h3c0cc987),
	.w7(32'h3be50c04),
	.w8(32'hbb0b212d),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee4383),
	.w1(32'hbb0694b1),
	.w2(32'hbc92d407),
	.w3(32'hbc2fbd1b),
	.w4(32'hbbce8d6e),
	.w5(32'hba81b7a4),
	.w6(32'hbb583c41),
	.w7(32'h3b9667f8),
	.w8(32'hbb123e76),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3711),
	.w1(32'h3b3a0544),
	.w2(32'h3b3f3a35),
	.w3(32'h3b1e22dc),
	.w4(32'h3ad8330f),
	.w5(32'hb9d379c8),
	.w6(32'h39cde733),
	.w7(32'hbb14e649),
	.w8(32'h3a8448ea),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad519ee),
	.w1(32'h3bac35db),
	.w2(32'hbbc18457),
	.w3(32'h3aa2f00f),
	.w4(32'h3b88dd22),
	.w5(32'hba6ebb5f),
	.w6(32'hbba1d83b),
	.w7(32'hbb1ea778),
	.w8(32'h391bb700),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0799b),
	.w1(32'h3c08588c),
	.w2(32'h3bbdaac8),
	.w3(32'h3bbd3055),
	.w4(32'h3bcb3789),
	.w5(32'h3c9a0e4b),
	.w6(32'h3ab871ba),
	.w7(32'h3b0f658b),
	.w8(32'hbc233f90),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b1dbd),
	.w1(32'h3b3f5478),
	.w2(32'hbb4c052b),
	.w3(32'h3c632020),
	.w4(32'h3c2c3630),
	.w5(32'hba03889b),
	.w6(32'hbc4ae8e9),
	.w7(32'hbc835122),
	.w8(32'hbb86e84e),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb038300),
	.w1(32'hbb2512da),
	.w2(32'h3aaea6ea),
	.w3(32'hbb2140dd),
	.w4(32'hba27ed6a),
	.w5(32'hbbb575d9),
	.w6(32'hbb481178),
	.w7(32'h39c14215),
	.w8(32'hbb7e5e06),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79239b),
	.w1(32'h3c28520b),
	.w2(32'h3bb119a4),
	.w3(32'hbc0520c8),
	.w4(32'hbb561429),
	.w5(32'hbc6eaeaf),
	.w6(32'hbc0360aa),
	.w7(32'hbbe698e3),
	.w8(32'h3c4c9c43),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc5c5c),
	.w1(32'h3baf5d2d),
	.w2(32'hbba36fcc),
	.w3(32'hbc2b79e9),
	.w4(32'h3b2a7154),
	.w5(32'hbbf9283b),
	.w6(32'hbb875293),
	.w7(32'hbbe7e832),
	.w8(32'hba2e7421),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1df037),
	.w1(32'h3b040e9f),
	.w2(32'hbae3eaeb),
	.w3(32'hbb60a6fc),
	.w4(32'h3b5794d4),
	.w5(32'hba76379f),
	.w6(32'hbc1c6449),
	.w7(32'hbc44a547),
	.w8(32'hbbc5cc38),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b96a3),
	.w1(32'hbb399313),
	.w2(32'h3b696a03),
	.w3(32'hbbb63139),
	.w4(32'hba6020e7),
	.w5(32'hbb992657),
	.w6(32'hbbbe20f6),
	.w7(32'hb9ab9c0c),
	.w8(32'hbaeac28d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc06e9e),
	.w1(32'h3b763316),
	.w2(32'hbbc86c3f),
	.w3(32'hbc2fe716),
	.w4(32'hbbc6c283),
	.w5(32'hbb878e27),
	.w6(32'hbb799660),
	.w7(32'h3b8798bb),
	.w8(32'hba35632b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28989),
	.w1(32'hbbc81063),
	.w2(32'hbba16790),
	.w3(32'hbbb950b8),
	.w4(32'hba4d4b95),
	.w5(32'hbbb90130),
	.w6(32'h3aef8dd3),
	.w7(32'h3b25a43a),
	.w8(32'h3a192f3f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a30f6),
	.w1(32'h39f9ccf3),
	.w2(32'h3c385491),
	.w3(32'hbb35f36c),
	.w4(32'hba3ec361),
	.w5(32'hbb446657),
	.w6(32'h3ae3b9ce),
	.w7(32'h3b7229a7),
	.w8(32'hb9d61359),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c288f42),
	.w1(32'hbaa98d23),
	.w2(32'hbae1bacb),
	.w3(32'hbbed08d1),
	.w4(32'h3a80f387),
	.w5(32'hbaf855d5),
	.w6(32'hbb6a9874),
	.w7(32'hbba78c2c),
	.w8(32'h3c46711a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf76242),
	.w1(32'h3c0f9a86),
	.w2(32'h3b227ce9),
	.w3(32'hbc8b2a39),
	.w4(32'hbc429c7d),
	.w5(32'hbad04bb3),
	.w6(32'hbbdfb7ce),
	.w7(32'hbbf103c0),
	.w8(32'h3bf97c51),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba65db9),
	.w1(32'h3b6308ef),
	.w2(32'hb9827dd3),
	.w3(32'hbc685688),
	.w4(32'hba90b7ba),
	.w5(32'hbb71488a),
	.w6(32'hb9d68815),
	.w7(32'h3b9a6258),
	.w8(32'h3c44298a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1c37b),
	.w1(32'hbacdf6c6),
	.w2(32'h3b5a3f2b),
	.w3(32'hbbf6e3ce),
	.w4(32'hbbfaeaa3),
	.w5(32'h3b1bc1ea),
	.w6(32'hbba06392),
	.w7(32'hba132cd4),
	.w8(32'h3b8356f2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe7137),
	.w1(32'h3b9db567),
	.w2(32'hbca525cc),
	.w3(32'hbc6d437a),
	.w4(32'hbb68a6b3),
	.w5(32'hbc49949b),
	.w6(32'hbb8b4f2b),
	.w7(32'h3c35fcde),
	.w8(32'hbb0f085b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b3550),
	.w1(32'hbaa3f75e),
	.w2(32'h3bd41fb4),
	.w3(32'hbb11d7bb),
	.w4(32'hbb505e80),
	.w5(32'hbb10437e),
	.w6(32'h3b7e77ca),
	.w7(32'h3ba34634),
	.w8(32'h3c47af6b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6216a),
	.w1(32'hbb8f2cf9),
	.w2(32'hba9c4a85),
	.w3(32'hbbfac694),
	.w4(32'hbc201ef9),
	.w5(32'h3c553982),
	.w6(32'h3c64a9de),
	.w7(32'h3c11e7ad),
	.w8(32'hbbb898d0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb68aae),
	.w1(32'h3b8be442),
	.w2(32'h3b9db398),
	.w3(32'h3b86dbd0),
	.w4(32'h3c9fa154),
	.w5(32'h3c9995f5),
	.w6(32'hbc67dfb5),
	.w7(32'h3c043e05),
	.w8(32'h3ca5600e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4ae65),
	.w1(32'hbbfeb6b9),
	.w2(32'hbc7ec34e),
	.w3(32'hbb809ef9),
	.w4(32'h3bed5d63),
	.w5(32'hbbe1556e),
	.w6(32'hbab7aff4),
	.w7(32'h3c487d85),
	.w8(32'hb9b2fb23),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc51fc0),
	.w1(32'h3b98fd72),
	.w2(32'hbb5f1084),
	.w3(32'h39e1abd4),
	.w4(32'h3b0e6768),
	.w5(32'h3b77be34),
	.w6(32'h3b96405f),
	.w7(32'h3c5dfd9f),
	.w8(32'h3aaac347),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01be4f),
	.w1(32'h3a68f6d1),
	.w2(32'hbb877e08),
	.w3(32'hbc08dc90),
	.w4(32'hbab95565),
	.w5(32'hbb7cb526),
	.w6(32'hbc225c0c),
	.w7(32'hbbd9552e),
	.w8(32'h3ab8b71d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3948f7),
	.w1(32'hbbebcdd8),
	.w2(32'h3c369894),
	.w3(32'hbc685c21),
	.w4(32'hbc4e91d3),
	.w5(32'hbc3e68cc),
	.w6(32'hba21bb21),
	.w7(32'hbbca2d9d),
	.w8(32'h3ba0f75b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006921),
	.w1(32'h3ab6b0b7),
	.w2(32'h3c3b45f6),
	.w3(32'hbc8e3768),
	.w4(32'hbc92a03b),
	.w5(32'hbc042195),
	.w6(32'h3c0dbc0c),
	.w7(32'h3be5f61d),
	.w8(32'hbba89ffc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dd8d1),
	.w1(32'h3c5db6d9),
	.w2(32'h3a2de936),
	.w3(32'hbc7b9d36),
	.w4(32'hbc4226b9),
	.w5(32'hba6833a5),
	.w6(32'hbac64a55),
	.w7(32'h3c1ac73d),
	.w8(32'hbc13b6fa),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b0995),
	.w1(32'hbba7d3bc),
	.w2(32'hbb001063),
	.w3(32'hba05f7db),
	.w4(32'h3b8c1dd6),
	.w5(32'hbc0d3525),
	.w6(32'hbc9c5ddc),
	.w7(32'hbc41fc30),
	.w8(32'h3ca0cef0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096845),
	.w1(32'h3c166c81),
	.w2(32'h3b48ac40),
	.w3(32'hbc95f34b),
	.w4(32'hbc2d109d),
	.w5(32'h3b3c31a0),
	.w6(32'h3b87c583),
	.w7(32'h3c70b5fe),
	.w8(32'hb99f3bdf),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1ffe),
	.w1(32'h3b84a044),
	.w2(32'h3b0d65ba),
	.w3(32'h3a6d16c7),
	.w4(32'h3a0f3792),
	.w5(32'h3c02925b),
	.w6(32'hbbf25b62),
	.w7(32'hbc30ed8a),
	.w8(32'h3bb6037f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9570a41),
	.w1(32'h3bdba328),
	.w2(32'h3bf8d210),
	.w3(32'hbbb09c99),
	.w4(32'h3c099ea8),
	.w5(32'h3cccb3d6),
	.w6(32'hbbd2b879),
	.w7(32'h3bff3155),
	.w8(32'hbcc1846e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabcebe6),
	.w1(32'hbbf593e5),
	.w2(32'hbc2828de),
	.w3(32'h3c9539e4),
	.w4(32'h3ca2d1b5),
	.w5(32'h3c47099b),
	.w6(32'hbcc129f8),
	.w7(32'hbc8e9a81),
	.w8(32'hbc103801),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2188d3),
	.w1(32'hbac309a4),
	.w2(32'h3b401c70),
	.w3(32'h3cdec498),
	.w4(32'h3cab5951),
	.w5(32'h3b3a886d),
	.w6(32'hbc6b0a9b),
	.w7(32'hbc6601c3),
	.w8(32'h3a5d8d04),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba44fa2),
	.w1(32'h3bd247a3),
	.w2(32'hbac06d0d),
	.w3(32'h39f261af),
	.w4(32'h390473f8),
	.w5(32'h3c231336),
	.w6(32'hbbca409c),
	.w7(32'h3b3cf73a),
	.w8(32'h3c5b98a3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b100),
	.w1(32'hbb98e7a9),
	.w2(32'hbc318347),
	.w3(32'h3a36dc4d),
	.w4(32'h3bd9a6a5),
	.w5(32'hbb1ada71),
	.w6(32'hbadebbe3),
	.w7(32'h3ad95ce3),
	.w8(32'h3bdd220f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5aa20),
	.w1(32'hbc0275e5),
	.w2(32'hba99c992),
	.w3(32'hbc0dc488),
	.w4(32'hbbcff507),
	.w5(32'h3890fd6b),
	.w6(32'h3c275a1a),
	.w7(32'h3c16e7d8),
	.w8(32'hba879495),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af43a29),
	.w1(32'hbaa3bca3),
	.w2(32'hbc016cc7),
	.w3(32'h3b340965),
	.w4(32'h3b26a548),
	.w5(32'hb9e0ef5c),
	.w6(32'hbb86b52c),
	.w7(32'h3ae99b5e),
	.w8(32'h3b462d89),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb637d13),
	.w1(32'hbba701e0),
	.w2(32'hbb072880),
	.w3(32'hb9c6c5a3),
	.w4(32'h3a7ac485),
	.w5(32'h3ad7d53c),
	.w6(32'hba833095),
	.w7(32'h3adda25b),
	.w8(32'hbb9f2bdf),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaca7a8),
	.w1(32'h3bdf7be8),
	.w2(32'h3abadb93),
	.w3(32'h3b6a0c47),
	.w4(32'h3ba3754a),
	.w5(32'hbc246979),
	.w6(32'hbbd60590),
	.w7(32'hbc1f390b),
	.w8(32'h3c1c9a93),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6811d),
	.w1(32'h3ba76d8a),
	.w2(32'hbaec21ab),
	.w3(32'hbc777fe7),
	.w4(32'hbb5842ce),
	.w5(32'h3c909194),
	.w6(32'h3b851b4c),
	.w7(32'h3b99d9a7),
	.w8(32'hbcaa805f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d169c),
	.w1(32'h39d9c4e4),
	.w2(32'h3c01bb10),
	.w3(32'h3c9de4b5),
	.w4(32'h3c6fb493),
	.w5(32'hbc902b2f),
	.w6(32'hbcf7a367),
	.w7(32'hbcc89817),
	.w8(32'h3c09fb06),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e17cc),
	.w1(32'h3b7efac2),
	.w2(32'h3bcaeffa),
	.w3(32'hbcca328f),
	.w4(32'hbc3edca3),
	.w5(32'hbb9d752c),
	.w6(32'h3acdfee0),
	.w7(32'h3bda59cc),
	.w8(32'h3c25c125),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd3964),
	.w1(32'h3b7ad6f7),
	.w2(32'hbc1e8c5f),
	.w3(32'hbc32ef0e),
	.w4(32'hbb8b6432),
	.w5(32'hbc32a4bf),
	.w6(32'h3c857c78),
	.w7(32'h3c497fda),
	.w8(32'h38aeb591),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307888),
	.w1(32'h3ae698b2),
	.w2(32'hba1f8200),
	.w3(32'hbb419940),
	.w4(32'hb9758bc1),
	.w5(32'h3bfaa531),
	.w6(32'h3bf2ae20),
	.w7(32'h3c47ce17),
	.w8(32'hbc9e17c9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c632f39),
	.w1(32'hb9c704f5),
	.w2(32'hbc68a0a7),
	.w3(32'h3b9b8b3f),
	.w4(32'h3c24a1a1),
	.w5(32'hba8a471b),
	.w6(32'hbc7dabf7),
	.w7(32'hbc51337e),
	.w8(32'hbc469ba2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89ff03),
	.w1(32'hbbdbd23a),
	.w2(32'hbb680e64),
	.w3(32'h3b743ba3),
	.w4(32'h3a6ca2e8),
	.w5(32'h3b730ca8),
	.w6(32'h3b4644d9),
	.w7(32'h3b107d21),
	.w8(32'hbaadde79),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13e1cf),
	.w1(32'hba213474),
	.w2(32'hbb9439cd),
	.w3(32'h3aed77f4),
	.w4(32'h3ad1bc22),
	.w5(32'hbabd15dd),
	.w6(32'hbae068b4),
	.w7(32'h3a350485),
	.w8(32'hbbac900f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9b969),
	.w1(32'hbb8712d0),
	.w2(32'hbc011d0c),
	.w3(32'hb8c435bb),
	.w4(32'hbaf760d9),
	.w5(32'hbbb9e6fe),
	.w6(32'hbba8d6ee),
	.w7(32'hbc170844),
	.w8(32'hb9f213e3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cafb8),
	.w1(32'hbbfb2730),
	.w2(32'hbbbdb7fe),
	.w3(32'hbbbb61d5),
	.w4(32'hbc00a8c9),
	.w5(32'h3c027246),
	.w6(32'h3a8bc9a2),
	.w7(32'h3a9afea0),
	.w8(32'hbce67483),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8f20),
	.w1(32'h3b91dc2c),
	.w2(32'hbc002f08),
	.w3(32'h3c766dc7),
	.w4(32'h3c45d12d),
	.w5(32'h3c7f21a0),
	.w6(32'hbd217a97),
	.w7(32'hbd1f339a),
	.w8(32'hbc807110),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba109d5c),
	.w1(32'hb9b473d1),
	.w2(32'h3c5c1ecb),
	.w3(32'h3cfa0e79),
	.w4(32'h3cb00a43),
	.w5(32'hbb03fb35),
	.w6(32'hbbb73f85),
	.w7(32'hbbc5a960),
	.w8(32'h3b61182a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc057d5),
	.w1(32'h3c014f59),
	.w2(32'h3a91d30c),
	.w3(32'hbc04f859),
	.w4(32'hbbf9671f),
	.w5(32'h3b41d901),
	.w6(32'h3b09bd56),
	.w7(32'h3c1d989e),
	.w8(32'h3a9d6665),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b997df5),
	.w1(32'h3b9d7d69),
	.w2(32'h3b1c0d99),
	.w3(32'h3bb70395),
	.w4(32'h3b9e58eb),
	.w5(32'h3b2f97f9),
	.w6(32'h3b897a5c),
	.w7(32'h3b4ad149),
	.w8(32'hba2295c6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6209fc),
	.w1(32'h3a311a09),
	.w2(32'h393a517a),
	.w3(32'h39aa043a),
	.w4(32'hbb045b09),
	.w5(32'hba43abbf),
	.w6(32'hba2b185b),
	.w7(32'hbb20d2a5),
	.w8(32'h3a19bf16),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a9662),
	.w1(32'hbc02e37c),
	.w2(32'h371a2cd3),
	.w3(32'h3a0e6c8b),
	.w4(32'h3b1fb82c),
	.w5(32'h3aa6580f),
	.w6(32'h3c133310),
	.w7(32'h3c425796),
	.w8(32'h3b2c5ff4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a1c6f),
	.w1(32'hbb897850),
	.w2(32'hbabe5c83),
	.w3(32'h3abd2b87),
	.w4(32'hbb037560),
	.w5(32'h3b943010),
	.w6(32'h3b068ae5),
	.w7(32'h3b548e4b),
	.w8(32'h3bf531c3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd6be),
	.w1(32'hbbf336f3),
	.w2(32'hbc559d8f),
	.w3(32'hbb0759d7),
	.w4(32'h3bf29dac),
	.w5(32'hbb4fd18d),
	.w6(32'h3c2babd1),
	.w7(32'h3ccc6138),
	.w8(32'hbc6ce3e4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3c0ab),
	.w1(32'hb99ecfca),
	.w2(32'hbbdbf765),
	.w3(32'h3b16b916),
	.w4(32'h3ba84253),
	.w5(32'h3a61a97a),
	.w6(32'h3c10c7d5),
	.w7(32'h3b3980fa),
	.w8(32'hbb0f6265),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5799dd),
	.w1(32'hbb64f9d5),
	.w2(32'h3bd74b14),
	.w3(32'hbc484b0e),
	.w4(32'hba29fe4a),
	.w5(32'hbaf757dd),
	.w6(32'hbbe74b05),
	.w7(32'h3b6fcc0d),
	.w8(32'h3b34eb13),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule