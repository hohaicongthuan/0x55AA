module layer_8_featuremap_154(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16f690),
	.w1(32'h3a2afa0a),
	.w2(32'hbbce8596),
	.w3(32'h3b2930a9),
	.w4(32'h3b1758fa),
	.w5(32'h39765c7b),
	.w6(32'h3b2a8619),
	.w7(32'h3b9c95b0),
	.w8(32'hba19c84d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd831e3),
	.w1(32'hbba304d7),
	.w2(32'h3b03c4a3),
	.w3(32'hbb9aebd5),
	.w4(32'h3b240b32),
	.w5(32'h3bdd6bd2),
	.w6(32'hbaafda6b),
	.w7(32'h3b337443),
	.w8(32'h3b95693c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b782d7f),
	.w1(32'hbb6ad518),
	.w2(32'hbb01eb94),
	.w3(32'hbb1f17d5),
	.w4(32'hbabb32e7),
	.w5(32'h3bc19725),
	.w6(32'hbb868314),
	.w7(32'hbb306779),
	.w8(32'h3a3b50e3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28f205),
	.w1(32'hba8ec5c6),
	.w2(32'h3b6b4dd4),
	.w3(32'h3b413ac2),
	.w4(32'hbad5e9af),
	.w5(32'h3a72b730),
	.w6(32'hb92665ee),
	.w7(32'h3b788b0a),
	.w8(32'h3bdcff1d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c108762),
	.w1(32'h3b08c84b),
	.w2(32'hbae30d6d),
	.w3(32'h3c05256e),
	.w4(32'h3ba7fcc1),
	.w5(32'hbb14667e),
	.w6(32'h3c31a041),
	.w7(32'h3aa9e90d),
	.w8(32'hbb9f0ddc),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb820d5d),
	.w1(32'h3b0d58d3),
	.w2(32'h3be60373),
	.w3(32'hbbae2ec8),
	.w4(32'hbb3536c1),
	.w5(32'hba77961d),
	.w6(32'hbabff290),
	.w7(32'hbb3088c9),
	.w8(32'h3bcf1ac5),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3f35),
	.w1(32'hbadd39fd),
	.w2(32'h3b4bffe5),
	.w3(32'h3c0277a1),
	.w4(32'hba956358),
	.w5(32'h3add5741),
	.w6(32'h3beea4c8),
	.w7(32'hbaca1dd9),
	.w8(32'h3b4a7da8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab82516),
	.w1(32'h39273a03),
	.w2(32'hbba671e3),
	.w3(32'h3afb0c3a),
	.w4(32'hbc36c480),
	.w5(32'hbbb2b7a6),
	.w6(32'h399375aa),
	.w7(32'hbb9e2656),
	.w8(32'hbb2f58ea),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc72afe),
	.w1(32'hbc3f9edb),
	.w2(32'h3bb2994f),
	.w3(32'hba5ea8b7),
	.w4(32'h3bd073bc),
	.w5(32'h3bf475cc),
	.w6(32'hbbd5c985),
	.w7(32'h3c48ffac),
	.w8(32'h3c8ed4ea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23d778),
	.w1(32'h3bab14a3),
	.w2(32'h3c072208),
	.w3(32'h3c67844b),
	.w4(32'h3a89d7ef),
	.w5(32'h3acac547),
	.w6(32'h3c9ce125),
	.w7(32'h3be90ccc),
	.w8(32'h3bfb348b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67b8be),
	.w1(32'h3b98bc91),
	.w2(32'h3b6a234d),
	.w3(32'h3b5f4c47),
	.w4(32'h3ae06b97),
	.w5(32'hb89513c9),
	.w6(32'h3c076eef),
	.w7(32'h3b0b8799),
	.w8(32'hbb87b470),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36e75b),
	.w1(32'hbbc68e7b),
	.w2(32'h3946f196),
	.w3(32'h3a8d4ebc),
	.w4(32'hbabe7c32),
	.w5(32'h3b4c7a5a),
	.w6(32'hbb306de0),
	.w7(32'hbaacb79e),
	.w8(32'hbb89d95c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb68e),
	.w1(32'hbc1579a1),
	.w2(32'hba45c1a6),
	.w3(32'hbbae5254),
	.w4(32'hba87a257),
	.w5(32'h3911a6af),
	.w6(32'hbc30f4b5),
	.w7(32'hbba56e66),
	.w8(32'h3aae5bc4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28e2b3),
	.w1(32'h3bcc82df),
	.w2(32'hbae051d3),
	.w3(32'h3b1be1a5),
	.w4(32'h3b13de41),
	.w5(32'h3a8eafb0),
	.w6(32'h3b964dc7),
	.w7(32'hbb9eb30a),
	.w8(32'hbbe53e7c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf947b2),
	.w1(32'h3aef32d5),
	.w2(32'h3b337ae1),
	.w3(32'h3b5ee588),
	.w4(32'h3b8cd1bc),
	.w5(32'h3adc76b6),
	.w6(32'h3a717513),
	.w7(32'h3a4afd4e),
	.w8(32'hbbc4bd67),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac76aac),
	.w1(32'h3c03bc6f),
	.w2(32'hbb93651f),
	.w3(32'h3ba118eb),
	.w4(32'h3ad5d4d8),
	.w5(32'h3b87704a),
	.w6(32'h396e464c),
	.w7(32'h3bfd7bfa),
	.w8(32'hbc98e41c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa52b8a),
	.w1(32'hb9cd4882),
	.w2(32'hbae99b1d),
	.w3(32'h39f674e2),
	.w4(32'hbbbf6c31),
	.w5(32'hbc4b1d5c),
	.w6(32'hbba4efa8),
	.w7(32'h3bb67e3d),
	.w8(32'h3c0c98a2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb72342),
	.w1(32'hbc21b355),
	.w2(32'hbc2d187a),
	.w3(32'h3bf03770),
	.w4(32'h3afcad8f),
	.w5(32'hbc784c0f),
	.w6(32'hbc55ec8b),
	.w7(32'h3c4fb6ee),
	.w8(32'hbc664026),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29154b),
	.w1(32'hbb894e91),
	.w2(32'hbc5941d9),
	.w3(32'h3c921d7a),
	.w4(32'hbc0d7195),
	.w5(32'hbc76cea0),
	.w6(32'hbaae26a8),
	.w7(32'h3c3212db),
	.w8(32'hbbf57422),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4fcae),
	.w1(32'hbcdab639),
	.w2(32'hbc6a3843),
	.w3(32'h3c294fc4),
	.w4(32'hbaf503c8),
	.w5(32'hbc64f7a0),
	.w6(32'hbc939852),
	.w7(32'hbb5c874e),
	.w8(32'hbc3592f3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4509),
	.w1(32'h3bff9d5e),
	.w2(32'hbc56722d),
	.w3(32'h3bf9d2a0),
	.w4(32'hbcdaf83e),
	.w5(32'h3d32cbc2),
	.w6(32'hbbce8aea),
	.w7(32'h3d0c6f51),
	.w8(32'hbda934d8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c862efd),
	.w1(32'hbc9aa3c8),
	.w2(32'hbba6d60e),
	.w3(32'hbcc868ac),
	.w4(32'h3b3fa6ee),
	.w5(32'hbbd7c45a),
	.w6(32'h3d45f183),
	.w7(32'h3b0cf4e7),
	.w8(32'hbb54942c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c778c9f),
	.w1(32'hbb7c38eb),
	.w2(32'hbace47bc),
	.w3(32'hbc6cafcb),
	.w4(32'hbc08d4e2),
	.w5(32'h3b2e79fb),
	.w6(32'hbc6b2024),
	.w7(32'h3c0dc81b),
	.w8(32'hbd5045ed),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b061),
	.w1(32'h38b0cb7f),
	.w2(32'hbb8b1f5e),
	.w3(32'h3b2114fe),
	.w4(32'h3c1abcf7),
	.w5(32'h3a8dd27a),
	.w6(32'h3c21215d),
	.w7(32'h3b8d8e04),
	.w8(32'h3c544856),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf7b13),
	.w1(32'h3be4d601),
	.w2(32'h3b42f62a),
	.w3(32'h3a0dbcaa),
	.w4(32'hbbff4e07),
	.w5(32'hbbb260d5),
	.w6(32'hbbb922b4),
	.w7(32'hbb62623c),
	.w8(32'hbcbf587e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b417461),
	.w1(32'hbbc2752f),
	.w2(32'hbc4d9d96),
	.w3(32'h3b027696),
	.w4(32'h3afdfd19),
	.w5(32'h3bde5d40),
	.w6(32'h3c044822),
	.w7(32'h3af4bd05),
	.w8(32'h3ceb8b1e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca12fb2),
	.w1(32'h3b8d2f27),
	.w2(32'h3b8f0f27),
	.w3(32'h3c3f4f3b),
	.w4(32'hba67bf7a),
	.w5(32'h3c3329c8),
	.w6(32'hbbb1eb0b),
	.w7(32'hbb996be5),
	.w8(32'h3bb2d337),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159454),
	.w1(32'hbc418e4d),
	.w2(32'hbb544d1f),
	.w3(32'h3c216092),
	.w4(32'h37ca996d),
	.w5(32'hb890ba45),
	.w6(32'h3c2768b4),
	.w7(32'hbc8b6a52),
	.w8(32'hbb7cb40f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0cad5),
	.w1(32'h3bf51c1e),
	.w2(32'hbc1c9dd4),
	.w3(32'hbbf22af9),
	.w4(32'h3b2d634e),
	.w5(32'hbccf59aa),
	.w6(32'hbbaf5f09),
	.w7(32'hbc902b22),
	.w8(32'h3cc89207),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad96455),
	.w1(32'hbc0f2f4d),
	.w2(32'hbc7c97fe),
	.w3(32'h3c39ee93),
	.w4(32'hbc4c0e36),
	.w5(32'h3c44bbf7),
	.w6(32'hbcb5c3fc),
	.w7(32'h3cf2cdd2),
	.w8(32'hbd3bd711),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3be5d0),
	.w1(32'hbb92ce15),
	.w2(32'h3c2c8852),
	.w3(32'h3af9faad),
	.w4(32'h3c6d1018),
	.w5(32'h3c0383d4),
	.w6(32'h3d0326e9),
	.w7(32'h3bc9ae50),
	.w8(32'h3b080ccc),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a09e2),
	.w1(32'h3af39686),
	.w2(32'hbc515a3c),
	.w3(32'h3b13de50),
	.w4(32'h3ad4d9ac),
	.w5(32'hba8449ff),
	.w6(32'hbb96439a),
	.w7(32'hbb148753),
	.w8(32'hbd208087),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95fe82),
	.w1(32'hbc0e728e),
	.w2(32'h3c4836b1),
	.w3(32'hbc043e59),
	.w4(32'hbc2c071d),
	.w5(32'h3b26c61c),
	.w6(32'hb910ceff),
	.w7(32'hbbb73923),
	.w8(32'h3c6f5f38),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccff764),
	.w1(32'hbb953baf),
	.w2(32'hbc15f06a),
	.w3(32'h3bfd22a0),
	.w4(32'hbad1c649),
	.w5(32'h3c3008b5),
	.w6(32'h3c11cc49),
	.w7(32'h3c5ef9ab),
	.w8(32'hbd46b198),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c1237),
	.w1(32'h3bdae820),
	.w2(32'hba36b4f8),
	.w3(32'hbc8ef37c),
	.w4(32'h3a8f0c10),
	.w5(32'h3b959b51),
	.w6(32'h3c17320f),
	.w7(32'h3beab0de),
	.w8(32'hbc2788c8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3bab),
	.w1(32'h3b611d81),
	.w2(32'hbc3a1267),
	.w3(32'h3a940d96),
	.w4(32'hbbcba3a0),
	.w5(32'hbc95d8f7),
	.w6(32'h3c335c28),
	.w7(32'h3cd44b59),
	.w8(32'h3c1c15bd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b765a),
	.w1(32'h3c314d98),
	.w2(32'hbb8374c1),
	.w3(32'hba6ee6b9),
	.w4(32'h3bcb6ecf),
	.w5(32'hbc4b224b),
	.w6(32'hbc366543),
	.w7(32'hbc3d6f3d),
	.w8(32'h3c11bec5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229d7c),
	.w1(32'hbb889101),
	.w2(32'h3c3ac86d),
	.w3(32'h3c1048bb),
	.w4(32'h3c5ca10c),
	.w5(32'hbb9809e4),
	.w6(32'hbc813787),
	.w7(32'h3a6ac013),
	.w8(32'h3c28029f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb60fd3),
	.w1(32'h3bd31108),
	.w2(32'hbce0532c),
	.w3(32'h3bfd7abf),
	.w4(32'hbb3780ff),
	.w5(32'hbc706f8f),
	.w6(32'h3c295dd7),
	.w7(32'hbb82d0e5),
	.w8(32'hbc1736ed),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c897ec9),
	.w1(32'h37b19cd7),
	.w2(32'h3b12cc1a),
	.w3(32'hbc077614),
	.w4(32'h3c2600f7),
	.w5(32'h3bc0e0af),
	.w6(32'hbd0c6212),
	.w7(32'h3b8844df),
	.w8(32'hbbded45a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d90d5),
	.w1(32'hbbe34b51),
	.w2(32'hbc2642bc),
	.w3(32'h3be41b23),
	.w4(32'hbbbc8d7c),
	.w5(32'hbbb2c8df),
	.w6(32'h3bf38b05),
	.w7(32'h3c3e4d4a),
	.w8(32'hbc96ec34),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9ae94),
	.w1(32'hbb390399),
	.w2(32'hbbc20e9f),
	.w3(32'h3bd40903),
	.w4(32'hbbed04c4),
	.w5(32'hbc1df529),
	.w6(32'hbbd9e504),
	.w7(32'h3c89a700),
	.w8(32'hbcd6dcfd),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f9216),
	.w1(32'hbbad4772),
	.w2(32'h3b9b8e97),
	.w3(32'h3cbd96b8),
	.w4(32'hbcdca0a9),
	.w5(32'hbb3c65e4),
	.w6(32'hb9e19792),
	.w7(32'h3c67bfcd),
	.w8(32'hbca7e1d9),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40da13),
	.w1(32'h3c5b41c5),
	.w2(32'hba810de6),
	.w3(32'hbb07aa85),
	.w4(32'hb9fb167d),
	.w5(32'h38239a75),
	.w6(32'h3c118ce3),
	.w7(32'hbc041cf8),
	.w8(32'h3b3eab13),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d895e),
	.w1(32'h3c1c89dc),
	.w2(32'hbcb6ca47),
	.w3(32'h3c0827f8),
	.w4(32'h3bb68fa8),
	.w5(32'hbcaf4f66),
	.w6(32'h3c406230),
	.w7(32'hbbf8558d),
	.w8(32'h3d126e00),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2c283),
	.w1(32'h3ae830fb),
	.w2(32'hb8735488),
	.w3(32'h3ba16f33),
	.w4(32'h3c9812f4),
	.w5(32'hbd1470ae),
	.w6(32'hbbf329f6),
	.w7(32'hbc1b9425),
	.w8(32'h3d266d45),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccad62),
	.w1(32'h3bb47b86),
	.w2(32'h3bdf0e59),
	.w3(32'h3c29cd50),
	.w4(32'hbc47e04e),
	.w5(32'h3c141c27),
	.w6(32'hbcafc446),
	.w7(32'hbbe046b0),
	.w8(32'h3c815354),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa6b7c),
	.w1(32'h3b9a7fa2),
	.w2(32'hbd0a5c3b),
	.w3(32'hbc766386),
	.w4(32'h3b94e57a),
	.w5(32'hbcf9b320),
	.w6(32'h3c26517a),
	.w7(32'hbb4c5e92),
	.w8(32'h3d5eaa35),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af571e8),
	.w1(32'h3c77f2c9),
	.w2(32'h3c07c1bc),
	.w3(32'hbbcc045d),
	.w4(32'hbb325004),
	.w5(32'h3c410098),
	.w6(32'h3986a462),
	.w7(32'hbc402a77),
	.w8(32'hbbc35c93),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91cb9c),
	.w1(32'hb967a7f2),
	.w2(32'hbc0ce576),
	.w3(32'hbbae2338),
	.w4(32'hbb29959f),
	.w5(32'hbc537276),
	.w6(32'h3c9b9bce),
	.w7(32'hbb754fd1),
	.w8(32'h3a5176ab),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ce557),
	.w1(32'hbc2a9f5b),
	.w2(32'hbba27ec4),
	.w3(32'hbc8b39f8),
	.w4(32'h3b6a0b63),
	.w5(32'hbce61022),
	.w6(32'hbc7c3660),
	.w7(32'hbcff5a24),
	.w8(32'h3cc9fb06),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688239),
	.w1(32'hbcd32c52),
	.w2(32'h3bcaa303),
	.w3(32'h3bf15772),
	.w4(32'hbc65b8f9),
	.w5(32'h3bd313fa),
	.w6(32'hbcf41ff2),
	.w7(32'hbb89b04f),
	.w8(32'hba5b0454),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d68d1),
	.w1(32'hbc50d81a),
	.w2(32'hbadf94e8),
	.w3(32'hba2688d9),
	.w4(32'hbc7179fe),
	.w5(32'h3bd47dd9),
	.w6(32'h3c6d9c9f),
	.w7(32'hbc36d086),
	.w8(32'hbc8dc2ba),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc271950),
	.w1(32'hbb0f47c0),
	.w2(32'hbb37f404),
	.w3(32'h3b871260),
	.w4(32'h3acbe1e8),
	.w5(32'hba692479),
	.w6(32'h3c29e6c0),
	.w7(32'hbbe226b5),
	.w8(32'hba0e74b3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a1ed2),
	.w1(32'h3bd9c090),
	.w2(32'hba5ade54),
	.w3(32'h3ab6d509),
	.w4(32'h3b59ddeb),
	.w5(32'hbc662265),
	.w6(32'h39205dec),
	.w7(32'hbccc15a1),
	.w8(32'h3d4a7af5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8afad),
	.w1(32'hbb8dad25),
	.w2(32'hbc0db57e),
	.w3(32'h3bacbef3),
	.w4(32'hbb998588),
	.w5(32'hbc2e3851),
	.w6(32'hbc810f67),
	.w7(32'hbc385611),
	.w8(32'h3cb85779),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72a71b),
	.w1(32'hbbe8f242),
	.w2(32'h3bcb59d5),
	.w3(32'hbc11188a),
	.w4(32'h3a5fc587),
	.w5(32'hba81f9e5),
	.w6(32'hbc9038ef),
	.w7(32'hbb85c1ab),
	.w8(32'hbc0ecb34),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb998533),
	.w1(32'h3b8d4501),
	.w2(32'hbc6bf56d),
	.w3(32'h3bcb51c4),
	.w4(32'h3b1d6c47),
	.w5(32'hbba14d3e),
	.w6(32'h3b83e7b3),
	.w7(32'h3caecac9),
	.w8(32'hbbc9d413),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d16b3b4),
	.w1(32'hbc5a3d10),
	.w2(32'h39f93af5),
	.w3(32'hbb3e3a88),
	.w4(32'h3b04dab1),
	.w5(32'h3ada82bf),
	.w6(32'hbc7918f5),
	.w7(32'hbbc782b5),
	.w8(32'h3bcaf004),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6eb0e),
	.w1(32'h3c08c92b),
	.w2(32'hbbe76f01),
	.w3(32'h3b58c2b4),
	.w4(32'hbc638551),
	.w5(32'h3b7e3c50),
	.w6(32'h3ad380b6),
	.w7(32'hbadce71f),
	.w8(32'h3cd44dcb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b2086),
	.w1(32'h3c526ff5),
	.w2(32'hbcaf370d),
	.w3(32'h3bf25924),
	.w4(32'hbbd0b472),
	.w5(32'hbcf7e25c),
	.w6(32'hbabe3a53),
	.w7(32'h3c03d644),
	.w8(32'hbd5217bb),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d41e8fd),
	.w1(32'hbcdce2e1),
	.w2(32'h3ae2526b),
	.w3(32'h3c96e509),
	.w4(32'hbb833666),
	.w5(32'h3ab2b48b),
	.w6(32'h3ca81a58),
	.w7(32'hbc130b69),
	.w8(32'hb97288c9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba225d),
	.w1(32'hbbd66061),
	.w2(32'h3bd0972e),
	.w3(32'h3a0bc12b),
	.w4(32'hbc7bb432),
	.w5(32'hbc1cf18c),
	.w6(32'h3b26eace),
	.w7(32'hbd10112d),
	.w8(32'h3be59ca3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fc077),
	.w1(32'hba4e4023),
	.w2(32'h3b29967d),
	.w3(32'hbcd5696a),
	.w4(32'hba6ea482),
	.w5(32'hbbd7f6c7),
	.w6(32'h3c27aa46),
	.w7(32'hbc0b7d5a),
	.w8(32'hbc388b9e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a940cd5),
	.w1(32'h3adf9603),
	.w2(32'h3c02be0c),
	.w3(32'hbb621eca),
	.w4(32'hbabf121e),
	.w5(32'h3ad5c47d),
	.w6(32'hbbe12736),
	.w7(32'hbc10a016),
	.w8(32'hbc8fda22),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ea260),
	.w1(32'h399544b3),
	.w2(32'h3badc9db),
	.w3(32'h3b62cf3e),
	.w4(32'hbaae71a6),
	.w5(32'hbb3c75a0),
	.w6(32'hbb8bc9c9),
	.w7(32'h3c01517d),
	.w8(32'hbc974c5d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77edd6),
	.w1(32'hbc655e86),
	.w2(32'hbb29845f),
	.w3(32'hbb76e5f3),
	.w4(32'hbb96f9ac),
	.w5(32'hbc3fa4d7),
	.w6(32'hbbf0314d),
	.w7(32'hbcd8168a),
	.w8(32'h3b61b536),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba43d25f),
	.w1(32'hbbb6e8de),
	.w2(32'h39423b4f),
	.w3(32'hbcbcabdd),
	.w4(32'hbbdb2f3d),
	.w5(32'h3c4e71e8),
	.w6(32'hbc85e594),
	.w7(32'h3c9bac83),
	.w8(32'hbd4b5ebc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8495b),
	.w1(32'hbbfc1e67),
	.w2(32'hbb0f883e),
	.w3(32'h3abeec8b),
	.w4(32'h3a4d7254),
	.w5(32'hbab32b19),
	.w6(32'h3d0e51e0),
	.w7(32'hbbdc68dc),
	.w8(32'hb9909117),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7ab3d),
	.w1(32'hbca1262a),
	.w2(32'hbbfe399a),
	.w3(32'hbbfece2c),
	.w4(32'hbc89528f),
	.w5(32'h3c489a07),
	.w6(32'hbc178cd8),
	.w7(32'h3c516773),
	.w8(32'hbd0303d5),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c20f1),
	.w1(32'hbc293ff1),
	.w2(32'h3c218396),
	.w3(32'h3c141e53),
	.w4(32'hbb916a6d),
	.w5(32'h3aa0531f),
	.w6(32'h3c8595a0),
	.w7(32'h3c9c9717),
	.w8(32'hbc8e6049),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fb951),
	.w1(32'hbb243b06),
	.w2(32'hbc1c7325),
	.w3(32'h3bcf7966),
	.w4(32'h3b8dc5cc),
	.w5(32'h3bcd2ee3),
	.w6(32'h3ca66243),
	.w7(32'hba94956b),
	.w8(32'hbc633fd1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf90622),
	.w1(32'h3a22c2b0),
	.w2(32'h3c4e0ec5),
	.w3(32'h3b03025a),
	.w4(32'h3c3dbe0c),
	.w5(32'h3ae5c36d),
	.w6(32'hbc0897bb),
	.w7(32'h3b804b4d),
	.w8(32'hbb69c437),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9d40),
	.w1(32'hba88cd8f),
	.w2(32'h3c4ab26c),
	.w3(32'hba26b5c6),
	.w4(32'hbc98bc92),
	.w5(32'h3cb3e4ec),
	.w6(32'h39c52330),
	.w7(32'hbc45ecf4),
	.w8(32'h39794c01),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd704cf6),
	.w1(32'h3cb528cd),
	.w2(32'hbb319e1e),
	.w3(32'hbc20fddb),
	.w4(32'hbbf5590d),
	.w5(32'hbc9b1d3b),
	.w6(32'hbc3c073e),
	.w7(32'hbc7db77d),
	.w8(32'h3bf140ae),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fcaec),
	.w1(32'hbb0e8913),
	.w2(32'hbb60c342),
	.w3(32'hbcb5464b),
	.w4(32'hbbb96648),
	.w5(32'hbc347d58),
	.w6(32'hbc76f8c8),
	.w7(32'hbc0bc550),
	.w8(32'hbc91f0c1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16cc73),
	.w1(32'hbb752967),
	.w2(32'h39d1e3bc),
	.w3(32'h3a9f8168),
	.w4(32'h3a9b2b2d),
	.w5(32'h3a0c6451),
	.w6(32'hbbd0f822),
	.w7(32'h3aa30bda),
	.w8(32'hb96f6821),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e46ee),
	.w1(32'hb9e1b986),
	.w2(32'hbb8a7b3b),
	.w3(32'h3b2076f4),
	.w4(32'hbb6bdb28),
	.w5(32'hbba3f219),
	.w6(32'h3b34091b),
	.w7(32'hbad5bf0e),
	.w8(32'hbb927355),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3db815),
	.w1(32'h380768b8),
	.w2(32'hbb2cf3d0),
	.w3(32'h3a1608d2),
	.w4(32'hbb8d7a14),
	.w5(32'hbb2aaca2),
	.w6(32'hbaa91071),
	.w7(32'hbb5e2e1a),
	.w8(32'hbb74dd7b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97feb4),
	.w1(32'hbb5d6d60),
	.w2(32'hbb814a15),
	.w3(32'hbb6d54f4),
	.w4(32'hbac93e8d),
	.w5(32'hba283e5f),
	.w6(32'hbb4bce32),
	.w7(32'hbabfc3b9),
	.w8(32'hbb0eaebb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add441b),
	.w1(32'h3b23aa57),
	.w2(32'hbbdb3a4d),
	.w3(32'h3ba43d23),
	.w4(32'hbbac3b80),
	.w5(32'hbc0a508f),
	.w6(32'h3bd16705),
	.w7(32'hbc0218e5),
	.w8(32'hbc278398),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda1b0c),
	.w1(32'hbbd30576),
	.w2(32'hbb92d0bb),
	.w3(32'hbbe32dc9),
	.w4(32'h3b3d6a21),
	.w5(32'h3c43d924),
	.w6(32'hbbcbfb32),
	.w7(32'h3b6363db),
	.w8(32'h3c6a636d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21a31e),
	.w1(32'h3c44f753),
	.w2(32'h3a0aeecb),
	.w3(32'h3c0911b1),
	.w4(32'h3a231fab),
	.w5(32'h3be29dbc),
	.w6(32'h3c9f3383),
	.w7(32'h3bc98e71),
	.w8(32'h3a2a8f45),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef3230),
	.w1(32'h3b999b14),
	.w2(32'hbaa424e6),
	.w3(32'h3c652730),
	.w4(32'h3c106fa9),
	.w5(32'hb96b3600),
	.w6(32'h3c31aaaa),
	.w7(32'h3c1f6dca),
	.w8(32'h3c16522f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0774b),
	.w1(32'hbb63d124),
	.w2(32'hbbd431d7),
	.w3(32'hba9e861b),
	.w4(32'hbaae970d),
	.w5(32'hbc2d92fa),
	.w6(32'h3b609cb5),
	.w7(32'hbc331779),
	.w8(32'hbc89a11c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f4b25),
	.w1(32'h3add0d76),
	.w2(32'hb9fa70e7),
	.w3(32'h3bd2d26e),
	.w4(32'hbb33f6ff),
	.w5(32'hbb7aff03),
	.w6(32'hba8ef19a),
	.w7(32'hb9d62166),
	.w8(32'h3bcb8969),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14c1e1),
	.w1(32'h3b95221b),
	.w2(32'h3aaf6349),
	.w3(32'hb95263be),
	.w4(32'hbbb5232f),
	.w5(32'hbb06605c),
	.w6(32'h39257342),
	.w7(32'h3a66f4a7),
	.w8(32'h3aab0e91),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c677b),
	.w1(32'hbbb639a4),
	.w2(32'h3b754c78),
	.w3(32'hbb89967e),
	.w4(32'h3b9a4775),
	.w5(32'h3b50a315),
	.w6(32'hbb21b106),
	.w7(32'h3b89d8ee),
	.w8(32'h3b5e1108),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9cb6),
	.w1(32'h3b741aac),
	.w2(32'hbb1a9efb),
	.w3(32'h3ad51d7e),
	.w4(32'hb9936414),
	.w5(32'h3a5b9257),
	.w6(32'h3b1feb9b),
	.w7(32'hbb078e52),
	.w8(32'h3a74f5a7),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990f810),
	.w1(32'hb8c55ae0),
	.w2(32'h3aaf642d),
	.w3(32'h3b43797d),
	.w4(32'h3ac95764),
	.w5(32'hbb7e361f),
	.w6(32'h3a894b10),
	.w7(32'h3bc36402),
	.w8(32'h3b7b3a58),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd43443),
	.w1(32'h3b4b70f4),
	.w2(32'h3a4d5ca5),
	.w3(32'hbaf413ca),
	.w4(32'h3b476425),
	.w5(32'hbacd9309),
	.w6(32'h3a1d3f38),
	.w7(32'hbb0e7499),
	.w8(32'hbbc32dbe),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81b6e),
	.w1(32'hbab4da2d),
	.w2(32'hbb05224b),
	.w3(32'h3ae88e1b),
	.w4(32'hb9cab6c2),
	.w5(32'hbbd5eee3),
	.w6(32'hbbdbf767),
	.w7(32'hbbf7f8ad),
	.w8(32'hbc976c54),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d6b21),
	.w1(32'hbc4da3cc),
	.w2(32'hba5bf637),
	.w3(32'hbc0a01f7),
	.w4(32'h3b536fb2),
	.w5(32'hba9b7628),
	.w6(32'hbc42bf7d),
	.w7(32'h3bb4b648),
	.w8(32'hb9fbbcb6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b2b21),
	.w1(32'h3bb63c29),
	.w2(32'h3ae8ec17),
	.w3(32'h3acac173),
	.w4(32'h3a8d2609),
	.w5(32'hbace3164),
	.w6(32'h3c3c99ec),
	.w7(32'h3c069e6f),
	.w8(32'h3bfc37e3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac834b),
	.w1(32'hbb25fa15),
	.w2(32'h3ba8ef9d),
	.w3(32'h3b10aa05),
	.w4(32'h3b39d477),
	.w5(32'h3ba808ba),
	.w6(32'h3b39d63a),
	.w7(32'h3c1fa61b),
	.w8(32'h3c27d507),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd3cf0),
	.w1(32'hba36e448),
	.w2(32'hbb08d635),
	.w3(32'hbb24f7cf),
	.w4(32'hbc0569bd),
	.w5(32'hbc09e9c1),
	.w6(32'hb9a027fe),
	.w7(32'hbb7a6d67),
	.w8(32'hbc08271e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a1b8d1),
	.w1(32'h3b9159b1),
	.w2(32'hbc009430),
	.w3(32'hbb6dfa12),
	.w4(32'hbc39b670),
	.w5(32'hbc108b90),
	.w6(32'h3abd7ed7),
	.w7(32'hbc06f365),
	.w8(32'hbb73fb5f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820192),
	.w1(32'h3b5add43),
	.w2(32'hbbe50f63),
	.w3(32'hbb647d38),
	.w4(32'hbb599159),
	.w5(32'hbb887284),
	.w6(32'hbad7e57f),
	.w7(32'hbbb9c764),
	.w8(32'hbb0d983c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc4893),
	.w1(32'hbbeeaabb),
	.w2(32'h3b0c6de1),
	.w3(32'hbb85b935),
	.w4(32'h3b9d17b8),
	.w5(32'h3bae53c4),
	.w6(32'hbbaf8482),
	.w7(32'h3b2b03dc),
	.w8(32'h3b8e571f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69149f),
	.w1(32'h3ba1579f),
	.w2(32'hbb82c3c7),
	.w3(32'h3bca4d20),
	.w4(32'hbb38ce11),
	.w5(32'hba9334b2),
	.w6(32'h3b89d417),
	.w7(32'hba5ab43d),
	.w8(32'h3b6f0e9b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa34546),
	.w1(32'h3a08b908),
	.w2(32'hbc0b325f),
	.w3(32'hba0d5f2d),
	.w4(32'hbc4fd996),
	.w5(32'hbc30d5e6),
	.w6(32'h3b8df864),
	.w7(32'hbc67fd4a),
	.w8(32'hbc1e0ea0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc637a0d),
	.w1(32'hbc886195),
	.w2(32'hbb57ae05),
	.w3(32'hbbf14b93),
	.w4(32'hbbe540c9),
	.w5(32'hbc032dd3),
	.w6(32'hbb9c70ea),
	.w7(32'h3afb424a),
	.w8(32'hb894e108),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31dd08),
	.w1(32'hbaf8f4a3),
	.w2(32'hbb831a22),
	.w3(32'hbb411059),
	.w4(32'hbba26544),
	.w5(32'hbae54832),
	.w6(32'hbc629401),
	.w7(32'hbc132fa1),
	.w8(32'h3ad33c2c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1454),
	.w1(32'h3bf8aa64),
	.w2(32'h39de277b),
	.w3(32'hb952f2d5),
	.w4(32'hbbd24a45),
	.w5(32'hbb9ca62e),
	.w6(32'h3c1b4465),
	.w7(32'h3b4d05c5),
	.w8(32'h3b40ef1e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad64c04),
	.w1(32'h3ae78631),
	.w2(32'h3b74c2f1),
	.w3(32'h3b120af3),
	.w4(32'h3a7bf281),
	.w5(32'h3b6b17f6),
	.w6(32'h3bed633b),
	.w7(32'h3c30fee5),
	.w8(32'h3bc00b2f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01bd5),
	.w1(32'h3a127239),
	.w2(32'hbb98ceab),
	.w3(32'hbaf55370),
	.w4(32'hbbabef07),
	.w5(32'hbc252881),
	.w6(32'hbb5f4f9e),
	.w7(32'hbc06847e),
	.w8(32'hbb9e0b9b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2eaa5),
	.w1(32'h395dac0e),
	.w2(32'h3b4c7a02),
	.w3(32'h3b031862),
	.w4(32'h3a03f933),
	.w5(32'h3b1947b3),
	.w6(32'h3b8fff18),
	.w7(32'h384a4f51),
	.w8(32'hbb7917e0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc875eda),
	.w1(32'hbc199463),
	.w2(32'hbb896691),
	.w3(32'hb92ab0dc),
	.w4(32'hbad040dd),
	.w5(32'hbb21d150),
	.w6(32'hbb9e2177),
	.w7(32'h3b1e716f),
	.w8(32'h3a95809c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3b3e),
	.w1(32'h3c1483c7),
	.w2(32'h3c0a4030),
	.w3(32'h3c15acd1),
	.w4(32'h3c22621e),
	.w5(32'h3b2bcbc7),
	.w6(32'h3c24edd2),
	.w7(32'h3c1beb89),
	.w8(32'h3ba66791),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba981b6),
	.w1(32'h3b693bdd),
	.w2(32'hbaaa1368),
	.w3(32'hbc12bd87),
	.w4(32'h3ba5fb47),
	.w5(32'h39e531dc),
	.w6(32'hbb178201),
	.w7(32'h3bdfd8f3),
	.w8(32'h3b8b3f8d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d5967),
	.w1(32'hbae7bea5),
	.w2(32'hbbfdc062),
	.w3(32'hba40029d),
	.w4(32'hbb3a0fbf),
	.w5(32'hbb887574),
	.w6(32'hbba234ee),
	.w7(32'hb959284d),
	.w8(32'h3b5e8b39),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd3e9),
	.w1(32'h3a504ca7),
	.w2(32'hbc201b16),
	.w3(32'hba4585b0),
	.w4(32'h3ab13ddc),
	.w5(32'hbc0cf0b0),
	.w6(32'h38b81500),
	.w7(32'h3ac89d86),
	.w8(32'hba8a43d5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e65c),
	.w1(32'h3b2894d6),
	.w2(32'h3b424ea3),
	.w3(32'hbb46ae69),
	.w4(32'h3ba7a0ee),
	.w5(32'h3babb65d),
	.w6(32'hbbb17b86),
	.w7(32'h39a9055d),
	.w8(32'h3b70b075),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad7147),
	.w1(32'h3beb46bd),
	.w2(32'hbc0d8ca3),
	.w3(32'h3bbb3e69),
	.w4(32'hbc7db261),
	.w5(32'hbb93ae96),
	.w6(32'h3c063bec),
	.w7(32'hbc165e06),
	.w8(32'h3acc1fb6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d3466),
	.w1(32'hbac41593),
	.w2(32'h3b5d4cd7),
	.w3(32'hbbdd84a3),
	.w4(32'h3b8edac3),
	.w5(32'h396ad2f2),
	.w6(32'h3b8ec4c9),
	.w7(32'h3c25e8d6),
	.w8(32'h3c37697b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b4141),
	.w1(32'h3bc57573),
	.w2(32'hbafd7ad5),
	.w3(32'hbb7633b4),
	.w4(32'h3b18a782),
	.w5(32'hba826579),
	.w6(32'h3a9cc6d7),
	.w7(32'h3aef83aa),
	.w8(32'h3bb2142e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f8860),
	.w1(32'h39ad170b),
	.w2(32'hbb766273),
	.w3(32'hbaa1c321),
	.w4(32'hb99d893f),
	.w5(32'hbbc8819a),
	.w6(32'hb8d19477),
	.w7(32'h3b2196e3),
	.w8(32'hbb7c23b0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb655c78),
	.w1(32'h3b970cd0),
	.w2(32'hbaae6a27),
	.w3(32'hbadcbcde),
	.w4(32'hba4febd2),
	.w5(32'hbaa2eeee),
	.w6(32'h3b083eb9),
	.w7(32'h3a054391),
	.w8(32'hb9e285c1),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcb25d),
	.w1(32'h3af932ad),
	.w2(32'h3bc28edd),
	.w3(32'h3aaa729d),
	.w4(32'h3b7c4b8d),
	.w5(32'h3b0276d8),
	.w6(32'h3b143e80),
	.w7(32'h3c0e5ee2),
	.w8(32'h3b05ae99),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b927820),
	.w1(32'h3b2aa8a3),
	.w2(32'h3b8b1cab),
	.w3(32'h3c3d5fe6),
	.w4(32'h3a967d13),
	.w5(32'h3bacad60),
	.w6(32'h3b876be1),
	.w7(32'h3b787ac4),
	.w8(32'hbadee075),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24f063),
	.w1(32'h3b793a02),
	.w2(32'hbafb831c),
	.w3(32'h3b813a24),
	.w4(32'hbb610c21),
	.w5(32'hbbb0e61c),
	.w6(32'h3b72dc55),
	.w7(32'hbba703d4),
	.w8(32'hbbb41d1f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3899),
	.w1(32'h3b880bbf),
	.w2(32'hbacab7ca),
	.w3(32'h38a52cab),
	.w4(32'h3bba4356),
	.w5(32'h3ae5be00),
	.w6(32'h3b2a2301),
	.w7(32'h3b637783),
	.w8(32'hba2c2fe0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba613ea),
	.w1(32'hbac20770),
	.w2(32'h3b0b942f),
	.w3(32'h3a845a87),
	.w4(32'h3a717bed),
	.w5(32'h3a877096),
	.w6(32'hbb2abb63),
	.w7(32'h3abba6ce),
	.w8(32'h3ab9eb7c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6edad3),
	.w1(32'h3bc95ab9),
	.w2(32'h3b209eda),
	.w3(32'h3b122846),
	.w4(32'h3c3fb7a5),
	.w5(32'h3be70ae0),
	.w6(32'h3b61488a),
	.w7(32'h3a8fc139),
	.w8(32'hbad932a6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6cfcf),
	.w1(32'hbb9d5348),
	.w2(32'h3aad75ff),
	.w3(32'h3b3a9d67),
	.w4(32'h399ac35a),
	.w5(32'hbb1424fd),
	.w6(32'h3bd478c1),
	.w7(32'h3b0082e5),
	.w8(32'h3c17de9e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8aa48),
	.w1(32'h3b660bd1),
	.w2(32'hbbab8951),
	.w3(32'hbae207e8),
	.w4(32'hbb5d8741),
	.w5(32'hbaaf94fd),
	.w6(32'h3ae97dab),
	.w7(32'hbbad3c24),
	.w8(32'hbba1c191),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d2622),
	.w1(32'hbbc71e43),
	.w2(32'h3bfff0da),
	.w3(32'hb8f47059),
	.w4(32'h395d6a70),
	.w5(32'h3bc95c4a),
	.w6(32'hbbe8fac9),
	.w7(32'h3bd0b64d),
	.w8(32'hbaac9532),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9edc),
	.w1(32'h3a4a9023),
	.w2(32'h3b93ed1a),
	.w3(32'h3bc95a79),
	.w4(32'h3af5a64e),
	.w5(32'hbaf0ac63),
	.w6(32'h3b917255),
	.w7(32'h3b9deedf),
	.w8(32'h3a80190b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule