module layer_8_featuremap_115(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f995e),
	.w1(32'hbb27bd46),
	.w2(32'hbbf12162),
	.w3(32'hbac890c4),
	.w4(32'hbb755c50),
	.w5(32'hbbcf4156),
	.w6(32'hbb7f4070),
	.w7(32'hbb8c6b7c),
	.w8(32'hbc24b486),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc234ab7),
	.w1(32'hbb555cdf),
	.w2(32'h3b681da6),
	.w3(32'hbb04bac2),
	.w4(32'h3bc99aba),
	.w5(32'h3c979b64),
	.w6(32'hbb76c088),
	.w7(32'h3ba1a2a0),
	.w8(32'h3c707b28),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67a435),
	.w1(32'h3c040a41),
	.w2(32'hbbce5108),
	.w3(32'h3c915a3d),
	.w4(32'hbbcab269),
	.w5(32'h3aa750f1),
	.w6(32'h3c7a7fd3),
	.w7(32'hbbb1925b),
	.w8(32'hbb01058b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8ed4f),
	.w1(32'h3b70a697),
	.w2(32'h3be73fba),
	.w3(32'hbaafb772),
	.w4(32'hbbbb98b1),
	.w5(32'hbc60e0d0),
	.w6(32'h3b72cb9c),
	.w7(32'hbc28ce78),
	.w8(32'hbc8e84c1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf80304),
	.w1(32'hbc70ccff),
	.w2(32'h3b273d8f),
	.w3(32'hbb1e348d),
	.w4(32'h3b2ecb37),
	.w5(32'h3b53c875),
	.w6(32'hbc288145),
	.w7(32'hbb1b8c9c),
	.w8(32'hba8c3308),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baa75e),
	.w1(32'hbb7c7fbe),
	.w2(32'h3b3f651a),
	.w3(32'h3b9498f9),
	.w4(32'h3ba19282),
	.w5(32'hbbd63b1d),
	.w6(32'h3a826ed2),
	.w7(32'h3b25d25d),
	.w8(32'hbc1f04d7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb040cdc),
	.w1(32'hbc8d3702),
	.w2(32'hba37ccb1),
	.w3(32'hbc0dd9b9),
	.w4(32'hbb530823),
	.w5(32'hbbe017fa),
	.w6(32'hbc1e6e73),
	.w7(32'hbba29faa),
	.w8(32'hbc0cee5b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38224c),
	.w1(32'hbc26e38a),
	.w2(32'hbad41278),
	.w3(32'h3bbe9acb),
	.w4(32'hbb831db3),
	.w5(32'h3a433aa7),
	.w6(32'hbbc30ff0),
	.w7(32'h3acdb200),
	.w8(32'h3b003711),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906a7ef),
	.w1(32'hbbff70ce),
	.w2(32'h3a112a6a),
	.w3(32'hbbb1408d),
	.w4(32'hbb47a3f4),
	.w5(32'hbbd42526),
	.w6(32'hbc0d9819),
	.w7(32'hbb8452a1),
	.w8(32'hbb8b020a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9d45c),
	.w1(32'hbbfa35ed),
	.w2(32'h39912e58),
	.w3(32'h3ae83137),
	.w4(32'h3b75bfd1),
	.w5(32'hb9b65a62),
	.w6(32'hbb538ab3),
	.w7(32'hbb029acb),
	.w8(32'hbba2c168),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac4a6),
	.w1(32'hbb11dff2),
	.w2(32'h3c079544),
	.w3(32'h3c40c57a),
	.w4(32'h3b303bbd),
	.w5(32'h3b42b299),
	.w6(32'h3c2ab98e),
	.w7(32'h3c16c299),
	.w8(32'h3c7102b0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37c6c3),
	.w1(32'h3abddb69),
	.w2(32'hbbb019be),
	.w3(32'hbb5000a6),
	.w4(32'h39cd9f4c),
	.w5(32'hbc1f0c2e),
	.w6(32'hbb21bc14),
	.w7(32'hbbc5612e),
	.w8(32'hbbd339b3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee6348),
	.w1(32'hbb9db64a),
	.w2(32'hbab488b6),
	.w3(32'hbbe22549),
	.w4(32'hb8585217),
	.w5(32'hbad45254),
	.w6(32'hbbee66ef),
	.w7(32'hba815620),
	.w8(32'hb9c3a3fa),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba972016),
	.w1(32'hba765097),
	.w2(32'hbb558c75),
	.w3(32'hba693ef6),
	.w4(32'hbb8aa02e),
	.w5(32'hbad75276),
	.w6(32'hba3d807c),
	.w7(32'hbb6147a2),
	.w8(32'hbacec311),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3701b9),
	.w1(32'hbb835a61),
	.w2(32'h3aaa86f2),
	.w3(32'hbb4c4c21),
	.w4(32'hba584c83),
	.w5(32'hba7e5c7e),
	.w6(32'hbae12ecd),
	.w7(32'hb8b2546c),
	.w8(32'hb920065a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9540c75),
	.w1(32'hbb547670),
	.w2(32'h3b89b90f),
	.w3(32'hbad73f59),
	.w4(32'hba225896),
	.w5(32'h3b3e96c8),
	.w6(32'hbaa73735),
	.w7(32'h3a089809),
	.w8(32'h3a6f65a8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95dd5e),
	.w1(32'hbb80a6c1),
	.w2(32'h3b78f055),
	.w3(32'h3b9c853f),
	.w4(32'h3bd6540f),
	.w5(32'h3cca2186),
	.w6(32'hb96d3836),
	.w7(32'h3b4c33e7),
	.w8(32'h3c7bbdc4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcab580),
	.w1(32'h3b105784),
	.w2(32'h3b6363e0),
	.w3(32'h3c0c41d8),
	.w4(32'hbb5eacec),
	.w5(32'hbbf9f527),
	.w6(32'h3b7856ae),
	.w7(32'h3aa5f948),
	.w8(32'hb9e5a9ed),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7592f3),
	.w1(32'hbbb06410),
	.w2(32'hba9c9c57),
	.w3(32'hbb9aa1ac),
	.w4(32'hbb14d058),
	.w5(32'h3b3746bd),
	.w6(32'hbbd0320f),
	.w7(32'hbb230b49),
	.w8(32'h3bd5621b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c313c48),
	.w1(32'h3a9b74a6),
	.w2(32'h3b7e2c70),
	.w3(32'hbbf03515),
	.w4(32'h3b8236ad),
	.w5(32'h3b100273),
	.w6(32'hbc144fa6),
	.w7(32'h3baeab2d),
	.w8(32'h3b84a707),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6ff8),
	.w1(32'hbb416e88),
	.w2(32'hbbbe0b54),
	.w3(32'hbba32e4b),
	.w4(32'hbc06c758),
	.w5(32'hbc0f3675),
	.w6(32'h3b50850f),
	.w7(32'hbc24f061),
	.w8(32'hbc14b80b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1da2a5),
	.w1(32'hbb406d82),
	.w2(32'hbb5e4cbd),
	.w3(32'hbaa5ce79),
	.w4(32'hbbbba1de),
	.w5(32'hbb9aeb1f),
	.w6(32'h3b9ad272),
	.w7(32'hbc04b38f),
	.w8(32'hbb22cd2e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0cd7d),
	.w1(32'hbbc6642c),
	.w2(32'h39e1dc80),
	.w3(32'hbc4397d9),
	.w4(32'hbbfbe917),
	.w5(32'hbc418f2d),
	.w6(32'hbc2d11c7),
	.w7(32'hbb94a5a4),
	.w8(32'hbc1243dc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e292),
	.w1(32'hbb2ec22a),
	.w2(32'h3c7dd411),
	.w3(32'hbbab31b9),
	.w4(32'h3bf4c970),
	.w5(32'h3c43c5fd),
	.w6(32'hbbc1d6a4),
	.w7(32'h3c6b372f),
	.w8(32'h3cb28ed2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd35155),
	.w1(32'hbc0b66bf),
	.w2(32'hbb780ab7),
	.w3(32'hbadedb03),
	.w4(32'hbbf0d320),
	.w5(32'hbbfd8c89),
	.w6(32'hbbaba5c4),
	.w7(32'hb9c328e2),
	.w8(32'hba732ca6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06f7d6),
	.w1(32'hb9fef5d6),
	.w2(32'hbb493c61),
	.w3(32'hba3bfdf7),
	.w4(32'hbb0e8860),
	.w5(32'h3bdbea81),
	.w6(32'h3bdd5e89),
	.w7(32'hb986eee4),
	.w8(32'h3ba48fbb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b004110),
	.w1(32'h3b7a8218),
	.w2(32'hbb86d54b),
	.w3(32'hbb3539bc),
	.w4(32'hbbbcbe0a),
	.w5(32'hbb75db33),
	.w6(32'h388a758f),
	.w7(32'hbb40b49d),
	.w8(32'hbb866d71),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed8d3),
	.w1(32'hbb48317b),
	.w2(32'hbaf22366),
	.w3(32'hbbaddc4b),
	.w4(32'hbb937289),
	.w5(32'h3acad166),
	.w6(32'hbbe0f8fd),
	.w7(32'hbc32879d),
	.w8(32'hbbba1a1f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4965fc),
	.w1(32'hb3be8dbb),
	.w2(32'h3b8ecc4c),
	.w3(32'hbc3dc602),
	.w4(32'h3b1e331f),
	.w5(32'hbc1895e6),
	.w6(32'hbb97d45a),
	.w7(32'h3b06b023),
	.w8(32'h3ba5f818),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a8b5e),
	.w1(32'h3c33de43),
	.w2(32'hbbd39b6d),
	.w3(32'hbc0a432e),
	.w4(32'h3acf8ff5),
	.w5(32'h3af2a12f),
	.w6(32'h3c6958fe),
	.w7(32'hbab0a6ac),
	.w8(32'hba1a14a1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb24d31),
	.w1(32'hba955916),
	.w2(32'hb7807708),
	.w3(32'h3bc94b98),
	.w4(32'hb98b52eb),
	.w5(32'hbb96486f),
	.w6(32'h3bcd2321),
	.w7(32'hb98069a8),
	.w8(32'hbb9c5c83),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5dc2),
	.w1(32'hbb0423a5),
	.w2(32'h3bd1fe8f),
	.w3(32'hbb2b9e47),
	.w4(32'hbb12c42c),
	.w5(32'hbb816620),
	.w6(32'hbb18806c),
	.w7(32'hb99d62cf),
	.w8(32'hbbb4eeab),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b672257),
	.w1(32'hbb3aeb3e),
	.w2(32'hbb4abd40),
	.w3(32'hbb399fb2),
	.w4(32'h3ac93a47),
	.w5(32'hbbf55971),
	.w6(32'h3a5805c1),
	.w7(32'hbb4e8fd5),
	.w8(32'hbb3d9256),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8cc67),
	.w1(32'hbb4d61b0),
	.w2(32'hbb86959f),
	.w3(32'hbbecbaff),
	.w4(32'h3b826612),
	.w5(32'h3bfe54aa),
	.w6(32'hbc50c209),
	.w7(32'hbaab960b),
	.w8(32'hbaa69db5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28bfff),
	.w1(32'h3a582d79),
	.w2(32'hbaf6ac96),
	.w3(32'h3c8b5035),
	.w4(32'hb93dfbbe),
	.w5(32'h3bc70321),
	.w6(32'h3b676555),
	.w7(32'hbb88cf2d),
	.w8(32'h3aff4c4a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02b2ff),
	.w1(32'h3a6ccdb0),
	.w2(32'hbbea5c6d),
	.w3(32'h3a5c8379),
	.w4(32'hbc0a423a),
	.w5(32'hbc07ff8b),
	.w6(32'h3a94ca16),
	.w7(32'hbc25755d),
	.w8(32'hbb6a5a48),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ed8f1),
	.w1(32'h3bb36c6d),
	.w2(32'hbb2a27a7),
	.w3(32'hbc0d1a31),
	.w4(32'hbb986e70),
	.w5(32'hbc3b0e00),
	.w6(32'hbb4c5964),
	.w7(32'h3c00244c),
	.w8(32'h3c6cdcb3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3538d2),
	.w1(32'h3c5f18cd),
	.w2(32'h3b449b4b),
	.w3(32'hbc2a2d1f),
	.w4(32'h3b94f2e6),
	.w5(32'hbc370595),
	.w6(32'h3bcaef9c),
	.w7(32'h3b3d80a6),
	.w8(32'hbc1a908f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc293b43),
	.w1(32'h39479342),
	.w2(32'h3c099185),
	.w3(32'hbb83ea1d),
	.w4(32'h3bafda4b),
	.w5(32'h3bf8f0e3),
	.w6(32'hbb90b108),
	.w7(32'h3b9cedca),
	.w8(32'h3b80c0ac),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa182a),
	.w1(32'h3c2ad837),
	.w2(32'hba6ad5a3),
	.w3(32'h3b8bfa70),
	.w4(32'hbb619768),
	.w5(32'hbae72cd7),
	.w6(32'h3befc7b5),
	.w7(32'hbba1f1b7),
	.w8(32'hbbfd83d5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7001),
	.w1(32'hbb19f10f),
	.w2(32'hba08b0c7),
	.w3(32'h3b7efceb),
	.w4(32'h3b5af32e),
	.w5(32'h3b172bfd),
	.w6(32'hbbb9d51d),
	.w7(32'hb981f2bf),
	.w8(32'h3adcdf82),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbea6e2),
	.w1(32'h39a44442),
	.w2(32'h3b47d2da),
	.w3(32'hbae111d1),
	.w4(32'hbb756597),
	.w5(32'hbb122721),
	.w6(32'hbc1e01c5),
	.w7(32'hbb1f8e7b),
	.w8(32'hbb952574),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20368),
	.w1(32'h3bbba91c),
	.w2(32'hbc27bb00),
	.w3(32'h3c4042ac),
	.w4(32'h3a11e835),
	.w5(32'hbb9ce07d),
	.w6(32'h3b004bb5),
	.w7(32'hbc1028a6),
	.w8(32'hbb5b79e3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e3052),
	.w1(32'h3b6b6835),
	.w2(32'hbadc0a6b),
	.w3(32'hbbb5926d),
	.w4(32'h3987dff5),
	.w5(32'h393e8b84),
	.w6(32'hbbb81414),
	.w7(32'hbadee572),
	.w8(32'h3a66dd5b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0c6f5),
	.w1(32'hba166ef0),
	.w2(32'h3a3ae7f3),
	.w3(32'hb9c6f467),
	.w4(32'h3b4bf938),
	.w5(32'h3b99633c),
	.w6(32'h3a25fb83),
	.w7(32'hbaa6db8d),
	.w8(32'hbb2e6ea4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7a6f0),
	.w1(32'hbaa88234),
	.w2(32'h3c5c3e06),
	.w3(32'hbaffd749),
	.w4(32'h38828d92),
	.w5(32'hbb507c24),
	.w6(32'hbb48b361),
	.w7(32'h3bff4bd0),
	.w8(32'h3a98db01),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814fdc),
	.w1(32'h3c3baf9b),
	.w2(32'h3a5a50c3),
	.w3(32'h3c1235c6),
	.w4(32'hba221ed7),
	.w5(32'hbaa80656),
	.w6(32'h3c2bc72c),
	.w7(32'hbb73fcd0),
	.w8(32'hba3b9da5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e265e),
	.w1(32'h3b01bf96),
	.w2(32'h3bd46746),
	.w3(32'hbbc463fa),
	.w4(32'h3b549c72),
	.w5(32'hba0c7512),
	.w6(32'h3b95ae95),
	.w7(32'hbb1ff9f1),
	.w8(32'hba8405d9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37eebe),
	.w1(32'h3b8a9342),
	.w2(32'h3bfb9fde),
	.w3(32'hba21a57f),
	.w4(32'h3b075273),
	.w5(32'h3b5c586c),
	.w6(32'hbad4afba),
	.w7(32'h3abdab2a),
	.w8(32'hb97690a9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5367b),
	.w1(32'hbb77d065),
	.w2(32'h3c142b11),
	.w3(32'h3ab8e033),
	.w4(32'hb8d09542),
	.w5(32'h3b4b806b),
	.w6(32'hba225abe),
	.w7(32'h3bc1dc4f),
	.w8(32'h3c06f57d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5a4d9),
	.w1(32'hb9edc194),
	.w2(32'h3c36a995),
	.w3(32'hbb1dbbee),
	.w4(32'h3c2aec05),
	.w5(32'h3c094259),
	.w6(32'h3b58884d),
	.w7(32'h3c0e86a1),
	.w8(32'h3ae6b4ea),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c225a24),
	.w1(32'hbb10cd45),
	.w2(32'h3bbaa970),
	.w3(32'h3c2a237d),
	.w4(32'hbb26e3c1),
	.w5(32'h3b947a47),
	.w6(32'h3b404625),
	.w7(32'hbb477c4b),
	.w8(32'hbb65b463),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc5571),
	.w1(32'h3a46bd61),
	.w2(32'h3b54b666),
	.w3(32'h3c6ba642),
	.w4(32'hbb0d31b3),
	.w5(32'h39a49053),
	.w6(32'h3b8ffcff),
	.w7(32'hb840b2bd),
	.w8(32'hbab674f5),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa9c46),
	.w1(32'hbbc9babf),
	.w2(32'hbb106fac),
	.w3(32'hbbde32b0),
	.w4(32'hba93f512),
	.w5(32'h38e0bdc4),
	.w6(32'hbb4ad4d6),
	.w7(32'hbb2190ce),
	.w8(32'h3a4939dc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0a29c),
	.w1(32'hba4e4173),
	.w2(32'hbba0d2c4),
	.w3(32'hba831d6e),
	.w4(32'hbb49544b),
	.w5(32'hbc0ab839),
	.w6(32'h3a2730e3),
	.w7(32'hba9136a4),
	.w8(32'hbaf066a8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff7aad),
	.w1(32'hbabb62ed),
	.w2(32'h3b933050),
	.w3(32'hbb4cf6b7),
	.w4(32'h38ae0e2a),
	.w5(32'hba5f05be),
	.w6(32'hbadc635c),
	.w7(32'h38c36fbb),
	.w8(32'h3b8739ef),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbbb9b),
	.w1(32'h39af1b67),
	.w2(32'h3a1e5fe7),
	.w3(32'hbc17d543),
	.w4(32'hb9a2c694),
	.w5(32'h3a7e0f82),
	.w6(32'hbb8d32f3),
	.w7(32'hb9ac7153),
	.w8(32'hbadd2c70),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae00758),
	.w1(32'hba95b1fa),
	.w2(32'hbb2a1184),
	.w3(32'h3b050506),
	.w4(32'h3c4258db),
	.w5(32'h3b69cc01),
	.w6(32'hbab6cd45),
	.w7(32'h3bbb0767),
	.w8(32'h3b355d17),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02e22f),
	.w1(32'h3c0837e0),
	.w2(32'hbb096e3d),
	.w3(32'hbb1ada8e),
	.w4(32'h392a41e9),
	.w5(32'h38884964),
	.w6(32'h3b17e4cf),
	.w7(32'hbb093355),
	.w8(32'h3a18bad6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d24ea),
	.w1(32'hb9f5e2f5),
	.w2(32'h3c0c193e),
	.w3(32'hb9815ea2),
	.w4(32'h3bc2d766),
	.w5(32'h3b4c38ca),
	.w6(32'h3a0bf50e),
	.w7(32'h3aec0ef0),
	.w8(32'h3b879fa1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3c599),
	.w1(32'hbac6b05b),
	.w2(32'hb8add9e7),
	.w3(32'hbc0c985f),
	.w4(32'hbbc1063c),
	.w5(32'hbc11456a),
	.w6(32'hbb1ad2d7),
	.w7(32'hbb75ad07),
	.w8(32'hbc025bd2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae32476),
	.w1(32'hbbf37538),
	.w2(32'h3c12c3d7),
	.w3(32'hbbf8367d),
	.w4(32'h3c85f923),
	.w5(32'h3c8383fb),
	.w6(32'hbc88a833),
	.w7(32'h3ca9c64d),
	.w8(32'h3ccc24cd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4181),
	.w1(32'h3c3021e5),
	.w2(32'hbbd9ef8b),
	.w3(32'h3bfd97bb),
	.w4(32'hbb80b9e2),
	.w5(32'hbc0911db),
	.w6(32'h3cb71ff2),
	.w7(32'hbb85b3c0),
	.w8(32'hbb09c77b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937c241),
	.w1(32'hbc11618a),
	.w2(32'h3ae89da1),
	.w3(32'hbc8387d2),
	.w4(32'hba92c2ef),
	.w5(32'hbbbce3b1),
	.w6(32'hbc89138c),
	.w7(32'h3a0ce654),
	.w8(32'hba22851d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b82f3),
	.w1(32'h3b68cc7b),
	.w2(32'h39decd8b),
	.w3(32'hbbf23750),
	.w4(32'h3a302b5e),
	.w5(32'hbb344a62),
	.w6(32'h3b39bb18),
	.w7(32'h3bc90c9a),
	.w8(32'h3c1059bb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b321870),
	.w1(32'h3c1c0999),
	.w2(32'h39ea9b60),
	.w3(32'hbb133c58),
	.w4(32'h3b46dbce),
	.w5(32'h3c63ae01),
	.w6(32'h3c83f30a),
	.w7(32'h3ad4233b),
	.w8(32'h3c485138),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bfba3),
	.w1(32'hbb047e64),
	.w2(32'h3c6afec9),
	.w3(32'h3be3ea95),
	.w4(32'h3c191eda),
	.w5(32'h3b72c567),
	.w6(32'h3a913027),
	.w7(32'h3c4cf356),
	.w8(32'h3b819dbc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7da2),
	.w1(32'h3c2092a2),
	.w2(32'hbb05e72e),
	.w3(32'h3ba2e016),
	.w4(32'h3a79adf5),
	.w5(32'hba087cbb),
	.w6(32'h3c48f1c4),
	.w7(32'hbaeda3ee),
	.w8(32'hbc0b0a91),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205e28),
	.w1(32'hbbe8be3f),
	.w2(32'h3b190f01),
	.w3(32'h3c25d497),
	.w4(32'hbb3c96bc),
	.w5(32'h39e806a8),
	.w6(32'h3af6cd28),
	.w7(32'hbb98dd13),
	.w8(32'hb997c643),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c2f48),
	.w1(32'hba75c79a),
	.w2(32'hbc1079ef),
	.w3(32'hbaa5ef8d),
	.w4(32'hbbd10260),
	.w5(32'hbc2c59a8),
	.w6(32'hb8b59a61),
	.w7(32'hbbf09681),
	.w8(32'hbc25c857),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd51628),
	.w1(32'hbc4de7f3),
	.w2(32'hbb25792a),
	.w3(32'hbb8f11ef),
	.w4(32'hbb4c0ada),
	.w5(32'hba8178eb),
	.w6(32'hbb8fc254),
	.w7(32'hbb4ad69b),
	.w8(32'hbc0fabd2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe60ab3),
	.w1(32'hbb9f1424),
	.w2(32'h3ad39b6a),
	.w3(32'h3c1fcbdf),
	.w4(32'h3bbebdb7),
	.w5(32'h3b3b914a),
	.w6(32'hbb4747da),
	.w7(32'h3b0894a3),
	.w8(32'hba8f2f86),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a70e8),
	.w1(32'hbbd2fe2c),
	.w2(32'h3b8b7b1a),
	.w3(32'hbbe43699),
	.w4(32'h39f2fcf6),
	.w5(32'hbb0a2d43),
	.w6(32'hbc1df24f),
	.w7(32'h3c336038),
	.w8(32'h3c16d4b7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3244e0),
	.w1(32'h3bbe24f8),
	.w2(32'hbb20e82f),
	.w3(32'h38bc4bed),
	.w4(32'hbac7cf5f),
	.w5(32'h3bcfb59f),
	.w6(32'h3c8d9df0),
	.w7(32'h3b008fb3),
	.w8(32'hbb6d1d08),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97bd88),
	.w1(32'hbba358ad),
	.w2(32'h3b305fb3),
	.w3(32'h3c52e346),
	.w4(32'h3a2724bd),
	.w5(32'hbb7b3f69),
	.w6(32'h39d10bb0),
	.w7(32'h3b7e5f95),
	.w8(32'h3ae9ffc0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c130672),
	.w1(32'h3b8a9e1b),
	.w2(32'h3bd47878),
	.w3(32'hbb269b68),
	.w4(32'h39170a39),
	.w5(32'h3bbe94f1),
	.w6(32'hbb0b8b6c),
	.w7(32'h3b32d950),
	.w8(32'h3b6aee6e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b734489),
	.w1(32'hbb294464),
	.w2(32'hbb3b12ac),
	.w3(32'hbb0d4c09),
	.w4(32'h3aeb03e2),
	.w5(32'h3b784b81),
	.w6(32'h3b3227f6),
	.w7(32'hbb617356),
	.w8(32'h3c37ce37),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14536c),
	.w1(32'h3b73bb50),
	.w2(32'hbb8e4fe8),
	.w3(32'h3af21ff3),
	.w4(32'hbb1c1167),
	.w5(32'h3a22de1c),
	.w6(32'h3af2029b),
	.w7(32'hbbf7a524),
	.w8(32'h3b421236),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c02a9),
	.w1(32'h392afc34),
	.w2(32'hbba01074),
	.w3(32'h3ba70dfe),
	.w4(32'hbb45b44f),
	.w5(32'hbb18197c),
	.w6(32'h3afd8022),
	.w7(32'hbb9161c8),
	.w8(32'hbb162339),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00c42c),
	.w1(32'h3be5af11),
	.w2(32'h3a1159fb),
	.w3(32'h3b5e3686),
	.w4(32'hba5b16e9),
	.w5(32'h3b9e49a8),
	.w6(32'h3b8b3c39),
	.w7(32'h3c24e395),
	.w8(32'hb9efaef0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8893cc),
	.w1(32'h3a86d5ed),
	.w2(32'hbc3ce1bd),
	.w3(32'hbbd39c98),
	.w4(32'hbc126868),
	.w5(32'h3baf3b1b),
	.w6(32'h3bf1e85a),
	.w7(32'h3b9a63cb),
	.w8(32'h3cf6ac75),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836ff2),
	.w1(32'hbc8510dc),
	.w2(32'hbbf968a7),
	.w3(32'hbc20980d),
	.w4(32'hbbc43d21),
	.w5(32'hb9c05a87),
	.w6(32'hbb951583),
	.w7(32'hbb110a4f),
	.w8(32'h3bb4be5c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8ca8),
	.w1(32'h3bd3b8a4),
	.w2(32'h3c52fda9),
	.w3(32'hba3e1f3c),
	.w4(32'h3bf343c5),
	.w5(32'h3b9f0a03),
	.w6(32'h39744e04),
	.w7(32'h3cdc5ab6),
	.w8(32'h3c400e8c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9854b),
	.w1(32'hbb16a15a),
	.w2(32'h3b3a0c7d),
	.w3(32'h3a0d99ca),
	.w4(32'hbb9e5b29),
	.w5(32'h3c1f4d15),
	.w6(32'hbc4e797d),
	.w7(32'hba3f9416),
	.w8(32'hba90c7a3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc124cf3),
	.w1(32'hbc0bf380),
	.w2(32'h3c12011c),
	.w3(32'h3aa4d458),
	.w4(32'h3c901de9),
	.w5(32'hbcfa384c),
	.w6(32'h3c10517d),
	.w7(32'h3cbb72e7),
	.w8(32'hbdb8cb22),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04cac6),
	.w1(32'h3cd5833e),
	.w2(32'hbcacd0d0),
	.w3(32'h3bfb48f7),
	.w4(32'hbb2d11a8),
	.w5(32'h3ba69c36),
	.w6(32'h3d11738b),
	.w7(32'hbcaab254),
	.w8(32'h3ca73ead),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86ff16),
	.w1(32'hbc20fc2c),
	.w2(32'h3a67c3c2),
	.w3(32'hbb21866f),
	.w4(32'hbb43a331),
	.w5(32'h3be89f4f),
	.w6(32'hbb1f9338),
	.w7(32'h3b1804c0),
	.w8(32'h3baceb27),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43839),
	.w1(32'h3bbb95eb),
	.w2(32'h3a7b2649),
	.w3(32'hba61e3e3),
	.w4(32'h3b0d69e1),
	.w5(32'hbb415b58),
	.w6(32'h3c029623),
	.w7(32'hba7772b2),
	.w8(32'h3c37c7d7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf29186),
	.w1(32'h3b8549c5),
	.w2(32'h3b96dab5),
	.w3(32'h3b5439df),
	.w4(32'hbae347f1),
	.w5(32'hba996d15),
	.w6(32'h3c2ae274),
	.w7(32'h3a8eed00),
	.w8(32'hbc24b504),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba48e6),
	.w1(32'hb89de20c),
	.w2(32'h3b0fb120),
	.w3(32'h3c0fb4b1),
	.w4(32'hbc2582f9),
	.w5(32'h3c347048),
	.w6(32'h3bc5b05a),
	.w7(32'hbc1aa1ae),
	.w8(32'h3b13edd5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e76f2),
	.w1(32'h3bd17cc3),
	.w2(32'h3b47d70d),
	.w3(32'h39970147),
	.w4(32'h3b0e8653),
	.w5(32'h3c0ac332),
	.w6(32'h3c80c055),
	.w7(32'h3badc4f4),
	.w8(32'hbb768c54),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb465a9c),
	.w1(32'hbbe13684),
	.w2(32'h3b1d4ed5),
	.w3(32'hbbbdb7fd),
	.w4(32'hbc2f0cf1),
	.w5(32'h3c458d6f),
	.w6(32'hbb110be4),
	.w7(32'hbb2574f8),
	.w8(32'hbc6c50c9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2870f),
	.w1(32'hbbca16ed),
	.w2(32'h3c99d313),
	.w3(32'h3a4f83e2),
	.w4(32'h3aa9f350),
	.w5(32'h3cb89bcd),
	.w6(32'h3aed3c61),
	.w7(32'hba735051),
	.w8(32'h3be27570),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b1300),
	.w1(32'h3c8a3ee8),
	.w2(32'h3b145f46),
	.w3(32'hb983d45f),
	.w4(32'h3bff5465),
	.w5(32'hbd0553e1),
	.w6(32'hbca41875),
	.w7(32'h3be76f32),
	.w8(32'hbd3f5e06),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6994),
	.w1(32'h3bea7731),
	.w2(32'hb9c19260),
	.w3(32'h3b77acda),
	.w4(32'hbacf551c),
	.w5(32'h3b5c434f),
	.w6(32'h3ce52521),
	.w7(32'hbb6266f7),
	.w8(32'h3bb3acbd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d4bf),
	.w1(32'h3ba21014),
	.w2(32'h3938a3a4),
	.w3(32'hba864b2c),
	.w4(32'hbb9d853b),
	.w5(32'h3c1cb7bd),
	.w6(32'h3991bc26),
	.w7(32'h3a9d562a),
	.w8(32'hbab985a7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf12e17),
	.w1(32'h3bca7af5),
	.w2(32'hbc777e9c),
	.w3(32'h3b2e0bd1),
	.w4(32'h3c2103e9),
	.w5(32'hbc55e9ab),
	.w6(32'h3c208a57),
	.w7(32'h3a8237d1),
	.w8(32'h3c8792ea),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c068689),
	.w1(32'hbba9bfd8),
	.w2(32'hbc36b509),
	.w3(32'h3c330a1b),
	.w4(32'hbb854427),
	.w5(32'hbcd046d9),
	.w6(32'h399c956e),
	.w7(32'hbca47d49),
	.w8(32'hbcb53ef9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce59df),
	.w1(32'h3b887c21),
	.w2(32'h3c7c2257),
	.w3(32'hbc95605f),
	.w4(32'h3c44ec90),
	.w5(32'hbc4429c2),
	.w6(32'hbbdf0bc0),
	.w7(32'h3c400efd),
	.w8(32'hbcabfcff),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be0b4),
	.w1(32'h3ba99e6c),
	.w2(32'hbb65b92a),
	.w3(32'h3b87ee03),
	.w4(32'h3c3fe50a),
	.w5(32'hbc2e0885),
	.w6(32'h3b97cb42),
	.w7(32'h3c8e94dd),
	.w8(32'hbb4acd42),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86d7be),
	.w1(32'hbcfdbec5),
	.w2(32'h3c506458),
	.w3(32'hbc08cd16),
	.w4(32'h3b84366d),
	.w5(32'hbbebe674),
	.w6(32'hbd00b8bc),
	.w7(32'h39b9005b),
	.w8(32'hbadb562a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23845e),
	.w1(32'hba544323),
	.w2(32'hbba66326),
	.w3(32'hbc32fb46),
	.w4(32'hbc28b410),
	.w5(32'h3b86ec34),
	.w6(32'hbc469834),
	.w7(32'hb9fbf142),
	.w8(32'h3d015c6c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c486397),
	.w1(32'hbb98b9fb),
	.w2(32'hbb9a92a7),
	.w3(32'hbc8a9146),
	.w4(32'h39a41230),
	.w5(32'hba972450),
	.w6(32'hbbcedd14),
	.w7(32'h3aa0fddc),
	.w8(32'hbcd5fa3a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b79d7),
	.w1(32'h3c5fb48d),
	.w2(32'hbc01a843),
	.w3(32'hbca29ecf),
	.w4(32'hba694b45),
	.w5(32'hbbac71d5),
	.w6(32'hbc834522),
	.w7(32'h3a4d2311),
	.w8(32'hbbff8979),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9610d),
	.w1(32'h3bc4974c),
	.w2(32'h3bb9336c),
	.w3(32'hba28726c),
	.w4(32'h3b92ed94),
	.w5(32'h3c0b6a0b),
	.w6(32'h3b9e68df),
	.w7(32'hbbc3abc2),
	.w8(32'hbbb2a28a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82c575),
	.w1(32'h3b689730),
	.w2(32'h3c6ec86e),
	.w3(32'hbaa247d9),
	.w4(32'h3c473230),
	.w5(32'hbcb32b75),
	.w6(32'h3ac56308),
	.w7(32'h3c9a8eca),
	.w8(32'hbd0f4008),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b34c),
	.w1(32'h3c35401b),
	.w2(32'h3a3b9e92),
	.w3(32'h3c53f219),
	.w4(32'h3c8a3953),
	.w5(32'hbc8ddfa3),
	.w6(32'h3bec4dfe),
	.w7(32'h3c331e72),
	.w8(32'h3caceeac),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8498dd),
	.w1(32'hbb0c3987),
	.w2(32'hbb84b4dc),
	.w3(32'h3b5160dc),
	.w4(32'hba92db95),
	.w5(32'h3aeffc8e),
	.w6(32'hbbed60d1),
	.w7(32'hbbdf3f8a),
	.w8(32'h3c6e66a7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c747369),
	.w1(32'h3b980e8c),
	.w2(32'hbb9fb006),
	.w3(32'h3ac1d01a),
	.w4(32'h3b23c27c),
	.w5(32'hbca3cae0),
	.w6(32'h3b7eb8e0),
	.w7(32'hbbe3bac7),
	.w8(32'hbb654751),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce8aee),
	.w1(32'hbc467bd8),
	.w2(32'hbb1ec1fb),
	.w3(32'hbba199cd),
	.w4(32'hbc7eb194),
	.w5(32'h3be188da),
	.w6(32'hbcea9db5),
	.w7(32'hbc9b784b),
	.w8(32'h3cdacffb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b190a5d),
	.w1(32'hbc41bfdc),
	.w2(32'h3c0abc8b),
	.w3(32'hbc0ffc5f),
	.w4(32'h3bc6f86e),
	.w5(32'hb9960c3d),
	.w6(32'hbc4bc159),
	.w7(32'hb9dc009f),
	.w8(32'hbca0070d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ded38),
	.w1(32'h3bd9c826),
	.w2(32'hba85e818),
	.w3(32'h3c737039),
	.w4(32'hbbd85fa9),
	.w5(32'h3bab969e),
	.w6(32'h3aaae087),
	.w7(32'hbba3e4a8),
	.w8(32'h3d98eae1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf0e3e0),
	.w1(32'hbd40367c),
	.w2(32'h3b6b8203),
	.w3(32'h3c39eaaa),
	.w4(32'hba1d6b26),
	.w5(32'hbb8dea0e),
	.w6(32'hbc19dd72),
	.w7(32'h3ba637e1),
	.w8(32'hbcd28867),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57029c),
	.w1(32'hbbb49950),
	.w2(32'hbcc449a7),
	.w3(32'hbc475471),
	.w4(32'hbca8334a),
	.w5(32'hbbd0f847),
	.w6(32'hbc047b10),
	.w7(32'hbca2da7f),
	.w8(32'h3bab7c4a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe32a47),
	.w1(32'hbc869667),
	.w2(32'hb9adc41a),
	.w3(32'hbcc85330),
	.w4(32'hbc94d0b8),
	.w5(32'h3cbb7ca7),
	.w6(32'hbc941db2),
	.w7(32'h3a94a093),
	.w8(32'h3d06bbe8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3e8f6),
	.w1(32'hbc9fdbf6),
	.w2(32'h3c8e71db),
	.w3(32'hbbb1f8f2),
	.w4(32'h3bc35deb),
	.w5(32'hbbf7df67),
	.w6(32'hba9f80d9),
	.w7(32'h3b3ba958),
	.w8(32'hbccebe1b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc880e99),
	.w1(32'h3c01fd18),
	.w2(32'hbbbc6a24),
	.w3(32'h3c9bfaac),
	.w4(32'hbb7a3c49),
	.w5(32'h3b3359fc),
	.w6(32'h3c6abcf3),
	.w7(32'hbbaf422d),
	.w8(32'hbca2c53b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993550),
	.w1(32'h3c5c42ce),
	.w2(32'hbb8d59c8),
	.w3(32'h3c1c9b4d),
	.w4(32'hba935d43),
	.w5(32'h3aee1a5c),
	.w6(32'h3b3a5533),
	.w7(32'hbbcb839d),
	.w8(32'h3c0ef214),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41d57f),
	.w1(32'hba655c4a),
	.w2(32'h3bff3b50),
	.w3(32'h37e871bb),
	.w4(32'h3c510cce),
	.w5(32'hbc5fd8d0),
	.w6(32'hbb13dda1),
	.w7(32'h3b3d5a1f),
	.w8(32'hbce35f00),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc51230),
	.w1(32'h3c6579d7),
	.w2(32'hbb9a4409),
	.w3(32'h3cac7bff),
	.w4(32'hbc88d01c),
	.w5(32'h3cbb90ff),
	.w6(32'h3ac129df),
	.w7(32'hbc15308e),
	.w8(32'h3d6c4807),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab3b69),
	.w1(32'hbca0f6d8),
	.w2(32'h3bbf574c),
	.w3(32'hbc87441e),
	.w4(32'h3c4ef7a4),
	.w5(32'h3a6b994e),
	.w6(32'hbc802001),
	.w7(32'h3c5ba5b7),
	.w8(32'hbb931776),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b416),
	.w1(32'h3ba03f04),
	.w2(32'h3b08919c),
	.w3(32'hbb093820),
	.w4(32'hbb550ea0),
	.w5(32'h3ca7c546),
	.w6(32'h3bb8f1e4),
	.w7(32'hbbe3f514),
	.w8(32'h3c9d8486),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a8db5),
	.w1(32'hbbbd4ef2),
	.w2(32'hbb738c71),
	.w3(32'hbaa52c99),
	.w4(32'hbb146571),
	.w5(32'h3aca55df),
	.w6(32'hbb33a7fd),
	.w7(32'hbbd8708a),
	.w8(32'h3c5ba43a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74a4cc),
	.w1(32'h3b0807fb),
	.w2(32'h3bab223f),
	.w3(32'h39fb6ced),
	.w4(32'hbc24295c),
	.w5(32'h3c9f3024),
	.w6(32'h3a79c46a),
	.w7(32'h3bc7d7e5),
	.w8(32'h3c33745c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840a08),
	.w1(32'hbc18d1c9),
	.w2(32'hbc6709a3),
	.w3(32'hbc8404c7),
	.w4(32'h3bdc977d),
	.w5(32'hbca7c85d),
	.w6(32'hbc574ce8),
	.w7(32'hbc2942c0),
	.w8(32'h3cbb4bba),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d447d0a),
	.w1(32'hbd0a11f1),
	.w2(32'hbacda021),
	.w3(32'hbc6abaed),
	.w4(32'hbaffe8de),
	.w5(32'hbb6a3183),
	.w6(32'hbc7e1b54),
	.w7(32'h39f8e9b9),
	.w8(32'h3b8b32b4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0e87c),
	.w1(32'h3a2b4522),
	.w2(32'hba613a84),
	.w3(32'h3aa6c7e6),
	.w4(32'hbc66729c),
	.w5(32'h3b733921),
	.w6(32'h3b9d3515),
	.w7(32'hbcaee7b1),
	.w8(32'h3cf0f801),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74dbc9),
	.w1(32'hbc556343),
	.w2(32'h3bb2c9c1),
	.w3(32'hbb90a061),
	.w4(32'h3b4b4167),
	.w5(32'h3b7d70c0),
	.w6(32'hbbf05f51),
	.w7(32'h3a14341e),
	.w8(32'h3aa9891a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule