module layer_10_featuremap_147(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb852a337),
	.w1(32'h39599ab6),
	.w2(32'h3a818ccf),
	.w3(32'h38390e5a),
	.w4(32'hb89038ce),
	.w5(32'h394e70bb),
	.w6(32'hb84ab412),
	.w7(32'hba0308b9),
	.w8(32'hba86d201),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cdee7),
	.w1(32'hbac68659),
	.w2(32'hba4a5772),
	.w3(32'hba16801e),
	.w4(32'hba5f23e9),
	.w5(32'hb97fdebb),
	.w6(32'hb8d26db8),
	.w7(32'h39848761),
	.w8(32'h3769f406),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb660bbda),
	.w1(32'h38b9428e),
	.w2(32'hb9bc2db3),
	.w3(32'hb85f6e85),
	.w4(32'h39802314),
	.w5(32'h399dc1f2),
	.w6(32'h398c844a),
	.w7(32'h398b963d),
	.w8(32'h39387bb6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca4102),
	.w1(32'hba1bd143),
	.w2(32'hb999ac11),
	.w3(32'h39d92f69),
	.w4(32'hb98d0f74),
	.w5(32'hb959ce65),
	.w6(32'hb9559b05),
	.w7(32'hb89a1400),
	.w8(32'h394886ac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7c96f),
	.w1(32'hb9ef4d1b),
	.w2(32'h3a48712c),
	.w3(32'h38fb5c1d),
	.w4(32'hba928c0b),
	.w5(32'hb89d75da),
	.w6(32'h39c228cf),
	.w7(32'h3a44db43),
	.w8(32'h39e8e16e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80952d5),
	.w1(32'h3897e066),
	.w2(32'h393a653e),
	.w3(32'h39b67eba),
	.w4(32'hb8f023bc),
	.w5(32'h39bc98a4),
	.w6(32'hb91c07a2),
	.w7(32'h391df671),
	.w8(32'h394a1f7b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac66ee8),
	.w1(32'h39fa0dcb),
	.w2(32'h3a25a84b),
	.w3(32'h3a12d7a7),
	.w4(32'h3a16f200),
	.w5(32'h39e3bb19),
	.w6(32'hba16c9db),
	.w7(32'h38168839),
	.w8(32'hb94afa31),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae077c9),
	.w1(32'h3a785a21),
	.w2(32'hb9ca794d),
	.w3(32'h3ace0929),
	.w4(32'hbaab70b7),
	.w5(32'hbae9da2e),
	.w6(32'h3aae0dc7),
	.w7(32'hba0a5455),
	.w8(32'h3a273e19),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93317c6),
	.w1(32'h3a17877e),
	.w2(32'h39753d7f),
	.w3(32'hb8d2009c),
	.w4(32'h39d17a2b),
	.w5(32'h3a7bec20),
	.w6(32'h39ac7f64),
	.w7(32'h39406be9),
	.w8(32'h3a2ed928),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1298ce),
	.w1(32'hba8f4871),
	.w2(32'h3a36d990),
	.w3(32'hbada39b7),
	.w4(32'hbac4f6af),
	.w5(32'h3a72dd98),
	.w6(32'h3a24e5be),
	.w7(32'hb93f7732),
	.w8(32'h3aaaaf92),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ebd166),
	.w1(32'hb9ae6a1f),
	.w2(32'hb9f42714),
	.w3(32'hb99c5046),
	.w4(32'hb9f60f9b),
	.w5(32'hba03d40a),
	.w6(32'hbab242d0),
	.w7(32'hba911c79),
	.w8(32'hba73b05c),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93d650),
	.w1(32'h3aa5fe47),
	.w2(32'h3a98e4dd),
	.w3(32'hba18d271),
	.w4(32'hb989edc1),
	.w5(32'h39cd3fac),
	.w6(32'hbaf72d9b),
	.w7(32'hbaea234a),
	.w8(32'hba9fd49f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036b91),
	.w1(32'hbafc5c96),
	.w2(32'hbb4c5b1c),
	.w3(32'hbb1eb256),
	.w4(32'hbb00c189),
	.w5(32'hbb684010),
	.w6(32'hbb482b10),
	.w7(32'hbb87cc21),
	.w8(32'hbb4ed54b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c7f1),
	.w1(32'hbab82e81),
	.w2(32'hbae59d39),
	.w3(32'hb9c66b46),
	.w4(32'hba89967f),
	.w5(32'hba97f906),
	.w6(32'hbae9b0c7),
	.w7(32'hba33ccf8),
	.w8(32'hba47c95d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf344a8),
	.w1(32'h388500a0),
	.w2(32'h3ae4dd68),
	.w3(32'hbad852c8),
	.w4(32'hbadb69ff),
	.w5(32'h3a419571),
	.w6(32'h3a9d0969),
	.w7(32'h36532862),
	.w8(32'h3a8a6683),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e04459),
	.w1(32'hba60edbc),
	.w2(32'hb8f93e94),
	.w3(32'h38151258),
	.w4(32'hba6b2fe5),
	.w5(32'h39b7a108),
	.w6(32'h3a58169b),
	.w7(32'h37c7b515),
	.w8(32'h3acfd6da),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397edae8),
	.w1(32'h395d3a98),
	.w2(32'hb9f4affc),
	.w3(32'hb78a7e87),
	.w4(32'h394d74dc),
	.w5(32'h3920c0ca),
	.w6(32'hb83685b8),
	.w7(32'h38978923),
	.w8(32'hba1e6a06),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f18af),
	.w1(32'h3b801ee1),
	.w2(32'h3acf342c),
	.w3(32'h3b39cdd5),
	.w4(32'h3b2686bd),
	.w5(32'hb8920f4f),
	.w6(32'h3b5a840e),
	.w7(32'h3a1fe158),
	.w8(32'h3a404be1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c2dff),
	.w1(32'h39026463),
	.w2(32'hbb01458f),
	.w3(32'hba33d63b),
	.w4(32'hba478fe8),
	.w5(32'hba9656d4),
	.w6(32'h39b6ac9f),
	.w7(32'hbab64578),
	.w8(32'hbaeb4e50),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c3aaf),
	.w1(32'h374e4252),
	.w2(32'hb9b35a4b),
	.w3(32'h39207bf7),
	.w4(32'hb9035061),
	.w5(32'hb8000a65),
	.w6(32'hb7fa5570),
	.w7(32'hb87222cc),
	.w8(32'hb8f0930e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab534b),
	.w1(32'hb895e909),
	.w2(32'h39500c16),
	.w3(32'hb90d7383),
	.w4(32'hb9e18b1e),
	.w5(32'hb9800585),
	.w6(32'hba2fad7e),
	.w7(32'hb9ca914e),
	.w8(32'hb9c3fadf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aaeeaf),
	.w1(32'hb8ebb4fb),
	.w2(32'hbaed507d),
	.w3(32'hba10f676),
	.w4(32'h396e135e),
	.w5(32'h388be3df),
	.w6(32'hb7e2d944),
	.w7(32'hb95bc35a),
	.w8(32'hb80399c9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1226aa),
	.w1(32'h3c159ed9),
	.w2(32'h3b77da6e),
	.w3(32'h3bb3646d),
	.w4(32'h3beadc1a),
	.w5(32'h3b8ecfa8),
	.w6(32'h3c5a4cc2),
	.w7(32'h3c105d41),
	.w8(32'h3c0860f3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac02c8),
	.w1(32'hbb046c73),
	.w2(32'hba383024),
	.w3(32'hbad654e9),
	.w4(32'hbb1e6391),
	.w5(32'hb96b65e9),
	.w6(32'hb9a2a30f),
	.w7(32'hba024e14),
	.w8(32'h3ad1ff9e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c22ea),
	.w1(32'hbaa2fb86),
	.w2(32'h395b2369),
	.w3(32'hbb530c94),
	.w4(32'hbb5b0117),
	.w5(32'hb9395a9c),
	.w6(32'hb82a56a2),
	.w7(32'hb89f5ea9),
	.w8(32'h3b1d30ba),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c8b6d),
	.w1(32'h39c72e83),
	.w2(32'h3883de2e),
	.w3(32'hb9614d38),
	.w4(32'h3882c10f),
	.w5(32'h3a29d7d9),
	.w6(32'h37adb830),
	.w7(32'h38575d72),
	.w8(32'h389befa9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1d5f8),
	.w1(32'hb98775d4),
	.w2(32'hb9b033f2),
	.w3(32'hb9bf6f7a),
	.w4(32'hb9d1818e),
	.w5(32'hb9418437),
	.w6(32'hb9daa11c),
	.w7(32'hb9b4553d),
	.w8(32'hb9b9055b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e3610),
	.w1(32'hba3ad112),
	.w2(32'h3a685a9c),
	.w3(32'hbab11c9b),
	.w4(32'hbac63e4e),
	.w5(32'h3a1820fc),
	.w6(32'hba8e280c),
	.w7(32'hbaac3441),
	.w8(32'hb8f3189b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381775d6),
	.w1(32'hb94b4ea8),
	.w2(32'h386e52b8),
	.w3(32'hba0b7259),
	.w4(32'hb9e4cb81),
	.w5(32'hb9e8fe41),
	.w6(32'hba7ff997),
	.w7(32'hba96b282),
	.w8(32'hba6a4675),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1065b1),
	.w1(32'hbae3f170),
	.w2(32'hba97615f),
	.w3(32'hbacf4a41),
	.w4(32'hbad88dd8),
	.w5(32'hb9270641),
	.w6(32'hb9b7da63),
	.w7(32'h36d2c8ce),
	.w8(32'h3b06af3c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba086be1),
	.w1(32'hb8fff9cc),
	.w2(32'h38c09628),
	.w3(32'hb9cfc9a9),
	.w4(32'hb9e5bb47),
	.w5(32'hb9abc8a8),
	.w6(32'hba03c201),
	.w7(32'hb93b4e46),
	.w8(32'hb9518a68),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a775f5),
	.w1(32'hb8d51a27),
	.w2(32'hb9292c8e),
	.w3(32'hb9ac1ce9),
	.w4(32'hb980f93c),
	.w5(32'hb8c8420e),
	.w6(32'hb981c17e),
	.w7(32'hb93986c5),
	.w8(32'hb8d12c43),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a802de2),
	.w1(32'hba361a7d),
	.w2(32'hb9654dc7),
	.w3(32'h396d651a),
	.w4(32'hb9e81980),
	.w5(32'h3a0d48b3),
	.w6(32'h3a3a42bf),
	.w7(32'h3a0018a8),
	.w8(32'h3a03f495),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab28289),
	.w1(32'hba9b946b),
	.w2(32'h399c7dbd),
	.w3(32'hb9f2f3ac),
	.w4(32'hba86674c),
	.w5(32'h3a39398c),
	.w6(32'hba05f42d),
	.w7(32'hb8f9be45),
	.w8(32'h3a7383b4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394a13be),
	.w1(32'h3a24e5be),
	.w2(32'h3a48364f),
	.w3(32'h39d941ca),
	.w4(32'h39b2aa3a),
	.w5(32'h39b10626),
	.w6(32'h389a9748),
	.w7(32'h398bc87c),
	.w8(32'h3897498f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89571a),
	.w1(32'h39d5f8b1),
	.w2(32'h39e54a4a),
	.w3(32'h39058071),
	.w4(32'hb99c1720),
	.w5(32'h36719da4),
	.w6(32'hb9839eea),
	.w7(32'hba061a03),
	.w8(32'hb9928ff7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78627d),
	.w1(32'h3b054d49),
	.w2(32'hb945d13c),
	.w3(32'h3a014bdb),
	.w4(32'h3a655c6f),
	.w5(32'h3a6b50ad),
	.w6(32'h3aafddf7),
	.w7(32'h3b410f93),
	.w8(32'h3b3b45bf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81c228),
	.w1(32'hbb89fcc9),
	.w2(32'h3aa22c72),
	.w3(32'hbbc2d0d5),
	.w4(32'hbba57b53),
	.w5(32'h3a932ef5),
	.w6(32'hbb3d153e),
	.w7(32'hbb397f4a),
	.w8(32'h3b57c8f8),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c2fe),
	.w1(32'hbb0ec7cf),
	.w2(32'h3a5f3dc5),
	.w3(32'hbb4d0e87),
	.w4(32'hbb1d3d51),
	.w5(32'h3a8aa214),
	.w6(32'hba7a1acf),
	.w7(32'hba33d919),
	.w8(32'h3ad911b5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e184d1),
	.w1(32'hba04eb35),
	.w2(32'h380edfb2),
	.w3(32'hba40c285),
	.w4(32'hbab2f5c9),
	.w5(32'hb9efc30b),
	.w6(32'hb97d2283),
	.w7(32'hb9f6538a),
	.w8(32'hba033412),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389ea998),
	.w1(32'hba262eb8),
	.w2(32'hbaa7b9fb),
	.w3(32'hb887dac6),
	.w4(32'hb99c1dfc),
	.w5(32'hba3daee1),
	.w6(32'hb9f2c15d),
	.w7(32'hba61204c),
	.w8(32'hb9bf376c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b4a76),
	.w1(32'hb9fc3a26),
	.w2(32'hb9e5d938),
	.w3(32'hba165a17),
	.w4(32'hba0dbd58),
	.w5(32'hb9c6c1be),
	.w6(32'h37daaaef),
	.w7(32'h38b1ed8b),
	.w8(32'h38f01618),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac9b4b),
	.w1(32'hba1891bb),
	.w2(32'h3a3a4278),
	.w3(32'hbac6e9e2),
	.w4(32'hba312879),
	.w5(32'h3a7da907),
	.w6(32'hba950ca9),
	.w7(32'hb9284a3f),
	.w8(32'h3a85dca2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53c363),
	.w1(32'hb8077556),
	.w2(32'h3a0fd186),
	.w3(32'h39271729),
	.w4(32'hba03b92e),
	.w5(32'h3aa2a3d3),
	.w6(32'h3b26094e),
	.w7(32'h39fe262c),
	.w8(32'h3ad4afe2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72168d),
	.w1(32'hba83750f),
	.w2(32'hb8b70a9b),
	.w3(32'hba817017),
	.w4(32'hba830afd),
	.w5(32'h3a121b44),
	.w6(32'h385bc52d),
	.w7(32'h3985810f),
	.w8(32'h3b0d89fa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba993cd5),
	.w1(32'hbaf4ddd6),
	.w2(32'hba5d8aee),
	.w3(32'hbae66a68),
	.w4(32'hbb0ef7d3),
	.w5(32'hba5657d0),
	.w6(32'h3a5b358e),
	.w7(32'h3877b808),
	.w8(32'h3b058f1a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac67824),
	.w1(32'hb9b9d4c3),
	.w2(32'h39fec863),
	.w3(32'h39e2e858),
	.w4(32'hbac8c1c5),
	.w5(32'hba0bdfdf),
	.w6(32'h3b10397f),
	.w7(32'h3aa90683),
	.w8(32'h3b0af644),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd435fa),
	.w1(32'h3b93b3d2),
	.w2(32'hb9952446),
	.w3(32'h3bc42f5e),
	.w4(32'h3ba453d6),
	.w5(32'h39f59bf7),
	.w6(32'h3bc65d61),
	.w7(32'h3b2b51b6),
	.w8(32'hbac413a8),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3bc41),
	.w1(32'hb96480ab),
	.w2(32'hba08bd0f),
	.w3(32'hb9b941f4),
	.w4(32'hb8c69e53),
	.w5(32'hb9011f86),
	.w6(32'hb7bbd871),
	.w7(32'hb97a8249),
	.w8(32'hb9363470),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374a5af2),
	.w1(32'hb9aefcf2),
	.w2(32'hb9befd8f),
	.w3(32'hb8ca6385),
	.w4(32'hba1ea430),
	.w5(32'hb92d8294),
	.w6(32'hb9d59ce8),
	.w7(32'hb98feb40),
	.w8(32'hb98920f1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f2bf3),
	.w1(32'hba9538cc),
	.w2(32'hba5cc4a8),
	.w3(32'hba28be6d),
	.w4(32'hba5d3f6a),
	.w5(32'hba559da7),
	.w6(32'hba398655),
	.w7(32'hba08a67a),
	.w8(32'hba27dd38),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d2211c),
	.w1(32'hba71f8e5),
	.w2(32'hbaa4fbd7),
	.w3(32'hba967606),
	.w4(32'hba60da0e),
	.w5(32'hba25bb2c),
	.w6(32'h39852f69),
	.w7(32'h362aaebc),
	.w8(32'h3aa6ba9b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d1152),
	.w1(32'h3a0e94fb),
	.w2(32'h39d53482),
	.w3(32'hb9a42765),
	.w4(32'h38c6eacd),
	.w5(32'h3a4bc902),
	.w6(32'h3a0d5dd0),
	.w7(32'h3a56dc64),
	.w8(32'h3a3a024a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b982c65),
	.w1(32'h3b72a794),
	.w2(32'h3b1b1cf3),
	.w3(32'h3b4b5e65),
	.w4(32'h3ac9ce17),
	.w5(32'h3ae714c1),
	.w6(32'h3b365076),
	.w7(32'h3b098428),
	.w8(32'h3b20df07),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39913c7d),
	.w1(32'h3a3efaf0),
	.w2(32'h3a44eae2),
	.w3(32'h3962032d),
	.w4(32'h39772012),
	.w5(32'h3a08e132),
	.w6(32'hb920201e),
	.w7(32'h36a7dd9e),
	.w8(32'h39e3858f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39846943),
	.w1(32'hba7ab8b7),
	.w2(32'hbaded9f7),
	.w3(32'h38deb0b9),
	.w4(32'hba66b0a3),
	.w5(32'hbaa5c2e4),
	.w6(32'hba69f182),
	.w7(32'hba7a26e3),
	.w8(32'hb59ecfa8),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13e189),
	.w1(32'hb9c89d72),
	.w2(32'hba49816c),
	.w3(32'hba14cede),
	.w4(32'hb9c635cf),
	.w5(32'hba2bcbe6),
	.w6(32'hba02d8de),
	.w7(32'hb9ede4eb),
	.w8(32'hba230f2c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb95a1),
	.w1(32'hbaa43f8e),
	.w2(32'h3661a56c),
	.w3(32'hba65b912),
	.w4(32'hba9d17d7),
	.w5(32'hba3a9fc0),
	.w6(32'hb98c297b),
	.w7(32'h380744e6),
	.w8(32'hb8c8c872),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd195c),
	.w1(32'hb9be9d4e),
	.w2(32'hb921346f),
	.w3(32'hb8fd58b1),
	.w4(32'hb9ddf760),
	.w5(32'hb67f2f61),
	.w6(32'hb9fb1b13),
	.w7(32'hb9384444),
	.w8(32'hb8fd37f1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb586c023),
	.w1(32'hb99919ee),
	.w2(32'hb9fe5c16),
	.w3(32'hb96743f9),
	.w4(32'hb9e67154),
	.w5(32'hb97449f2),
	.w6(32'hba1cfa81),
	.w7(32'hb9d6d38e),
	.w8(32'hb9008d01),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859f39d),
	.w1(32'h3a0b9bf0),
	.w2(32'hba018c3c),
	.w3(32'hba853eff),
	.w4(32'hba6d7804),
	.w5(32'hba820d74),
	.w6(32'hb9ca40c2),
	.w7(32'hbab154d9),
	.w8(32'hbaa3bf56),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102420),
	.w1(32'h3a80620b),
	.w2(32'h388e2182),
	.w3(32'h3ab60cf6),
	.w4(32'h39ec0f35),
	.w5(32'h397697ed),
	.w6(32'h3a6edc9d),
	.w7(32'h38c1e0c5),
	.w8(32'h3a9433f5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca4fc1),
	.w1(32'hb797f3d0),
	.w2(32'h39e96fd2),
	.w3(32'hb9e73611),
	.w4(32'h3a318c0b),
	.w5(32'h3a7dcef3),
	.w6(32'h3998a5aa),
	.w7(32'h3a091fb5),
	.w8(32'h3a1853f4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9068959),
	.w1(32'h3968fb9c),
	.w2(32'h3a0557b9),
	.w3(32'h3a24b9d3),
	.w4(32'h3a06e73e),
	.w5(32'h39ec5d15),
	.w6(32'h3927944e),
	.w7(32'h3977bcca),
	.w8(32'hb971aae6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df5b8a),
	.w1(32'h39cfdcad),
	.w2(32'hb9879c6f),
	.w3(32'h3921345b),
	.w4(32'h3a12a968),
	.w5(32'h39897680),
	.w6(32'h3999a53a),
	.w7(32'h3930fcf6),
	.w8(32'hb9ab6f4b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93cba5a),
	.w1(32'hba03c6ac),
	.w2(32'hb9f78f0a),
	.w3(32'h383b4f34),
	.w4(32'hb8bb8c87),
	.w5(32'h360ffb82),
	.w6(32'hb921db01),
	.w7(32'hb6b6a9c3),
	.w8(32'h39bc61a1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acacf58),
	.w1(32'hba52ebdf),
	.w2(32'hbb25af7c),
	.w3(32'h3af72f10),
	.w4(32'hb9a33b30),
	.w5(32'hb9b7a9f9),
	.w6(32'h3a114e09),
	.w7(32'hbab7a2a3),
	.w8(32'hba2a6a77),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bd34d0),
	.w1(32'hb8ef5b59),
	.w2(32'h3a02773e),
	.w3(32'hbada0da4),
	.w4(32'hba9c0c7a),
	.w5(32'hb98498dc),
	.w6(32'h3a4e85e4),
	.w7(32'hb8707b26),
	.w8(32'h3b09ad4b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b397c97),
	.w1(32'h3ad76ee6),
	.w2(32'h3b1d4a51),
	.w3(32'h3a1875c4),
	.w4(32'hb90edae9),
	.w5(32'h3a184db1),
	.w6(32'h3ac62eb1),
	.w7(32'h38e4f21c),
	.w8(32'h3aaafbc9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb286ae8),
	.w1(32'hbb842190),
	.w2(32'h3936ade7),
	.w3(32'hbb5d66ff),
	.w4(32'hbba1e3a2),
	.w5(32'hbaab458b),
	.w6(32'hbaa29294),
	.w7(32'h39b26195),
	.w8(32'h3b4471d7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c621c),
	.w1(32'hb884d7e2),
	.w2(32'hb99d6062),
	.w3(32'hba1e435b),
	.w4(32'h37dfb344),
	.w5(32'h3886da1c),
	.w6(32'hb882a9e8),
	.w7(32'h371966c6),
	.w8(32'h38925fd3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e4ddc0),
	.w1(32'hb984d788),
	.w2(32'hb9e334d9),
	.w3(32'h37d63420),
	.w4(32'hb9b7df5c),
	.w5(32'hb936fe85),
	.w6(32'hb9c481c6),
	.w7(32'hb986ae52),
	.w8(32'hb9690c9c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982d610),
	.w1(32'hb9c7ac14),
	.w2(32'hba20e0c2),
	.w3(32'hb8e14699),
	.w4(32'hb9c6d8ce),
	.w5(32'hb971dccc),
	.w6(32'hb9d604bd),
	.w7(32'hb9a61071),
	.w8(32'hb92c5b1d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d26cd),
	.w1(32'h391c594d),
	.w2(32'hb9d11c6d),
	.w3(32'h3a24a912),
	.w4(32'hba7fea80),
	.w5(32'hba5baeb5),
	.w6(32'hb9ebd1e0),
	.w7(32'hbad7eadc),
	.w8(32'hba6552fa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eba33e),
	.w1(32'h3935db3f),
	.w2(32'h38e51dbd),
	.w3(32'hb947c43e),
	.w4(32'h393817e6),
	.w5(32'h399e8ba9),
	.w6(32'hb6c6d5c4),
	.w7(32'h38ceedd7),
	.w8(32'hb8aef2f0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8617cb),
	.w1(32'h3aad637a),
	.w2(32'hba6c6eee),
	.w3(32'h3b556e92),
	.w4(32'h3ae933a7),
	.w5(32'hb80a8038),
	.w6(32'h3ad2f280),
	.w7(32'hb9f93dfd),
	.w8(32'hba438faf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b505525),
	.w1(32'h3b47ab6f),
	.w2(32'h39ccc6b0),
	.w3(32'h3b0c3a64),
	.w4(32'h3a782c60),
	.w5(32'hba1706ed),
	.w6(32'h3a9cfa9c),
	.w7(32'hba1fab43),
	.w8(32'h38ee755a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bac54),
	.w1(32'hbafeba65),
	.w2(32'hbad479f8),
	.w3(32'hbaa20735),
	.w4(32'hbac9c869),
	.w5(32'hba9648b8),
	.w6(32'hba6394c9),
	.w7(32'hbae52e14),
	.w8(32'hba6f540d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20609b),
	.w1(32'hb93ecb22),
	.w2(32'hb9530ada),
	.w3(32'h39ca177e),
	.w4(32'hb9b1585d),
	.w5(32'h39c27b7a),
	.w6(32'h3991f623),
	.w7(32'hb99dd0e9),
	.w8(32'h390ff479),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada9bb1),
	.w1(32'h399751e3),
	.w2(32'hb9b06129),
	.w3(32'h3aaf384f),
	.w4(32'hb70878b5),
	.w5(32'hb9f6c159),
	.w6(32'hba2ed1af),
	.w7(32'hb9c9571f),
	.w8(32'hb9cef1b0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb58ef),
	.w1(32'hba9ab1ec),
	.w2(32'hba20a6e0),
	.w3(32'hba864abd),
	.w4(32'hba7e3cbc),
	.w5(32'hb9a7fc4c),
	.w6(32'hb97be40e),
	.w7(32'hb9d44bd3),
	.w8(32'h3a715bf4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b193f1e),
	.w1(32'h3b057ddc),
	.w2(32'h38486538),
	.w3(32'h3ae5b248),
	.w4(32'h3abe2264),
	.w5(32'h39215caf),
	.w6(32'h3ae2f473),
	.w7(32'h3a90aa19),
	.w8(32'hba6bfcde),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9525f2d),
	.w1(32'hb91faebd),
	.w2(32'hb9e1ec67),
	.w3(32'hb9abc2e2),
	.w4(32'hb915cf5e),
	.w5(32'hb90ce2b7),
	.w6(32'hb955b324),
	.w7(32'hb91a4283),
	.w8(32'hb91fc481),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37940fc5),
	.w1(32'h38b6df0d),
	.w2(32'hb8a7dda1),
	.w3(32'hb9aeaab6),
	.w4(32'h37e5ddcf),
	.w5(32'h388d75e2),
	.w6(32'hb872d4e3),
	.w7(32'h38d627d8),
	.w8(32'h37b10be0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ac1457),
	.w1(32'hb917f7a8),
	.w2(32'hb9a86028),
	.w3(32'h37a17459),
	.w4(32'h3a0f81eb),
	.w5(32'hb904a654),
	.w6(32'hb9752d4a),
	.w7(32'hb96f7c37),
	.w8(32'h3913b160),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91705c0),
	.w1(32'hb98d2c2f),
	.w2(32'hba906159),
	.w3(32'h396316c0),
	.w4(32'hb9be3948),
	.w5(32'hba2f5e16),
	.w6(32'h3765b31d),
	.w7(32'hb966ab7a),
	.w8(32'hb95a2e20),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e0ff2e),
	.w1(32'hba0612c6),
	.w2(32'hb9b194a6),
	.w3(32'hbac0adad),
	.w4(32'hbabe4051),
	.w5(32'h3a490349),
	.w6(32'hba474cac),
	.w7(32'hba773b44),
	.w8(32'h3ad3864a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c0b52),
	.w1(32'h39709731),
	.w2(32'h39e5183b),
	.w3(32'hb76b4697),
	.w4(32'hba1a3263),
	.w5(32'hb9de225c),
	.w6(32'hb9785966),
	.w7(32'hb9a074fd),
	.w8(32'hb9b1e323),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8929c9),
	.w1(32'hb8839530),
	.w2(32'h37c000fe),
	.w3(32'hb99e61a5),
	.w4(32'hb8390740),
	.w5(32'h39c06602),
	.w6(32'h3a5a81bd),
	.w7(32'h3a9642df),
	.w8(32'h3a947269),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0a167),
	.w1(32'h3ba6f9be),
	.w2(32'h3b1706d3),
	.w3(32'h3bae7ddf),
	.w4(32'h3b38e057),
	.w5(32'hb9e82bb5),
	.w6(32'h3bd365b6),
	.w7(32'h3b4b56e6),
	.w8(32'h3a1fc4b0),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44acef),
	.w1(32'hb9e57611),
	.w2(32'h3afaadc0),
	.w3(32'hba9fd7a6),
	.w4(32'hba6c478b),
	.w5(32'h3aac5dcf),
	.w6(32'hba70543a),
	.w7(32'hba2414cc),
	.w8(32'h3a3db648),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62fa6),
	.w1(32'h39fda8be),
	.w2(32'h39829a95),
	.w3(32'h3a566eb4),
	.w4(32'h3acc2d47),
	.w5(32'h3adc80ec),
	.w6(32'h3b013b56),
	.w7(32'h3ae71a16),
	.w8(32'h3ac26708),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389fdb79),
	.w1(32'h3a98ef63),
	.w2(32'h39cf057a),
	.w3(32'hba5b58ef),
	.w4(32'h3a475b68),
	.w5(32'h39cf84a8),
	.w6(32'h39ab3c4a),
	.w7(32'h3aa01009),
	.w8(32'h3a616139),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac79fd5),
	.w1(32'h3a6e093b),
	.w2(32'h3b1b77af),
	.w3(32'hb95198bc),
	.w4(32'h3a2b8cd2),
	.w5(32'h3af42feb),
	.w6(32'hba85dd0b),
	.w7(32'h39e36bde),
	.w8(32'h3b276b8a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a753b),
	.w1(32'h39a2b70d),
	.w2(32'hb8cfea39),
	.w3(32'h397ba810),
	.w4(32'h3886fdd6),
	.w5(32'h39d10ec7),
	.w6(32'h3ab3bd29),
	.w7(32'h3aa37222),
	.w8(32'h3a9e09c2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0b6fd),
	.w1(32'hb936b5d5),
	.w2(32'hb675b5e7),
	.w3(32'hba6885fa),
	.w4(32'hba49aea2),
	.w5(32'h3a580667),
	.w6(32'hba2a0e26),
	.w7(32'hba885b70),
	.w8(32'h3a27af4f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eb64f),
	.w1(32'hb9313417),
	.w2(32'hba17baff),
	.w3(32'hb9b99605),
	.w4(32'h398ea23d),
	.w5(32'h3941e690),
	.w6(32'h39969eb1),
	.w7(32'h370f268c),
	.w8(32'h39c4cd68),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a3891),
	.w1(32'hb9539b1b),
	.w2(32'h3ae48de8),
	.w3(32'h3a3b6980),
	.w4(32'hb8d0bddc),
	.w5(32'h3b048067),
	.w6(32'h3ac8205c),
	.w7(32'h3a9115ca),
	.w8(32'h3b33c61c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9003a),
	.w1(32'h3a98c25c),
	.w2(32'h3a8031db),
	.w3(32'h39ac6ce0),
	.w4(32'hb9e760c2),
	.w5(32'h3a5e79e7),
	.w6(32'h3970f760),
	.w7(32'hb9a4500b),
	.w8(32'h3ac1063b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ca831),
	.w1(32'h3b43dea2),
	.w2(32'h3a4d0ca8),
	.w3(32'h3b7974f8),
	.w4(32'h3b10bf32),
	.w5(32'h39f77aad),
	.w6(32'h3bafd88c),
	.w7(32'h3b913dd8),
	.w8(32'h39f62f90),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69db0a),
	.w1(32'hbb5ffd4e),
	.w2(32'h3ba5d133),
	.w3(32'hbba1d1db),
	.w4(32'hbb68ae5b),
	.w5(32'h3ba4d852),
	.w6(32'hbb1503e7),
	.w7(32'hb9fbbc9e),
	.w8(32'h3bde5b22),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98862b),
	.w1(32'hbb2e67ef),
	.w2(32'hba197bb0),
	.w3(32'hba929bed),
	.w4(32'hba91127d),
	.w5(32'h39818943),
	.w6(32'h39aed7b4),
	.w7(32'h3a9bdc2e),
	.w8(32'h3b43ab91),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b272c91),
	.w1(32'h3a93f87f),
	.w2(32'h38d903c2),
	.w3(32'h3a0e82e4),
	.w4(32'h39a140e1),
	.w5(32'h3aa98b06),
	.w6(32'h3a7f8231),
	.w7(32'h3a4fc214),
	.w8(32'h3ac86058),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92d940),
	.w1(32'hba1411c2),
	.w2(32'hba34c977),
	.w3(32'hba4fb432),
	.w4(32'hba3c7493),
	.w5(32'hb9f9852f),
	.w6(32'hb987bc6c),
	.w7(32'hb9839347),
	.w8(32'hb9a7042b),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4a01d),
	.w1(32'h3bd3e86a),
	.w2(32'h3b3569a7),
	.w3(32'h3b9a9d62),
	.w4(32'h3b5d5579),
	.w5(32'h3b23e7e0),
	.w6(32'h3b3a5209),
	.w7(32'h3afdd8e7),
	.w8(32'hb97fb3ca),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba354082),
	.w1(32'hb9d04421),
	.w2(32'h3b06be12),
	.w3(32'hba9991b6),
	.w4(32'hba7fc9d7),
	.w5(32'h3aec9bf3),
	.w6(32'hbad9cdf3),
	.w7(32'hbab0576c),
	.w8(32'h3922fa1e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da1790),
	.w1(32'h3a043a5b),
	.w2(32'h36a37d71),
	.w3(32'hb9162186),
	.w4(32'h3a2214a4),
	.w5(32'h39fe07df),
	.w6(32'h39950002),
	.w7(32'h39ae4c81),
	.w8(32'h39870894),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c725b1),
	.w1(32'hb9d18cc1),
	.w2(32'h36d3078a),
	.w3(32'h3a3b702f),
	.w4(32'hb99ccd80),
	.w5(32'hb9ffcd59),
	.w6(32'h391abcc6),
	.w7(32'h3951c106),
	.w8(32'hb92e3b16),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a38a2),
	.w1(32'hbb16d00a),
	.w2(32'hbafd41ba),
	.w3(32'hba543c6c),
	.w4(32'hbaa5dca4),
	.w5(32'hba07d0b4),
	.w6(32'h3999d40d),
	.w7(32'hba065b8a),
	.w8(32'hb985737f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad04f34),
	.w1(32'hbb118cba),
	.w2(32'hbab5f55c),
	.w3(32'hbaed1753),
	.w4(32'hbb20255a),
	.w5(32'hba1fde97),
	.w6(32'hb9fdc366),
	.w7(32'hb9c4ec4e),
	.w8(32'h3a8c6bb1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbf271),
	.w1(32'hba2e666f),
	.w2(32'h38381d9b),
	.w3(32'hba7850ee),
	.w4(32'hba8f0a79),
	.w5(32'h3af0ca80),
	.w6(32'h3ae8271c),
	.w7(32'hb9796b52),
	.w8(32'h3b27fd02),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba448246),
	.w1(32'hba89e72a),
	.w2(32'hba1006ef),
	.w3(32'hba295f9a),
	.w4(32'hba98f481),
	.w5(32'hb8eb3680),
	.w6(32'h3aa0fffc),
	.w7(32'h3ab386fa),
	.w8(32'h3b0f24e9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995011e),
	.w1(32'h3a94f861),
	.w2(32'h3a71568d),
	.w3(32'h39977770),
	.w4(32'h39d50b94),
	.w5(32'h3970620a),
	.w6(32'hb84bba36),
	.w7(32'hb981eb5d),
	.w8(32'h39121195),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9badc),
	.w1(32'h39ebc010),
	.w2(32'h3a0ba074),
	.w3(32'h39fe9488),
	.w4(32'h38f804a1),
	.w5(32'h39b9ea1b),
	.w6(32'h39c992a6),
	.w7(32'h39354cc0),
	.w8(32'h39903e9e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a0955a),
	.w1(32'hbaaf853e),
	.w2(32'hba23ec2a),
	.w3(32'hb9e66ac3),
	.w4(32'hbab30f00),
	.w5(32'h3949f14f),
	.w6(32'hb9d24485),
	.w7(32'hb98c1dd0),
	.w8(32'h3a785680),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02c7ab),
	.w1(32'hba3d2fb5),
	.w2(32'hba6a8b86),
	.w3(32'hba0a6b8d),
	.w4(32'hba137be4),
	.w5(32'hb9c2f63e),
	.w6(32'hba62ec6d),
	.w7(32'hba430bcf),
	.w8(32'hba16231c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d6242),
	.w1(32'hb96559b9),
	.w2(32'hb9d120b4),
	.w3(32'hb9e40f3b),
	.w4(32'hb8ded5b7),
	.w5(32'hb80b2d7e),
	.w6(32'hb9db1979),
	.w7(32'hb999be3a),
	.w8(32'hb90c3dc2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87416be),
	.w1(32'hb8e896a0),
	.w2(32'hb90c80ec),
	.w3(32'h38b886f2),
	.w4(32'hb7a22c02),
	.w5(32'h3965a9a3),
	.w6(32'hb9bac5b3),
	.w7(32'hb93a375c),
	.w8(32'hb8732dbe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a86c2b),
	.w1(32'hb9810377),
	.w2(32'hbabbc806),
	.w3(32'h3a06a9ba),
	.w4(32'hb94465dd),
	.w5(32'hba21e16b),
	.w6(32'hb9550df7),
	.w7(32'hb94e096f),
	.w8(32'hb9f0e7dd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6f42f),
	.w1(32'hbab57bf6),
	.w2(32'hb987ed9e),
	.w3(32'hbacae4cc),
	.w4(32'hbaae2a63),
	.w5(32'hb76c3341),
	.w6(32'h391af9da),
	.w7(32'h39489e2d),
	.w8(32'h3abbeb8f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad5d17),
	.w1(32'hb91294d5),
	.w2(32'h3936d6ca),
	.w3(32'h39c88d56),
	.w4(32'hba2394c3),
	.w5(32'h384a66bf),
	.w6(32'hba1affed),
	.w7(32'hb8e92587),
	.w8(32'hb9398257),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a857a87),
	.w1(32'h3a87a049),
	.w2(32'h3a93549e),
	.w3(32'h3a3f9c61),
	.w4(32'h3a6a6d33),
	.w5(32'h39561a99),
	.w6(32'h39f2f076),
	.w7(32'h39d6efdb),
	.w8(32'hb98a3cf6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb6651),
	.w1(32'hbb5a68d4),
	.w2(32'hbb0fd14c),
	.w3(32'hbac1d65e),
	.w4(32'hbb2f7b50),
	.w5(32'hbaa5f84f),
	.w6(32'h3938f67b),
	.w7(32'hb9d093a1),
	.w8(32'h3a88b2cf),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdf352),
	.w1(32'hb9c3117b),
	.w2(32'hba8e22db),
	.w3(32'hb98f7974),
	.w4(32'h39e9b651),
	.w5(32'hb912955e),
	.w6(32'hba20b449),
	.w7(32'hba6f6fa2),
	.w8(32'hb93afe9b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf5ba7),
	.w1(32'h38b06a63),
	.w2(32'h38fd0d63),
	.w3(32'hba7be69d),
	.w4(32'hb90c7cff),
	.w5(32'h39c45c45),
	.w6(32'hb9e96633),
	.w7(32'h39c64d48),
	.w8(32'h38e9eb1c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c000e),
	.w1(32'h3965330e),
	.w2(32'h396f1a50),
	.w3(32'h39dc123e),
	.w4(32'hb9b473bc),
	.w5(32'hb9979f96),
	.w6(32'hb9e6eb3b),
	.w7(32'hb8f5801e),
	.w8(32'hb97bb872),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393000d3),
	.w1(32'hba8b3ab5),
	.w2(32'hba750fff),
	.w3(32'hb9be8234),
	.w4(32'hba3a8b0e),
	.w5(32'hba202621),
	.w6(32'hb96216b6),
	.w7(32'hba4f22a9),
	.w8(32'hb881005e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0085f0),
	.w1(32'h3a4313d5),
	.w2(32'h3a201db0),
	.w3(32'hba0e5585),
	.w4(32'hb80539b7),
	.w5(32'h38c33e41),
	.w6(32'h39b09941),
	.w7(32'hba3de425),
	.w8(32'hb9ced137),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a1abf),
	.w1(32'h39993003),
	.w2(32'h3a8655ed),
	.w3(32'h3972ddb3),
	.w4(32'h390d5852),
	.w5(32'h3a9a4a79),
	.w6(32'h399eee8b),
	.w7(32'h384c45d3),
	.w8(32'h3a23b8ae),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17ca6a),
	.w1(32'h3902d109),
	.w2(32'h3903fc3a),
	.w3(32'hba3e5b19),
	.w4(32'h3987ccc4),
	.w5(32'h393b2bd9),
	.w6(32'h39cfc8df),
	.w7(32'h3954edcf),
	.w8(32'h37aa423b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a129dd0),
	.w1(32'h37dc662b),
	.w2(32'h399bfa9a),
	.w3(32'hb8c38a7d),
	.w4(32'h37bdb801),
	.w5(32'hb9460232),
	.w6(32'h37860812),
	.w7(32'h396e5f07),
	.w8(32'h3a594131),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9672e7c),
	.w1(32'hbaaa14c7),
	.w2(32'h38439da9),
	.w3(32'h3842a154),
	.w4(32'hba8a546e),
	.w5(32'hb9ea969f),
	.w6(32'h39e8319b),
	.w7(32'h39c97a36),
	.w8(32'h3a739949),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98886f5),
	.w1(32'h3ab4c489),
	.w2(32'h3a5a3935),
	.w3(32'hba19c632),
	.w4(32'h3a26652d),
	.w5(32'h394f4f79),
	.w6(32'h3a8e10b9),
	.w7(32'hb896b944),
	.w8(32'h3a001f3c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e205f9),
	.w1(32'hb9b8731d),
	.w2(32'hb94b6954),
	.w3(32'h39d4345c),
	.w4(32'h3a041053),
	.w5(32'h399ed7d2),
	.w6(32'h3a267008),
	.w7(32'h398b1f60),
	.w8(32'hb8afca27),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b941f6c),
	.w1(32'h3b377f9a),
	.w2(32'h3ae81904),
	.w3(32'h3b362198),
	.w4(32'h3ad8c0e8),
	.w5(32'h3a9b9f89),
	.w6(32'h3b69843d),
	.w7(32'h3aada0be),
	.w8(32'h3a7b9dd7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b5944),
	.w1(32'hb9b21581),
	.w2(32'h39c923f9),
	.w3(32'hb97162ae),
	.w4(32'hb9b4b77e),
	.w5(32'h3a40f06a),
	.w6(32'h3aac4701),
	.w7(32'h3aaf62a1),
	.w8(32'h3adfa62a),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a168c7b),
	.w1(32'h3a9a8a22),
	.w2(32'h3a0e4816),
	.w3(32'hba138a75),
	.w4(32'h395747ac),
	.w5(32'h3a9cf132),
	.w6(32'h3a64509d),
	.w7(32'h38e7f53e),
	.w8(32'h3adda59a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e107),
	.w1(32'h3b668f57),
	.w2(32'h3aeb35f0),
	.w3(32'h3b5712d5),
	.w4(32'h3b8fb1ec),
	.w5(32'h3b0c766f),
	.w6(32'h3b5faea5),
	.w7(32'h3b5b487c),
	.w8(32'h3b1763fb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4581f5),
	.w1(32'hbae6e68a),
	.w2(32'hba6d8ab1),
	.w3(32'h3a8a3681),
	.w4(32'hbaa7a241),
	.w5(32'hba2ba8a3),
	.w6(32'h399fac0b),
	.w7(32'h3a7d5364),
	.w8(32'h3a4abe13),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79630a),
	.w1(32'h3a1485c5),
	.w2(32'h3a52e674),
	.w3(32'h39eb710c),
	.w4(32'h396bdff0),
	.w5(32'h399c1351),
	.w6(32'h3ae60f38),
	.w7(32'h3b0b2a2f),
	.w8(32'h3b28ec99),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb920cb4d),
	.w1(32'hba689b46),
	.w2(32'hba273829),
	.w3(32'hba665c67),
	.w4(32'hba5296d9),
	.w5(32'hba126a8b),
	.w6(32'hba49c317),
	.w7(32'hba586306),
	.w8(32'hb912bb31),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba077a29),
	.w1(32'hbb3a7292),
	.w2(32'hbae290a5),
	.w3(32'hbab9774b),
	.w4(32'hbb483f86),
	.w5(32'hba149314),
	.w6(32'h3ae0a1fc),
	.w7(32'h3aab854a),
	.w8(32'h3b101396),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a702014),
	.w1(32'h3a745bfc),
	.w2(32'h3b2438e3),
	.w3(32'h3a7b7da9),
	.w4(32'h393b481b),
	.w5(32'h3a03e846),
	.w6(32'h3aeb0284),
	.w7(32'h3a3b0b2c),
	.w8(32'h3a914974),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21f9fa),
	.w1(32'h3a068d1e),
	.w2(32'hb90cccd1),
	.w3(32'h38a212ab),
	.w4(32'h39eafcec),
	.w5(32'h38a38afc),
	.w6(32'h391f6517),
	.w7(32'hb9e8ed9c),
	.w8(32'hb9f08603),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba017589),
	.w1(32'h39ade848),
	.w2(32'h3a3dc658),
	.w3(32'hb9345d90),
	.w4(32'h39908b80),
	.w5(32'h3998708b),
	.w6(32'h3a2a6b51),
	.w7(32'h3a3820ab),
	.w8(32'h3a2e7e74),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e4339),
	.w1(32'hba13a071),
	.w2(32'h399aa734),
	.w3(32'hb983ef1a),
	.w4(32'hb9ce8925),
	.w5(32'h39926cb1),
	.w6(32'hba3a00ef),
	.w7(32'hba4fc44e),
	.w8(32'h3a09121f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67a702),
	.w1(32'h3991c9a4),
	.w2(32'h3a5e3f2e),
	.w3(32'h394a56de),
	.w4(32'hba4be0d3),
	.w5(32'h3a606b6c),
	.w6(32'h3abdc199),
	.w7(32'h3a0e3793),
	.w8(32'h3a4ce789),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b198f),
	.w1(32'hbb136076),
	.w2(32'hbb2c899b),
	.w3(32'hbae15f60),
	.w4(32'hbb1a431b),
	.w5(32'hbb56329e),
	.w6(32'hbaecc496),
	.w7(32'hbb8b911b),
	.w8(32'hbb41eb6f),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9878fd8),
	.w1(32'hba036810),
	.w2(32'hba6f14cc),
	.w3(32'hb92ced3e),
	.w4(32'hb987e6ee),
	.w5(32'hba04796b),
	.w6(32'hb99d77f0),
	.w7(32'hba12ee6d),
	.w8(32'hb86cc8f6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21bd28),
	.w1(32'hbb12ff72),
	.w2(32'hbaf68c75),
	.w3(32'hba30d0dc),
	.w4(32'hbab1dee8),
	.w5(32'hba134b33),
	.w6(32'hba9433c1),
	.w7(32'hbacf3ac9),
	.w8(32'h3827ed10),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20292d),
	.w1(32'h370d5109),
	.w2(32'h397ef9ba),
	.w3(32'hb9ebb0cc),
	.w4(32'h37b486c3),
	.w5(32'h3a5d74cb),
	.w6(32'h3ab26d88),
	.w7(32'h3abedc56),
	.w8(32'h3b1769a3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f57f6),
	.w1(32'h3a874df9),
	.w2(32'h39e9186f),
	.w3(32'h3b37831a),
	.w4(32'h3ac7c2ee),
	.w5(32'h39933193),
	.w6(32'h38a260ac),
	.w7(32'hb9ed9c13),
	.w8(32'hbab68692),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba149b4e),
	.w1(32'hba765ad4),
	.w2(32'h39299d70),
	.w3(32'hb9f20fb2),
	.w4(32'hbac29e55),
	.w5(32'hb95af4c9),
	.w6(32'h3a90abfd),
	.w7(32'h39cfd4f6),
	.w8(32'h3ac446e1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41c00a),
	.w1(32'hba2d10e6),
	.w2(32'hb7e9e9d2),
	.w3(32'hba3e0765),
	.w4(32'hba53dd24),
	.w5(32'hb9ecbe23),
	.w6(32'hb8ce5fa2),
	.w7(32'h3a8539f6),
	.w8(32'h3adbfdbf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80f423),
	.w1(32'hb9c072c3),
	.w2(32'hba289a24),
	.w3(32'hba392d10),
	.w4(32'hb97de4c0),
	.w5(32'hb9f3aa32),
	.w6(32'hb9c81597),
	.w7(32'hba0abf36),
	.w8(32'hb949605f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88bc2ea),
	.w1(32'hba8badd7),
	.w2(32'hb993cb66),
	.w3(32'hba2bea82),
	.w4(32'hba9c2acb),
	.w5(32'hb97044fb),
	.w6(32'hba8e765f),
	.w7(32'hb9af3552),
	.w8(32'h3a7ac114),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb231824),
	.w1(32'hba9b20fb),
	.w2(32'h3a04e92c),
	.w3(32'hbb1c01c7),
	.w4(32'hbaeeb270),
	.w5(32'h398c867a),
	.w6(32'hba9d01e8),
	.w7(32'hbafb1585),
	.w8(32'h3ac978e7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab5cb6),
	.w1(32'h3a431fb3),
	.w2(32'h3aab17f8),
	.w3(32'h38d47c2f),
	.w4(32'h38cea451),
	.w5(32'h3a63fc28),
	.w6(32'h3a1d35a9),
	.w7(32'h3a0a3a93),
	.w8(32'h3a51f2a0),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36c494),
	.w1(32'h3a8ff7a4),
	.w2(32'hb8f62073),
	.w3(32'h3b1509c5),
	.w4(32'h3a916b90),
	.w5(32'h39e153c2),
	.w6(32'h3a8b6531),
	.w7(32'h39f13d78),
	.w8(32'hb82b11ac),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931ab9b),
	.w1(32'hb9c4074b),
	.w2(32'hb9cc998c),
	.w3(32'h384231dd),
	.w4(32'hb981e356),
	.w5(32'hb9b53a16),
	.w6(32'hb9632a9e),
	.w7(32'hb99e4062),
	.w8(32'hb7c120ab),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a602f6c),
	.w1(32'h3a0d7298),
	.w2(32'h3ae576c2),
	.w3(32'h39c39a6e),
	.w4(32'h3a2021c0),
	.w5(32'h3a4c9e39),
	.w6(32'h3aab7c4e),
	.w7(32'h3a948831),
	.w8(32'h3ab31d03),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06cbc8),
	.w1(32'hb94ce7cd),
	.w2(32'hba2a3167),
	.w3(32'h39d0dbe0),
	.w4(32'h39848980),
	.w5(32'hb93a375f),
	.w6(32'hb94a9647),
	.w7(32'hba231bc6),
	.w8(32'h3abc8430),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac39fd4),
	.w1(32'hb796643f),
	.w2(32'hb8acc0f2),
	.w3(32'h396491da),
	.w4(32'h394e2a36),
	.w5(32'h3a69431d),
	.w6(32'h3992ca5e),
	.w7(32'h39a4b832),
	.w8(32'h3aee6752),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a188ac7),
	.w1(32'h38e129b7),
	.w2(32'h37b1e5f7),
	.w3(32'h3a4e5a06),
	.w4(32'hb8535cff),
	.w5(32'hb9c5cfec),
	.w6(32'hb91adff7),
	.w7(32'hb9896613),
	.w8(32'hb7b30ed7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cfdb6e),
	.w1(32'h3a57e29c),
	.w2(32'h39e3d4e2),
	.w3(32'hba8dccd1),
	.w4(32'hba9c6822),
	.w5(32'hbb04a96d),
	.w6(32'h3a1542f8),
	.w7(32'h3a3dd63b),
	.w8(32'hbadd3719),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b3c59),
	.w1(32'hb99f5ca3),
	.w2(32'hb9a01bd6),
	.w3(32'h3a34df19),
	.w4(32'h390800d2),
	.w5(32'hb7b54b12),
	.w6(32'h3584168f),
	.w7(32'hb8f2d26b),
	.w8(32'hb94927ce),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d8329),
	.w1(32'h3957decb),
	.w2(32'hb88310d2),
	.w3(32'h39256d78),
	.w4(32'h37c17ef1),
	.w5(32'hb900327c),
	.w6(32'h389fc433),
	.w7(32'hb9a2a870),
	.w8(32'hb9bdd353),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a144b),
	.w1(32'hbac0f85b),
	.w2(32'h399be11e),
	.w3(32'hba190745),
	.w4(32'hba964138),
	.w5(32'h3a3159d8),
	.w6(32'hb814f3ea),
	.w7(32'h37ef60e3),
	.w8(32'h3ae8d7a8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3132b3),
	.w1(32'h3b325998),
	.w2(32'h3ad73736),
	.w3(32'h3adb1421),
	.w4(32'h3b1a91b3),
	.w5(32'h3ae23edb),
	.w6(32'h3b8ad30e),
	.w7(32'h3b86062c),
	.w8(32'h3b8945d3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa4290),
	.w1(32'h39dae2b7),
	.w2(32'h3a7a9f9c),
	.w3(32'h3a86a3f9),
	.w4(32'h397673db),
	.w5(32'h39d65b6b),
	.w6(32'h39f754cd),
	.w7(32'h3a175bdd),
	.w8(32'h3a16961a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2be86),
	.w1(32'hbb03ac0f),
	.w2(32'hba61aaeb),
	.w3(32'hba278c67),
	.w4(32'hbb0cce03),
	.w5(32'hba306386),
	.w6(32'hb887834f),
	.w7(32'hb8a88c4e),
	.w8(32'h3a957eb3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959bc4d),
	.w1(32'h3902941a),
	.w2(32'hb9051f69),
	.w3(32'hb9979907),
	.w4(32'h3a965577),
	.w5(32'h3a4857e2),
	.w6(32'h3a50bb7f),
	.w7(32'h3a19daee),
	.w8(32'hb890338d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8718c),
	.w1(32'hbb3d534b),
	.w2(32'hb9eed826),
	.w3(32'hba869968),
	.w4(32'hbb58749b),
	.w5(32'hbaa465be),
	.w6(32'hbb6f66d0),
	.w7(32'hbba5b506),
	.w8(32'hbadf456c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891154a),
	.w1(32'hba0f5389),
	.w2(32'h391ecbf3),
	.w3(32'hb91c9557),
	.w4(32'hb945d630),
	.w5(32'h3a08a3bc),
	.w6(32'h386ce1ba),
	.w7(32'hb957ba12),
	.w8(32'h3ac3f3dd),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8c7c8),
	.w1(32'h3aafff54),
	.w2(32'h39b947ef),
	.w3(32'h3aa2909a),
	.w4(32'h3a509a5a),
	.w5(32'hb86dbba9),
	.w6(32'h3b30bc45),
	.w7(32'h3ac334e1),
	.w8(32'h3a7d8291),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee0857),
	.w1(32'h3a478c41),
	.w2(32'h397910f2),
	.w3(32'hb918ea4b),
	.w4(32'h3a7ba7be),
	.w5(32'h3a395c44),
	.w6(32'h3a9f8807),
	.w7(32'h3a4929f3),
	.w8(32'h3a48252f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab67d4a),
	.w1(32'h3a081a56),
	.w2(32'h3a20963d),
	.w3(32'h3a5edd60),
	.w4(32'h39d3b09f),
	.w5(32'h3a25743f),
	.w6(32'h36cbfcd2),
	.w7(32'h397ffe5c),
	.w8(32'h3a253e8f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9960390),
	.w1(32'hb9b87541),
	.w2(32'hb99dc0d6),
	.w3(32'hb97b5709),
	.w4(32'hba058390),
	.w5(32'hb9e70f86),
	.w6(32'hb920005b),
	.w7(32'hb974c7bb),
	.w8(32'hb9d23afe),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a86d22),
	.w1(32'hbad36a85),
	.w2(32'hbae19db4),
	.w3(32'hb9984295),
	.w4(32'hbac2f68d),
	.w5(32'hbadc1607),
	.w6(32'hb8dbfef3),
	.w7(32'hb98b8132),
	.w8(32'h395bbb53),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba311bda),
	.w1(32'h39b3ab36),
	.w2(32'hb9b0888b),
	.w3(32'hba40d6e4),
	.w4(32'h398c7bde),
	.w5(32'hb9b13750),
	.w6(32'h3a6b4983),
	.w7(32'h3a1f74d0),
	.w8(32'hba1fbbb9),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab207ee),
	.w1(32'hba25884d),
	.w2(32'hba135b7a),
	.w3(32'hba287edd),
	.w4(32'h37a114a6),
	.w5(32'hb8bafe67),
	.w6(32'hb96b742f),
	.w7(32'hba873c8d),
	.w8(32'hba4cbf78),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba146124),
	.w1(32'hb9d3273c),
	.w2(32'hb9297c45),
	.w3(32'hb98fe1d4),
	.w4(32'hb9f73604),
	.w5(32'hba33344c),
	.w6(32'hb8a4f180),
	.w7(32'hb9e13259),
	.w8(32'hb97df6d0),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816f12d),
	.w1(32'h39407511),
	.w2(32'h3a1087bd),
	.w3(32'hb92f2b15),
	.w4(32'h39a778d4),
	.w5(32'h39978900),
	.w6(32'h3a03c0ae),
	.w7(32'h3a2f6226),
	.w8(32'h3a2322cc),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dee0f),
	.w1(32'hb9177a1d),
	.w2(32'h3a04fc54),
	.w3(32'h3960ed85),
	.w4(32'hb8744b35),
	.w5(32'h39d773b3),
	.w6(32'h39dcc833),
	.w7(32'h3a31c4f9),
	.w8(32'h3aae7ffa),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0734ec),
	.w1(32'h3a9142c6),
	.w2(32'h3ab1e572),
	.w3(32'h3a212fc0),
	.w4(32'h3a3246fe),
	.w5(32'h3aaaa2a9),
	.w6(32'h3abbf3cf),
	.w7(32'h3ad593c1),
	.w8(32'h3b3a0473),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9ac10),
	.w1(32'h39e45fa4),
	.w2(32'h3986c0ed),
	.w3(32'h3ab39a6d),
	.w4(32'hb952dded),
	.w5(32'hb9a6a350),
	.w6(32'h39aab931),
	.w7(32'hb99a06a5),
	.w8(32'hb9f41953),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d4c9c),
	.w1(32'hb9a8d71b),
	.w2(32'hb9ba8c7b),
	.w3(32'hb92ce9a5),
	.w4(32'hb9974b86),
	.w5(32'hba24e065),
	.w6(32'h39994b28),
	.w7(32'hb9650bce),
	.w8(32'hba310201),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba334798),
	.w1(32'hbaa8ab84),
	.w2(32'hbb7f76ec),
	.w3(32'hbb7e9ec2),
	.w4(32'hbbcaefac),
	.w5(32'hbbb91a28),
	.w6(32'hbbf1039e),
	.w7(32'hbc477130),
	.w8(32'hbc04addd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2e539),
	.w1(32'hbb31cbc8),
	.w2(32'hbaa4ba9b),
	.w3(32'hba8462c9),
	.w4(32'hbb14e00a),
	.w5(32'hb9bfd853),
	.w6(32'hb9506038),
	.w7(32'hbae2a15e),
	.w8(32'h3a575aa3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26b33c),
	.w1(32'h39137802),
	.w2(32'h35a751af),
	.w3(32'h3a1e8e9f),
	.w4(32'h3983cc9d),
	.w5(32'h3990d6b2),
	.w6(32'hb9ae3a92),
	.w7(32'hb7636a6e),
	.w8(32'hb75c9b3c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99de17c),
	.w1(32'hba0c2826),
	.w2(32'h39b59334),
	.w3(32'hb9398063),
	.w4(32'h39d28670),
	.w5(32'hb903f1d8),
	.w6(32'hba04f476),
	.w7(32'hb9a0b713),
	.w8(32'h390a7cdf),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c73bd8),
	.w1(32'h37ed5e0e),
	.w2(32'h386aa1df),
	.w3(32'hb9224e40),
	.w4(32'h3a2f2197),
	.w5(32'h3a1b0c99),
	.w6(32'h39fbf6b2),
	.w7(32'h39e6a27f),
	.w8(32'h398849ba),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72fca08),
	.w1(32'hb98f0d74),
	.w2(32'h3949316d),
	.w3(32'h39bf8342),
	.w4(32'hb82431fe),
	.w5(32'hb8d0cd73),
	.w6(32'h391df79e),
	.w7(32'h3919a152),
	.w8(32'h392886a2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e47c2),
	.w1(32'hb90ecd14),
	.w2(32'h39fa8e07),
	.w3(32'h39a739e2),
	.w4(32'hb9bfc03d),
	.w5(32'h39717fb8),
	.w6(32'hb8c1dd2e),
	.w7(32'hb927839f),
	.w8(32'h3a39befa),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2ab75),
	.w1(32'h3acc8689),
	.w2(32'h3b220dc0),
	.w3(32'h3908d21d),
	.w4(32'hba50d8c1),
	.w5(32'h3774fade),
	.w6(32'h3aee103f),
	.w7(32'h3ae95500),
	.w8(32'h3b0d6f56),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a9a0b),
	.w1(32'h3935477d),
	.w2(32'hbab4414f),
	.w3(32'hba98384f),
	.w4(32'hbaa4058b),
	.w5(32'hba789ad6),
	.w6(32'h3765bb20),
	.w7(32'hbae698c2),
	.w8(32'h3aaeff27),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a901eeb),
	.w1(32'h3a36e8e4),
	.w2(32'h389f9bc7),
	.w3(32'h3a972ea8),
	.w4(32'h3a10fd5a),
	.w5(32'h37d0551d),
	.w6(32'h3a587667),
	.w7(32'h39a9c6f6),
	.w8(32'h39172140),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b7645d),
	.w1(32'hbb2fb862),
	.w2(32'hba937976),
	.w3(32'hba585549),
	.w4(32'hbaf5bd45),
	.w5(32'hbaa7d408),
	.w6(32'hb8598b8e),
	.w7(32'hba079032),
	.w8(32'hb9e9268e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6fb55),
	.w1(32'h38babf9a),
	.w2(32'h3a638a40),
	.w3(32'hb9b33ca0),
	.w4(32'h3809f2e6),
	.w5(32'h3a85a826),
	.w6(32'hba088f31),
	.w7(32'hb7362530),
	.w8(32'h3a6ae9d3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39560ff3),
	.w1(32'h38f9d946),
	.w2(32'h388b63a6),
	.w3(32'h39b6c83a),
	.w4(32'h3850ba1d),
	.w5(32'hb7d7188f),
	.w6(32'h3835acad),
	.w7(32'hb9aea6b4),
	.w8(32'hb9076e57),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a264d29),
	.w1(32'h3a6d8f62),
	.w2(32'h3802a1df),
	.w3(32'h39b3c387),
	.w4(32'h39f25488),
	.w5(32'h3935465f),
	.w6(32'h38cdb0cc),
	.w7(32'hb8ee42f6),
	.w8(32'hb91518f6),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad5703),
	.w1(32'hb947a35c),
	.w2(32'hb9ab6e68),
	.w3(32'hb96311f8),
	.w4(32'hb98de9f6),
	.w5(32'hb9e94f1c),
	.w6(32'hb9626532),
	.w7(32'hb9f695ea),
	.w8(32'hb9557aaf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997ef26),
	.w1(32'h3656e0c8),
	.w2(32'hba0e27e1),
	.w3(32'h3722abf1),
	.w4(32'hba862fdf),
	.w5(32'hbabe4d08),
	.w6(32'h3a8e536c),
	.w7(32'h39d288f5),
	.w8(32'h3a8f04c9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb28c3),
	.w1(32'hba240ee6),
	.w2(32'h3a0cd3c3),
	.w3(32'hbae44a15),
	.w4(32'hbafd15ca),
	.w5(32'hbabd1dba),
	.w6(32'h38e6be4d),
	.w7(32'h3a3fa09d),
	.w8(32'h3b1abe30),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3950589e),
	.w1(32'hba0b65d1),
	.w2(32'h37a15bc8),
	.w3(32'hba66a2b8),
	.w4(32'hb9f90f71),
	.w5(32'h3a3921c0),
	.w6(32'h3a75b144),
	.w7(32'h3a741c70),
	.w8(32'h3aedecc0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bb37a3),
	.w1(32'h39fa5366),
	.w2(32'h3a7e4f87),
	.w3(32'h397e7d4a),
	.w4(32'h3a31ded3),
	.w5(32'h3a829408),
	.w6(32'h3a623a2a),
	.w7(32'h39c2d958),
	.w8(32'h399e0a71),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11e9a6),
	.w1(32'hb9e28032),
	.w2(32'h3aeb326b),
	.w3(32'hba7a6268),
	.w4(32'hba02c708),
	.w5(32'h3abe1916),
	.w6(32'h3aaf0238),
	.w7(32'h3af6b625),
	.w8(32'h3b52685a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1992e),
	.w1(32'hb8d403f6),
	.w2(32'hb9c58e22),
	.w3(32'h3ab12b89),
	.w4(32'hb89d79ca),
	.w5(32'h391bc076),
	.w6(32'h3a66e642),
	.w7(32'h379404dc),
	.w8(32'h3a10fd7d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1ccd),
	.w1(32'hba7e2994),
	.w2(32'hbaedca47),
	.w3(32'hbb6d5b84),
	.w4(32'hbb363c12),
	.w5(32'hbb4e580d),
	.w6(32'hbb18a10e),
	.w7(32'hbb92e83f),
	.w8(32'hbb208f4a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804c97),
	.w1(32'h3a774e82),
	.w2(32'h3a95a0ea),
	.w3(32'h3a95131d),
	.w4(32'h3a30155c),
	.w5(32'h3a8fc27e),
	.w6(32'h3aa65b53),
	.w7(32'h3aa47303),
	.w8(32'h3aa6e819),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab079db),
	.w1(32'hb7f5b2aa),
	.w2(32'h38b1f016),
	.w3(32'h3a75579b),
	.w4(32'h380054e1),
	.w5(32'hb8f3cd1e),
	.w6(32'h39a3195e),
	.w7(32'h396c3ef8),
	.w8(32'h39c19a7c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9540848),
	.w1(32'h3a25196b),
	.w2(32'h3ab78b20),
	.w3(32'hba4d6f40),
	.w4(32'hb9cca450),
	.w5(32'h3a5705e2),
	.w6(32'h39877812),
	.w7(32'hb53523a8),
	.w8(32'h3ac9387b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3040ee),
	.w1(32'h3b686aee),
	.w2(32'h3b323859),
	.w3(32'h3a95f4a3),
	.w4(32'h3ae19eac),
	.w5(32'h3b0294e0),
	.w6(32'h3b67a236),
	.w7(32'h3b539cb6),
	.w8(32'h3b9a9d1c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a831061),
	.w1(32'hb817d579),
	.w2(32'h3a92e311),
	.w3(32'hb99a24a2),
	.w4(32'hb7afa5b2),
	.w5(32'h3aae4a18),
	.w6(32'h3af67349),
	.w7(32'h3b0128bd),
	.w8(32'h3b34b004),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ab0f5),
	.w1(32'hb68480b5),
	.w2(32'h3a0d597c),
	.w3(32'h3b116f2b),
	.w4(32'h38b00d3b),
	.w5(32'h398a11ef),
	.w6(32'h39527568),
	.w7(32'h3a0c26b0),
	.w8(32'h39f4ae85),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925e3cb),
	.w1(32'hb7f8e30b),
	.w2(32'hb9a9aafb),
	.w3(32'hb9315ec2),
	.w4(32'h38412f9b),
	.w5(32'hb8dfa58b),
	.w6(32'hb77177e1),
	.w7(32'hb9917459),
	.w8(32'h36e50be9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93be840),
	.w1(32'h39b22ff5),
	.w2(32'h39ce763d),
	.w3(32'hb924c816),
	.w4(32'h3978e17e),
	.w5(32'h396a0097),
	.w6(32'h39bddfee),
	.w7(32'h3a04ac58),
	.w8(32'h3a144e86),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac04883),
	.w1(32'h3ac6ba3e),
	.w2(32'h3a65d10c),
	.w3(32'h3a58a8c7),
	.w4(32'h3a9f6174),
	.w5(32'h39ea502b),
	.w6(32'h3a436173),
	.w7(32'h3a8bb5f6),
	.w8(32'hb9b00ddc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40ff3f),
	.w1(32'hba61e39f),
	.w2(32'hbb119a4a),
	.w3(32'hbacfca21),
	.w4(32'hbb7bf58c),
	.w5(32'hbb78db8f),
	.w6(32'hbb12cb0a),
	.w7(32'hbbbf8dd6),
	.w8(32'hbba67952),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e6a48),
	.w1(32'h3b62d5a5),
	.w2(32'h3aedcfb7),
	.w3(32'h3b964999),
	.w4(32'h3b986644),
	.w5(32'h3b29ac67),
	.w6(32'h3b85af61),
	.w7(32'h3b4826fa),
	.w8(32'h39ff6c2c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392754fa),
	.w1(32'hb8a07fe7),
	.w2(32'h3afb6b9d),
	.w3(32'hba07d2b9),
	.w4(32'hba19c02b),
	.w5(32'h3ad159a2),
	.w6(32'h38ba6923),
	.w7(32'h39da5f55),
	.w8(32'h3b051343),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f11fe1),
	.w1(32'hba4794b3),
	.w2(32'h39f09d4e),
	.w3(32'hba74cdf9),
	.w4(32'hbaad02dc),
	.w5(32'h39d0f898),
	.w6(32'hb9630feb),
	.w7(32'hb9e82708),
	.w8(32'h3b09f83d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17d37f),
	.w1(32'hb9bcf03a),
	.w2(32'h38995bfc),
	.w3(32'h3a48c7c3),
	.w4(32'hb8754d46),
	.w5(32'h38558c70),
	.w6(32'hb8e01a77),
	.w7(32'h38c939a9),
	.w8(32'h3973e426),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f6177),
	.w1(32'hbab20ead),
	.w2(32'hbaba4eaf),
	.w3(32'h39b9aab1),
	.w4(32'hbab205d3),
	.w5(32'hba9c19e9),
	.w6(32'hbad57815),
	.w7(32'hba9db949),
	.w8(32'hba99c3cc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa67050),
	.w1(32'h39f846f3),
	.w2(32'h399545ed),
	.w3(32'hba6c373b),
	.w4(32'h39acaabf),
	.w5(32'h387db82e),
	.w6(32'h39ae1c1c),
	.w7(32'h39811434),
	.w8(32'h3a47517e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0885e0),
	.w1(32'hbad91081),
	.w2(32'hba081813),
	.w3(32'h39983a1c),
	.w4(32'hba3d3f40),
	.w5(32'hb9fd538b),
	.w6(32'hbaa2987f),
	.w7(32'hb98b3e6d),
	.w8(32'h384b36f6),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb879ae46),
	.w1(32'h3a19c5f2),
	.w2(32'h3a962443),
	.w3(32'hb9874414),
	.w4(32'h39b00e54),
	.w5(32'h3a6a500c),
	.w6(32'h3a6763b6),
	.w7(32'h3a425a2e),
	.w8(32'h3a5a4e10),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afbe2fd),
	.w1(32'h3a16b75e),
	.w2(32'h3a74d92a),
	.w3(32'h3acf6a58),
	.w4(32'h3a8e44cd),
	.w5(32'h3ab6bd91),
	.w6(32'h3ad9167b),
	.w7(32'h3af972d8),
	.w8(32'h3b399541),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91383b5),
	.w1(32'hba8654a7),
	.w2(32'h3a2e4b30),
	.w3(32'hb9cbb4a2),
	.w4(32'hba98a87e),
	.w5(32'hb85da179),
	.w6(32'h3a9f3073),
	.w7(32'h3aa31042),
	.w8(32'h3b813e09),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1408f0),
	.w1(32'h39a989dd),
	.w2(32'hba815ca9),
	.w3(32'h3a98f645),
	.w4(32'hb92f8f27),
	.w5(32'hbaf28b6e),
	.w6(32'h397aef67),
	.w7(32'hb9bf518f),
	.w8(32'h395c3d4c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94ff96),
	.w1(32'h3b681ce1),
	.w2(32'h3b3becce),
	.w3(32'h3b638c32),
	.w4(32'h3b618ba4),
	.w5(32'h3b1ea300),
	.w6(32'h3b655dcc),
	.w7(32'h3b15bedb),
	.w8(32'h3a482dc8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d0572),
	.w1(32'h3a9a0a6d),
	.w2(32'h3a1d267b),
	.w3(32'h3a741276),
	.w4(32'h3a86c3e0),
	.w5(32'h3a05f0cd),
	.w6(32'h3a98ecb1),
	.w7(32'h3a062001),
	.w8(32'h393a8f14),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d32fc3),
	.w1(32'h39936840),
	.w2(32'h39bee505),
	.w3(32'h39e4f2e3),
	.w4(32'h39856679),
	.w5(32'h39f85efa),
	.w6(32'h394be6d3),
	.w7(32'h399fbf9a),
	.w8(32'h39b91d36),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5eadc),
	.w1(32'h3a5897ff),
	.w2(32'h3925650a),
	.w3(32'h3ab832b6),
	.w4(32'h3a6f15af),
	.w5(32'hb94d374a),
	.w6(32'h3a88e14c),
	.w7(32'h39c6a7c7),
	.w8(32'hb9aa11ac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9350b8b),
	.w1(32'h39628a9f),
	.w2(32'h398065ce),
	.w3(32'hb8d12fa4),
	.w4(32'h3a1fe4ab),
	.w5(32'h39f69dd4),
	.w6(32'h39eb9a03),
	.w7(32'h39b78791),
	.w8(32'h39e05c64),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bb95b),
	.w1(32'hb8eb24e6),
	.w2(32'hba11f2ee),
	.w3(32'h3a0b6d2b),
	.w4(32'hb6c2d59c),
	.w5(32'hb931450e),
	.w6(32'hb7d98a79),
	.w7(32'hb8d55ce1),
	.w8(32'hb7b7cb3a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986be8c),
	.w1(32'h393b0494),
	.w2(32'h39128033),
	.w3(32'hb88c9691),
	.w4(32'h3912e3fc),
	.w5(32'h39842489),
	.w6(32'h39362390),
	.w7(32'h38fea2ef),
	.w8(32'h386e909a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dafc04),
	.w1(32'hba9b5f03),
	.w2(32'hbaa118fe),
	.w3(32'h3915bd89),
	.w4(32'hba3f8305),
	.w5(32'hba9f5971),
	.w6(32'hba4ab76d),
	.w7(32'hba72ffbf),
	.w8(32'hba9785fb),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb180747),
	.w1(32'hba057a8e),
	.w2(32'hba002d78),
	.w3(32'hbb0bd2a0),
	.w4(32'hba4b1990),
	.w5(32'hba11d417),
	.w6(32'hba15ba87),
	.w7(32'hba5437f6),
	.w8(32'hb9bd38e9),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbabca),
	.w1(32'h3ac507f4),
	.w2(32'h3ae8e203),
	.w3(32'h3a4f73e9),
	.w4(32'h3ae77360),
	.w5(32'h3a9af930),
	.w6(32'h3b079727),
	.w7(32'h3afd0b59),
	.w8(32'h3a8f5385),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ccbf87),
	.w1(32'h3a517e40),
	.w2(32'h3a1d14d9),
	.w3(32'hb9db5250),
	.w4(32'h3a5c0a77),
	.w5(32'h3a2bae25),
	.w6(32'h3a0bbc51),
	.w7(32'h39f9ad27),
	.w8(32'h3a1cea32),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d7dd5),
	.w1(32'hba1329ef),
	.w2(32'hba72129a),
	.w3(32'hbaa2fa93),
	.w4(32'hbb005818),
	.w5(32'hbab08b4e),
	.w6(32'h38b2d948),
	.w7(32'hbae01960),
	.w8(32'hbaa9a3d4),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d8666),
	.w1(32'hb9979cfb),
	.w2(32'hb913ccbb),
	.w3(32'hba09e468),
	.w4(32'hb87ec207),
	.w5(32'hb94d31a5),
	.w6(32'hba224092),
	.w7(32'hba14165d),
	.w8(32'hb916d82e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5c4d1),
	.w1(32'h39239fd8),
	.w2(32'h39225f2b),
	.w3(32'hb8f7a204),
	.w4(32'h39007710),
	.w5(32'h399aac7c),
	.w6(32'h3934621b),
	.w7(32'h38a39640),
	.w8(32'hb7707c5d),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ccacf),
	.w1(32'h39c581b6),
	.w2(32'h39bba7f4),
	.w3(32'h39286b93),
	.w4(32'h39388973),
	.w5(32'h397a7867),
	.w6(32'h397f2a35),
	.w7(32'h38f68139),
	.w8(32'h38297caf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d637b),
	.w1(32'h39f34887),
	.w2(32'h39d609e1),
	.w3(32'h391a8697),
	.w4(32'h397a3d4f),
	.w5(32'h39ad1cfc),
	.w6(32'h39b870a5),
	.w7(32'h3955cc61),
	.w8(32'h367769f8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae66ffa),
	.w1(32'hba23417b),
	.w2(32'hb9f5d72e),
	.w3(32'h3ad1de89),
	.w4(32'h3a0bda49),
	.w5(32'h37d5bcc4),
	.w6(32'h396b2815),
	.w7(32'hb893e9c2),
	.w8(32'hb9b7cdc1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba905371),
	.w1(32'hba86fa14),
	.w2(32'hb99f979a),
	.w3(32'hba43917f),
	.w4(32'hba3c05aa),
	.w5(32'hb9d0852c),
	.w6(32'hba1780bd),
	.w7(32'hb99074af),
	.w8(32'h39ce2a12),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16654b),
	.w1(32'h3a338431),
	.w2(32'h38d0571f),
	.w3(32'h3a01366c),
	.w4(32'h39d4a1e2),
	.w5(32'h3980420c),
	.w6(32'h3a16ea0f),
	.w7(32'hb9c22a70),
	.w8(32'hb9b1ca29),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391710b3),
	.w1(32'h39ac6830),
	.w2(32'hb9aabfdc),
	.w3(32'h39d9aa9f),
	.w4(32'h381ca8f5),
	.w5(32'h390df250),
	.w6(32'hb9c9d42b),
	.w7(32'hba75a97b),
	.w8(32'hb9eb6267),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27f05),
	.w1(32'hb91b4df6),
	.w2(32'hb9a0d99c),
	.w3(32'hb7804b09),
	.w4(32'hb997d34d),
	.w5(32'hb9bc4332),
	.w6(32'hb92763a7),
	.w7(32'hb9e13c8d),
	.w8(32'hb9dc1a79),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba910ad5),
	.w1(32'hba439988),
	.w2(32'hbaf16404),
	.w3(32'hba43df68),
	.w4(32'hb7a6bbda),
	.w5(32'hba9019e3),
	.w6(32'hba837393),
	.w7(32'hbaf6215f),
	.w8(32'hba500ca8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994148),
	.w1(32'hb92d6354),
	.w2(32'hb9a631ff),
	.w3(32'hba5a1d2d),
	.w4(32'hb936e5e5),
	.w5(32'h393d544a),
	.w6(32'hba2a2fb1),
	.w7(32'hba3da911),
	.w8(32'hba0f62c4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2defa8),
	.w1(32'h3ab0c500),
	.w2(32'hba466b72),
	.w3(32'h3b0e3c4b),
	.w4(32'h3ac835a4),
	.w5(32'h38afc9b3),
	.w6(32'h3afe1025),
	.w7(32'h3a1b502a),
	.w8(32'h38c73652),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94c1e46),
	.w1(32'h37945763),
	.w2(32'h3817472b),
	.w3(32'hb7e088ea),
	.w4(32'h36adc13f),
	.w5(32'h3786b008),
	.w6(32'hb6fed2b1),
	.w7(32'h37585671),
	.w8(32'hb7ed7568),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36df849d),
	.w1(32'h39d2124c),
	.w2(32'h3aa7d96b),
	.w3(32'hba8a7c8e),
	.w4(32'hba777ac7),
	.w5(32'hba51785d),
	.w6(32'h3842b50c),
	.w7(32'hba3db22f),
	.w8(32'h3a60eae1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule