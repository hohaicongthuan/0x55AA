module layer_10_featuremap_94(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71ee307),
	.w1(32'h36a7b6f3),
	.w2(32'h37638aed),
	.w3(32'hb7b6ee7e),
	.w4(32'h36cec1f1),
	.w5(32'hb63e6a9b),
	.w6(32'hb7a5e196),
	.w7(32'hb5acab65),
	.w8(32'hb7869a67),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf5b81),
	.w1(32'hbab0c3aa),
	.w2(32'hbb22446a),
	.w3(32'h3aef121f),
	.w4(32'hbadde682),
	.w5(32'hbb29e3dc),
	.w6(32'h3b1158de),
	.w7(32'h3914574e),
	.w8(32'hba639dca),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34488916),
	.w1(32'h350b3f05),
	.w2(32'hb6c2904a),
	.w3(32'hb6d17413),
	.w4(32'hb5cc2232),
	.w5(32'hb6f0138b),
	.w6(32'h363d1cc4),
	.w7(32'h366cc46e),
	.w8(32'hb6acb145),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1786c6),
	.w1(32'hba290605),
	.w2(32'hba35080e),
	.w3(32'h3a730244),
	.w4(32'h3a6306a4),
	.w5(32'h3a42c32e),
	.w6(32'h3a0b2aaf),
	.w7(32'h39981901),
	.w8(32'h3a03146b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a2795b),
	.w1(32'h37c8b7e8),
	.w2(32'hb7645120),
	.w3(32'hb682c505),
	.w4(32'h3648d61e),
	.w5(32'hb81c8fa0),
	.w6(32'hb7265b1f),
	.w7(32'h36e5d906),
	.w8(32'hb7bc08d4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372d3ea6),
	.w1(32'h37925f3c),
	.w2(32'hb75c9b8d),
	.w3(32'hb65cb408),
	.w4(32'h3458e96e),
	.w5(32'hb7cfced5),
	.w6(32'hb7599014),
	.w7(32'h363fde1d),
	.w8(32'hb788d2ad),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f42ec),
	.w1(32'h3b6fd3fe),
	.w2(32'h3b8282e4),
	.w3(32'h3b12dd6b),
	.w4(32'h3bcb6a0e),
	.w5(32'h3bb84e19),
	.w6(32'h3a06c80a),
	.w7(32'h3b505b93),
	.w8(32'h3b411308),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b905781),
	.w1(32'h3b5dc88f),
	.w2(32'h3bb297af),
	.w3(32'h3c0ff147),
	.w4(32'h3bebf639),
	.w5(32'h3aed8e02),
	.w6(32'h3b814bae),
	.w7(32'h3c40e309),
	.w8(32'h3ba169cd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900a4e9),
	.w1(32'hb84db9f3),
	.w2(32'h37070fca),
	.w3(32'hb7861361),
	.w4(32'hb8921e21),
	.w5(32'hb8b05d06),
	.w6(32'hb9002598),
	.w7(32'hb8b10006),
	.w8(32'hb8ab9253),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00358e),
	.w1(32'hbae0e801),
	.w2(32'h3b2aa9bd),
	.w3(32'h3a6e2c5d),
	.w4(32'h3acf974f),
	.w5(32'h3b88b352),
	.w6(32'h3ace0df9),
	.w7(32'h3a25c51f),
	.w8(32'h3b20ecc4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d135cd),
	.w1(32'h387aad25),
	.w2(32'h3885ae58),
	.w3(32'h38941677),
	.w4(32'h37091128),
	.w5(32'h3880dcc6),
	.w6(32'h37e2e1d8),
	.w7(32'h376dafbe),
	.w8(32'h380efc80),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f7ddc),
	.w1(32'hba8842e0),
	.w2(32'h3af2e255),
	.w3(32'h3af0554f),
	.w4(32'h3b55bb21),
	.w5(32'h3b923b3f),
	.w6(32'hb910bacd),
	.w7(32'h3b03bf9b),
	.w8(32'h3b050798),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2ca6),
	.w1(32'h39a96a31),
	.w2(32'h3b849cb1),
	.w3(32'h3b228304),
	.w4(32'h3b89bd9f),
	.w5(32'h3bc56ad2),
	.w6(32'h3ab412b8),
	.w7(32'h3ae2b1d3),
	.w8(32'h3b8bc688),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab048eb),
	.w1(32'h390620ef),
	.w2(32'h3a619198),
	.w3(32'hba645ed9),
	.w4(32'hba042f11),
	.w5(32'h3a4f9dd3),
	.w6(32'hbac5d293),
	.w7(32'hb9b70ff8),
	.w8(32'h3a3e4bfa),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b7dfc),
	.w1(32'hbaf0e073),
	.w2(32'hbb13fa99),
	.w3(32'hba8cd3a9),
	.w4(32'hbb3f2282),
	.w5(32'hbb306d6a),
	.w6(32'hb9adc5f3),
	.w7(32'hbaa66b0c),
	.w8(32'hb9c9c429),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38798608),
	.w1(32'hbad1ab3f),
	.w2(32'h3b3ac66a),
	.w3(32'h3ac39a58),
	.w4(32'hba685305),
	.w5(32'h3a81f54f),
	.w6(32'h3bbc812d),
	.w7(32'h3a9a4b64),
	.w8(32'h39cd8140),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f40fb7),
	.w1(32'h38457707),
	.w2(32'h3855efd6),
	.w3(32'h36c8cc95),
	.w4(32'hb78bee65),
	.w5(32'hb664841e),
	.w6(32'h388fb823),
	.w7(32'h3761f863),
	.w8(32'hb7dfeccf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d77fe),
	.w1(32'h3b8fed4c),
	.w2(32'h3bf9f19f),
	.w3(32'h3bf23903),
	.w4(32'h3bd38fa7),
	.w5(32'h3bf40cb0),
	.w6(32'h3b8d52cd),
	.w7(32'h3b7e5980),
	.w8(32'h3b79f95b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d180d),
	.w1(32'h3ae3e726),
	.w2(32'h3b233d9f),
	.w3(32'h3b3dad86),
	.w4(32'h3b5bf09b),
	.w5(32'h3b7480a6),
	.w6(32'h3a9e409a),
	.w7(32'h3ad33e65),
	.w8(32'h3b04c157),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b14434),
	.w1(32'hb895e952),
	.w2(32'h3861adcf),
	.w3(32'h36eec452),
	.w4(32'hb956e3c3),
	.w5(32'hb888bc50),
	.w6(32'h3898c2c9),
	.w7(32'hb836e1bc),
	.w8(32'hb5bc20fd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3847d7f1),
	.w1(32'h38cf31ab),
	.w2(32'h391ec900),
	.w3(32'h3818df75),
	.w4(32'h38874743),
	.w5(32'h3948b809),
	.w6(32'h37fa839f),
	.w7(32'hb82ae2be),
	.w8(32'h385df599),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e5e79),
	.w1(32'hbaaab2e7),
	.w2(32'hba6c3a5d),
	.w3(32'hbb0084c2),
	.w4(32'hba4e6e19),
	.w5(32'h3738dbc6),
	.w6(32'hbacfe00d),
	.w7(32'hba34b3df),
	.w8(32'h39478a63),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b470808),
	.w1(32'h3ada851c),
	.w2(32'h3b82a441),
	.w3(32'h3b889b51),
	.w4(32'h3be30b12),
	.w5(32'h3c0d69d6),
	.w6(32'h3ba952c9),
	.w7(32'h3b2a33e4),
	.w8(32'h3bb55a39),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3948e1),
	.w1(32'hbb34c8e5),
	.w2(32'h3a3e92a8),
	.w3(32'hb9a48e00),
	.w4(32'hba20bc26),
	.w5(32'h3ae2f40c),
	.w6(32'hba2a765e),
	.w7(32'hbab709bf),
	.w8(32'h3ac2a3c6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadfd26),
	.w1(32'hbbb6db7d),
	.w2(32'hbbb72662),
	.w3(32'hbb1362fb),
	.w4(32'hbba52d69),
	.w5(32'hbba6ec11),
	.w6(32'hbab2456d),
	.w7(32'hbb7d5e1e),
	.w8(32'hbb2f285e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ea5190),
	.w1(32'h37a9b4ac),
	.w2(32'hb6664751),
	.w3(32'h358eeec0),
	.w4(32'h369fa8b8),
	.w5(32'hb7a970e3),
	.w6(32'hb72acdc8),
	.w7(32'h37af9ada),
	.w8(32'h3685268c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e66fac),
	.w1(32'h37856a61),
	.w2(32'hb847ada6),
	.w3(32'hb861f026),
	.w4(32'hb7a52549),
	.w5(32'hb8b74286),
	.w6(32'hb81c5d84),
	.w7(32'hb75c042c),
	.w8(32'hb89633e3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfc1cae),
	.w1(32'h3b994403),
	.w2(32'h3c02a457),
	.w3(32'hbc943760),
	.w4(32'h3c14e25a),
	.w5(32'h3c2b2c57),
	.w6(32'hbc968ea0),
	.w7(32'h3c195660),
	.w8(32'h3af251c1),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba058e5c),
	.w1(32'hba13dc43),
	.w2(32'h3a714465),
	.w3(32'hb9e6aac7),
	.w4(32'hba0916f4),
	.w5(32'h3ab9b326),
	.w6(32'hba59ce5c),
	.w7(32'hba40e267),
	.w8(32'h3a3d4db8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc2cd38),
	.w1(32'hbba3eb1e),
	.w2(32'hbb4b84ca),
	.w3(32'hbc51a677),
	.w4(32'h3a2c22d4),
	.w5(32'h3b6af989),
	.w6(32'hbc5ed193),
	.w7(32'hb89f9de0),
	.w8(32'h3b2a949e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb779fb5e),
	.w1(32'hb69c0793),
	.w2(32'hb6a98b83),
	.w3(32'hb7c4af50),
	.w4(32'hb7440c70),
	.w5(32'hb6c5b03a),
	.w6(32'hb7b49b08),
	.w7(32'hb71011e1),
	.w8(32'hb6b80215),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c26d40),
	.w1(32'h36fcf0f6),
	.w2(32'hb7d655cd),
	.w3(32'h366cf97f),
	.w4(32'hb7c1b261),
	.w5(32'hb831b052),
	.w6(32'hb6923b09),
	.w7(32'hb73d2686),
	.w8(32'hb68e7ed2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba413dc7),
	.w1(32'hba4f1d3a),
	.w2(32'h3a76aba2),
	.w3(32'h39ca333a),
	.w4(32'hb5f52576),
	.w5(32'h3aba06ef),
	.w6(32'h39035421),
	.w7(32'h39fddfff),
	.w8(32'h3a93e356),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a52b),
	.w1(32'hbb047464),
	.w2(32'hbaa8f4a4),
	.w3(32'h397a3c79),
	.w4(32'hbaef04de),
	.w5(32'hbac267f4),
	.w6(32'h39c78758),
	.w7(32'hba85b9f4),
	.w8(32'hba209040),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6785ba),
	.w1(32'hb90ba398),
	.w2(32'hba0f29e3),
	.w3(32'hb8aa5d48),
	.w4(32'h3a0aef5c),
	.w5(32'h3a2399f5),
	.w6(32'h3843ec08),
	.w7(32'h3a2fb54a),
	.w8(32'h39631e46),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376e68a6),
	.w1(32'h3af0bbfc),
	.w2(32'h3b2987f9),
	.w3(32'h3af99b7f),
	.w4(32'h3b6a22c2),
	.w5(32'h3b82ed60),
	.w6(32'h39947984),
	.w7(32'h3ad90874),
	.w8(32'h3ab3b933),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c291eba),
	.w1(32'hbbce559a),
	.w2(32'h3ac8a44b),
	.w3(32'h3ac3518c),
	.w4(32'hbc0f287a),
	.w5(32'hb8b4ef8d),
	.w6(32'h3b1ec43e),
	.w7(32'hbc048cdd),
	.w8(32'hbb3ced76),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc534761),
	.w1(32'hbb462766),
	.w2(32'hbacc90d9),
	.w3(32'hbc250964),
	.w4(32'hbb29fd0a),
	.w5(32'h3b040998),
	.w6(32'hbc014ab3),
	.w7(32'hbaa6fabd),
	.w8(32'h3bc1382f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc32359),
	.w1(32'h3ad447ba),
	.w2(32'h3a806afe),
	.w3(32'hbc9345a4),
	.w4(32'h3b9f37f6),
	.w5(32'h3c12c0aa),
	.w6(32'hbc8beff3),
	.w7(32'h3b3db44b),
	.w8(32'h3c1a05bc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d55b38),
	.w1(32'hba9b9d8b),
	.w2(32'hba503764),
	.w3(32'hb9c31a40),
	.w4(32'hba91e1e2),
	.w5(32'hb9953841),
	.w6(32'hb9a34a8f),
	.w7(32'hba57e94c),
	.w8(32'h399dbb47),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38369166),
	.w1(32'h389e8831),
	.w2(32'hb766c715),
	.w3(32'h37b6bbf8),
	.w4(32'h37ab6ae9),
	.w5(32'hb84efa36),
	.w6(32'hb704b812),
	.w7(32'h37d52c88),
	.w8(32'hb855976b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85695de),
	.w1(32'hb7396b61),
	.w2(32'hb842ace3),
	.w3(32'hb8d81514),
	.w4(32'hb899e12c),
	.w5(32'hb9258e3a),
	.w6(32'hb83fe386),
	.w7(32'hb7f579e8),
	.w8(32'hb8ca1f32),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5fb1c),
	.w1(32'hba58572b),
	.w2(32'h3a10bcd6),
	.w3(32'h3a00639d),
	.w4(32'hb9aae6d2),
	.w5(32'h3a959305),
	.w6(32'hb90c2cd0),
	.w7(32'hba00c976),
	.w8(32'h3a08e4c7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3d8f4),
	.w1(32'h3bb6e928),
	.w2(32'h3c0f1a51),
	.w3(32'h3b1b93a5),
	.w4(32'h3c02449e),
	.w5(32'h3c050f82),
	.w6(32'h3b2eb513),
	.w7(32'h3b67484a),
	.w8(32'h3b7bf314),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c9971),
	.w1(32'hbb714534),
	.w2(32'hbae1d10d),
	.w3(32'hbb0831c7),
	.w4(32'hbb1a40d1),
	.w5(32'hba3a9c33),
	.w6(32'hbb05e58a),
	.w7(32'hbadb435a),
	.w8(32'h3936a123),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb314181),
	.w1(32'hbb85964b),
	.w2(32'hbb08acc1),
	.w3(32'h3a43eade),
	.w4(32'hbaa42270),
	.w5(32'hba0d32d7),
	.w6(32'hb7e9f969),
	.w7(32'hbb27a59a),
	.w8(32'hbaf39e54),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb107bf2),
	.w1(32'hbb48f140),
	.w2(32'hba537790),
	.w3(32'hb91515bd),
	.w4(32'hba6da578),
	.w5(32'h3ad9320d),
	.w6(32'hb8be187b),
	.w7(32'h39a97f3e),
	.w8(32'h3a84cb88),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23ee5f),
	.w1(32'h3b19e97b),
	.w2(32'h3be74989),
	.w3(32'h3bbafd54),
	.w4(32'h3be2994a),
	.w5(32'h3c2cba33),
	.w6(32'h3a744e5c),
	.w7(32'h3b469a39),
	.w8(32'h3b9cb4ca),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87ec220),
	.w1(32'h36c60211),
	.w2(32'h35cee9c0),
	.w3(32'hb824606f),
	.w4(32'h36d2c87a),
	.w5(32'hb72ea391),
	.w6(32'hb863de14),
	.w7(32'h37f99db6),
	.w8(32'hb7259541),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb868b1f9),
	.w1(32'hb832aeb2),
	.w2(32'hb749f77e),
	.w3(32'h38e11236),
	.w4(32'h3916d65c),
	.w5(32'h38550834),
	.w6(32'h384808d2),
	.w7(32'h38e65d24),
	.w8(32'h383442ff),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37336526),
	.w1(32'hb61d3c30),
	.w2(32'h378ed958),
	.w3(32'hb821828a),
	.w4(32'h3770c6f8),
	.w5(32'h37f5c495),
	.w6(32'h380f10ba),
	.w7(32'h388c2d89),
	.w8(32'h3839fd13),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0164f9),
	.w1(32'h3a512bd4),
	.w2(32'h3a38adef),
	.w3(32'h39a63932),
	.w4(32'h3aee7fe1),
	.w5(32'h3ad61202),
	.w6(32'h3997ca27),
	.w7(32'h3b02ae40),
	.w8(32'h3a3c6575),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea3652),
	.w1(32'hb9a418a7),
	.w2(32'h3a8e831b),
	.w3(32'h39b163d5),
	.w4(32'h3a10f43d),
	.w5(32'h3a920c03),
	.w6(32'hb91036e9),
	.w7(32'h39bac248),
	.w8(32'h3a598687),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63c6a8),
	.w1(32'h3b7b8678),
	.w2(32'h3bb9a158),
	.w3(32'h3bbb330c),
	.w4(32'h3bbdd7f7),
	.w5(32'h3c0661b9),
	.w6(32'h3b09ad70),
	.w7(32'h3b90db71),
	.w8(32'h3b88b48c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cd20b),
	.w1(32'h3b185a4e),
	.w2(32'h3adb6e5c),
	.w3(32'h3a8a6bb2),
	.w4(32'h3b197671),
	.w5(32'h3aae6244),
	.w6(32'hb9c92ac8),
	.w7(32'h39fc6c0f),
	.w8(32'h3a3cbaa7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d0e39),
	.w1(32'hb9f6305b),
	.w2(32'hba1ef60c),
	.w3(32'hb8a289fb),
	.w4(32'hba28d417),
	.w5(32'hba4adb11),
	.w6(32'h37d96bef),
	.w7(32'hb9eaa04f),
	.w8(32'hb9f5f497),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7989432),
	.w1(32'hb80719e0),
	.w2(32'hb7c950ce),
	.w3(32'hb7751f09),
	.w4(32'hb844e326),
	.w5(32'hb81be98c),
	.w6(32'hb794cec5),
	.w7(32'hb7d0702e),
	.w8(32'hb73b8a28),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a3fa),
	.w1(32'hb93da97f),
	.w2(32'h39865ae0),
	.w3(32'hba167db0),
	.w4(32'h392edf47),
	.w5(32'h3a2309f2),
	.w6(32'hba1db140),
	.w7(32'hb804765e),
	.w8(32'h39e3dfe2),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59b547),
	.w1(32'hba37f34b),
	.w2(32'hb884aa94),
	.w3(32'hb9d8bb6b),
	.w4(32'hb99b42cc),
	.w5(32'h3a0f2c39),
	.w6(32'hba0afcc7),
	.w7(32'hb9057ccc),
	.w8(32'h3a0982fe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba251737),
	.w1(32'h38d142db),
	.w2(32'hba148d52),
	.w3(32'h391c978b),
	.w4(32'h3a4d8977),
	.w5(32'h39a894cb),
	.w6(32'hb94b4c30),
	.w7(32'h3a224044),
	.w8(32'h398906cb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dee3b4),
	.w1(32'h3ac97411),
	.w2(32'h3b3ed740),
	.w3(32'h3ae43b9c),
	.w4(32'h3b1b5cb2),
	.w5(32'h3b60ecb7),
	.w6(32'h3a92748e),
	.w7(32'h39de04d1),
	.w8(32'h3b0e8df5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c2fa7),
	.w1(32'h3ba3af66),
	.w2(32'h3b6c0ee0),
	.w3(32'hba676f1a),
	.w4(32'h3bd0250c),
	.w5(32'h3b22f2be),
	.w6(32'h39c59978),
	.w7(32'h3b70e5ac),
	.w8(32'hb91460f5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787b667),
	.w1(32'h36f98e5f),
	.w2(32'hb7d952a1),
	.w3(32'h375e9550),
	.w4(32'h36810425),
	.w5(32'hb868e854),
	.w6(32'h3791d2a8),
	.w7(32'h37cd19d3),
	.w8(32'hb81a6772),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7935ede),
	.w1(32'h3740cab5),
	.w2(32'hb7e6d85d),
	.w3(32'hb780b064),
	.w4(32'h36e480b5),
	.w5(32'hb7fecfe9),
	.w6(32'hb775b270),
	.w7(32'h3718ec2c),
	.w8(32'hb7ba3e66),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369ecd77),
	.w1(32'h371c2b2d),
	.w2(32'hb786cc4c),
	.w3(32'hb79ee61d),
	.w4(32'hb7aba965),
	.w5(32'hb80be45b),
	.w6(32'hb7aae756),
	.w7(32'hb789b9b1),
	.w8(32'hb80ade96),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b2198b),
	.w1(32'h373ec899),
	.w2(32'hb800522a),
	.w3(32'hb8201850),
	.w4(32'h3369476e),
	.w5(32'hb875f8ec),
	.w6(32'hb7fe83e4),
	.w7(32'h3781b63b),
	.w8(32'hb824f719),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40a413),
	.w1(32'h3a9b53c5),
	.w2(32'h3b9f53dd),
	.w3(32'h3b696efc),
	.w4(32'h3bbf46d0),
	.w5(32'h3bccde95),
	.w6(32'h3bcb1bb2),
	.w7(32'h3be7c877),
	.w8(32'h3b92016a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4efb),
	.w1(32'hbb261d21),
	.w2(32'h396dc93e),
	.w3(32'h3b3cd835),
	.w4(32'h3b01b7d0),
	.w5(32'h3b5e55c2),
	.w6(32'h3aeac6cc),
	.w7(32'h39b86373),
	.w8(32'h3ae47450),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d0b3dd),
	.w1(32'h398ccccd),
	.w2(32'h3bb7e25d),
	.w3(32'h3b3d38bc),
	.w4(32'h3b1ca93e),
	.w5(32'h3ba1df64),
	.w6(32'h3b4f645e),
	.w7(32'hb9bf4a30),
	.w8(32'h3aa5d0b5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc592fa6),
	.w1(32'hbbca3d12),
	.w2(32'hbba12d6b),
	.w3(32'hbbd25dbf),
	.w4(32'hbbab04eb),
	.w5(32'hbb79f394),
	.w6(32'hbb90a650),
	.w7(32'hbb3bca16),
	.w8(32'h398b93e4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c62d9),
	.w1(32'h384ccbf4),
	.w2(32'hb7b6ead9),
	.w3(32'h37d5c2c6),
	.w4(32'h36f0853b),
	.w5(32'hb89455eb),
	.w6(32'h3809fae8),
	.w7(32'h3792c70b),
	.w8(32'hb8609431),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a519d),
	.w1(32'h38386087),
	.w2(32'hb887845a),
	.w3(32'hb7925625),
	.w4(32'hb7464412),
	.w5(32'hb8f9cd02),
	.w6(32'h346b5c00),
	.w7(32'h374ca0a3),
	.w8(32'hb8c57143),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38051e4c),
	.w1(32'h38d22f01),
	.w2(32'hb7d3dcee),
	.w3(32'hb792e75a),
	.w4(32'h38448cf0),
	.w5(32'hb892a2ac),
	.w6(32'h37604ed0),
	.w7(32'h3886ab2a),
	.w8(32'hb88a2de9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a125eba),
	.w1(32'h3a88b68f),
	.w2(32'h3ab649db),
	.w3(32'h3ab57a5d),
	.w4(32'h3ac47a59),
	.w5(32'h3ae273b9),
	.w6(32'h3a994805),
	.w7(32'h3a976a92),
	.w8(32'h3a828968),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d2171c),
	.w1(32'h36e3f06f),
	.w2(32'hb7bb03a3),
	.w3(32'hb7e4bfc9),
	.w4(32'h37bc27ab),
	.w5(32'hb828ff88),
	.w6(32'hb6eefbbc),
	.w7(32'h37bbac06),
	.w8(32'hb827af6d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae931f5),
	.w1(32'h3a640a29),
	.w2(32'h3ac290da),
	.w3(32'h3ada3a38),
	.w4(32'h3b75f2af),
	.w5(32'h3b8370f3),
	.w6(32'h3a8c4cbf),
	.w7(32'h3b48f364),
	.w8(32'h3b0b0a9f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51a007),
	.w1(32'hb871717e),
	.w2(32'h3b376c88),
	.w3(32'h3b057c59),
	.w4(32'h3af0106c),
	.w5(32'h3b804587),
	.w6(32'h3a88841d),
	.w7(32'h3b81e361),
	.w8(32'h3b7ae80f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d7c51),
	.w1(32'hbb08f2fc),
	.w2(32'hbb425422),
	.w3(32'hb94f9d9b),
	.w4(32'hbace25c3),
	.w5(32'hbb0fd346),
	.w6(32'hba9959ac),
	.w7(32'hba109791),
	.w8(32'hba170116),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb985a715),
	.w1(32'hba4117c4),
	.w2(32'h3b0f31db),
	.w3(32'h3a787ade),
	.w4(32'h38fe64c9),
	.w5(32'h3af67796),
	.w6(32'h3ac20c05),
	.w7(32'hb89871fd),
	.w8(32'h3a5f8b82),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85747f),
	.w1(32'hba0abb8f),
	.w2(32'hba55c06c),
	.w3(32'h3aaf079f),
	.w4(32'h3a6d572b),
	.w5(32'h3b10dbc8),
	.w6(32'h3b0e5871),
	.w7(32'h3b6fdcda),
	.w8(32'h3a9fe0f4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8b36b),
	.w1(32'hb9e1c555),
	.w2(32'h3a74897c),
	.w3(32'hba6e5c77),
	.w4(32'hb9d670d0),
	.w5(32'hb992f782),
	.w6(32'hb9d14645),
	.w7(32'hb92c7ef8),
	.w8(32'hb99d7fb6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94eb52),
	.w1(32'h3a4de2f7),
	.w2(32'h3b23dd46),
	.w3(32'h3b0bcbe4),
	.w4(32'h3b39a1a5),
	.w5(32'h3b8045b1),
	.w6(32'h3aa753f5),
	.w7(32'h3a8b771c),
	.w8(32'h3af7b065),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f9a75d),
	.w1(32'h3733d481),
	.w2(32'h352e33ad),
	.w3(32'hb5cb1de0),
	.w4(32'h36d7f875),
	.w5(32'hb6ad78d0),
	.w6(32'h35ed2ede),
	.w7(32'h374ce6ea),
	.w8(32'h360a6258),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3855f772),
	.w1(32'h387da2b3),
	.w2(32'h383526e1),
	.w3(32'h36be1f8c),
	.w4(32'h37003088),
	.w5(32'hb60eb367),
	.w6(32'h38bddf1d),
	.w7(32'h381a5bf6),
	.w8(32'hb7b7cc83),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a47139),
	.w1(32'h36dc5331),
	.w2(32'hb8367726),
	.w3(32'hb80f50da),
	.w4(32'h320f3a3b),
	.w5(32'hb8144841),
	.w6(32'hb792f13d),
	.w7(32'h384abe04),
	.w8(32'hb5b97708),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944e61),
	.w1(32'hb992916b),
	.w2(32'hb8855cbb),
	.w3(32'hba26413c),
	.w4(32'h39090208),
	.w5(32'h3a3f3008),
	.w6(32'hba8066b6),
	.w7(32'h382c3bf4),
	.w8(32'h3a40d097),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983f860),
	.w1(32'hbb0599dc),
	.w2(32'hba7ba6fb),
	.w3(32'h3b0aa113),
	.w4(32'hbb268416),
	.w5(32'hbad3f53a),
	.w6(32'h3b09a87d),
	.w7(32'hbabbb5f7),
	.w8(32'hb9e15205),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f375bc),
	.w1(32'hba4d19fd),
	.w2(32'hb97dbd9c),
	.w3(32'h35ec77fd),
	.w4(32'hb9b4e3e8),
	.w5(32'h39942eb3),
	.w6(32'h37e8109c),
	.w7(32'hb995ef39),
	.w8(32'h3913986b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08ebb0),
	.w1(32'hbb02c439),
	.w2(32'hbb5a330f),
	.w3(32'h3aba03c4),
	.w4(32'hbac13f2a),
	.w5(32'hbb89045f),
	.w6(32'h3a3a803e),
	.w7(32'hbab3f46f),
	.w8(32'hbb33e0d2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a95051f),
	.w1(32'h3affcba3),
	.w2(32'h3b3e04ed),
	.w3(32'h3b4eb4fc),
	.w4(32'h3b55db90),
	.w5(32'h3b91f611),
	.w6(32'h3b3099b3),
	.w7(32'h3b2f137b),
	.w8(32'h3b415a91),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2679a1),
	.w1(32'hba8432db),
	.w2(32'hb8dd7518),
	.w3(32'hbbeffd4a),
	.w4(32'h3b080337),
	.w5(32'h3bace046),
	.w6(32'hbbf0b39b),
	.w7(32'h3a327c7a),
	.w8(32'h3b9b6f05),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db6f9),
	.w1(32'h3984421e),
	.w2(32'h3b38aaba),
	.w3(32'h3b4231a6),
	.w4(32'h3b6c8904),
	.w5(32'h3ba90d0f),
	.w6(32'h3b8e34cf),
	.w7(32'h3b9c0b6e),
	.w8(32'h3b04f481),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50a686),
	.w1(32'hba80ddc9),
	.w2(32'h3a81a63c),
	.w3(32'hb9f2699a),
	.w4(32'h39c5d14d),
	.w5(32'h3b48fe6c),
	.w6(32'hbab49405),
	.w7(32'h39816a08),
	.w8(32'h3b275add),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a0db0),
	.w1(32'hbb247a49),
	.w2(32'h3b5cd797),
	.w3(32'h39cca28a),
	.w4(32'hbae21d77),
	.w5(32'h3a08b1f2),
	.w6(32'h3b678b10),
	.w7(32'h3a65bd38),
	.w8(32'hba3fd86d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba417f2f),
	.w1(32'hbaf0481c),
	.w2(32'hbb3b091d),
	.w3(32'h397db60f),
	.w4(32'hba65d996),
	.w5(32'hbafcc254),
	.w6(32'h3ac851fb),
	.w7(32'h3abbd01f),
	.w8(32'hbaacc9a7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119565),
	.w1(32'hbb23b9d5),
	.w2(32'hbb3ca997),
	.w3(32'hbbc50665),
	.w4(32'hba93771d),
	.w5(32'h3a9ec380),
	.w6(32'hbb9584a0),
	.w7(32'hba59a7df),
	.w8(32'h3b02eaa1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907df8c),
	.w1(32'hb800a222),
	.w2(32'hb75721e8),
	.w3(32'hb749659f),
	.w4(32'h387509ee),
	.w5(32'hb79e83b2),
	.w6(32'hb853eadc),
	.w7(32'hb84ad188),
	.w8(32'hb8c263a8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6fe3a0),
	.w1(32'h39f1ff5b),
	.w2(32'h3b4ace59),
	.w3(32'h3b175950),
	.w4(32'h3b329cc9),
	.w5(32'h3b9585c3),
	.w6(32'h3a9b27e7),
	.w7(32'h3b0a08b9),
	.w8(32'h3b541f66),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a61e2),
	.w1(32'h3a311812),
	.w2(32'h3a429390),
	.w3(32'h3a4f7ad4),
	.w4(32'h3b5e9868),
	.w5(32'h3b814172),
	.w6(32'h3a9352e3),
	.w7(32'h3b860035),
	.w8(32'h3b54743b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c0482),
	.w1(32'hbb4d36fa),
	.w2(32'h3b3ff6d2),
	.w3(32'h3b81db82),
	.w4(32'h39819180),
	.w5(32'h3ba8a352),
	.w6(32'h3bf619ab),
	.w7(32'hbac57f29),
	.w8(32'hb9bd3e1c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfd351),
	.w1(32'hbb2b84ad),
	.w2(32'h3aceb997),
	.w3(32'hbbb3376c),
	.w4(32'hba8d9de3),
	.w5(32'h3b966a7e),
	.w6(32'hbb2c7f37),
	.w7(32'hb8d04e8e),
	.w8(32'h3b8c0c70),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaf92e),
	.w1(32'hbb888736),
	.w2(32'hbb462cf9),
	.w3(32'hba72fcb3),
	.w4(32'hbaf38349),
	.w5(32'hbb3cd429),
	.w6(32'hbac005f5),
	.w7(32'hbb40c317),
	.w8(32'hbad4d101),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f32a6),
	.w1(32'hbb6a08e0),
	.w2(32'h3b181e6f),
	.w3(32'h3a3b0789),
	.w4(32'hba9aa077),
	.w5(32'h3b7345d7),
	.w6(32'h39dd76db),
	.w7(32'hbb4d7001),
	.w8(32'hbab00d3a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c977fd),
	.w1(32'hb92b5562),
	.w2(32'hb91b6274),
	.w3(32'hb9438770),
	.w4(32'hb702be7f),
	.w5(32'h36ba69cd),
	.w6(32'hb93e9678),
	.w7(32'h390b3ac6),
	.w8(32'hb895b6cb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd09b30),
	.w1(32'hbbc4aa99),
	.w2(32'h3b84d650),
	.w3(32'h3ba09679),
	.w4(32'hbb239ee5),
	.w5(32'h3b9d304a),
	.w6(32'h3bb58f5d),
	.w7(32'hbb0981b2),
	.w8(32'hb9080273),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4af950),
	.w1(32'h38f79148),
	.w2(32'h3b6c0300),
	.w3(32'h3a7fc6e9),
	.w4(32'h3b79d8d4),
	.w5(32'h3bbce4c3),
	.w6(32'h39d07920),
	.w7(32'h3b521bcf),
	.w8(32'h3b8affb7),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f55cc),
	.w1(32'h38509bc5),
	.w2(32'h38ddf555),
	.w3(32'hba3bfb7b),
	.w4(32'hb756331f),
	.w5(32'h39183b4f),
	.w6(32'hba38a686),
	.w7(32'hb6851661),
	.w8(32'h3893226c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a458c6),
	.w1(32'hba0811fb),
	.w2(32'hba1fa0d4),
	.w3(32'h3a35a633),
	.w4(32'hb9b9d734),
	.w5(32'hbacf9c66),
	.w6(32'h3adf0e3f),
	.w7(32'h3a27524c),
	.w8(32'hbafcc72c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac09278),
	.w1(32'hb95913c6),
	.w2(32'h3b2c2344),
	.w3(32'h3a204fcb),
	.w4(32'h3b0bc138),
	.w5(32'h3b9217c3),
	.w6(32'h3956f05f),
	.w7(32'h39d0a61c),
	.w8(32'h3b1b163b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94a6e7),
	.w1(32'hbb3e2c62),
	.w2(32'hbac4786a),
	.w3(32'hbaf998b7),
	.w4(32'hba88980a),
	.w5(32'hba1c0cb4),
	.w6(32'hbb0ba08f),
	.w7(32'hbae978b5),
	.w8(32'hba0d40ba),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf2b1b),
	.w1(32'h3afe684f),
	.w2(32'hbaa64eaf),
	.w3(32'hbbc1b9e4),
	.w4(32'h39d6d3d0),
	.w5(32'h38773968),
	.w6(32'hbbf63b4c),
	.w7(32'h3a1474bc),
	.w8(32'h3ab83c9b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f46e8),
	.w1(32'hbb26ff2b),
	.w2(32'hbb281001),
	.w3(32'hbad54744),
	.w4(32'hbb1f6a4a),
	.w5(32'hbb3979fb),
	.w6(32'hbaa23b87),
	.w7(32'hba84dd13),
	.w8(32'hba2780f9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8107f6),
	.w1(32'h39dccd66),
	.w2(32'hbb7da4fd),
	.w3(32'h3b6f4775),
	.w4(32'h3b34f484),
	.w5(32'hbb0fcc06),
	.w6(32'h3a96f93e),
	.w7(32'h39d863be),
	.w8(32'hbb68218c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4438e4),
	.w1(32'hba1a7514),
	.w2(32'h3b0ec182),
	.w3(32'h3b1f3d67),
	.w4(32'hba2d881a),
	.w5(32'hb8a65698),
	.w6(32'h3bc24481),
	.w7(32'h3b3a4ad2),
	.w8(32'hb9052f47),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0c63b),
	.w1(32'hbac87b63),
	.w2(32'hb9daf0a8),
	.w3(32'hb9c7ed65),
	.w4(32'hb9ee61cb),
	.w5(32'h396fc900),
	.w6(32'hba0e1c8c),
	.w7(32'hba337901),
	.w8(32'h399b6940),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dc31fe),
	.w1(32'h38267cb4),
	.w2(32'h37b3c749),
	.w3(32'h3894cb7f),
	.w4(32'h37f4ba98),
	.w5(32'h3618a7a6),
	.w6(32'h3914e4a9),
	.w7(32'h38cb2be5),
	.w8(32'h37f7efd8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c8cd4),
	.w1(32'hb9a022be),
	.w2(32'hba1d0c02),
	.w3(32'h3a26626b),
	.w4(32'hb908f735),
	.w5(32'hba75a2c2),
	.w6(32'h3a87e604),
	.w7(32'h397e6672),
	.w8(32'hba0380d9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a62a06),
	.w1(32'hb8066312),
	.w2(32'hb8160e19),
	.w3(32'h3784c6fa),
	.w4(32'hb71dbf9c),
	.w5(32'hb78aa04d),
	.w6(32'hb71fcd96),
	.w7(32'hb73c94a3),
	.w8(32'hb700b213),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d5c319),
	.w1(32'h381dcef0),
	.w2(32'h352eb8fa),
	.w3(32'h35026376),
	.w4(32'h37a466be),
	.w5(32'hb7c19bee),
	.w6(32'hb60385f8),
	.w7(32'h3788c680),
	.w8(32'hb8211c52),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb246ded),
	.w1(32'hbafb8072),
	.w2(32'hba68b355),
	.w3(32'hba144477),
	.w4(32'hba51258a),
	.w5(32'hba17e122),
	.w6(32'hba5509e8),
	.w7(32'hbab5171d),
	.w8(32'hba0cd2d8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378841fc),
	.w1(32'hb89a778c),
	.w2(32'hb8cbe428),
	.w3(32'h38bfdf09),
	.w4(32'h378e49f0),
	.w5(32'h38f31049),
	.w6(32'hb9327404),
	.w7(32'h383c11f5),
	.w8(32'h397143ff),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ace2b),
	.w1(32'h3a865b7e),
	.w2(32'h3b104e97),
	.w3(32'h3a9a0d91),
	.w4(32'h3b0fc5df),
	.w5(32'h3b4cf0fe),
	.w6(32'h39898564),
	.w7(32'h3a885a38),
	.w8(32'h3acd51bf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc91268),
	.w1(32'hbb2a568e),
	.w2(32'hbb7c0780),
	.w3(32'hbbaf96de),
	.w4(32'hbb367bbd),
	.w5(32'hbb5e87c5),
	.w6(32'hbb86609f),
	.w7(32'hba6fe56a),
	.w8(32'hb94b1c1c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a89905),
	.w1(32'h36d3e2ba),
	.w2(32'hb81cb00f),
	.w3(32'hb8af77c8),
	.w4(32'hb851cfbe),
	.w5(32'hb89ba2bf),
	.w6(32'hb8ac8961),
	.w7(32'hb8551a21),
	.w8(32'hb8ad1c63),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377aa6f8),
	.w1(32'h3782d2b2),
	.w2(32'h3795f695),
	.w3(32'hb74ac759),
	.w4(32'hb6d07b19),
	.w5(32'h36f4328a),
	.w6(32'hb7c7e225),
	.w7(32'hb7450a8e),
	.w8(32'hb57c00a3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ce7d34),
	.w1(32'h366f36a3),
	.w2(32'h367b046c),
	.w3(32'hb72ee1aa),
	.w4(32'hb7287ce5),
	.w5(32'hb707f71d),
	.w6(32'h36680353),
	.w7(32'h36b8cbaa),
	.w8(32'h3693ed1e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c201c4),
	.w1(32'hbaad2df3),
	.w2(32'hbb04c667),
	.w3(32'hb8d6e286),
	.w4(32'hba1bdf85),
	.w5(32'hba1ef992),
	.w6(32'h3ae6ffc5),
	.w7(32'h3b0c2244),
	.w8(32'hb9843d7b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada9bad),
	.w1(32'h3b648bd0),
	.w2(32'h3af0b440),
	.w3(32'h3bc3a87f),
	.w4(32'h3bb839fa),
	.w5(32'h3af20b04),
	.w6(32'hbb0553a3),
	.w7(32'h3b123a6d),
	.w8(32'h3ae1d0b4),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaf32f),
	.w1(32'h3adaef2e),
	.w2(32'h3b62aa08),
	.w3(32'h3b4a5a93),
	.w4(32'h3bf0af99),
	.w5(32'h3b1f66c1),
	.w6(32'hbb840601),
	.w7(32'h3a6d160b),
	.w8(32'hba1af0fb),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4658),
	.w1(32'h3ad9fdd4),
	.w2(32'h3b1a60b1),
	.w3(32'hba8ecb88),
	.w4(32'h3aaa8d08),
	.w5(32'h3afc0400),
	.w6(32'hb82cf9d3),
	.w7(32'h3a52f795),
	.w8(32'h39f87d5f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a48d1),
	.w1(32'h3b761509),
	.w2(32'h3b7d1f2f),
	.w3(32'h3b1bbc17),
	.w4(32'hbaacbb83),
	.w5(32'hbb0ac7ae),
	.w6(32'hb8150aa5),
	.w7(32'h3a2de709),
	.w8(32'h3aa72be3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c2f73),
	.w1(32'hbb36d345),
	.w2(32'hbbf43183),
	.w3(32'hbb486a04),
	.w4(32'hbb2a85dc),
	.w5(32'hba8c9774),
	.w6(32'h38abfe5a),
	.w7(32'h3ad13ed9),
	.w8(32'h3af9f28a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139673),
	.w1(32'hba063e5f),
	.w2(32'h3aff89df),
	.w3(32'hb9a2a5d6),
	.w4(32'hbab73be2),
	.w5(32'hba75a028),
	.w6(32'h3b0a1b4a),
	.w7(32'h3a0cc70f),
	.w8(32'hb93c16a6),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6d8a6),
	.w1(32'h3b1d7210),
	.w2(32'h3a8da43b),
	.w3(32'h398b2214),
	.w4(32'hb9de3bd6),
	.w5(32'hb9f4b150),
	.w6(32'hba9ec202),
	.w7(32'hbb403e39),
	.w8(32'hbba41ec3),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446846),
	.w1(32'h3bab9113),
	.w2(32'h3bf70140),
	.w3(32'h3bb56930),
	.w4(32'h3bfa82e2),
	.w5(32'h3c0bc0f6),
	.w6(32'h3b658e72),
	.w7(32'h3ba84f74),
	.w8(32'h3b9e7e3c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba45a2e7),
	.w1(32'hba984cbf),
	.w2(32'hbaebbee4),
	.w3(32'h39e7d374),
	.w4(32'hbaff8e4d),
	.w5(32'hba1aa161),
	.w6(32'hbb163b12),
	.w7(32'hbb223468),
	.w8(32'hbafd26ad),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af10be0),
	.w1(32'hba56b2c9),
	.w2(32'hba1ba7b8),
	.w3(32'h3aedb101),
	.w4(32'hb8f0ea9c),
	.w5(32'hbabfa769),
	.w6(32'h3b490eba),
	.w7(32'h3a7b6d6f),
	.w8(32'hba9897f9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a960b1c),
	.w1(32'h3b8deb3a),
	.w2(32'h3aa24e9b),
	.w3(32'h3b75b96b),
	.w4(32'h3c0a64f2),
	.w5(32'h3bae60c6),
	.w6(32'hbb887872),
	.w7(32'hbbb3b873),
	.w8(32'hbbaf0f52),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e40b4),
	.w1(32'h3c55ee84),
	.w2(32'h3c348fed),
	.w3(32'h3b370947),
	.w4(32'hbbf0ca46),
	.w5(32'hbc0262e8),
	.w6(32'hba23e21e),
	.w7(32'hbb35ccc4),
	.w8(32'hbb72f21b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c683468),
	.w1(32'hbb38a1fe),
	.w2(32'hba953c9f),
	.w3(32'hbbbe6ce2),
	.w4(32'h3b534941),
	.w5(32'h3bb9c638),
	.w6(32'h3a1d7167),
	.w7(32'h3abc6d6c),
	.w8(32'h3af83377),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23c814),
	.w1(32'hba54ebbd),
	.w2(32'hb9a13ea9),
	.w3(32'h3adfe4e8),
	.w4(32'hba4447d0),
	.w5(32'h397fe891),
	.w6(32'h394a012b),
	.w7(32'h38cbb1da),
	.w8(32'hba6a57cc),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe0401),
	.w1(32'h3b072adf),
	.w2(32'hbae8c470),
	.w3(32'hbc8805cc),
	.w4(32'h3b99b394),
	.w5(32'h3b9e1891),
	.w6(32'hbca6c745),
	.w7(32'h3ab46a37),
	.w8(32'h3b340cdd),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b140e2e),
	.w1(32'hbbb9eb24),
	.w2(32'hbbd312f3),
	.w3(32'h3b586ab8),
	.w4(32'hbb0b8ab5),
	.w5(32'hb99bc8dc),
	.w6(32'h3a1e9754),
	.w7(32'hbb10fa03),
	.w8(32'hbb31a134),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2c47),
	.w1(32'h38a8fbfc),
	.w2(32'hb9795e34),
	.w3(32'h3a851f38),
	.w4(32'h394e7483),
	.w5(32'hb9b91906),
	.w6(32'h38d474ca),
	.w7(32'h3a3a815a),
	.w8(32'h37d0c47d),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8824),
	.w1(32'h3c234a04),
	.w2(32'h3b9c26fb),
	.w3(32'hba4532ec),
	.w4(32'h3badeba4),
	.w5(32'h3a63c4bb),
	.w6(32'h3b89a4e1),
	.w7(32'h3b04d1f0),
	.w8(32'hbad52fd3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ad41c),
	.w1(32'h3b019b42),
	.w2(32'h3b58a532),
	.w3(32'hbb39970b),
	.w4(32'h3b20f048),
	.w5(32'h3b174d00),
	.w6(32'h38e861db),
	.w7(32'hba54ead9),
	.w8(32'h3aa65bc1),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02001a),
	.w1(32'hbad0e6f9),
	.w2(32'hbb74a3b3),
	.w3(32'h3b592d28),
	.w4(32'hbb334066),
	.w5(32'hbb5201c7),
	.w6(32'h3ae19456),
	.w7(32'hbb072a6a),
	.w8(32'hb9b49afb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3030e7),
	.w1(32'hbad07102),
	.w2(32'hb918b525),
	.w3(32'h3a9fa941),
	.w4(32'h3ad3853f),
	.w5(32'h3b3068e9),
	.w6(32'h39c04e64),
	.w7(32'h39a2d602),
	.w8(32'h3acc584e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2b01),
	.w1(32'h3a7d7ee0),
	.w2(32'hb8718e75),
	.w3(32'hb9e61ba1),
	.w4(32'hb9d0de33),
	.w5(32'hb9477095),
	.w6(32'h3b1bba03),
	.w7(32'h3b14902e),
	.w8(32'h3a1fc0d6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a567e0e),
	.w1(32'hbad23cf1),
	.w2(32'hb897ba17),
	.w3(32'h3ad4631b),
	.w4(32'h3b29babc),
	.w5(32'h3b9061d0),
	.w6(32'h3a4ad072),
	.w7(32'h3b950325),
	.w8(32'h3b5f4c49),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1d3ce),
	.w1(32'h39eefffd),
	.w2(32'h3b8b53e8),
	.w3(32'hbb63c968),
	.w4(32'hbb504812),
	.w5(32'h3af147c0),
	.w6(32'h3bd7d236),
	.w7(32'h3c0b543f),
	.w8(32'h3c03eab0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c257e66),
	.w1(32'h3abdeaa8),
	.w2(32'h3b704874),
	.w3(32'h3b5bf7f3),
	.w4(32'h3aecb6f1),
	.w5(32'h3b89b59c),
	.w6(32'h3a8caf07),
	.w7(32'h39858439),
	.w8(32'hbac19669),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91eb88),
	.w1(32'h3b58c067),
	.w2(32'hb96a99a4),
	.w3(32'hbc5981df),
	.w4(32'h3b0c9351),
	.w5(32'h3a8546bd),
	.w6(32'hbc642e70),
	.w7(32'h38bde59c),
	.w8(32'h3b877101),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3dc6b),
	.w1(32'h3b45da5b),
	.w2(32'h3b245721),
	.w3(32'hba3073e8),
	.w4(32'hb9a90ed6),
	.w5(32'hb92d7564),
	.w6(32'h391f1f27),
	.w7(32'hbb3ff976),
	.w8(32'hbbc87ecb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd6ac1),
	.w1(32'hb9b8cdd6),
	.w2(32'hba1cbb26),
	.w3(32'hbb9fa9b5),
	.w4(32'h3a46f52c),
	.w5(32'h39a8a49b),
	.w6(32'h397a798f),
	.w7(32'h3a877609),
	.w8(32'hba4f5f81),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9b61e),
	.w1(32'hbb9b83d8),
	.w2(32'hbba6c1af),
	.w3(32'hbb4e831e),
	.w4(32'hbb7a7886),
	.w5(32'hbb98a2eb),
	.w6(32'hbb879fcf),
	.w7(32'hbb4c6d58),
	.w8(32'hb9c8f90b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfc20a),
	.w1(32'h3b9c85d7),
	.w2(32'h3c2891f6),
	.w3(32'hbb3d5b29),
	.w4(32'hbbf021ed),
	.w5(32'hbb130686),
	.w6(32'hba0dd333),
	.w7(32'h3a777027),
	.w8(32'h3b14f2ff),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cd62c),
	.w1(32'h3b6756a4),
	.w2(32'h3adac335),
	.w3(32'hbb7dd7b1),
	.w4(32'h3b49c9f1),
	.w5(32'h3ad5255e),
	.w6(32'h3b4c736b),
	.w7(32'h3a07399b),
	.w8(32'h3b892d71),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5c4de),
	.w1(32'h3a6f5ed2),
	.w2(32'h3adfcf74),
	.w3(32'h3b163389),
	.w4(32'h3aa7c26a),
	.w5(32'h3ad70f40),
	.w6(32'h3b03530c),
	.w7(32'h3b080980),
	.w8(32'h3a5fdb21),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8f7f4),
	.w1(32'h39f4d8a3),
	.w2(32'h3a817c1e),
	.w3(32'h39aa9a72),
	.w4(32'hb9dabf5d),
	.w5(32'hb8edd0ca),
	.w6(32'h39e6f175),
	.w7(32'h3a33da19),
	.w8(32'hbab0e902),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6686),
	.w1(32'h3b8a6d6e),
	.w2(32'h3ae701bb),
	.w3(32'hb9035ab9),
	.w4(32'h3b829d5c),
	.w5(32'hb922acea),
	.w6(32'h3b577fbc),
	.w7(32'h3b2651f6),
	.w8(32'h3a87e023),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e882f),
	.w1(32'hbad25934),
	.w2(32'h3a5381fe),
	.w3(32'hba3f433b),
	.w4(32'h3ae9d973),
	.w5(32'h3b8ff5cc),
	.w6(32'h3ada700d),
	.w7(32'h3bb38b10),
	.w8(32'hb8b0f83b),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e755f),
	.w1(32'h3b6b4219),
	.w2(32'hba366507),
	.w3(32'hbba284a2),
	.w4(32'h3baaec23),
	.w5(32'h39d70085),
	.w6(32'hbb81eaaf),
	.w7(32'hbb44c3d4),
	.w8(32'hbb0b0ef0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa90730),
	.w1(32'h38cb2dc3),
	.w2(32'h3a49159d),
	.w3(32'h3ae5519d),
	.w4(32'hb9cf7e42),
	.w5(32'hba2f5fcf),
	.w6(32'hb931c3be),
	.w7(32'h3a9d8834),
	.w8(32'hba4be50d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae11088),
	.w1(32'h3b06d09a),
	.w2(32'h3b59aba6),
	.w3(32'h36b70f3d),
	.w4(32'h3b7e12ff),
	.w5(32'h3bb67d4b),
	.w6(32'hb9bed8c5),
	.w7(32'h3a5a3798),
	.w8(32'h3b16d0e8),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393a2081),
	.w1(32'h3b1aa8d9),
	.w2(32'h3b03a8f9),
	.w3(32'h3a969f38),
	.w4(32'h3b17745c),
	.w5(32'h3b0fcaac),
	.w6(32'h3a7b086c),
	.w7(32'h3af1b32e),
	.w8(32'h3a86f263),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f6509),
	.w1(32'h3ab2090d),
	.w2(32'h3b0803fa),
	.w3(32'h3af84ebf),
	.w4(32'hb8ead27b),
	.w5(32'h3a368c4e),
	.w6(32'h38eaa3df),
	.w7(32'h3a536de6),
	.w8(32'hb9e4c09f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba945be7),
	.w1(32'hba1cced2),
	.w2(32'hb9c43c3f),
	.w3(32'hba9b3f91),
	.w4(32'hb9b84578),
	.w5(32'h3a63a6ea),
	.w6(32'hba87eec2),
	.w7(32'hba13065c),
	.w8(32'h399389b2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0191a2),
	.w1(32'hbb274773),
	.w2(32'h3b006f2f),
	.w3(32'h3b07900f),
	.w4(32'h3be45b5d),
	.w5(32'h3c0c316a),
	.w6(32'h3c09632b),
	.w7(32'h3bdebe07),
	.w8(32'h3c2f6a1b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd08f8),
	.w1(32'hb9afdcb4),
	.w2(32'h3a444673),
	.w3(32'h3af5d502),
	.w4(32'hbb523ae5),
	.w5(32'hbae4ecb0),
	.w6(32'hb9aaf3bb),
	.w7(32'h390ace12),
	.w8(32'h3a1166a4),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaefb91),
	.w1(32'hbb3617c0),
	.w2(32'hbb1c8766),
	.w3(32'hbb8a5d72),
	.w4(32'hba9d454b),
	.w5(32'hb9980dd4),
	.w6(32'hbadaa833),
	.w7(32'h38b229b5),
	.w8(32'hbaae92b0),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf45bbd),
	.w1(32'h3b4912a5),
	.w2(32'h3984d8ad),
	.w3(32'hbba4b362),
	.w4(32'h3bc3f24d),
	.w5(32'h3af6680d),
	.w6(32'hbc67cc8b),
	.w7(32'hbc3068c8),
	.w8(32'hbc594853),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b09ad),
	.w1(32'h3b43af37),
	.w2(32'h3b11b20d),
	.w3(32'h3aa1139b),
	.w4(32'h3bc5cdb4),
	.w5(32'h3b5708ac),
	.w6(32'h39394ae7),
	.w7(32'h3aa2a416),
	.w8(32'h3b3939e7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a517d88),
	.w1(32'hbaaf574e),
	.w2(32'h3a1a7b9e),
	.w3(32'h3a7b924c),
	.w4(32'h3a1e201c),
	.w5(32'h3af37fad),
	.w6(32'h3a8f7d79),
	.w7(32'h3a575a20),
	.w8(32'h3b7ae420),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1281f4),
	.w1(32'hba07a237),
	.w2(32'h3ac5c7ce),
	.w3(32'h3b2a8c4f),
	.w4(32'h3b0f999e),
	.w5(32'h3ba94abb),
	.w6(32'h3b6f8955),
	.w7(32'h3adec48f),
	.w8(32'h3b382fcc),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93f466),
	.w1(32'h3c2705e1),
	.w2(32'h3c309f0e),
	.w3(32'h3ab3f5ac),
	.w4(32'hbadc993e),
	.w5(32'h3a36b783),
	.w6(32'h3b62ffee),
	.w7(32'h3bbe688a),
	.w8(32'h3b13f9a9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38ecae),
	.w1(32'hbab397bd),
	.w2(32'hb973691c),
	.w3(32'hbb0c64c1),
	.w4(32'h398a51cd),
	.w5(32'h3a3955bd),
	.w6(32'hba922f30),
	.w7(32'h39e26418),
	.w8(32'hbb604e5b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca523),
	.w1(32'h3a7c5e0a),
	.w2(32'h3ae6e4cc),
	.w3(32'hbaaa1c39),
	.w4(32'hb9f1b45f),
	.w5(32'h39e9bbcf),
	.w6(32'hba9b5c69),
	.w7(32'hba4ea176),
	.w8(32'hbb042530),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ec0c1),
	.w1(32'h3a9d68aa),
	.w2(32'h3b3b42b1),
	.w3(32'h3a1e2b2b),
	.w4(32'h3b0e33c7),
	.w5(32'h3add8a31),
	.w6(32'hbaee33fe),
	.w7(32'hb89afba7),
	.w8(32'hb8b7bb49),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b706f),
	.w1(32'h39fc9dae),
	.w2(32'hbb84d1e6),
	.w3(32'h3aec419b),
	.w4(32'h3ae71a73),
	.w5(32'hbb550b70),
	.w6(32'hbb0265be),
	.w7(32'hbac81a65),
	.w8(32'h399ebf51),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1687b4),
	.w1(32'h3a9b4850),
	.w2(32'h3b57f5fc),
	.w3(32'hb78923d4),
	.w4(32'h391390e4),
	.w5(32'h3b137eca),
	.w6(32'h3b53a9e5),
	.w7(32'h3a935767),
	.w8(32'hbb192dbc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffff49),
	.w1(32'h38183aa6),
	.w2(32'h3b00610b),
	.w3(32'hba843550),
	.w4(32'h39641183),
	.w5(32'h39e339f9),
	.w6(32'h3aa64b5d),
	.w7(32'h3a9401e6),
	.w8(32'hba6eb920),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4b543),
	.w1(32'h3a14ed7a),
	.w2(32'hbaad4396),
	.w3(32'h39d34639),
	.w4(32'h3aed4ba5),
	.w5(32'hb8a4e1b4),
	.w6(32'h3ac90748),
	.w7(32'h3a8c3a6d),
	.w8(32'hbb5e3fd9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0436fd),
	.w1(32'hbb1e2a9d),
	.w2(32'h3ace7880),
	.w3(32'hbbabda89),
	.w4(32'h3b24bf88),
	.w5(32'h3b71a095),
	.w6(32'h3b6d930b),
	.w7(32'h3c065465),
	.w8(32'h3bb585d3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab813fc),
	.w1(32'hbb846281),
	.w2(32'h3aada87a),
	.w3(32'h3b6efdd6),
	.w4(32'hbb14b447),
	.w5(32'h3b176eed),
	.w6(32'h3b8f5a59),
	.w7(32'h3a07d3bb),
	.w8(32'h39a5fc56),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b757fef),
	.w1(32'h3b05305d),
	.w2(32'h3bb70682),
	.w3(32'h3b9b1ba4),
	.w4(32'h3b1929a5),
	.w5(32'h3b73d002),
	.w6(32'h3b02d2f0),
	.w7(32'h3ae1975c),
	.w8(32'h3b42d31f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31e62c),
	.w1(32'h3aeec8a9),
	.w2(32'h3a2f9b5a),
	.w3(32'h3acd462d),
	.w4(32'h3abc689e),
	.w5(32'h3a26fdc2),
	.w6(32'h38daf253),
	.w7(32'h39e311bd),
	.w8(32'h3a017669),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f64d5),
	.w1(32'h3b96a607),
	.w2(32'h3c253eaf),
	.w3(32'h3c1bc4c3),
	.w4(32'h3bf328ac),
	.w5(32'h3c292e23),
	.w6(32'h3b80f9d5),
	.w7(32'h3ab1bddd),
	.w8(32'h3b9be9a0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc407e80),
	.w1(32'hba2adb72),
	.w2(32'hba6ed063),
	.w3(32'hbc07baef),
	.w4(32'h39df685e),
	.w5(32'hbaaca228),
	.w6(32'hbbe7f172),
	.w7(32'h3ad8fa80),
	.w8(32'hbae0499f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98117e2),
	.w1(32'h3a91ba04),
	.w2(32'h3aaf4637),
	.w3(32'hb9997b91),
	.w4(32'h3aeda92b),
	.w5(32'h3a9b0b7e),
	.w6(32'hb94f92be),
	.w7(32'h3b0933c4),
	.w8(32'h3a6c6bf8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7b625),
	.w1(32'h3b637dfb),
	.w2(32'hb9f79877),
	.w3(32'h39c32a5d),
	.w4(32'h3b6213db),
	.w5(32'hbac24a44),
	.w6(32'h3b72380f),
	.w7(32'h3ad29dc7),
	.w8(32'h3a0c85b0),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78a193),
	.w1(32'h3ae2e0c3),
	.w2(32'hba0c2aca),
	.w3(32'hb9c8e320),
	.w4(32'h3b4e32bf),
	.w5(32'h397c4247),
	.w6(32'hbbf48f9b),
	.w7(32'hbc0176b0),
	.w8(32'hbc06cbbd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbb742),
	.w1(32'hbaf2efa2),
	.w2(32'hbb3689a6),
	.w3(32'h39750960),
	.w4(32'hbb10a10c),
	.w5(32'hbafdf5ea),
	.w6(32'hbb1537a7),
	.w7(32'hbb169c37),
	.w8(32'hba4b9086),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865f0b3),
	.w1(32'h3ae353cc),
	.w2(32'h3b0cfe17),
	.w3(32'h39a8c90d),
	.w4(32'h3b120eb7),
	.w5(32'h3ac19c3b),
	.w6(32'h3ae34dfd),
	.w7(32'h3b63c702),
	.w8(32'h3b1860d2),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a4280),
	.w1(32'hba5116f0),
	.w2(32'h3b43e94a),
	.w3(32'h3901165e),
	.w4(32'h3b866618),
	.w5(32'h3bbae10c),
	.w6(32'h3b8d9ecf),
	.w7(32'h3ba76950),
	.w8(32'h3bfca66e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a2670),
	.w1(32'hbb755a3d),
	.w2(32'h3b0f5484),
	.w3(32'h3bd2c0eb),
	.w4(32'hbb4acc3d),
	.w5(32'h3b26ef8e),
	.w6(32'h3c2ec92d),
	.w7(32'h3c476c0a),
	.w8(32'h3c0c6529),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4ef73),
	.w1(32'h3adac6b1),
	.w2(32'h3abd93b8),
	.w3(32'h3b53fabc),
	.w4(32'h37d20731),
	.w5(32'h3a81d731),
	.w6(32'h394b6fdd),
	.w7(32'h3aa69b56),
	.w8(32'h371bb478),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c943),
	.w1(32'h396c8b8c),
	.w2(32'h3b2ad9ab),
	.w3(32'h3ae8bede),
	.w4(32'h3ad296c1),
	.w5(32'h3b52c922),
	.w6(32'hba754aaf),
	.w7(32'hbb151f16),
	.w8(32'h395c52d6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29b212),
	.w1(32'h3b309d76),
	.w2(32'h3b4cdd56),
	.w3(32'h3a98e52c),
	.w4(32'h3b2511a8),
	.w5(32'h3b2e1627),
	.w6(32'h3abd8a01),
	.w7(32'h3a1083c6),
	.w8(32'h3a7eb80f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f08b0),
	.w1(32'h3a082e3f),
	.w2(32'h3adb4182),
	.w3(32'h3aabc64b),
	.w4(32'hb9f268a5),
	.w5(32'h3a2d9996),
	.w6(32'h3918d3d9),
	.w7(32'h3a72dace),
	.w8(32'hba75feb4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2718),
	.w1(32'h3a15e016),
	.w2(32'h3b93cc4f),
	.w3(32'h3a4a5aac),
	.w4(32'hba639181),
	.w5(32'h3ac761a8),
	.w6(32'h3aca1153),
	.w7(32'h390eb8dd),
	.w8(32'hb9faffa2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aded219),
	.w1(32'h3b1982f9),
	.w2(32'h3b31fc3c),
	.w3(32'h3a31f9c1),
	.w4(32'hba05ec0a),
	.w5(32'hb95f0248),
	.w6(32'hb972c38c),
	.w7(32'h3a2f5845),
	.w8(32'hbabc90db),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83252d7),
	.w1(32'hb9da80ef),
	.w2(32'h3afe00d8),
	.w3(32'hba9b1b97),
	.w4(32'hb9218bbf),
	.w5(32'h3a87c050),
	.w6(32'hbadeb7eb),
	.w7(32'hba130ea0),
	.w8(32'h3b0d226b),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd9fa9),
	.w1(32'hbb8f0b8f),
	.w2(32'hbb90774d),
	.w3(32'hbb19bbe0),
	.w4(32'hb9ffb964),
	.w5(32'hbb1f443e),
	.w6(32'h39b268f4),
	.w7(32'hbb2c8ad8),
	.w8(32'hbb7cd53b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf56c3c),
	.w1(32'hba07d1e4),
	.w2(32'h39e920b0),
	.w3(32'hbbafc520),
	.w4(32'hba2ebdaf),
	.w5(32'h3a5f3e76),
	.w6(32'hbb978c8e),
	.w7(32'hbbabdd0c),
	.w8(32'hbb99556a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab59a5c),
	.w1(32'h3a674a84),
	.w2(32'h39b4d7fe),
	.w3(32'h3a842e23),
	.w4(32'h3a9533fa),
	.w5(32'hb802a385),
	.w6(32'h3a931c58),
	.w7(32'h3a8498d3),
	.w8(32'h3b6ff02c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f7171),
	.w1(32'h3baf2a8b),
	.w2(32'h3a3f997a),
	.w3(32'hbaacf907),
	.w4(32'h3b4ecfcb),
	.w5(32'hb74bda9d),
	.w6(32'h3a735645),
	.w7(32'h3b0a181a),
	.w8(32'hbb575d72),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bcfb7),
	.w1(32'hb9dc20cb),
	.w2(32'h3aacf456),
	.w3(32'hbb8aec46),
	.w4(32'hb979367e),
	.w5(32'h3aa2810d),
	.w6(32'h3b65cac5),
	.w7(32'h3b49565d),
	.w8(32'h3a76a665),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9888cee),
	.w1(32'hbbf47178),
	.w2(32'h3b57a028),
	.w3(32'h3b1e1429),
	.w4(32'h3972b3b5),
	.w5(32'h3bf48369),
	.w6(32'h3c1ae2f0),
	.w7(32'h3c6d1054),
	.w8(32'h3c5353d1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0fbd0),
	.w1(32'h3ad9437e),
	.w2(32'h3ac53715),
	.w3(32'h3b7e39e6),
	.w4(32'h3a3801de),
	.w5(32'hb9b59427),
	.w6(32'h3a2a16d8),
	.w7(32'h3a99359c),
	.w8(32'h3b01c1e8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08423f),
	.w1(32'h3bbd91c7),
	.w2(32'h3bb25bd7),
	.w3(32'h3a06c084),
	.w4(32'h3918e0be),
	.w5(32'h3a2511a1),
	.w6(32'h3aaede64),
	.w7(32'h3b466b22),
	.w8(32'h3a925e74),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b537382),
	.w1(32'hba8e324a),
	.w2(32'h3a815af3),
	.w3(32'hb9d59926),
	.w4(32'h3b06d13e),
	.w5(32'h3b49e454),
	.w6(32'h3a1749ce),
	.w7(32'hb9db1422),
	.w8(32'h38f8bb72),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4bca3),
	.w1(32'h3a064b51),
	.w2(32'h3c2065ff),
	.w3(32'h3b1a2b33),
	.w4(32'hbb079486),
	.w5(32'h3c12ba57),
	.w6(32'h3ba5b10d),
	.w7(32'h3c55dfa8),
	.w8(32'h3c357138),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14764d),
	.w1(32'hbacfdb10),
	.w2(32'h3ae58959),
	.w3(32'h3b6a8946),
	.w4(32'h39df462c),
	.w5(32'h3a1a279d),
	.w6(32'h3b31d901),
	.w7(32'h3b079074),
	.w8(32'h3b191850),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc7260),
	.w1(32'hbacd4c22),
	.w2(32'hbb19c60b),
	.w3(32'h3bdb8364),
	.w4(32'h3b639af0),
	.w5(32'h3ae57108),
	.w6(32'hba7b78af),
	.w7(32'h3b0274ba),
	.w8(32'hba4876e4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ddb54),
	.w1(32'h3acd57e5),
	.w2(32'h3b156c10),
	.w3(32'h3a4e8186),
	.w4(32'hb98d09ee),
	.w5(32'h3a45e146),
	.w6(32'h3ac08d02),
	.w7(32'h3b0169d7),
	.w8(32'h3a3fe95c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d220),
	.w1(32'hb9487c41),
	.w2(32'hba4f8164),
	.w3(32'h3a330277),
	.w4(32'h3a99360b),
	.w5(32'h396075bc),
	.w6(32'h3b1c1786),
	.w7(32'h3aeafdf6),
	.w8(32'hbb0b510e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f9028),
	.w1(32'h3b880e32),
	.w2(32'h3ba30cde),
	.w3(32'h3ac5a7a3),
	.w4(32'h3bcb317a),
	.w5(32'h3bf818dd),
	.w6(32'h3ba1e083),
	.w7(32'h3bd0a041),
	.w8(32'h3b9f0f52),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0086),
	.w1(32'h3bd1bf66),
	.w2(32'h3c0fd2ce),
	.w3(32'h3b9d3841),
	.w4(32'h3b6a8393),
	.w5(32'h3ba7cbd0),
	.w6(32'h3b1cbbb6),
	.w7(32'h3b156ba0),
	.w8(32'h3b7d0289),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053d2e),
	.w1(32'h380661b1),
	.w2(32'h3b96950f),
	.w3(32'h3afa550e),
	.w4(32'h3bbe8927),
	.w5(32'h3bf7db70),
	.w6(32'h3a9c0af6),
	.w7(32'hbaa93e80),
	.w8(32'hba0046c7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe11723),
	.w1(32'hb9c241e7),
	.w2(32'hba9c215b),
	.w3(32'hbb3a750c),
	.w4(32'h3a040f15),
	.w5(32'h3a8d851d),
	.w6(32'hbb12c952),
	.w7(32'h39aa6cd1),
	.w8(32'h3ae31411),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bee4),
	.w1(32'hbc4aeb85),
	.w2(32'hba54a5ad),
	.w3(32'hbb8daf29),
	.w4(32'hbbcaf185),
	.w5(32'h3b016139),
	.w6(32'h3b39fd2c),
	.w7(32'h3c31983b),
	.w8(32'h3c25bdad),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2340ef),
	.w1(32'h3b136b37),
	.w2(32'h3b3bcbf4),
	.w3(32'h3b24e9c3),
	.w4(32'hba9e41e7),
	.w5(32'hb9cc96bc),
	.w6(32'hba9773db),
	.w7(32'hb83dfa84),
	.w8(32'hba4f1cb9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa53a1),
	.w1(32'hbabe9529),
	.w2(32'hba6456b9),
	.w3(32'hba8c07af),
	.w4(32'hba394ace),
	.w5(32'hbab45030),
	.w6(32'hbb07b6cf),
	.w7(32'hbb38c719),
	.w8(32'hbb4f465e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4c9a5),
	.w1(32'hbb734a93),
	.w2(32'h38091e6c),
	.w3(32'h3a8dd98c),
	.w4(32'hbb0bcf28),
	.w5(32'h3b0eeab5),
	.w6(32'h3abb9ef5),
	.w7(32'h3ba99ef0),
	.w8(32'h3b07d88a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94972af),
	.w1(32'h3b1156ad),
	.w2(32'h3a53f021),
	.w3(32'hbaeaf755),
	.w4(32'hba7d1832),
	.w5(32'hbb1ec22c),
	.w6(32'h3a2fd0d0),
	.w7(32'hb74bbbc6),
	.w8(32'hba14ce17),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395bc1f3),
	.w1(32'h38607a1b),
	.w2(32'h3aa80510),
	.w3(32'h3a3f4672),
	.w4(32'h3a745f41),
	.w5(32'h3a90df1d),
	.w6(32'h3856bc3b),
	.w7(32'h3b1a41b9),
	.w8(32'h3b4fa2f3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a66fff8),
	.w1(32'h3ad24733),
	.w2(32'h3b399329),
	.w3(32'h3a9e1fb2),
	.w4(32'h3a30926f),
	.w5(32'h3af797bf),
	.w6(32'hb96747c4),
	.w7(32'h3a7f2ba3),
	.w8(32'h3a51b86b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0428f9),
	.w1(32'hb880f530),
	.w2(32'h3acdc430),
	.w3(32'hba48151e),
	.w4(32'hb96dabe9),
	.w5(32'h3b35cce2),
	.w6(32'h3a8be829),
	.w7(32'h3b14ffa0),
	.w8(32'hbb1890b3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb287e50),
	.w1(32'hbacb4656),
	.w2(32'hbb576cfd),
	.w3(32'hbafb7db1),
	.w4(32'h3aae55b4),
	.w5(32'h3ad4390e),
	.w6(32'h3af81ac2),
	.w7(32'hba0f777f),
	.w8(32'h3a6cc534),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0e617),
	.w1(32'h3a801a91),
	.w2(32'h3c0597dd),
	.w3(32'h3b978b74),
	.w4(32'h3b140ee6),
	.w5(32'h3c11ec66),
	.w6(32'hbb1d9981),
	.w7(32'hbbdb33af),
	.w8(32'hbbdfd16a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b737c58),
	.w1(32'h3b0239f4),
	.w2(32'h3b32a310),
	.w3(32'h3b668ed9),
	.w4(32'h3a74f9b7),
	.w5(32'h3b1f01fd),
	.w6(32'h3b1d556a),
	.w7(32'h3b3f39ae),
	.w8(32'h3a98538b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff2395),
	.w1(32'h3acc08ca),
	.w2(32'h3a915b8b),
	.w3(32'h3a6b1f21),
	.w4(32'h3a0081db),
	.w5(32'h39b9ed0e),
	.w6(32'hbb4954a4),
	.w7(32'hbb60eb45),
	.w8(32'hbb8dbb61),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02dad5),
	.w1(32'h3af508ff),
	.w2(32'h3ab92c07),
	.w3(32'h3b147d53),
	.w4(32'h3b4ee20a),
	.w5(32'h3b2f18cc),
	.w6(32'h3ac5b90d),
	.w7(32'h3b40c84f),
	.w8(32'h3adae154),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04b69e),
	.w1(32'h3b4d8298),
	.w2(32'h3b460c19),
	.w3(32'hba7163b5),
	.w4(32'hbac50915),
	.w5(32'hbac62a65),
	.w6(32'hba8e5df9),
	.w7(32'hb6bb110d),
	.w8(32'h3a1fda39),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b748832),
	.w1(32'h3b957549),
	.w2(32'h3b74b54a),
	.w3(32'hbadf9f3a),
	.w4(32'hba4211ff),
	.w5(32'hb9c37437),
	.w6(32'h3ab934d1),
	.w7(32'h3a9313da),
	.w8(32'hb9f32db4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2bbdb),
	.w1(32'h3ac31b06),
	.w2(32'h3a835ac6),
	.w3(32'hb91aa2bb),
	.w4(32'h3a25e5ad),
	.w5(32'h3a0d4c48),
	.w6(32'hbb3bd73b),
	.w7(32'hbb540c5d),
	.w8(32'hbb8b3155),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8b722),
	.w1(32'h3a2603a8),
	.w2(32'h3b420fae),
	.w3(32'h3a715bb3),
	.w4(32'h3ae26403),
	.w5(32'h3af8bef0),
	.w6(32'hba71da2d),
	.w7(32'h3a83ed47),
	.w8(32'h3a9d5f7b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06efb1),
	.w1(32'hba319cdd),
	.w2(32'hb97fd3e4),
	.w3(32'h3aadd52a),
	.w4(32'h372421c7),
	.w5(32'h3a11d7d6),
	.w6(32'hba23c290),
	.w7(32'h3ab73d12),
	.w8(32'h3adad9ac),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba0a27),
	.w1(32'hb90d5bcd),
	.w2(32'h3b602a75),
	.w3(32'h3aaae2a0),
	.w4(32'h3b9034c9),
	.w5(32'h3a826273),
	.w6(32'h3b1108ea),
	.w7(32'h3b5e262f),
	.w8(32'h3b53c33b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998ba1e),
	.w1(32'h3b5997e7),
	.w2(32'h3baa00b9),
	.w3(32'h3b3a5ab4),
	.w4(32'h3af804c3),
	.w5(32'h3b822c0a),
	.w6(32'h3a16179f),
	.w7(32'h3b2673b3),
	.w8(32'h3b4d5443),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855405),
	.w1(32'h3a9e2feb),
	.w2(32'h3b36da60),
	.w3(32'h3ae78256),
	.w4(32'h3b8561e6),
	.w5(32'h3b2f2dce),
	.w6(32'hb87eb60a),
	.w7(32'h3a86f01b),
	.w8(32'h3a801b08),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ad8c87),
	.w1(32'hba56a7e9),
	.w2(32'hba9e2ca2),
	.w3(32'hba919ccb),
	.w4(32'hba2a0dc8),
	.w5(32'hbab9552e),
	.w6(32'h3a445865),
	.w7(32'h3a5f727d),
	.w8(32'hbaac5ee0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718b87),
	.w1(32'h3b0f1c9a),
	.w2(32'h3aae5d78),
	.w3(32'hbb157a70),
	.w4(32'h3a5942cf),
	.w5(32'h39dbf23c),
	.w6(32'hbb8ee577),
	.w7(32'hbb99c3ae),
	.w8(32'hbbcdb729),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07349e),
	.w1(32'h3aace8d1),
	.w2(32'h3a8ff71e),
	.w3(32'h3ab573ef),
	.w4(32'h3925bf21),
	.w5(32'h398be52e),
	.w6(32'hbabca61d),
	.w7(32'hbb0818ba),
	.w8(32'hbb3db4a7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9427a1),
	.w1(32'h3af3cb34),
	.w2(32'h3aa0d064),
	.w3(32'h3a0a713a),
	.w4(32'h393f3ac7),
	.w5(32'h38bd09a8),
	.w6(32'hbb152053),
	.w7(32'hbb480caa),
	.w8(32'hbb7a0a2f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf80f6),
	.w1(32'hb9a60ca7),
	.w2(32'h3a112333),
	.w3(32'h39f757c4),
	.w4(32'h39786edb),
	.w5(32'h3aa12e7e),
	.w6(32'hba05a943),
	.w7(32'h3974deb6),
	.w8(32'hb97973a4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a1d3e),
	.w1(32'hbaa5bd37),
	.w2(32'hbabac783),
	.w3(32'hbaa8280b),
	.w4(32'hbb15f507),
	.w5(32'hba975f38),
	.w6(32'h39d93271),
	.w7(32'h3ab0e27d),
	.w8(32'h38296e5b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba620cf4),
	.w1(32'hbaa34ec1),
	.w2(32'h3a9e3c31),
	.w3(32'hbac681a8),
	.w4(32'hba77f739),
	.w5(32'h3adb8bce),
	.w6(32'hbacf0f05),
	.w7(32'hb89f641a),
	.w8(32'hba6944c7),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38943bf4),
	.w1(32'h39635800),
	.w2(32'h3b220375),
	.w3(32'h3a5ae6a6),
	.w4(32'h3a6d6d70),
	.w5(32'h3b09e63a),
	.w6(32'hba95171e),
	.w7(32'h38d4f8d7),
	.w8(32'hb7b1675d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cb0c5),
	.w1(32'h3a879b1b),
	.w2(32'h3ac05edf),
	.w3(32'hba9b6b22),
	.w4(32'hb8f5e6dd),
	.w5(32'h3a06f384),
	.w6(32'hba691d38),
	.w7(32'hba0d121f),
	.w8(32'hbada14f8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96951c),
	.w1(32'hbb4c4669),
	.w2(32'hbb9e3056),
	.w3(32'h3a827222),
	.w4(32'h3babd43d),
	.w5(32'h3b07f680),
	.w6(32'h3996f9ae),
	.w7(32'h3a637d88),
	.w8(32'h3a92be63),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04c3b9),
	.w1(32'h3b301a23),
	.w2(32'h3b6824f5),
	.w3(32'h3a88ccb0),
	.w4(32'hba0963a2),
	.w5(32'h39bc3d97),
	.w6(32'hba4597c9),
	.w7(32'hba2832c0),
	.w8(32'hbb73b649),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72b7b1),
	.w1(32'h3ba5039b),
	.w2(32'h3c04712a),
	.w3(32'hba2630f1),
	.w4(32'h3a93fa49),
	.w5(32'h3a38c334),
	.w6(32'h3baa88e5),
	.w7(32'h3b985b8a),
	.w8(32'hbb9a03ef),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d668d),
	.w1(32'h3a949936),
	.w2(32'hb9c549d5),
	.w3(32'h3a0e123b),
	.w4(32'h3ab02e80),
	.w5(32'h39758523),
	.w6(32'h3aa2d97b),
	.w7(32'hb923629f),
	.w8(32'hb9718d33),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b79c1d),
	.w1(32'hbb0f8392),
	.w2(32'hbb7d5a0c),
	.w3(32'h3b2c6c2a),
	.w4(32'hb95e457b),
	.w5(32'hbb44a9ca),
	.w6(32'h3b170be0),
	.w7(32'hbb6f4c4d),
	.w8(32'hbb61df5b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule