module layer_10_featuremap_499(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840b81),
	.w1(32'h3afcc8d0),
	.w2(32'h3a07a59e),
	.w3(32'hba8993b2),
	.w4(32'h3c696dc4),
	.w5(32'h3b269369),
	.w6(32'h3c690f27),
	.w7(32'h3b75764a),
	.w8(32'h3b5d7a39),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb940386),
	.w1(32'h3ac9d89f),
	.w2(32'hb998c533),
	.w3(32'hbc147e7a),
	.w4(32'h3bb8c90e),
	.w5(32'h3bd453f6),
	.w6(32'hbc016a52),
	.w7(32'hba9e1e93),
	.w8(32'h3baf1e10),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b7e75),
	.w1(32'h3abeaba2),
	.w2(32'hbbcec101),
	.w3(32'h3b429de1),
	.w4(32'h3b790166),
	.w5(32'h390a0967),
	.w6(32'h3bc6c6b8),
	.w7(32'hbc05ae87),
	.w8(32'h3b37b33f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa3a78),
	.w1(32'hbb7a4a33),
	.w2(32'h3be25ba4),
	.w3(32'hbc374947),
	.w4(32'hbbdf46a5),
	.w5(32'h3ce9da9d),
	.w6(32'hbac0fd6f),
	.w7(32'h3b4905f6),
	.w8(32'hbb528f12),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49b2ed),
	.w1(32'hbbe4dcec),
	.w2(32'hbc266a07),
	.w3(32'h3b8dafb0),
	.w4(32'hbbf6e2a3),
	.w5(32'hbc8490d8),
	.w6(32'hbbac31b5),
	.w7(32'h3b9c5d3f),
	.w8(32'hbc15e59b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb932306),
	.w1(32'hbb6e203f),
	.w2(32'h3b56ddc9),
	.w3(32'hbc22a061),
	.w4(32'hbc6ce34f),
	.w5(32'hbc193618),
	.w6(32'hbbfb3509),
	.w7(32'hba803b30),
	.w8(32'hbb105b2e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc31501),
	.w1(32'h3c3903ee),
	.w2(32'hb899c6d0),
	.w3(32'h3bc1b1a5),
	.w4(32'h3a9c6a00),
	.w5(32'hbbf92b8e),
	.w6(32'h3b11005e),
	.w7(32'hbb0df88f),
	.w8(32'hb9c7df21),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92fb18),
	.w1(32'h3c00e6cf),
	.w2(32'hbb7d6a3a),
	.w3(32'hbbe3145e),
	.w4(32'h3b1ab172),
	.w5(32'hbaed770d),
	.w6(32'h3b15c0f9),
	.w7(32'h3b2f2f69),
	.w8(32'h3b6e6fba),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86c7bcc),
	.w1(32'hb94978fc),
	.w2(32'hbb2ee9b8),
	.w3(32'h3ba11a6d),
	.w4(32'hb9498829),
	.w5(32'h3c71d0d8),
	.w6(32'h3be74975),
	.w7(32'hbba01067),
	.w8(32'h39bc6286),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb788f22),
	.w1(32'hbc39f45a),
	.w2(32'h3b2457be),
	.w3(32'h3ae355f2),
	.w4(32'hbbedbd29),
	.w5(32'h3a984340),
	.w6(32'hbba0cd04),
	.w7(32'h3c21d057),
	.w8(32'h3aaf7a79),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbec1a),
	.w1(32'h38497faf),
	.w2(32'hb92e7800),
	.w3(32'hbadf8369),
	.w4(32'h3c0e573c),
	.w5(32'hbc0f00b1),
	.w6(32'h3b18e6d5),
	.w7(32'h3c23a008),
	.w8(32'hb9bb6f7a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f0505),
	.w1(32'h3b7bd4ae),
	.w2(32'hbc278e73),
	.w3(32'hbc187206),
	.w4(32'h3a96f618),
	.w5(32'hbca206b4),
	.w6(32'hb804183f),
	.w7(32'h3bd134f3),
	.w8(32'hbc65dbe7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf68d69),
	.w1(32'hba9c13da),
	.w2(32'hb9e20a1b),
	.w3(32'hbc3613f3),
	.w4(32'h3bb0c145),
	.w5(32'h3c57d8f7),
	.w6(32'hbbd85888),
	.w7(32'hb987a254),
	.w8(32'hbb88f9a0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27cc2c),
	.w1(32'h39ffb028),
	.w2(32'hbb6fbbe8),
	.w3(32'h3bdd9d4a),
	.w4(32'h3b445809),
	.w5(32'hb9f723a4),
	.w6(32'hba87d28c),
	.w7(32'h3b2075b8),
	.w8(32'h3a308ab2),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb83e60),
	.w1(32'hb9e831c0),
	.w2(32'hbc81a2c6),
	.w3(32'hbb01d88f),
	.w4(32'hbb0d137f),
	.w5(32'hbc657ee8),
	.w6(32'hbb978160),
	.w7(32'h3c1989ab),
	.w8(32'hbc039f06),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc240acc),
	.w1(32'h3b8af987),
	.w2(32'hbb84aa99),
	.w3(32'hbc7616df),
	.w4(32'h3c5a4630),
	.w5(32'hbb2781a5),
	.w6(32'hbba93f32),
	.w7(32'h3bff03ff),
	.w8(32'hbb5b6106),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166309),
	.w1(32'h3b47b760),
	.w2(32'hbafd8c87),
	.w3(32'hbc052c4d),
	.w4(32'h3b186978),
	.w5(32'hbbc0dfb2),
	.w6(32'hbb606523),
	.w7(32'h3b3e9451),
	.w8(32'hbb18d610),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f9d7),
	.w1(32'h3c3b684b),
	.w2(32'h3c6641a8),
	.w3(32'hbb8659a9),
	.w4(32'h3cf794ed),
	.w5(32'h3c99d67a),
	.w6(32'hbba436e9),
	.w7(32'h3c1dc774),
	.w8(32'h3c514990),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb670fe),
	.w1(32'hbb1eaeaf),
	.w2(32'hbc9b9744),
	.w3(32'hbc698f6d),
	.w4(32'hbc3b0269),
	.w5(32'hbcaaf3a1),
	.w6(32'hbc38a1d0),
	.w7(32'hbb461bc4),
	.w8(32'hbca0d653),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a792a),
	.w1(32'hbb1b35b9),
	.w2(32'hbbc2966c),
	.w3(32'hbc909100),
	.w4(32'h3bc3299e),
	.w5(32'hbba91570),
	.w6(32'hbc4984ab),
	.w7(32'h3b77938c),
	.w8(32'hbb946ef6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8c8e2),
	.w1(32'hbc5aab67),
	.w2(32'hbc82c594),
	.w3(32'hbbccb9b1),
	.w4(32'hbc9f328f),
	.w5(32'hbc85e8cd),
	.w6(32'hbb5be8b5),
	.w7(32'hbc61802f),
	.w8(32'hbc8aa075),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac8ba9),
	.w1(32'hbbb43acf),
	.w2(32'hbbfd4e2f),
	.w3(32'hbb710a48),
	.w4(32'hbc477374),
	.w5(32'hbc183ab8),
	.w6(32'h3ac077ea),
	.w7(32'hbbbcc312),
	.w8(32'hbb827740),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc409f39),
	.w1(32'hbc0c9254),
	.w2(32'h3c09b656),
	.w3(32'hbcb0e992),
	.w4(32'hbc32e7cb),
	.w5(32'h3b264ead),
	.w6(32'hbc4a6d17),
	.w7(32'hbae000e9),
	.w8(32'h3b2f24cc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f812),
	.w1(32'hbbf2d542),
	.w2(32'h3ae754b5),
	.w3(32'hbb8d84c5),
	.w4(32'hbb4c244a),
	.w5(32'h3a76279e),
	.w6(32'hbb71f77a),
	.w7(32'h3a8c79d2),
	.w8(32'h3bc0c98c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c0cc),
	.w1(32'h3a64ca80),
	.w2(32'hbc038c91),
	.w3(32'h397f0961),
	.w4(32'h3c5e1d9e),
	.w5(32'h3c149856),
	.w6(32'h39a46dcc),
	.w7(32'h3a9f0a19),
	.w8(32'hbbb316ed),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1c0b4),
	.w1(32'hbc787186),
	.w2(32'h3a84f7d3),
	.w3(32'hbb588ef1),
	.w4(32'hbcad15da),
	.w5(32'h3c185e8c),
	.w6(32'hbb07c658),
	.w7(32'hbc41a9dc),
	.w8(32'h3b06437e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e848d),
	.w1(32'h3c2e0775),
	.w2(32'hbc005d33),
	.w3(32'h3cb324e2),
	.w4(32'hbbd02f45),
	.w5(32'hbc211d24),
	.w6(32'h3c2baa20),
	.w7(32'hbc0a6527),
	.w8(32'hbc1348b8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81b9ba),
	.w1(32'h3b18c4df),
	.w2(32'h3bf694dd),
	.w3(32'hbab47963),
	.w4(32'h3b863639),
	.w5(32'h3ca08650),
	.w6(32'h3b8e05f4),
	.w7(32'h3b4efa2a),
	.w8(32'h3c158c3e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f80a5),
	.w1(32'h3b581500),
	.w2(32'h3bd9f284),
	.w3(32'h3b12c3af),
	.w4(32'h3c7db064),
	.w5(32'h3b72abc6),
	.w6(32'h3abaedc1),
	.w7(32'h3b1a6676),
	.w8(32'h3a332fea),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78466dd),
	.w1(32'h3aabe6d3),
	.w2(32'hbc82a92e),
	.w3(32'hbbffdca9),
	.w4(32'hbafad53d),
	.w5(32'hbc8814a9),
	.w6(32'h387a979e),
	.w7(32'h3ac72bf1),
	.w8(32'hbc279087),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6553a4),
	.w1(32'hbb808f31),
	.w2(32'h3bc13ecd),
	.w3(32'hbb48deb4),
	.w4(32'h3c15c195),
	.w5(32'h3adb889a),
	.w6(32'hba9b5480),
	.w7(32'h3c01db14),
	.w8(32'h3c119bd4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64945c),
	.w1(32'h3b19ddc4),
	.w2(32'h3c5aaa5f),
	.w3(32'hbb8da7cc),
	.w4(32'h3c1567f2),
	.w5(32'h3d14bfaa),
	.w6(32'hbbd21e6c),
	.w7(32'h3b8327b7),
	.w8(32'h3c69b34b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac460b6),
	.w1(32'h3c0cdb58),
	.w2(32'h3bf28a51),
	.w3(32'h3bf9cc64),
	.w4(32'h3bf5648f),
	.w5(32'h3b47ea68),
	.w6(32'h3aab5dc4),
	.w7(32'hbbd1537d),
	.w8(32'hbc23cc3a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b515637),
	.w1(32'hbbb9be77),
	.w2(32'hbbbfb536),
	.w3(32'h3bcd0751),
	.w4(32'hbba3dc6f),
	.w5(32'hb956e9ea),
	.w6(32'h3b2f5dea),
	.w7(32'hbaa82adc),
	.w8(32'h3b100a1f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974775),
	.w1(32'hb8f2974b),
	.w2(32'hbc1a3216),
	.w3(32'h3bd17270),
	.w4(32'h3b476026),
	.w5(32'hbbfe58a1),
	.w6(32'h3c386035),
	.w7(32'h3bc381cf),
	.w8(32'hbc17295c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3ad54),
	.w1(32'h3aa9b3fa),
	.w2(32'h3bee0f3b),
	.w3(32'h3b41f1c3),
	.w4(32'h3c200fcf),
	.w5(32'h3cc06fb5),
	.w6(32'hbb5ee0ef),
	.w7(32'h3afa1d00),
	.w8(32'h3c5b1aa9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42559f),
	.w1(32'hb9ebda38),
	.w2(32'h3aa3a972),
	.w3(32'h3bb4edbf),
	.w4(32'h3ba39ef4),
	.w5(32'hb8cc857e),
	.w6(32'h3b8c92a4),
	.w7(32'h3c08198c),
	.w8(32'hbb565e65),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0aeb),
	.w1(32'h3ad21257),
	.w2(32'h3bb7178d),
	.w3(32'hb9e9bb3f),
	.w4(32'h3b7eaeb7),
	.w5(32'h3cd1e2a4),
	.w6(32'hba804027),
	.w7(32'hbac81272),
	.w8(32'h3c51317a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb399d9),
	.w1(32'h3b001223),
	.w2(32'hbaa2bd8f),
	.w3(32'hba5b97f6),
	.w4(32'h3c4fe1e4),
	.w5(32'hbb3c4f7c),
	.w6(32'hbbb8e2c9),
	.w7(32'h3c49af84),
	.w8(32'h3b188305),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb1071),
	.w1(32'hbafbeff2),
	.w2(32'hb9bdcb10),
	.w3(32'h3acfa6ed),
	.w4(32'hbb187ba3),
	.w5(32'h3c999893),
	.w6(32'hbaf37cf9),
	.w7(32'hbb082897),
	.w8(32'h3a1e8b99),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb660d2d),
	.w1(32'hbbead70e),
	.w2(32'hbc0fd41b),
	.w3(32'h3b848bfe),
	.w4(32'hbc21f9fe),
	.w5(32'hbb38b93f),
	.w6(32'hbaafc744),
	.w7(32'hbc8384aa),
	.w8(32'hbc145acd),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2291b),
	.w1(32'hbbc09f03),
	.w2(32'hbbe7f24c),
	.w3(32'h3c324f1b),
	.w4(32'hbc7470bf),
	.w5(32'hbbdc4c08),
	.w6(32'hbc0fda6c),
	.w7(32'hbc2ce91a),
	.w8(32'hbc15afe4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09486b),
	.w1(32'hbb1737db),
	.w2(32'h3bf68d29),
	.w3(32'hbc67c2ee),
	.w4(32'h39a7bb80),
	.w5(32'h3cfddfe1),
	.w6(32'hbbc0b549),
	.w7(32'h3a9be044),
	.w8(32'h3a3a3bab),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec60fc),
	.w1(32'hbc0e0199),
	.w2(32'hbc47d049),
	.w3(32'h3b5edd26),
	.w4(32'h3aaa4297),
	.w5(32'hbac5e85f),
	.w6(32'hbac48a9a),
	.w7(32'hbb2badef),
	.w8(32'hbb80f108),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f81ca),
	.w1(32'hba7f76a0),
	.w2(32'hba8f363a),
	.w3(32'h3bef1692),
	.w4(32'h393ebf3f),
	.w5(32'h3ba23b7a),
	.w6(32'hbbd371ed),
	.w7(32'h38e0d08e),
	.w8(32'h3bb6a518),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a954d2a),
	.w1(32'h3c0adf2c),
	.w2(32'h3ab6d4f0),
	.w3(32'h3b13354e),
	.w4(32'h3c585c5e),
	.w5(32'h3b57571c),
	.w6(32'h3c0c6d81),
	.w7(32'h3c40400b),
	.w8(32'hbaca9b0a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc227585),
	.w1(32'hbabd46d8),
	.w2(32'hbaea8de3),
	.w3(32'hbc9e3937),
	.w4(32'hbb5a6644),
	.w5(32'h39db30d3),
	.w6(32'hbc1621d6),
	.w7(32'h3a0c9f88),
	.w8(32'hbafe9848),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beda3f5),
	.w1(32'h3bff384d),
	.w2(32'h3b90b64d),
	.w3(32'h3bc4579b),
	.w4(32'h3c16c0c7),
	.w5(32'h3c6335aa),
	.w6(32'h3beabf51),
	.w7(32'h3c102f38),
	.w8(32'h3c264cda),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b433080),
	.w1(32'hbc53d6d5),
	.w2(32'hbc80edee),
	.w3(32'h39f9ebc9),
	.w4(32'hbcd7013d),
	.w5(32'hbcb476aa),
	.w6(32'hbb0d3e0f),
	.w7(32'hbcacd727),
	.w8(32'hbc9e235e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6211fb),
	.w1(32'hbae449d3),
	.w2(32'h3c57fd07),
	.w3(32'hbbc399b3),
	.w4(32'hba3f6b8a),
	.w5(32'h3c2c0273),
	.w6(32'hbbebc2a6),
	.w7(32'hbb1065ba),
	.w8(32'h3be15adc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc45d10),
	.w1(32'h3c1ec198),
	.w2(32'hbaa01ed6),
	.w3(32'h3c9ec7aa),
	.w4(32'h3c70576c),
	.w5(32'hbbe02cbd),
	.w6(32'hbaa3d97b),
	.w7(32'h3c47d78c),
	.w8(32'hbb5382ca),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70e8fd),
	.w1(32'hbaa6a14d),
	.w2(32'hbb8656e1),
	.w3(32'hbb6a3f56),
	.w4(32'hba721181),
	.w5(32'h38b9e52d),
	.w6(32'hbb229385),
	.w7(32'h3ba4d8d4),
	.w8(32'h3b0342ee),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab202c),
	.w1(32'hbb310919),
	.w2(32'h3c151e69),
	.w3(32'h3c16cc4a),
	.w4(32'hbbecf5e7),
	.w5(32'h3b35363b),
	.w6(32'h3b96e1d8),
	.w7(32'hbb124ff4),
	.w8(32'h3c0f57cd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afdfd76),
	.w1(32'h3b116054),
	.w2(32'hbb45a657),
	.w3(32'h3b13e625),
	.w4(32'h3bbf8009),
	.w5(32'h3c5515ff),
	.w6(32'h3c17f15b),
	.w7(32'h3b8a97dc),
	.w8(32'h3c07b448),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3ce14),
	.w1(32'h3bd007d2),
	.w2(32'hba8894dc),
	.w3(32'h3952e7cb),
	.w4(32'h3c7bb8ea),
	.w5(32'h3c4bdd71),
	.w6(32'h3b6893eb),
	.w7(32'h3bf597ec),
	.w8(32'hbb1e8a39),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59adb3),
	.w1(32'h3b836c1e),
	.w2(32'hbb3dc736),
	.w3(32'hbbb8c436),
	.w4(32'h3c116b1d),
	.w5(32'h3c8e869b),
	.w6(32'hbb77797a),
	.w7(32'hbb23dc22),
	.w8(32'h3a239ae9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad998d),
	.w1(32'h3bde767f),
	.w2(32'hb9847652),
	.w3(32'h3b6b4252),
	.w4(32'h3b0e8111),
	.w5(32'hbbe9e1af),
	.w6(32'h3a09b38a),
	.w7(32'h3b4787d6),
	.w8(32'hbb29a50a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55e14d),
	.w1(32'hbbf3f108),
	.w2(32'hbb6d31d6),
	.w3(32'hba746f8c),
	.w4(32'hbc1108cb),
	.w5(32'hbb3b4d22),
	.w6(32'h3acae182),
	.w7(32'hbc2ded8d),
	.w8(32'hbc0bb033),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28da29),
	.w1(32'hbba858e2),
	.w2(32'hbcc84ee2),
	.w3(32'h3ba81a9d),
	.w4(32'h3a96c508),
	.w5(32'hbce23957),
	.w6(32'h3af40a14),
	.w7(32'h3b41325c),
	.w8(32'hbce96c4c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc352281),
	.w1(32'h3a16f5a8),
	.w2(32'hba57346f),
	.w3(32'hbc7d5db9),
	.w4(32'hbb89f54c),
	.w5(32'h3c8704db),
	.w6(32'hbc1e744a),
	.w7(32'h3a89cf3b),
	.w8(32'hbb35ff0a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a4752),
	.w1(32'hbacbc495),
	.w2(32'hb8d30aa9),
	.w3(32'h3c49fc10),
	.w4(32'hbc1f1e56),
	.w5(32'h3ae146af),
	.w6(32'h3c451c15),
	.w7(32'hbb607dbd),
	.w8(32'h3a819b0f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d02a7),
	.w1(32'h3b85c92e),
	.w2(32'hbb6df3e0),
	.w3(32'h3c11ffbb),
	.w4(32'hba15f35f),
	.w5(32'hbc683110),
	.w6(32'h3abae7c0),
	.w7(32'h3b8ecdf4),
	.w8(32'hbb9f1da9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a21ce),
	.w1(32'hbb1b5c14),
	.w2(32'h3bfcbda6),
	.w3(32'hbc30a4e1),
	.w4(32'h3bfa1d3e),
	.w5(32'h3d24e347),
	.w6(32'hba724b6c),
	.w7(32'hbb2b0257),
	.w8(32'hba14ea21),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe0473),
	.w1(32'h3bb6b4bd),
	.w2(32'hbba16fb9),
	.w3(32'h3bbdcb7b),
	.w4(32'h3ba96dcc),
	.w5(32'hbc61154c),
	.w6(32'hbb451633),
	.w7(32'h3b9a6ae9),
	.w8(32'hbb3f66aa),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7689b3),
	.w1(32'h3b7862f7),
	.w2(32'h3b9fe217),
	.w3(32'hbbcfde6a),
	.w4(32'h3a86900d),
	.w5(32'h3c2e0e60),
	.w6(32'h3ac19d1a),
	.w7(32'h3b861a27),
	.w8(32'h3bb94d0e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d967e),
	.w1(32'hbb24a23e),
	.w2(32'hbb1bf6b4),
	.w3(32'h3bce796e),
	.w4(32'hbc02cc32),
	.w5(32'hbc2a2e2b),
	.w6(32'h3b63c28c),
	.w7(32'hbb93f573),
	.w8(32'hbb83969e),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb104e40),
	.w1(32'hbba2d5cf),
	.w2(32'hbad20f07),
	.w3(32'hbba54479),
	.w4(32'hbb6ebe7d),
	.w5(32'h3a057d87),
	.w6(32'hb9366b9a),
	.w7(32'hbb8f7f32),
	.w8(32'h38923958),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac49e2c),
	.w1(32'h3bb591af),
	.w2(32'h3ab18071),
	.w3(32'hbb1d4415),
	.w4(32'h3c030a44),
	.w5(32'h3bba82de),
	.w6(32'h3b7a10e8),
	.w7(32'h3c867e96),
	.w8(32'h3aea5119),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd888b6),
	.w1(32'h3c3fb61b),
	.w2(32'hba994fda),
	.w3(32'hbc8262c0),
	.w4(32'h3cc9e92d),
	.w5(32'h3c16e2ee),
	.w6(32'hbc282efe),
	.w7(32'h3bea449d),
	.w8(32'h3b6c1e6e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb775d54),
	.w1(32'h3b68acbc),
	.w2(32'h3abfb3b3),
	.w3(32'hb9c38b10),
	.w4(32'h3b32d5cc),
	.w5(32'h3c448690),
	.w6(32'h3a917a24),
	.w7(32'h3ad7ea76),
	.w8(32'h3be3aa5c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b6612),
	.w1(32'h3a2f220e),
	.w2(32'h3ae7bc8a),
	.w3(32'hbc239602),
	.w4(32'h39f1ad7b),
	.w5(32'hb98892a5),
	.w6(32'hbbe55f59),
	.w7(32'h3a5366a2),
	.w8(32'h3827eb09),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e4096),
	.w1(32'h3b17b743),
	.w2(32'h3b3e64f5),
	.w3(32'h3a4e347c),
	.w4(32'h3b6cc0a4),
	.w5(32'hb830a431),
	.w6(32'h3a9d7c69),
	.w7(32'h3ba9f1c7),
	.w8(32'h3ab3969f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f1f9a),
	.w1(32'h3bb7d525),
	.w2(32'h3a1e8d92),
	.w3(32'hbb595664),
	.w4(32'h3a8783bb),
	.w5(32'h3bd8296d),
	.w6(32'hbab4ee9e),
	.w7(32'h398781fe),
	.w8(32'h392a08ef),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8053e2),
	.w1(32'hb8a4aa75),
	.w2(32'h3b683704),
	.w3(32'hbc0c8963),
	.w4(32'h3a00dde1),
	.w5(32'h3b976e69),
	.w6(32'hba9bbc3d),
	.w7(32'hb87d67b3),
	.w8(32'h3a9ae063),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc87dd),
	.w1(32'hbb87e9ce),
	.w2(32'hbb640202),
	.w3(32'h3b01b952),
	.w4(32'hbbb4d3e4),
	.w5(32'hbb0a18f4),
	.w6(32'h3a30088d),
	.w7(32'hbc02978b),
	.w8(32'hbbd38f13),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48e1d0),
	.w1(32'hbb74f97d),
	.w2(32'hbaa4b8ce),
	.w3(32'hbab77f7e),
	.w4(32'hbb22badd),
	.w5(32'hbb06c6cb),
	.w6(32'hb9ca573b),
	.w7(32'hbaf029b6),
	.w8(32'hbab1d41f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cf17a),
	.w1(32'h3bb92a88),
	.w2(32'hbae361b5),
	.w3(32'hba280502),
	.w4(32'h3bb2e918),
	.w5(32'h3b327e01),
	.w6(32'hba8074c6),
	.w7(32'h3b5dbecc),
	.w8(32'h3afe1adf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8f48),
	.w1(32'hba1b2a39),
	.w2(32'hbb81e32b),
	.w3(32'h3be70eac),
	.w4(32'h3ae0ab9b),
	.w5(32'hbb7c69b4),
	.w6(32'h3bbd4e40),
	.w7(32'h3bce02a5),
	.w8(32'hba50cae7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d885),
	.w1(32'hbb3666b0),
	.w2(32'hbbf70a3a),
	.w3(32'hbaa657e9),
	.w4(32'h3ad3d418),
	.w5(32'hbc18825f),
	.w6(32'hbbcd54d5),
	.w7(32'h3aa5de88),
	.w8(32'hbc1ba630),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840936),
	.w1(32'h396197f7),
	.w2(32'h3a965d65),
	.w3(32'hbb07f338),
	.w4(32'hbb846ae1),
	.w5(32'hbad9e5c6),
	.w6(32'hbb5b4b28),
	.w7(32'hbbc843c7),
	.w8(32'hba02069d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831ebf7),
	.w1(32'h3c52f5ab),
	.w2(32'h3c1684e6),
	.w3(32'h39440d31),
	.w4(32'h3c8389ec),
	.w5(32'h3c265570),
	.w6(32'hba24120a),
	.w7(32'h3c4abb94),
	.w8(32'h3c22aed7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30108c),
	.w1(32'hba7dcc98),
	.w2(32'h3af1173f),
	.w3(32'h3c6eda73),
	.w4(32'hbaa093e9),
	.w5(32'hb9a9759e),
	.w6(32'h3c316b35),
	.w7(32'h3a6b8fb8),
	.w8(32'h3914b88e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5ea68),
	.w1(32'hbb61aaa4),
	.w2(32'hbb08340d),
	.w3(32'h3b9d8fe6),
	.w4(32'hbb207a6c),
	.w5(32'hba4ec1c4),
	.w6(32'h3b650b21),
	.w7(32'hbb063998),
	.w8(32'hbae09bc4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03de21),
	.w1(32'hb9459add),
	.w2(32'h3ac68988),
	.w3(32'h3b05adbb),
	.w4(32'h3b75b6c3),
	.w5(32'h3bc124cd),
	.w6(32'h3aebb8c6),
	.w7(32'h3b8d9de5),
	.w8(32'h3b921998),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8050f5),
	.w1(32'hba864459),
	.w2(32'h3a335782),
	.w3(32'h3baf5303),
	.w4(32'hba9de5c2),
	.w5(32'hbb227024),
	.w6(32'h3b999f50),
	.w7(32'hbaeb2b9d),
	.w8(32'hbbcad3d3),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc76b6),
	.w1(32'hba2e6a26),
	.w2(32'h3a1fc0b6),
	.w3(32'hba32356c),
	.w4(32'h3b6230bc),
	.w5(32'h3baea18f),
	.w6(32'hba9fe479),
	.w7(32'h3bc64085),
	.w8(32'hba8264c1),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa8df1),
	.w1(32'h3b421d1f),
	.w2(32'h3b868357),
	.w3(32'hbb70010a),
	.w4(32'h3c08ccac),
	.w5(32'h3b28a1a9),
	.w6(32'hbbbf5b0f),
	.w7(32'h3b481b8a),
	.w8(32'h3bc6ae67),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3a441),
	.w1(32'hbafc3f97),
	.w2(32'hbb8d0e69),
	.w3(32'hba9e2285),
	.w4(32'h39fce56e),
	.w5(32'hbb6650d3),
	.w6(32'hb93b9c19),
	.w7(32'h3ab45f17),
	.w8(32'hbb04259d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7610f7),
	.w1(32'h3832757a),
	.w2(32'hbac8093c),
	.w3(32'hbb38400b),
	.w4(32'h3a6cce0e),
	.w5(32'h3a258536),
	.w6(32'hbb3f2dab),
	.w7(32'hbbc2c9a3),
	.w8(32'hba9ff64c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb665e18),
	.w1(32'hbb0cfba7),
	.w2(32'hbaf9f08d),
	.w3(32'hb7d431f9),
	.w4(32'h3a2eb0db),
	.w5(32'hba8605f7),
	.w6(32'hbab325ef),
	.w7(32'h3ad05513),
	.w8(32'hb8d8b4af),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c51b8),
	.w1(32'hbb4905eb),
	.w2(32'h3adc45c8),
	.w3(32'h3aeff705),
	.w4(32'hba72cd07),
	.w5(32'hb8028a79),
	.w6(32'h3b1d431c),
	.w7(32'hbb8c6ea1),
	.w8(32'h3a41a70f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3baec),
	.w1(32'h3adfd365),
	.w2(32'hba3b7116),
	.w3(32'hbbbc63c0),
	.w4(32'h3b0bcf58),
	.w5(32'h3b24f5cf),
	.w6(32'hbbaf98fd),
	.w7(32'h3a4b8006),
	.w8(32'h3b8009e7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8aa8ab),
	.w1(32'hbb57f942),
	.w2(32'hbb29e6fa),
	.w3(32'hbac493d1),
	.w4(32'hbaa33db2),
	.w5(32'hbabf1234),
	.w6(32'h3aa2243e),
	.w7(32'hbb48e631),
	.w8(32'hbb03afa7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae292f4),
	.w1(32'hb9f0e2e8),
	.w2(32'hbb7c2198),
	.w3(32'hbafd66f8),
	.w4(32'h3b079673),
	.w5(32'hbae9dd65),
	.w6(32'h3ac1ca46),
	.w7(32'h3ab49569),
	.w8(32'hb9cc9783),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38a771),
	.w1(32'hb6a21a79),
	.w2(32'hbb56b319),
	.w3(32'hbab99ab7),
	.w4(32'hbb23548c),
	.w5(32'hbacf5533),
	.w6(32'hba3f0caa),
	.w7(32'hbbc3d6c2),
	.w8(32'hbb60ab82),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc29fff),
	.w1(32'h3a74ad4d),
	.w2(32'h393efd9b),
	.w3(32'hbbacc057),
	.w4(32'hbbb0c205),
	.w5(32'h3b8f77ae),
	.w6(32'hbbb9dd1d),
	.w7(32'hbb5434d9),
	.w8(32'h3b4b9e2c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb871c7c),
	.w1(32'hba23f1ec),
	.w2(32'hbbca0c3f),
	.w3(32'hb9fa9952),
	.w4(32'h3af82651),
	.w5(32'hbafde893),
	.w6(32'hba35919f),
	.w7(32'hb9584538),
	.w8(32'hbb99cc9a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11ea79),
	.w1(32'hbb99eca6),
	.w2(32'hbbd0004a),
	.w3(32'hbbb45310),
	.w4(32'hbac4b8c1),
	.w5(32'hbb8e1c71),
	.w6(32'hbbd73a33),
	.w7(32'h3acfbbd1),
	.w8(32'hbb2e273b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4100b5),
	.w1(32'hb88f3403),
	.w2(32'h3c1293c0),
	.w3(32'h3a7872b7),
	.w4(32'hb903c27d),
	.w5(32'h3bfa5f65),
	.w6(32'h3aba077b),
	.w7(32'hba8905d8),
	.w8(32'h3bcc7c57),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8889db),
	.w1(32'hbac6d252),
	.w2(32'hb99bf776),
	.w3(32'h3c2d93e0),
	.w4(32'h3b15b02c),
	.w5(32'h3a63b75b),
	.w6(32'h3b790135),
	.w7(32'h3bc0cb9e),
	.w8(32'hbac8c99e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f69d),
	.w1(32'hbafa5c8d),
	.w2(32'h389f78d9),
	.w3(32'hbbf9b37a),
	.w4(32'h3b127c54),
	.w5(32'hb92ff04d),
	.w6(32'hbc14938e),
	.w7(32'hb9a4b993),
	.w8(32'hbab6a7a0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc288258),
	.w1(32'hbbcca4ec),
	.w2(32'hbc09e3c4),
	.w3(32'hbbe6f99a),
	.w4(32'hbb7545b2),
	.w5(32'hbbe1be71),
	.w6(32'hbbc9e012),
	.w7(32'hbba50a9f),
	.w8(32'hbc07b497),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26c41),
	.w1(32'hbb99774d),
	.w2(32'hbc00afe6),
	.w3(32'hbaf095c2),
	.w4(32'hbbcf75a6),
	.w5(32'hbc293506),
	.w6(32'hbb4f007b),
	.w7(32'hbb7134c7),
	.w8(32'hbba9d4ad),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb761e62),
	.w1(32'hbabbf416),
	.w2(32'hbbbad6ea),
	.w3(32'hbaf2f801),
	.w4(32'h3b224474),
	.w5(32'hbbcb9147),
	.w6(32'hb8d0a9f1),
	.w7(32'h3b9d679d),
	.w8(32'hbbc5ec88),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba8eb1),
	.w1(32'hb8d08592),
	.w2(32'hba90ea1e),
	.w3(32'hbb868a61),
	.w4(32'h3ba3b52f),
	.w5(32'h3beaf032),
	.w6(32'hbb90f46a),
	.w7(32'h3a6ff0ec),
	.w8(32'hba2032f7),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1a176),
	.w1(32'hbb8fc646),
	.w2(32'hbb439688),
	.w3(32'h3be881c6),
	.w4(32'hbb77fee0),
	.w5(32'hba970121),
	.w6(32'h3bbb0f51),
	.w7(32'hbb87821d),
	.w8(32'hbb4661f1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd70bb),
	.w1(32'hb9d08665),
	.w2(32'h3a3f6d37),
	.w3(32'hbb015b19),
	.w4(32'h39c8f740),
	.w5(32'hbb024b37),
	.w6(32'hbb23220f),
	.w7(32'h3b64fb9e),
	.w8(32'hbb2b42f0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa40c88),
	.w1(32'h3b4351c9),
	.w2(32'h3bf8f107),
	.w3(32'hba258b61),
	.w4(32'h3b582f4b),
	.w5(32'h3c626992),
	.w6(32'hbac1cc59),
	.w7(32'hbabaf00f),
	.w8(32'h3bf2bfd0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6d0e),
	.w1(32'hbb22cde4),
	.w2(32'hbb3c77ee),
	.w3(32'hbb7da2ab),
	.w4(32'h3b40e047),
	.w5(32'h3a72c08b),
	.w6(32'hbaeb4828),
	.w7(32'h3b57cab0),
	.w8(32'h392731f3),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9f27c),
	.w1(32'h3bee6813),
	.w2(32'hbb292a9e),
	.w3(32'h3abbd3f4),
	.w4(32'h3b8515a7),
	.w5(32'h3b80de4e),
	.w6(32'h3afb4ae1),
	.w7(32'hbb1b0ac2),
	.w8(32'h3b1a3687),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3b591),
	.w1(32'hbb767b54),
	.w2(32'h3a5637fe),
	.w3(32'hbb7c1c8c),
	.w4(32'hba55ed11),
	.w5(32'h3b09c954),
	.w6(32'hbb42a716),
	.w7(32'hbb27b9b3),
	.w8(32'hb9bd7620),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828478),
	.w1(32'hbb83c49a),
	.w2(32'hbb4c2eea),
	.w3(32'hbb0974c7),
	.w4(32'hbb21f598),
	.w5(32'hbb004044),
	.w6(32'hbb6eeb21),
	.w7(32'hbab63b9f),
	.w8(32'hbb34a2d7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc7205),
	.w1(32'h3accd769),
	.w2(32'hbb292fa3),
	.w3(32'hbb790883),
	.w4(32'h39ad76b9),
	.w5(32'hb90211a7),
	.w6(32'hbb91991e),
	.w7(32'h3b266bd9),
	.w8(32'hb80fe7bf),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b06c),
	.w1(32'hbada4c21),
	.w2(32'hbbc1175a),
	.w3(32'h3b03c8b2),
	.w4(32'h3a9cf7fb),
	.w5(32'hbbeac1f3),
	.w6(32'h3b3351ff),
	.w7(32'hbad7974b),
	.w8(32'hbba34246),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95830e),
	.w1(32'h3b0f232c),
	.w2(32'hbb871bd7),
	.w3(32'hbb41913c),
	.w4(32'h3ba1aa55),
	.w5(32'hbb722fa4),
	.w6(32'hbba6f6db),
	.w7(32'h3b846e5b),
	.w8(32'hb9b8ca24),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b690974),
	.w1(32'hbaa2dd94),
	.w2(32'hba1aea02),
	.w3(32'h3a17cc32),
	.w4(32'hbaaf3fc6),
	.w5(32'h389d53e7),
	.w6(32'h3b950181),
	.w7(32'hb9f17a1c),
	.w8(32'h39fe3f83),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d798d),
	.w1(32'hb93614c0),
	.w2(32'hbbcbc4ec),
	.w3(32'h3b0c24fa),
	.w4(32'hba700f67),
	.w5(32'hbc02774e),
	.w6(32'h3b118a8e),
	.w7(32'hbb08b289),
	.w8(32'hbba9df10),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f9923),
	.w1(32'hbb19f15b),
	.w2(32'hbb252e30),
	.w3(32'hba9a204f),
	.w4(32'hbb091e2e),
	.w5(32'hbba4aaff),
	.w6(32'hbb3019a9),
	.w7(32'hbb9650ad),
	.w8(32'hbc096255),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4aa26),
	.w1(32'hbbc1f8b6),
	.w2(32'hbb3d2a9e),
	.w3(32'hbb82959a),
	.w4(32'hbbc348bf),
	.w5(32'hbb8b149f),
	.w6(32'hbbe6e83c),
	.w7(32'hbbc8dfb3),
	.w8(32'hbb95718a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23943a),
	.w1(32'hbab5a18b),
	.w2(32'hbc03e213),
	.w3(32'hbb41fe55),
	.w4(32'hbb0f1b52),
	.w5(32'hbb205fb8),
	.w6(32'hbbb5d6c6),
	.w7(32'hbbd639a5),
	.w8(32'h39b6b7e2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdb44f),
	.w1(32'h3babdccb),
	.w2(32'h3b8a5680),
	.w3(32'hbbc02708),
	.w4(32'h3b6f93c3),
	.w5(32'h3b8a0bc0),
	.w6(32'hbb6ccdd0),
	.w7(32'h3afea06e),
	.w8(32'h3ac3ca19),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baedf50),
	.w1(32'h3b0078c7),
	.w2(32'h3b9bc9b7),
	.w3(32'h3b44c2ee),
	.w4(32'h3bafef81),
	.w5(32'h3c0554a8),
	.w6(32'h3bcda378),
	.w7(32'h3b9abdfd),
	.w8(32'h3bbd7190),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb486901),
	.w1(32'hbb2832d1),
	.w2(32'hbbbc31b2),
	.w3(32'hbb9225c2),
	.w4(32'h3a9011b2),
	.w5(32'hba3e1c37),
	.w6(32'hbbec7827),
	.w7(32'h3ae348f7),
	.w8(32'hb8aebced),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1650c),
	.w1(32'hbbdbf06a),
	.w2(32'hb98d5a7f),
	.w3(32'h3a822a62),
	.w4(32'hbbc0bfcb),
	.w5(32'h39ab5c1a),
	.w6(32'h3a1c89f5),
	.w7(32'hbb8248cd),
	.w8(32'hba3cdc8b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2207c),
	.w1(32'h3b8d0e3e),
	.w2(32'h3b4f7e7c),
	.w3(32'h3c083aa4),
	.w4(32'h3bf7f68b),
	.w5(32'hbab3397a),
	.w6(32'h3b990fda),
	.w7(32'h3c1557ca),
	.w8(32'hbb06eb00),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5759),
	.w1(32'hbbad6e13),
	.w2(32'hbaad2114),
	.w3(32'hbba71bf5),
	.w4(32'hbb760ce7),
	.w5(32'hbac61ccf),
	.w6(32'hbafd31a8),
	.w7(32'hbbce4d11),
	.w8(32'hbbaf909c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf3d27),
	.w1(32'hbc0be03b),
	.w2(32'hbbfd112c),
	.w3(32'hbaa5df5d),
	.w4(32'hbc59f174),
	.w5(32'hbc4a2bda),
	.w6(32'hbb4fa07e),
	.w7(32'hbc0642a5),
	.w8(32'hbc17fa39),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2972c8),
	.w1(32'hbb13114e),
	.w2(32'hbafd85d3),
	.w3(32'hbc07ad0a),
	.w4(32'hba68cf66),
	.w5(32'h3aad4926),
	.w6(32'hbc142581),
	.w7(32'h3a13b604),
	.w8(32'h3aa1469c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b3b4e),
	.w1(32'h3b3a44df),
	.w2(32'h3a8816a1),
	.w3(32'h3bd8445c),
	.w4(32'h3a4b63fb),
	.w5(32'hb8beb21d),
	.w6(32'h3b6591c4),
	.w7(32'hbb0e56f9),
	.w8(32'h3ac4a940),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31641c),
	.w1(32'hbaa83378),
	.w2(32'h38b2f531),
	.w3(32'h3a666949),
	.w4(32'h3af7d9de),
	.w5(32'h3a319fae),
	.w6(32'h39a2e3f8),
	.w7(32'h3b14dac5),
	.w8(32'h3ac6f345),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80c32),
	.w1(32'h3aeabc45),
	.w2(32'hbbc0db3c),
	.w3(32'hb9b075fe),
	.w4(32'h3b4eadc3),
	.w5(32'hbbe0e2cc),
	.w6(32'h3886127d),
	.w7(32'hbaa503de),
	.w8(32'hbba953cb),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9bad20),
	.w1(32'h3aaffbbc),
	.w2(32'h3b26e640),
	.w3(32'hbbc478b9),
	.w4(32'h3b811265),
	.w5(32'hb80502f7),
	.w6(32'hbbc20241),
	.w7(32'h398d117b),
	.w8(32'h3805d9ac),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea5dd),
	.w1(32'hbb851156),
	.w2(32'hbac49eb5),
	.w3(32'hba9aacad),
	.w4(32'hbb8b3d4f),
	.w5(32'hbad3312f),
	.w6(32'hba506efc),
	.w7(32'hbb8b1b5e),
	.w8(32'hbb7cb597),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b09a5),
	.w1(32'hbb240390),
	.w2(32'hbb99fa5e),
	.w3(32'hbaae77c6),
	.w4(32'hbb16c865),
	.w5(32'hbb80a931),
	.w6(32'hbb87beac),
	.w7(32'h3b09bc12),
	.w8(32'hbb34d57d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5a3c5),
	.w1(32'hbba11db7),
	.w2(32'hbb953d8e),
	.w3(32'h3b31d766),
	.w4(32'h3b005fc4),
	.w5(32'h3a8089f2),
	.w6(32'h3a5b3984),
	.w7(32'h3b6c90c7),
	.w8(32'h3b42a2d8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb928d79),
	.w1(32'hbb9bd0cc),
	.w2(32'hbaca1109),
	.w3(32'hba3c1a45),
	.w4(32'hba876cb6),
	.w5(32'hb94778a0),
	.w6(32'h39b3fa1a),
	.w7(32'h3ac16917),
	.w8(32'h3b01aa14),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1179),
	.w1(32'hbbc4448c),
	.w2(32'hbbb907aa),
	.w3(32'hbb3d3311),
	.w4(32'hbb866151),
	.w5(32'hbb8b06da),
	.w6(32'hbbd889cb),
	.w7(32'hbbae9161),
	.w8(32'hbbf15569),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4486a5),
	.w1(32'hbb964641),
	.w2(32'hbb865518),
	.w3(32'hbc285593),
	.w4(32'hba4a8f2c),
	.w5(32'hb9b3f8de),
	.w6(32'hbc3923a4),
	.w7(32'h3b1b97a8),
	.w8(32'h3abfa468),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5925),
	.w1(32'hb9c6183b),
	.w2(32'hbb1878fa),
	.w3(32'hbb54b740),
	.w4(32'h3a6916e6),
	.w5(32'hbb23e382),
	.w6(32'hbb313edc),
	.w7(32'h3bc8c08d),
	.w8(32'h3b5323ae),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d64fa),
	.w1(32'hbb5e963e),
	.w2(32'hbb88f720),
	.w3(32'hbb0561ca),
	.w4(32'hbb323a86),
	.w5(32'hbbb72a87),
	.w6(32'h3b0614fa),
	.w7(32'hbb42696c),
	.w8(32'hbb885d77),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38009720),
	.w1(32'hbb1a7527),
	.w2(32'h3a259c4d),
	.w3(32'hbabbc570),
	.w4(32'h394def00),
	.w5(32'hb87de3f2),
	.w6(32'hb9d448e8),
	.w7(32'h3a697689),
	.w8(32'hbb06a62c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39114ed7),
	.w1(32'hbb8a2889),
	.w2(32'hbbd3d8fd),
	.w3(32'h3a77e340),
	.w4(32'hbb74c01b),
	.w5(32'hbbbccf27),
	.w6(32'hbad56c63),
	.w7(32'hbb8aeb45),
	.w8(32'hbb889581),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c4719),
	.w1(32'h3779f130),
	.w2(32'h3b13f71e),
	.w3(32'hbb7edb9a),
	.w4(32'h3b2dd8b5),
	.w5(32'hbaad7a58),
	.w6(32'h38e794e9),
	.w7(32'h3b6766f2),
	.w8(32'hbae2ad29),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b5946),
	.w1(32'h3c0a2916),
	.w2(32'h3b6bad12),
	.w3(32'h3b05cab3),
	.w4(32'h3bd07569),
	.w5(32'h3a8e786d),
	.w6(32'h3b227899),
	.w7(32'h3bc98889),
	.w8(32'h3b2d528b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873ebf),
	.w1(32'h3a6dd7c6),
	.w2(32'h3ad764be),
	.w3(32'h3ac66792),
	.w4(32'h39f858ae),
	.w5(32'h39c071fc),
	.w6(32'h3b37e316),
	.w7(32'hba2d0e71),
	.w8(32'hb92bf667),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc6d60),
	.w1(32'h3b802ca7),
	.w2(32'h3ba75d58),
	.w3(32'h3b32b9ac),
	.w4(32'h3ba478e8),
	.w5(32'h390c072c),
	.w6(32'h3b07f584),
	.w7(32'h3b855320),
	.w8(32'h3ab7fe13),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95008),
	.w1(32'hbb6cb216),
	.w2(32'hbb788692),
	.w3(32'h3b13ea7f),
	.w4(32'hbb124ea2),
	.w5(32'hbb8adaf2),
	.w6(32'h39a8e6f9),
	.w7(32'hbb46a573),
	.w8(32'hbbc9bd4b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399da844),
	.w1(32'h3b5d7206),
	.w2(32'h3a4177c5),
	.w3(32'hba131143),
	.w4(32'h3c1012d2),
	.w5(32'hbb168238),
	.w6(32'hbb0c707d),
	.w7(32'h3be31969),
	.w8(32'hba4a4970),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78fff6),
	.w1(32'h3b078b8e),
	.w2(32'h3a6d2bab),
	.w3(32'h3a9ae642),
	.w4(32'h3a9e3fb7),
	.w5(32'hba9b8140),
	.w6(32'h3ad5fad4),
	.w7(32'h3b6e2142),
	.w8(32'hba0ab6ae),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31c49e),
	.w1(32'hba70b1ad),
	.w2(32'hbb9c204f),
	.w3(32'h3b6ec7af),
	.w4(32'h3a6ac86b),
	.w5(32'hbbbce41b),
	.w6(32'h3afb6d33),
	.w7(32'h3ba580e1),
	.w8(32'hbb497494),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab139f3),
	.w1(32'hbbad1ad7),
	.w2(32'hbba792f7),
	.w3(32'h3a8c8a1f),
	.w4(32'hbb3614fa),
	.w5(32'hba556dd4),
	.w6(32'h3af60eef),
	.w7(32'h38b623e3),
	.w8(32'h3af523d2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9392a6),
	.w1(32'h3bf500fc),
	.w2(32'hbb832a08),
	.w3(32'hbb884d89),
	.w4(32'h3c41537d),
	.w5(32'h39859be4),
	.w6(32'h3a6b3c0d),
	.w7(32'h3c041e06),
	.w8(32'hbaf1df24),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1885d),
	.w1(32'h3c25627c),
	.w2(32'hba1a4f8e),
	.w3(32'hbb5a79da),
	.w4(32'h3bf2da39),
	.w5(32'h3b61c851),
	.w6(32'hbb919462),
	.w7(32'h3bac4338),
	.w8(32'h3c2296a4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe0aff),
	.w1(32'hbb4f9a7c),
	.w2(32'h3acfc64c),
	.w3(32'hbc1f9e4f),
	.w4(32'hbb7ebc4e),
	.w5(32'hb98a7245),
	.w6(32'hbba4fa9b),
	.w7(32'h3931c4bc),
	.w8(32'h3b0a826f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e0059),
	.w1(32'h3ba5187c),
	.w2(32'hbbe8e84b),
	.w3(32'hbb8aa775),
	.w4(32'hb88ce45e),
	.w5(32'hbc0ec9e5),
	.w6(32'h3a85b25b),
	.w7(32'hbb747a1b),
	.w8(32'hbc034fbb),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f8bea),
	.w1(32'h3b71c5da),
	.w2(32'h3c2f090b),
	.w3(32'hbc06d279),
	.w4(32'h3bc22c96),
	.w5(32'h3c903a34),
	.w6(32'hbc313f45),
	.w7(32'h3bf6b807),
	.w8(32'h3c890201),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368ec2),
	.w1(32'hbbcf5085),
	.w2(32'hbb8e1f2e),
	.w3(32'h3a194af2),
	.w4(32'hbc34d53b),
	.w5(32'hbb8b6b6b),
	.w6(32'h3b6b5256),
	.w7(32'hbbe45f86),
	.w8(32'h3a516759),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963ed3),
	.w1(32'hbbe25c0a),
	.w2(32'hbada7ef8),
	.w3(32'hba273c67),
	.w4(32'hbc08f63a),
	.w5(32'hbbc95d5f),
	.w6(32'h39aad350),
	.w7(32'hbbd46c7d),
	.w8(32'hbbc39c6f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9d3fc),
	.w1(32'h3b957eb3),
	.w2(32'h3b88cb13),
	.w3(32'hb99c35a1),
	.w4(32'h3b8d588d),
	.w5(32'hb929bbd3),
	.w6(32'hbaffb772),
	.w7(32'h3b3aaf56),
	.w8(32'h3a01ccd2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b358bca),
	.w1(32'hbb7499ea),
	.w2(32'hbbb2f3d0),
	.w3(32'hbab2fb08),
	.w4(32'hbb5ce52f),
	.w5(32'hbb7666ec),
	.w6(32'hbac2917a),
	.w7(32'hbb459ddc),
	.w8(32'hbb04e446),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05ed7),
	.w1(32'h3b173f2f),
	.w2(32'hbb8d2248),
	.w3(32'hbbc1bb89),
	.w4(32'h3b5e6c3c),
	.w5(32'hbb60c076),
	.w6(32'hbbbeed0b),
	.w7(32'h3b7c5c00),
	.w8(32'hb901e01b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fe7e0),
	.w1(32'hbbdb5259),
	.w2(32'hbb95a309),
	.w3(32'hb99a95da),
	.w4(32'hbb94fe77),
	.w5(32'h3a015b60),
	.w6(32'h3a85cc37),
	.w7(32'h3abd874a),
	.w8(32'h3af2fc6f),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc009042),
	.w1(32'hbb3e0827),
	.w2(32'hbb1dc982),
	.w3(32'hbba272fb),
	.w4(32'hbaff523d),
	.w5(32'hbb955fb8),
	.w6(32'hbb3e6c4b),
	.w7(32'h3a8dd736),
	.w8(32'h3a22243b),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4929a5),
	.w1(32'h3bc3fde5),
	.w2(32'h3b352ad2),
	.w3(32'hbb97f42c),
	.w4(32'h3c0db7d3),
	.w5(32'hba4792a9),
	.w6(32'hbb6b630d),
	.w7(32'h3bbd0d19),
	.w8(32'hba94a2a1),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a419992),
	.w1(32'hbc00b060),
	.w2(32'hbc35a796),
	.w3(32'hb867c758),
	.w4(32'hbb8f27cd),
	.w5(32'hbbfd6bb4),
	.w6(32'hba26f8d3),
	.w7(32'hbbb26090),
	.w8(32'hbbe61e90),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5c2a),
	.w1(32'hba13b85c),
	.w2(32'h39baee8f),
	.w3(32'hb923f526),
	.w4(32'h3b6647cf),
	.w5(32'h3b2202fe),
	.w6(32'h3a109bb6),
	.w7(32'h3aa4237e),
	.w8(32'h3b407242),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba445ac),
	.w1(32'h3b97854d),
	.w2(32'h3c0085d7),
	.w3(32'h3bb21077),
	.w4(32'hbb8375fd),
	.w5(32'h3c46bba2),
	.w6(32'h3b65d203),
	.w7(32'hbbbf7d0f),
	.w8(32'h3bfc280b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90498f),
	.w1(32'h3a327d14),
	.w2(32'h3bac5479),
	.w3(32'hba23a9af),
	.w4(32'h3b1984dd),
	.w5(32'h3bff2af9),
	.w6(32'h3a06416f),
	.w7(32'hba9b2808),
	.w8(32'h3bffc014),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88ea17),
	.w1(32'hbc22053f),
	.w2(32'hbc2a85bf),
	.w3(32'hbba621e5),
	.w4(32'hbc56744d),
	.w5(32'hbbe3d493),
	.w6(32'hba9ea550),
	.w7(32'hbc39daa6),
	.w8(32'hbbcf6962),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6db0a),
	.w1(32'hbbb68c15),
	.w2(32'hbbe7d172),
	.w3(32'hbb187645),
	.w4(32'hbb6b397f),
	.w5(32'hbb9d4e9e),
	.w6(32'hbb8b7532),
	.w7(32'hbbbec75f),
	.w8(32'hbbc75d15),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c798d),
	.w1(32'hbc29e396),
	.w2(32'hbc137f45),
	.w3(32'hbb13d8ab),
	.w4(32'hbbe70410),
	.w5(32'hbc229f05),
	.w6(32'hbaae1efe),
	.w7(32'hbbe6e0d2),
	.w8(32'hbc172356),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14ce63),
	.w1(32'h3ac00bd8),
	.w2(32'h39a86456),
	.w3(32'hbb55b315),
	.w4(32'hba2868bb),
	.w5(32'h3b5de2e5),
	.w6(32'hbb54ac9a),
	.w7(32'h3a88da65),
	.w8(32'h3c2b4f45),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf05da),
	.w1(32'h3b21dd21),
	.w2(32'hba9c9cb3),
	.w3(32'hbb20327f),
	.w4(32'h3b4a58bf),
	.w5(32'h3b80fb58),
	.w6(32'hbad22b17),
	.w7(32'h3b5d3ae7),
	.w8(32'h3b882a38),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe812a),
	.w1(32'h3bdbf4c4),
	.w2(32'h3ba31e64),
	.w3(32'hbacff6be),
	.w4(32'h3b9d72fa),
	.w5(32'h3b018fba),
	.w6(32'h3b1c4be3),
	.w7(32'h3bba1e5f),
	.w8(32'h3baca72d),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f3e9db),
	.w1(32'hbb2beb36),
	.w2(32'hbbc5b7a4),
	.w3(32'hbaa7356b),
	.w4(32'h3b0c42bb),
	.w5(32'h3a54997d),
	.w6(32'h3b056633),
	.w7(32'hbb3a2c30),
	.w8(32'hbb848db9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb3d7c),
	.w1(32'h3befee08),
	.w2(32'h3c3660dc),
	.w3(32'hbb8c92ec),
	.w4(32'h3b5077d0),
	.w5(32'h3c82af39),
	.w6(32'hbb2212b1),
	.w7(32'h3bb48d34),
	.w8(32'h3c404b6f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4f0cb),
	.w1(32'hbb422669),
	.w2(32'hbb2c06f9),
	.w3(32'h3b391bf1),
	.w4(32'hbb3fdd77),
	.w5(32'hbb9b1f51),
	.w6(32'h3bb368f7),
	.w7(32'hbb2a8945),
	.w8(32'hbb07ecdd),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99f3f10),
	.w1(32'hbae8dde4),
	.w2(32'hbbdf3c72),
	.w3(32'hbac719e2),
	.w4(32'hbb419949),
	.w5(32'hbbc32362),
	.w6(32'hbb3e03ec),
	.w7(32'hbb8b37e2),
	.w8(32'hbb91d3f9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb65183),
	.w1(32'hbae7ba37),
	.w2(32'hba76575c),
	.w3(32'hbb95547c),
	.w4(32'hba70e53d),
	.w5(32'hb95ea65f),
	.w6(32'hbbdb68d4),
	.w7(32'h396e9b28),
	.w8(32'h3a09299e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecfa50),
	.w1(32'h3b88ea89),
	.w2(32'hbbaeaf87),
	.w3(32'h3a671255),
	.w4(32'h3ba3bd18),
	.w5(32'hbbade4cf),
	.w6(32'h3a818af3),
	.w7(32'h3b913603),
	.w8(32'hbbc212e3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc21628),
	.w1(32'hbbc49db5),
	.w2(32'hba489a7a),
	.w3(32'hbba1a2eb),
	.w4(32'hbb9d2b69),
	.w5(32'hbb727fa4),
	.w6(32'hbbb206ab),
	.w7(32'hba182178),
	.w8(32'hba3f4a91),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b401617),
	.w1(32'hba8d347c),
	.w2(32'hbb1b0b9b),
	.w3(32'h3a8d34a2),
	.w4(32'h3bde94ed),
	.w5(32'hbb4dabcd),
	.w6(32'h38bcf27f),
	.w7(32'h3c2397a3),
	.w8(32'h3ae957e8),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24a582),
	.w1(32'hbbe1f05d),
	.w2(32'hba89b2a3),
	.w3(32'hbacc4cd7),
	.w4(32'hbbcc7b3a),
	.w5(32'hbae2ef25),
	.w6(32'hbafd2149),
	.w7(32'hbc499782),
	.w8(32'hbb253525),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5d6ae),
	.w1(32'hbb7268b0),
	.w2(32'hbba69be0),
	.w3(32'hb80ee2a5),
	.w4(32'hba0107ae),
	.w5(32'hbbf46442),
	.w6(32'hbb6e83bc),
	.w7(32'hbacf4533),
	.w8(32'hbbda1b55),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb2dda),
	.w1(32'hba5ca6b9),
	.w2(32'hbb2560bb),
	.w3(32'hbb9615c7),
	.w4(32'h397281a5),
	.w5(32'hbb17bed2),
	.w6(32'hbbbc7241),
	.w7(32'hb9c31ff9),
	.w8(32'hbb4ca57b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb3cf),
	.w1(32'hba567c0c),
	.w2(32'h3b974559),
	.w3(32'hba12dd60),
	.w4(32'hbb0a7275),
	.w5(32'h3b30ee34),
	.w6(32'hbb0a4ac7),
	.w7(32'h3a96253e),
	.w8(32'h3ade4350),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae2895),
	.w1(32'h3b08e67d),
	.w2(32'hbb322a80),
	.w3(32'hbb265b7e),
	.w4(32'h3b7753b9),
	.w5(32'hbab39cc2),
	.w6(32'hb9ff0cce),
	.w7(32'h3b7d7cac),
	.w8(32'hb97b787b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb468d),
	.w1(32'hbaf38f76),
	.w2(32'hbb7df9d2),
	.w3(32'h3a0a6224),
	.w4(32'h3b161eb0),
	.w5(32'h3c4abbc5),
	.w6(32'h3b188e94),
	.w7(32'hb97c4e87),
	.w8(32'h3c0ad2fd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2fa2),
	.w1(32'h3b6aa36a),
	.w2(32'h3c0b8503),
	.w3(32'hbbec3d9c),
	.w4(32'h3a98b0d7),
	.w5(32'h3c165d10),
	.w6(32'hba952b6f),
	.w7(32'hbb508df3),
	.w8(32'h3b269edd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6090c),
	.w1(32'h3a7cc338),
	.w2(32'hb8adfe00),
	.w3(32'h3b30e0ed),
	.w4(32'hba42a811),
	.w5(32'hba004cb6),
	.w6(32'h3990d31b),
	.w7(32'hbb0eeb49),
	.w8(32'hbac37b8e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b132587),
	.w1(32'h3c154a46),
	.w2(32'h3b07a0e6),
	.w3(32'h3b81d8a6),
	.w4(32'h3c217d92),
	.w5(32'h3a854489),
	.w6(32'h3b6d51eb),
	.w7(32'h3b72d923),
	.w8(32'h3b66c701),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0abc68),
	.w1(32'hbb4f04b1),
	.w2(32'hbb1262e7),
	.w3(32'hbb0ecdf6),
	.w4(32'hba2b6b54),
	.w5(32'hbaa82212),
	.w6(32'hba41d1dc),
	.w7(32'hbae2b8ee),
	.w8(32'hbb2a1c2a),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad69cec),
	.w1(32'h3bbb041f),
	.w2(32'h3ba5091d),
	.w3(32'hbadc5871),
	.w4(32'h3bc4dda0),
	.w5(32'h3b78cac7),
	.w6(32'hbab76cd0),
	.w7(32'h3b128430),
	.w8(32'h3a8fdb09),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c1bf),
	.w1(32'hba7c0b44),
	.w2(32'h3ac02332),
	.w3(32'h3b5be471),
	.w4(32'hbb940bdb),
	.w5(32'h3b656567),
	.w6(32'hb9972e62),
	.w7(32'hbb69ddef),
	.w8(32'h3b6b56e5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52e49e),
	.w1(32'h3bf0eda1),
	.w2(32'h3c3ac453),
	.w3(32'h3bcddf5a),
	.w4(32'h3b9e13c6),
	.w5(32'h3c33bcad),
	.w6(32'h3bdaf470),
	.w7(32'h3bc73169),
	.w8(32'h3bf05bc9),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29d742),
	.w1(32'hb9d12c1a),
	.w2(32'hba8d8521),
	.w3(32'h3c1e7b3d),
	.w4(32'hbb78e61c),
	.w5(32'hbb11028d),
	.w6(32'h3c101263),
	.w7(32'hbab7a75e),
	.w8(32'hba2240c2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b9b4),
	.w1(32'h3b2a3372),
	.w2(32'h3bd58d5d),
	.w3(32'h3c08da7c),
	.w4(32'h36a62eec),
	.w5(32'h3c3bc054),
	.w6(32'h3b1c65bc),
	.w7(32'hb89317a7),
	.w8(32'h3c3e3400),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93c64),
	.w1(32'hbc12f303),
	.w2(32'hbb24c028),
	.w3(32'h3ad31014),
	.w4(32'hbb880953),
	.w5(32'hbb780728),
	.w6(32'h3b7c89ac),
	.w7(32'h3a9aa5cd),
	.w8(32'hbc2c508c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba17bac),
	.w1(32'hbc1a8228),
	.w2(32'hbc75e013),
	.w3(32'hbc29dd11),
	.w4(32'hbc85c97d),
	.w5(32'hbc0bf333),
	.w6(32'hbb162687),
	.w7(32'hbbc5e492),
	.w8(32'hbc2e7891),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc340372),
	.w1(32'hbc04efbf),
	.w2(32'hbc009d7b),
	.w3(32'hbbb5ba4b),
	.w4(32'hbba9a154),
	.w5(32'hbbb0c2e7),
	.w6(32'hbc39e0d9),
	.w7(32'hbc32851a),
	.w8(32'hbc668bbb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb7a21),
	.w1(32'hbb61beef),
	.w2(32'h3c0b42fd),
	.w3(32'hbbe1e5df),
	.w4(32'hbbc3f730),
	.w5(32'h3c68d56b),
	.w6(32'hbc17f181),
	.w7(32'h39ee1ec1),
	.w8(32'h3bdd0a60),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1d795),
	.w1(32'h3b4ff6f5),
	.w2(32'h39f5b663),
	.w3(32'hbbf00de1),
	.w4(32'h3b06ed94),
	.w5(32'h3bc1a092),
	.w6(32'h3a961e54),
	.w7(32'h3b3a978e),
	.w8(32'h3bf338ac),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e1bd9),
	.w1(32'hbb9b781d),
	.w2(32'hbba4c7d9),
	.w3(32'h3b570ba1),
	.w4(32'hbb94a956),
	.w5(32'h3c2f517e),
	.w6(32'h3bdfd694),
	.w7(32'hbbb0981a),
	.w8(32'hbc037040),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70c4aa),
	.w1(32'h3b690fd6),
	.w2(32'h3bb26d83),
	.w3(32'h38ca5c74),
	.w4(32'h3bb753cf),
	.w5(32'h3c1fdffe),
	.w6(32'hbbfcd3cf),
	.w7(32'h3b42ea4b),
	.w8(32'h3c164f62),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081815),
	.w1(32'hbba8824b),
	.w2(32'hbbe1b1b9),
	.w3(32'h3b802db6),
	.w4(32'h3bae491e),
	.w5(32'h3b441924),
	.w6(32'h3bd1a897),
	.w7(32'hbb9f1558),
	.w8(32'hb9900085),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7fc11),
	.w1(32'hba038629),
	.w2(32'hbb1d680a),
	.w3(32'hbbf13187),
	.w4(32'h3bc05b42),
	.w5(32'hbb656bb0),
	.w6(32'hbb83bd30),
	.w7(32'h3bd512d8),
	.w8(32'hbb8ad851),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a5c00),
	.w1(32'hbb4bd2f5),
	.w2(32'hbadfa45a),
	.w3(32'hbbead4bb),
	.w4(32'h39f6f9aa),
	.w5(32'hbb5a839b),
	.w6(32'hbc1cd2f8),
	.w7(32'hbb7dd2f4),
	.w8(32'hba7d0a58),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f51d88),
	.w1(32'h3b971c11),
	.w2(32'hbc431a9c),
	.w3(32'h3b88dcd0),
	.w4(32'h3c648364),
	.w5(32'h3c900813),
	.w6(32'hbbe672c4),
	.w7(32'hbb7791a8),
	.w8(32'h3a6255d8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedcfba),
	.w1(32'h3b84a33f),
	.w2(32'h3b21c52d),
	.w3(32'hbb7face6),
	.w4(32'hb99004f0),
	.w5(32'hbc1f5f25),
	.w6(32'h3b408e6b),
	.w7(32'h3b4a736a),
	.w8(32'h3b3b339c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6bbf4),
	.w1(32'h39b104be),
	.w2(32'hba0dcbf2),
	.w3(32'hbabb6e1a),
	.w4(32'hbafa85b2),
	.w5(32'hbc051135),
	.w6(32'h3b60d09b),
	.w7(32'h3b6059f7),
	.w8(32'hbb2b50e7),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85b50e),
	.w1(32'hbaeb35c2),
	.w2(32'hbbd24e6c),
	.w3(32'hbba3f509),
	.w4(32'h39c7fea9),
	.w5(32'h3bae7896),
	.w6(32'hbbd9762d),
	.w7(32'h3b2d72eb),
	.w8(32'h3b7c98cc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e7532),
	.w1(32'hba8b1bad),
	.w2(32'hbc0b1d0d),
	.w3(32'h3bc52d4a),
	.w4(32'hbb8f9752),
	.w5(32'h3b7e0830),
	.w6(32'h3ac8d3db),
	.w7(32'hbbb9cedb),
	.w8(32'hbb5d5d25),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d97f7),
	.w1(32'hbb576800),
	.w2(32'hbb4d0e29),
	.w3(32'h3beba0f2),
	.w4(32'hbc1073bb),
	.w5(32'hbaf09809),
	.w6(32'hbc4a148c),
	.w7(32'hbbc50e27),
	.w8(32'hbb7fdbe5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff4d00),
	.w1(32'hbbd4ce81),
	.w2(32'hbbb9f33f),
	.w3(32'hbbfb8f73),
	.w4(32'h3c6402ce),
	.w5(32'h3cad0485),
	.w6(32'hbc01e0cc),
	.w7(32'h3bf461a4),
	.w8(32'h3be204f4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd61653),
	.w1(32'h3c41d0d4),
	.w2(32'h3b1745b1),
	.w3(32'hbb68785e),
	.w4(32'h3b8d650c),
	.w5(32'h3c8587c1),
	.w6(32'hbb33e0d2),
	.w7(32'hbb3e93a6),
	.w8(32'hbb171307),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a904),
	.w1(32'h3c34e5c2),
	.w2(32'h399f3f29),
	.w3(32'h3bdc48e9),
	.w4(32'h3c2b2233),
	.w5(32'h3c997fc9),
	.w6(32'h3bb8a064),
	.w7(32'h3bbac3f3),
	.w8(32'hbb50a005),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ad680),
	.w1(32'hbb22b83e),
	.w2(32'hbb9bfd20),
	.w3(32'h3b9c9cba),
	.w4(32'hba2c6403),
	.w5(32'hbaf512e5),
	.w6(32'h3b791a38),
	.w7(32'hbb85c01b),
	.w8(32'hba0fe526),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdaa35d),
	.w1(32'h3a8fbc31),
	.w2(32'h3b97b840),
	.w3(32'h3b3c5cbe),
	.w4(32'h3b795199),
	.w5(32'hbb4834cc),
	.w6(32'hbc265f6e),
	.w7(32'h3bf0bd28),
	.w8(32'hbc0d01fc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec1d18),
	.w1(32'hbbaa7d80),
	.w2(32'hbbb15fdf),
	.w3(32'h3b729b83),
	.w4(32'hbb378729),
	.w5(32'hbbb21d93),
	.w6(32'hbb46c671),
	.w7(32'hbb17b6f0),
	.w8(32'hbb860487),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d85560),
	.w1(32'hb8601cd5),
	.w2(32'hbb38427c),
	.w3(32'hb982250d),
	.w4(32'hb80fac74),
	.w5(32'h3c1572e8),
	.w6(32'hba999f43),
	.w7(32'hba9b8c3d),
	.w8(32'hbc32a9d7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0ac52),
	.w1(32'hba6e1663),
	.w2(32'hbbb7e550),
	.w3(32'h3b8834f9),
	.w4(32'h3bdbcaf6),
	.w5(32'h3b220758),
	.w6(32'hbb0401cd),
	.w7(32'h3b5325ba),
	.w8(32'h39f16ae1),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae32d7),
	.w1(32'h3a737c32),
	.w2(32'h3b798343),
	.w3(32'hba08ac06),
	.w4(32'h3b0ea9c5),
	.w5(32'hbb122dcd),
	.w6(32'h3b2ea8f0),
	.w7(32'hbb383029),
	.w8(32'h3a460fb8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23b081),
	.w1(32'hbc0a851e),
	.w2(32'hbc7f2100),
	.w3(32'hbad510e3),
	.w4(32'hbb006b2f),
	.w5(32'h3ce60cbe),
	.w6(32'h3b727885),
	.w7(32'hbad0c739),
	.w8(32'hbb44e8f4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87aedc),
	.w1(32'h3b711f09),
	.w2(32'hbb944667),
	.w3(32'hbb08f565),
	.w4(32'h3c0662fe),
	.w5(32'h3b9c38cf),
	.w6(32'h3b5ff918),
	.w7(32'h3a21241b),
	.w8(32'h3b8e6a41),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc269981),
	.w1(32'hb97b3635),
	.w2(32'hbc05f2f7),
	.w3(32'hbc019e8c),
	.w4(32'hbaafd7c9),
	.w5(32'h3ac9fdaf),
	.w6(32'h3bb3378e),
	.w7(32'hbb8980ab),
	.w8(32'hbbf23274),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f35e7),
	.w1(32'hbc0e19d3),
	.w2(32'hbc3b3a7b),
	.w3(32'h3ace137b),
	.w4(32'h39908bd4),
	.w5(32'hbbf53d26),
	.w6(32'hbbb51d71),
	.w7(32'hbbb1f314),
	.w8(32'h3b075cc4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2458a),
	.w1(32'h3a9ebf10),
	.w2(32'h3c07410e),
	.w3(32'hbc07ed68),
	.w4(32'hbb123354),
	.w5(32'hbbb34cf8),
	.w6(32'hbbd45e3d),
	.w7(32'h3b142ce3),
	.w8(32'h3b2741e7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b619cfe),
	.w1(32'hbb762f51),
	.w2(32'hbb8ce326),
	.w3(32'hba38e699),
	.w4(32'hba951a76),
	.w5(32'hbca3fb13),
	.w6(32'hbb8b3258),
	.w7(32'hbb4ffbb3),
	.w8(32'hbb6c31bf),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17c888),
	.w1(32'h3911f04c),
	.w2(32'hbc370f17),
	.w3(32'hbb236e76),
	.w4(32'h3b64e0a9),
	.w5(32'h3c5c8237),
	.w6(32'hbc0a35f3),
	.w7(32'hbbbf36e4),
	.w8(32'hbb866137),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb636343),
	.w1(32'h3abb3359),
	.w2(32'hba8e6ca0),
	.w3(32'h3abed653),
	.w4(32'h3c366ab8),
	.w5(32'hba4f8865),
	.w6(32'hbae5e8e5),
	.w7(32'h3c6c22f8),
	.w8(32'h3bc0fe0d),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c024bee),
	.w1(32'h3b808f0f),
	.w2(32'hbc138fef),
	.w3(32'h3b2a9213),
	.w4(32'h3bcd4243),
	.w5(32'h3b94e1bb),
	.w6(32'h39f1e3d5),
	.w7(32'h3b8a72c9),
	.w8(32'hbbc75dd6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca5933),
	.w1(32'h395515fa),
	.w2(32'hbb12c7e0),
	.w3(32'h3bf8c485),
	.w4(32'h3c27696b),
	.w5(32'h3b62085e),
	.w6(32'hbb8b0168),
	.w7(32'h3bd87edf),
	.w8(32'h3ae72791),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73b5b7),
	.w1(32'h3a2c2187),
	.w2(32'hbb2bda56),
	.w3(32'hbb07d22b),
	.w4(32'hbb835447),
	.w5(32'h3c9a7257),
	.w6(32'hbc03cdd7),
	.w7(32'hb8f237eb),
	.w8(32'hba829ade),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93e22a),
	.w1(32'h3b1ed174),
	.w2(32'hb94564c0),
	.w3(32'h3bfb6ef7),
	.w4(32'hb99fa968),
	.w5(32'hbae9198a),
	.w6(32'h3a6d01ee),
	.w7(32'h3870f57e),
	.w8(32'hbb43fce8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a18d4),
	.w1(32'h3b27cbd5),
	.w2(32'hbbb6019e),
	.w3(32'hb99526e0),
	.w4(32'h3c025e20),
	.w5(32'hbbc12ee9),
	.w6(32'hbb6fe8c5),
	.w7(32'h3c4c94d4),
	.w8(32'h3b1541ce),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa792c3),
	.w1(32'h3bdc1bb5),
	.w2(32'h3c8acc4e),
	.w3(32'h39c7e143),
	.w4(32'hbba2bdd0),
	.w5(32'hbba8c95d),
	.w6(32'hba8ce68f),
	.w7(32'hbb0e1688),
	.w8(32'hbb5c5448),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b076e),
	.w1(32'hbb580134),
	.w2(32'hbb00fa4d),
	.w3(32'h3be7aba6),
	.w4(32'hbad1c0fe),
	.w5(32'hbbf78ae4),
	.w6(32'h3c187037),
	.w7(32'h3bfe14c8),
	.w8(32'h3b2bc8e5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd8e6),
	.w1(32'h3b5bbcb2),
	.w2(32'hbb4b684a),
	.w3(32'hbbbb54f0),
	.w4(32'hba837ad7),
	.w5(32'h3cb3f81f),
	.w6(32'h3bb10b82),
	.w7(32'hbbc29b65),
	.w8(32'hbacf2add),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb923e88),
	.w1(32'h3a39b371),
	.w2(32'h3cbb26c8),
	.w3(32'h3a927009),
	.w4(32'h38edc040),
	.w5(32'h3b49f2c1),
	.w6(32'hbb699213),
	.w7(32'h3a944401),
	.w8(32'h3ab51f4d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0852dc),
	.w1(32'hbb8fdc1f),
	.w2(32'hbb59b46c),
	.w3(32'h3ac5601a),
	.w4(32'hb8dd1c43),
	.w5(32'h3b6332a7),
	.w6(32'hba5cb303),
	.w7(32'h3bc92c57),
	.w8(32'h3aebb878),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06f096),
	.w1(32'h3b55deea),
	.w2(32'hbbea2a4d),
	.w3(32'h3b84acb9),
	.w4(32'h375cd545),
	.w5(32'hbb1140eb),
	.w6(32'hbb378ff0),
	.w7(32'h3bda95f7),
	.w8(32'h3bb71f63),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5404),
	.w1(32'hbb9b9660),
	.w2(32'hbba4055f),
	.w3(32'hbb97e12a),
	.w4(32'h39f5d3b6),
	.w5(32'h3a49bd46),
	.w6(32'hbbbd1e37),
	.w7(32'h3ae43917),
	.w8(32'hba2681c3),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0229f),
	.w1(32'h3b59357a),
	.w2(32'hbbf3ad44),
	.w3(32'h3b013f34),
	.w4(32'h3bff9835),
	.w5(32'hbb74e54c),
	.w6(32'hba3225f2),
	.w7(32'hbb053242),
	.w8(32'h3b8a7d59),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8caff4),
	.w1(32'hbbda4c73),
	.w2(32'hbbbfbcdc),
	.w3(32'h3b76e565),
	.w4(32'hbc32cc80),
	.w5(32'hbbda826c),
	.w6(32'h3b832c8f),
	.w7(32'hbc0c4c57),
	.w8(32'hbb5e3586),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95d079),
	.w1(32'h3ba253a7),
	.w2(32'hbc3f06e7),
	.w3(32'hbadd8f36),
	.w4(32'h3c4806fa),
	.w5(32'h3bed68eb),
	.w6(32'h3a82f42f),
	.w7(32'h3b9f400f),
	.w8(32'h3b6179c7),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae96766),
	.w1(32'h3ab209d5),
	.w2(32'h3ba938ca),
	.w3(32'h3b70bec9),
	.w4(32'h3bb4490a),
	.w5(32'hbc33bacd),
	.w6(32'h3c05d18c),
	.w7(32'h3b8807f0),
	.w8(32'h3b0c6186),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878f17),
	.w1(32'h3bac77d1),
	.w2(32'hbbc12d02),
	.w3(32'hbadd25dd),
	.w4(32'h3b152342),
	.w5(32'h3bd78456),
	.w6(32'h3be80754),
	.w7(32'h3b435290),
	.w8(32'h3b07601c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a925468),
	.w1(32'hbb84ded2),
	.w2(32'h3afcf97f),
	.w3(32'h3982cd3a),
	.w4(32'hbb098d82),
	.w5(32'h3b824714),
	.w6(32'h3bd1383d),
	.w7(32'h38e5c206),
	.w8(32'hbb082d51),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5998),
	.w1(32'hbbc51591),
	.w2(32'hbb15d181),
	.w3(32'h3b652053),
	.w4(32'hbb858a65),
	.w5(32'hb8ed646e),
	.w6(32'hbadaa84d),
	.w7(32'hbc007eba),
	.w8(32'hbb159f9a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba28b63),
	.w1(32'hbb68bd49),
	.w2(32'hbb530f08),
	.w3(32'hbb68554b),
	.w4(32'h36d30ce0),
	.w5(32'hbc41a8e7),
	.w6(32'hbbd665db),
	.w7(32'h3b6a3f01),
	.w8(32'hbb405a3a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eb7a2),
	.w1(32'h3b9faffd),
	.w2(32'hbc0efd9e),
	.w3(32'hba97d030),
	.w4(32'hb9d75ea4),
	.w5(32'h3bff5b00),
	.w6(32'h3c00b518),
	.w7(32'h3a8a1937),
	.w8(32'hbb9cd05b),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba526cf2),
	.w1(32'hba413e53),
	.w2(32'hbba1c891),
	.w3(32'h39fb3a55),
	.w4(32'h3b8653c5),
	.w5(32'hbb9f6f6e),
	.w6(32'hbb795f95),
	.w7(32'h3ba12141),
	.w8(32'hbb4888cc),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33b0e6),
	.w1(32'hba840a8f),
	.w2(32'hbad87599),
	.w3(32'h3a865b83),
	.w4(32'h3be8df6c),
	.w5(32'hbad1b650),
	.w6(32'hbb950a70),
	.w7(32'h3ba4a769),
	.w8(32'h3b901507),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcde2b),
	.w1(32'hba09f7eb),
	.w2(32'hbb100186),
	.w3(32'hbbcfe264),
	.w4(32'h3ac7f29d),
	.w5(32'h3b6048a0),
	.w6(32'h3a8fd8eb),
	.w7(32'hbb0cddc2),
	.w8(32'hbb8e1ebb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e254c),
	.w1(32'h3be650c4),
	.w2(32'h3b4a800a),
	.w3(32'h3b421c76),
	.w4(32'h3c136fd7),
	.w5(32'h3bba5234),
	.w6(32'hbb25aac0),
	.w7(32'h3b10415a),
	.w8(32'h3ba9ba6f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b3a16),
	.w1(32'hbbff1eef),
	.w2(32'hbbf22248),
	.w3(32'h3bdf513e),
	.w4(32'hba5b0adb),
	.w5(32'h3c182248),
	.w6(32'hbc142ede),
	.w7(32'h3b3978dd),
	.w8(32'h3b1867e7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule