module layer_6_featuremap_62(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce74128),
	.w1(32'hbaebd5c0),
	.w2(32'h3c33c525),
	.w3(32'hbbd36598),
	.w4(32'h3a59ac9b),
	.w5(32'hbbab5f68),
	.w6(32'h3853c376),
	.w7(32'h3c7b6f90),
	.w8(32'h3bd47e65),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd038b8),
	.w1(32'h3aff9d73),
	.w2(32'hbb26c681),
	.w3(32'h39fe48c1),
	.w4(32'h3b5f89ae),
	.w5(32'hb9c793fa),
	.w6(32'h3b866cc7),
	.w7(32'hbb3ac6df),
	.w8(32'h3982dc97),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf521f4),
	.w1(32'hbc8ee024),
	.w2(32'hbc8b8a87),
	.w3(32'h3c207153),
	.w4(32'hbc9d3aca),
	.w5(32'hbc94054c),
	.w6(32'h3c904734),
	.w7(32'h3c17c20b),
	.w8(32'hbb39a04f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd451e4),
	.w1(32'h3bb192da),
	.w2(32'h3a9de9f0),
	.w3(32'hbb8db1a7),
	.w4(32'hbc046971),
	.w5(32'hbb97a8cb),
	.w6(32'hbace01dd),
	.w7(32'hbc252267),
	.w8(32'hbc1f98ce),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5579fc),
	.w1(32'hbbf4aa43),
	.w2(32'h3cbeabf4),
	.w3(32'hbc94d1fd),
	.w4(32'h3c080d9a),
	.w5(32'hbc21f4b4),
	.w6(32'h3b988425),
	.w7(32'h3d931371),
	.w8(32'h3d28d7fd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bd42b),
	.w1(32'h3c6ead1e),
	.w2(32'h3cc2de79),
	.w3(32'h3c185bb1),
	.w4(32'h3c7f2b2f),
	.w5(32'h3c65d4b4),
	.w6(32'h3ca62254),
	.w7(32'h3d029654),
	.w8(32'h3ce3d3d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d163d51),
	.w1(32'hbbcc9af4),
	.w2(32'hbca18a98),
	.w3(32'hbbebd882),
	.w4(32'hbca7f7cb),
	.w5(32'hbc4c6eb4),
	.w6(32'hbca8e3f3),
	.w7(32'hbd26d2fa),
	.w8(32'hbcdf0d61),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b3b3e),
	.w1(32'h3c4e60c6),
	.w2(32'h3bd6c1d5),
	.w3(32'h3bd8f0a8),
	.w4(32'hbc30ef05),
	.w5(32'hb9083976),
	.w6(32'h3c2aa28d),
	.w7(32'hbc928a41),
	.w8(32'hbb42d0b9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41dce1),
	.w1(32'hbc996a5b),
	.w2(32'hbc8d0149),
	.w3(32'hbbbff0ca),
	.w4(32'hbbfef994),
	.w5(32'hbb4014c5),
	.w6(32'hbad3a420),
	.w7(32'h3c2ece6c),
	.w8(32'h3c217825),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93f335),
	.w1(32'h3c18ed2e),
	.w2(32'h3c7365d8),
	.w3(32'h3c3dfe0a),
	.w4(32'h3cbe61ca),
	.w5(32'h3c49db46),
	.w6(32'h3c761b96),
	.w7(32'h3cd248f7),
	.w8(32'h3c5434b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd4ec),
	.w1(32'hbadf4b62),
	.w2(32'h3b9ff23f),
	.w3(32'hbb428caa),
	.w4(32'hbc34334d),
	.w5(32'hbb1e1d7c),
	.w6(32'h3c0a1373),
	.w7(32'hba0dc7d9),
	.w8(32'h3c79a4f3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf72f0),
	.w1(32'hbc815fe8),
	.w2(32'hbb6bb0fb),
	.w3(32'hbb95fa5a),
	.w4(32'h3bb14167),
	.w5(32'hbbb7afb2),
	.w6(32'hbb3794ee),
	.w7(32'h3c0e3bf9),
	.w8(32'h3ba95c71),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75be90),
	.w1(32'hbbd7fdb3),
	.w2(32'h3bf6116e),
	.w3(32'h3a73fab7),
	.w4(32'h3c80055b),
	.w5(32'h3a22b5ee),
	.w6(32'hb9ecf09e),
	.w7(32'h3c43c0ec),
	.w8(32'h3a5e8bb3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3281d2),
	.w1(32'hbc59d504),
	.w2(32'hbbeddbfb),
	.w3(32'hbb14ed6e),
	.w4(32'hbd2de0a9),
	.w5(32'hbce77b9b),
	.w6(32'hbb4da057),
	.w7(32'hbc4568b8),
	.w8(32'hbbb2bbc0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9b952),
	.w1(32'h3b880b68),
	.w2(32'h3bdcf5fa),
	.w3(32'h3bd9c72d),
	.w4(32'h3c25453d),
	.w5(32'h3be287a2),
	.w6(32'h3a95ef6d),
	.w7(32'h3ba5f238),
	.w8(32'hbbaac045),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6eab13),
	.w1(32'h389f6caf),
	.w2(32'h3c14fc77),
	.w3(32'hbc04bd77),
	.w4(32'hbbd76a64),
	.w5(32'hbb293d7c),
	.w6(32'hbb77fed9),
	.w7(32'hba52a25c),
	.w8(32'h3c1179f8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9b5fb),
	.w1(32'hbb05c4c6),
	.w2(32'hbb11c6f5),
	.w3(32'hba3dacc2),
	.w4(32'hbd2dd27c),
	.w5(32'hbd0e7b39),
	.w6(32'h3c850057),
	.w7(32'hbc84247c),
	.w8(32'hbcd52b0e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc065b19),
	.w1(32'hbb99562c),
	.w2(32'h3b95c3dd),
	.w3(32'hb93be672),
	.w4(32'h3c48c7d9),
	.w5(32'h3c112d6b),
	.w6(32'hbb093be7),
	.w7(32'h3bf807b9),
	.w8(32'h3bfe0798),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8554),
	.w1(32'h3bb3f652),
	.w2(32'h3b2c728b),
	.w3(32'h398649fc),
	.w4(32'hbb8b19ee),
	.w5(32'hbb0aac4a),
	.w6(32'h39024cf8),
	.w7(32'hbbaf9a58),
	.w8(32'hbb9bcab8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe19a58),
	.w1(32'hbbd5ab00),
	.w2(32'hbc1dac5b),
	.w3(32'hbbca4e13),
	.w4(32'hbba13de7),
	.w5(32'hbc16db86),
	.w6(32'hbc0879c0),
	.w7(32'h3a31754e),
	.w8(32'hbc180445),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc249a27),
	.w1(32'hbacf908a),
	.w2(32'hbbd8dfd6),
	.w3(32'hbb746aa2),
	.w4(32'hbbd12acc),
	.w5(32'h3819ec9b),
	.w6(32'hbb95feb2),
	.w7(32'hbc1d43f8),
	.w8(32'hbb84755a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01de1a),
	.w1(32'hbc936b43),
	.w2(32'hbae4e07e),
	.w3(32'hbc27279f),
	.w4(32'hbd036d23),
	.w5(32'hbc8129a9),
	.w6(32'h3be1e524),
	.w7(32'h3ad5ad30),
	.w8(32'h3b4049a9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b152a3a),
	.w1(32'h3c5c6272),
	.w2(32'h3c4af14a),
	.w3(32'h3b376db2),
	.w4(32'h3a85f027),
	.w5(32'hbd1164a9),
	.w6(32'h3ce36cf2),
	.w7(32'h3c65a69f),
	.w8(32'hbd2f9bef),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7dd3c7),
	.w1(32'hbd44462f),
	.w2(32'hbd83adeb),
	.w3(32'hbc10aa77),
	.w4(32'hbd1c6d79),
	.w5(32'hbd4cff7a),
	.w6(32'hbcf89748),
	.w7(32'hbd411487),
	.w8(32'hbd48cf75),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9b0cf1),
	.w1(32'hbcaba711),
	.w2(32'hbcd396db),
	.w3(32'hbd3df596),
	.w4(32'hbd99a299),
	.w5(32'hbd4a3bda),
	.w6(32'h3c0cac61),
	.w7(32'hbc83a0d4),
	.w8(32'hbcd8f194),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc347218),
	.w1(32'h3c012f70),
	.w2(32'h3c9def0c),
	.w3(32'h3aa5c490),
	.w4(32'h3a9be02c),
	.w5(32'h3b137a41),
	.w6(32'h3c2dcd50),
	.w7(32'h3c1e0639),
	.w8(32'hbb4fca09),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba788e),
	.w1(32'hbc32479d),
	.w2(32'h3c0ef045),
	.w3(32'hbbeac353),
	.w4(32'hbca8a673),
	.w5(32'hbcf9d213),
	.w6(32'hbc49fbc9),
	.w7(32'h3c00f280),
	.w8(32'h3a56bb51),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4b93),
	.w1(32'hbc278efd),
	.w2(32'hbc8c24bf),
	.w3(32'hbc2f0b55),
	.w4(32'hbcad3ffa),
	.w5(32'hbbb39d7e),
	.w6(32'hbc5b2b9e),
	.w7(32'hbce0eaa0),
	.w8(32'hbc63ba21),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4ffd2),
	.w1(32'h3a7c803f),
	.w2(32'hbad4e247),
	.w3(32'h3b6177ea),
	.w4(32'h3a141a3a),
	.w5(32'h3b9c3754),
	.w6(32'h3a8867ea),
	.w7(32'hbad684bf),
	.w8(32'h3ab54060),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4e7a),
	.w1(32'h3b2ea588),
	.w2(32'h3c4d1a10),
	.w3(32'h3ac0611a),
	.w4(32'h3d986e89),
	.w5(32'h3d8659b4),
	.w6(32'h3cf6136f),
	.w7(32'hbcc4ec45),
	.w8(32'hbcccee77),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9461e6),
	.w1(32'h3c6cf7d3),
	.w2(32'h3d04860c),
	.w3(32'hbc80f3bd),
	.w4(32'hbd04c396),
	.w5(32'hbca9e06b),
	.w6(32'hbc64e3b3),
	.w7(32'hbc9c020b),
	.w8(32'hbc87c21a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c886d2d),
	.w1(32'hbc241dbf),
	.w2(32'h3c5ba6ad),
	.w3(32'hbc61b852),
	.w4(32'h3c27a63e),
	.w5(32'hbb6f0dbe),
	.w6(32'h3b164923),
	.w7(32'h3d026665),
	.w8(32'h3cc58a88),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80d1cf),
	.w1(32'hbc14f69d),
	.w2(32'hbaa99b67),
	.w3(32'hbb731cdd),
	.w4(32'h3ae2d220),
	.w5(32'hbc340ed0),
	.w6(32'hbbb54b7b),
	.w7(32'h3b914597),
	.w8(32'hbc108ab8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5eb3a6),
	.w1(32'h3b5c15d0),
	.w2(32'h3c31633f),
	.w3(32'h3bd7138e),
	.w4(32'hbb2045f8),
	.w5(32'hbc333fed),
	.w6(32'h3c2b4016),
	.w7(32'h3b967399),
	.w8(32'hbc27d122),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b4bd),
	.w1(32'h3c01629f),
	.w2(32'h3c49be16),
	.w3(32'h3be758b2),
	.w4(32'h3c3f8fa5),
	.w5(32'h3bd74eca),
	.w6(32'h3c81cff3),
	.w7(32'h3ca87f73),
	.w8(32'h3c567c82),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74499d),
	.w1(32'h3be42684),
	.w2(32'h3c830db1),
	.w3(32'h3b2154d5),
	.w4(32'h3b93093f),
	.w5(32'h3c74ba86),
	.w6(32'h39d7c2e4),
	.w7(32'hbb98691b),
	.w8(32'hbc4da6af),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90aa63),
	.w1(32'hbacb5b5a),
	.w2(32'h3c3c1120),
	.w3(32'hbc09cb38),
	.w4(32'hbb957cf2),
	.w5(32'hbbc60486),
	.w6(32'hba091572),
	.w7(32'h3c6e2cbc),
	.w8(32'h3b8f38dc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1161c8),
	.w1(32'hb99bfeb9),
	.w2(32'hbb79e917),
	.w3(32'hbc078ef4),
	.w4(32'hbb42c8d3),
	.w5(32'h3be73721),
	.w6(32'hbb7f7e22),
	.w7(32'hbc7f2543),
	.w8(32'hbbf3f28d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbea04),
	.w1(32'h3af5f7ec),
	.w2(32'hbbcea918),
	.w3(32'hbb82156b),
	.w4(32'hbc46031c),
	.w5(32'hbbb1a0ab),
	.w6(32'hbc44a618),
	.w7(32'hbbd7ec84),
	.w8(32'hbb5669a9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd55cc62),
	.w1(32'hbd434520),
	.w2(32'h3c64cbe5),
	.w3(32'hbc1648ac),
	.w4(32'hbd44a961),
	.w5(32'hbc9a64a7),
	.w6(32'hb99cc788),
	.w7(32'h3c44f119),
	.w8(32'h3d2bc948),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d012641),
	.w1(32'h3c91c780),
	.w2(32'h3c3c330f),
	.w3(32'hbc6ea8d1),
	.w4(32'hbb3f4734),
	.w5(32'h3cc836f8),
	.w6(32'hba98ac60),
	.w7(32'hbbba3d70),
	.w8(32'hbc861093),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8d12d),
	.w1(32'h3c11b5b8),
	.w2(32'h3b697b9c),
	.w3(32'hbbe08de5),
	.w4(32'hbb6f593f),
	.w5(32'h3b2f8a91),
	.w6(32'hbc1b3401),
	.w7(32'hbcbb4b16),
	.w8(32'hbc513b3c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb638d3d),
	.w1(32'h3a83d924),
	.w2(32'h3c30922b),
	.w3(32'hbb565ff1),
	.w4(32'h3b9d3d57),
	.w5(32'h3b64c599),
	.w6(32'h3a5deccd),
	.w7(32'h3c7dfa95),
	.w8(32'h3c06cb57),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d74a658),
	.w1(32'h3d2e9a32),
	.w2(32'h3d0f83b7),
	.w3(32'h3c736f9d),
	.w4(32'h3d5967f5),
	.w5(32'h3d99308a),
	.w6(32'h3d2838aa),
	.w7(32'hbd055e4f),
	.w8(32'hbc9fd1f0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca7eca3),
	.w1(32'hbcdf811a),
	.w2(32'hbc140a73),
	.w3(32'h3b926aea),
	.w4(32'hbcc0ee8a),
	.w5(32'hbc205364),
	.w6(32'h3c0f3859),
	.w7(32'h3b9d93ea),
	.w8(32'h3c29ee3f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7978c2),
	.w1(32'h3c216ca5),
	.w2(32'h3b4fbca7),
	.w3(32'hbc8c19c4),
	.w4(32'hbb85788e),
	.w5(32'hbb2bf8a8),
	.w6(32'hbb394bf2),
	.w7(32'h3c4ef67d),
	.w8(32'h3b2e03d7),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1792de),
	.w1(32'h3c8e789c),
	.w2(32'h3ab079dd),
	.w3(32'h3b5e58c6),
	.w4(32'h3c4ca09f),
	.w5(32'h3c8275c9),
	.w6(32'h3c05ad17),
	.w7(32'hbc02e458),
	.w8(32'hbb2c1134),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd91f99),
	.w1(32'hbd365c1c),
	.w2(32'hbd16c769),
	.w3(32'hbd266778),
	.w4(32'hbd60752b),
	.w5(32'hbd541b02),
	.w6(32'hbcd1ebd1),
	.w7(32'hbd125f31),
	.w8(32'hbd1f1203),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e4427),
	.w1(32'h3bb4808c),
	.w2(32'h3b4fbba3),
	.w3(32'h3b79f4e1),
	.w4(32'h3b2ead17),
	.w5(32'h3bc0600f),
	.w6(32'h3b5b0842),
	.w7(32'h3a5c123c),
	.w8(32'h3b7cc328),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b9bd3),
	.w1(32'hbcc073b5),
	.w2(32'hbbe38ea9),
	.w3(32'hbc77e82b),
	.w4(32'hbd33e8c4),
	.w5(32'hbd78606f),
	.w6(32'hba8c60a5),
	.w7(32'h3b3208f0),
	.w8(32'hbc9bcdfa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cfb3e),
	.w1(32'h3bc21dea),
	.w2(32'h3b0f13f0),
	.w3(32'h3b720914),
	.w4(32'hbabf1c5d),
	.w5(32'h3ae0255d),
	.w6(32'h3bcaaa52),
	.w7(32'hbc30e0b4),
	.w8(32'hbc0524a1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c569f8e),
	.w1(32'h3d22cca8),
	.w2(32'h3b812e6a),
	.w3(32'h3cc5bb98),
	.w4(32'hbab92b52),
	.w5(32'h3b8684e4),
	.w6(32'h3ca9ff17),
	.w7(32'hbc685edf),
	.w8(32'hbc41d2ab),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2072a3),
	.w1(32'hbcb8d673),
	.w2(32'hbc9cbb9a),
	.w3(32'hba821a86),
	.w4(32'hbd4b64e0),
	.w5(32'hbcf00749),
	.w6(32'h3b0fe555),
	.w7(32'hbcc9e8fa),
	.w8(32'hbc0e26a4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a34b8),
	.w1(32'hbcd400a0),
	.w2(32'hbd2f2c00),
	.w3(32'hbcf1c803),
	.w4(32'hbd16b466),
	.w5(32'hbccb55d2),
	.w6(32'hbcffa2f1),
	.w7(32'hbd3e91d4),
	.w8(32'hbd189189),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdefa62),
	.w1(32'hbb9db56c),
	.w2(32'hbc3bd00c),
	.w3(32'h3c04d943),
	.w4(32'h3bc7e266),
	.w5(32'h3b96c74e),
	.w6(32'h3ad13703),
	.w7(32'hbc2f76ad),
	.w8(32'hbc0901f6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b2136),
	.w1(32'h3c97bac4),
	.w2(32'h3c5f93b2),
	.w3(32'hbc507e56),
	.w4(32'hbc8c70cf),
	.w5(32'hb9f217b7),
	.w6(32'h3b3a58d7),
	.w7(32'hbc9a6b88),
	.w8(32'hbc86a236),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55ab42),
	.w1(32'hbba81bc3),
	.w2(32'hbbcd48b8),
	.w3(32'hbc02d28d),
	.w4(32'h39f6a065),
	.w5(32'h3bba45a3),
	.w6(32'hbc0fec0f),
	.w7(32'hbb881cbd),
	.w8(32'h3c0ddfac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a894bcf),
	.w1(32'h3c2393f0),
	.w2(32'h3c9c7214),
	.w3(32'hb8fb2b62),
	.w4(32'hbbba636e),
	.w5(32'hbb1c3d19),
	.w6(32'h3c7bda48),
	.w7(32'h3b3429eb),
	.w8(32'hbd021390),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf0826),
	.w1(32'hbb581ee9),
	.w2(32'hbb5cdeaf),
	.w3(32'hbb501be4),
	.w4(32'hbb405c57),
	.w5(32'hbaf761f1),
	.w6(32'hbb0c1ce1),
	.w7(32'hbb808b75),
	.w8(32'hbb1aa904),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd20bf35),
	.w1(32'hbc420d8d),
	.w2(32'hbc067c9e),
	.w3(32'hbc2994eb),
	.w4(32'hbd3c67a8),
	.w5(32'hbcdddcb8),
	.w6(32'h3d161578),
	.w7(32'h3cb1513e),
	.w8(32'h3c800505),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85b5eb),
	.w1(32'hbbea68ee),
	.w2(32'hbaeacaf6),
	.w3(32'hbadc5704),
	.w4(32'hbc018a20),
	.w5(32'hbc67ae3e),
	.w6(32'hba6d1c8f),
	.w7(32'hbab2acac),
	.w8(32'hbc676838),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc892464),
	.w1(32'hbbf3b733),
	.w2(32'hbd114afc),
	.w3(32'hbcf7ab47),
	.w4(32'hbd86e612),
	.w5(32'hbcb42b96),
	.w6(32'hbc735a19),
	.w7(32'hbd43f7cb),
	.w8(32'hbd08ab7e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96c706),
	.w1(32'hbd3f2c6d),
	.w2(32'hbd9d54f3),
	.w3(32'h3c0cc56a),
	.w4(32'h3d563857),
	.w5(32'h3d13aa17),
	.w6(32'hbccd5975),
	.w7(32'h3ab61872),
	.w8(32'h3d8530fc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf014f8),
	.w1(32'hbc858aa6),
	.w2(32'h3b9c94b0),
	.w3(32'hba1a4120),
	.w4(32'h3b34b4e5),
	.w5(32'hbc043360),
	.w6(32'hbae0985f),
	.w7(32'h3c6f261b),
	.w8(32'hbab51882),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule