module layer_8_featuremap_56(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bea2c5),
	.w1(32'hb812297b),
	.w2(32'h38d927ea),
	.w3(32'h38fff556),
	.w4(32'h38ed41a8),
	.w5(32'hb6b277c8),
	.w6(32'hb8a35989),
	.w7(32'hb8fda83d),
	.w8(32'hb9dc3984),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd2642),
	.w1(32'h38c157dd),
	.w2(32'h38deb254),
	.w3(32'h3959ae34),
	.w4(32'h3896a13e),
	.w5(32'h38b2c3ca),
	.w6(32'h395180b2),
	.w7(32'h388bf551),
	.w8(32'hb4edf96e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3832738d),
	.w1(32'h38a92fa2),
	.w2(32'h3950596b),
	.w3(32'h396a7261),
	.w4(32'h3909df7f),
	.w5(32'h38cc7fa8),
	.w6(32'h39007fb6),
	.w7(32'h378be4f4),
	.w8(32'h3718a767),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba795a),
	.w1(32'h39790f61),
	.w2(32'h399fa444),
	.w3(32'h38a33d27),
	.w4(32'h3883b988),
	.w5(32'hb6f930b6),
	.w6(32'h39a65e03),
	.w7(32'h396164e5),
	.w8(32'h3841f032),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922dfac),
	.w1(32'h391347e7),
	.w2(32'h393546a4),
	.w3(32'h38fd1df0),
	.w4(32'h38b4b14e),
	.w5(32'hb70a6f69),
	.w6(32'h3984c7f2),
	.w7(32'h39307456),
	.w8(32'hb8c0dffe),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bc93f),
	.w1(32'h399b495c),
	.w2(32'h392fcd55),
	.w3(32'hb8aacee6),
	.w4(32'hb96a12fe),
	.w5(32'hb98b38f5),
	.w6(32'h39420c2f),
	.w7(32'hb91bdbc2),
	.w8(32'hb9b50326),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70d3876),
	.w1(32'hb5d41949),
	.w2(32'hb5fbbbcb),
	.w3(32'hb6dc54fd),
	.w4(32'h34abdbc1),
	.w5(32'hb452110e),
	.w6(32'hb6f31b38),
	.w7(32'hb56999d2),
	.w8(32'hb512d36c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391733bb),
	.w1(32'hb9092d08),
	.w2(32'hb802a610),
	.w3(32'h39c04761),
	.w4(32'hb8c9a799),
	.w5(32'hb99452ed),
	.w6(32'h39a5ab04),
	.w7(32'h37895c73),
	.w8(32'hb9537b8a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c372b1),
	.w1(32'h38396a4a),
	.w2(32'h38855052),
	.w3(32'hb870d54e),
	.w4(32'hb8da4974),
	.w5(32'hb9403e77),
	.w6(32'h3920677d),
	.w7(32'hb910be9f),
	.w8(32'hb9b1b760),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cdff44),
	.w1(32'h383bc38c),
	.w2(32'h384b4a4a),
	.w3(32'h39da0f8f),
	.w4(32'h39ab0c24),
	.w5(32'h39491599),
	.w6(32'h3934abd7),
	.w7(32'h389552d6),
	.w8(32'hb997bcd1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386da784),
	.w1(32'hb828043b),
	.w2(32'h3958c6e0),
	.w3(32'h3855c368),
	.w4(32'hb905224d),
	.w5(32'hb90f0fc8),
	.w6(32'h3873cc4d),
	.w7(32'hb883c9ea),
	.w8(32'hb9b6256d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1d0d6),
	.w1(32'h395635c8),
	.w2(32'h38e74b4b),
	.w3(32'h3a0d397a),
	.w4(32'h393cb903),
	.w5(32'h39529d42),
	.w6(32'h39a3e437),
	.w7(32'h385be6dd),
	.w8(32'hb74949ee),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcf9e6),
	.w1(32'h39811beb),
	.w2(32'h399e79a0),
	.w3(32'h399024a7),
	.w4(32'h39169a1a),
	.w5(32'h395b3a2c),
	.w6(32'h398d2050),
	.w7(32'h389cb860),
	.w8(32'h38d1e24c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c9c036),
	.w1(32'hb5e82f94),
	.w2(32'hb5cea1e3),
	.w3(32'hb6478d7a),
	.w4(32'h35f7de8f),
	.w5(32'hb427109f),
	.w6(32'hb619189e),
	.w7(32'h3614010b),
	.w8(32'hb4b333a8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6afa205),
	.w1(32'hb3a37dd4),
	.w2(32'hb5266fab),
	.w3(32'hb661cd6b),
	.w4(32'h35d21380),
	.w5(32'h35543ad1),
	.w6(32'hb6494bb6),
	.w7(32'h3599fe16),
	.w8(32'h344f3c72),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35a3f5dc),
	.w1(32'hb7b5b1ce),
	.w2(32'hb6bb855c),
	.w3(32'h36460076),
	.w4(32'hb7e54447),
	.w5(32'hb68d2e42),
	.w6(32'hb86039a3),
	.w7(32'hb872335f),
	.w8(32'hb87eefeb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8115afc),
	.w1(32'hb8b8e29f),
	.w2(32'hb8b7dcfa),
	.w3(32'hb81e6e06),
	.w4(32'hb8e119b1),
	.w5(32'hb89ed412),
	.w6(32'h36379256),
	.w7(32'hb88366e6),
	.w8(32'hb866a35f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae3a5a),
	.w1(32'h39ae32f3),
	.w2(32'h39938b5b),
	.w3(32'h39efb20b),
	.w4(32'h39f825f3),
	.w5(32'h3a1ecaea),
	.w6(32'h39cb7cb7),
	.w7(32'h3948f556),
	.w8(32'h39c91d58),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997baf2),
	.w1(32'hb9c4f53f),
	.w2(32'h39631eb3),
	.w3(32'h3a127634),
	.w4(32'hb8daeb0a),
	.w5(32'hb9e9bea8),
	.w6(32'hb91cf6f7),
	.w7(32'hba05fa53),
	.w8(32'hba3a1071),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2abe7),
	.w1(32'h380d6fd0),
	.w2(32'h39d9a63b),
	.w3(32'h388839b9),
	.w4(32'hb9aa5e93),
	.w5(32'hb9c5b511),
	.w6(32'hb62b810b),
	.w7(32'hb9507383),
	.w8(32'hb98e5532),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38313c2f),
	.w1(32'hb9b4fa6d),
	.w2(32'hb9edaf7e),
	.w3(32'hb8ee762b),
	.w4(32'hba0e9a46),
	.w5(32'hba2f6fa1),
	.w6(32'hb892e07a),
	.w7(32'hb9a21628),
	.w8(32'hba0e1911),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1d760),
	.w1(32'h38cb8b3f),
	.w2(32'h394888cc),
	.w3(32'hb81ef251),
	.w4(32'hb8af5eaf),
	.w5(32'hb8aee1f5),
	.w6(32'h3841305f),
	.w7(32'h37fc85dc),
	.w8(32'h3821ccd9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c08f8),
	.w1(32'hb9c7399f),
	.w2(32'hb93e8770),
	.w3(32'hb9461437),
	.w4(32'hb989fa4e),
	.w5(32'hba106b2c),
	.w6(32'hb9b95d31),
	.w7(32'hb9d23ed1),
	.w8(32'hba84738f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ccbb2),
	.w1(32'hb847cbfd),
	.w2(32'hb717382c),
	.w3(32'hb885961b),
	.w4(32'hb83f0bc9),
	.w5(32'h361accf0),
	.w6(32'hb784f98b),
	.w7(32'hb904d262),
	.w8(32'hb90bf2d9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b037be),
	.w1(32'hb6fee554),
	.w2(32'h36a245b0),
	.w3(32'hb6d8b044),
	.w4(32'hb7cb00b2),
	.w5(32'hb76c86c3),
	.w6(32'h368d6f55),
	.w7(32'hb6320f52),
	.w8(32'h366d23bb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a8a18),
	.w1(32'hb917ee0b),
	.w2(32'hb9aeef6a),
	.w3(32'h39e87ceb),
	.w4(32'hb89df26a),
	.w5(32'hb9ac41d8),
	.w6(32'h39c5f9b3),
	.w7(32'hb88c80ed),
	.w8(32'hb9a83e25),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362c7090),
	.w1(32'h369ea574),
	.w2(32'h37072d66),
	.w3(32'h35805773),
	.w4(32'h36823f94),
	.w5(32'h37082741),
	.w6(32'h365f6eb3),
	.w7(32'h36a0e4b8),
	.w8(32'h3710c726),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9499d9f),
	.w1(32'hbb88c96e),
	.w2(32'hbb592147),
	.w3(32'h3accb089),
	.w4(32'hbb2f3476),
	.w5(32'hbb388198),
	.w6(32'h39d4a30e),
	.w7(32'hb9fc7ce3),
	.w8(32'h39ccb082),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394ffe58),
	.w1(32'hb88fc0be),
	.w2(32'h35d93819),
	.w3(32'h39437b00),
	.w4(32'h3736aa4e),
	.w5(32'hb84313da),
	.w6(32'h393d30b8),
	.w7(32'hb904bdbc),
	.w8(32'hb95e2839),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901e7cb),
	.w1(32'h3884d9a4),
	.w2(32'h38b4a0f5),
	.w3(32'h3870df5b),
	.w4(32'hb79ad374),
	.w5(32'hb615f0fa),
	.w6(32'h3902d601),
	.w7(32'h37cdede1),
	.w8(32'h355c8e84),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dacac1),
	.w1(32'h38a3907c),
	.w2(32'h38c36b6d),
	.w3(32'h37c3a05e),
	.w4(32'hb74ce25c),
	.w5(32'h38cbbc2a),
	.w6(32'h37ba0c9d),
	.w7(32'h3719e458),
	.w8(32'h388792db),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39480adc),
	.w1(32'hb738d1ff),
	.w2(32'h36e0773f),
	.w3(32'hb7ba45ad),
	.w4(32'hb984b6bd),
	.w5(32'hb9c88a1a),
	.w6(32'h3797cf1c),
	.w7(32'hb957631c),
	.w8(32'hb999a067),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb789ac8f),
	.w1(32'hb694c31b),
	.w2(32'hb62bbdb3),
	.w3(32'hb769bde5),
	.w4(32'hb63db3f9),
	.w5(32'hb49d67c3),
	.w6(32'hb732b864),
	.w7(32'hb61a5764),
	.w8(32'hb5df4bc6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7846241),
	.w1(32'hb714d140),
	.w2(32'hb6ec3d87),
	.w3(32'hb74c2d03),
	.w4(32'hb6d9b1ea),
	.w5(32'hb67706c0),
	.w6(32'hb74bf6df),
	.w7(32'hb6ce1c33),
	.w8(32'hb68833fd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395753cf),
	.w1(32'h39717b86),
	.w2(32'h398a309c),
	.w3(32'hb8b900d7),
	.w4(32'h37d27871),
	.w5(32'h38bcd6e8),
	.w6(32'h38ea38c9),
	.w7(32'h397534db),
	.w8(32'h39848370),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34ba8eaa),
	.w1(32'hb9acefd7),
	.w2(32'hb9951796),
	.w3(32'h3999c026),
	.w4(32'hb7f50748),
	.w5(32'hb9695d2d),
	.w6(32'h3921ff63),
	.w7(32'hb735051e),
	.w8(32'hb92d64f6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb52c61a8),
	.w1(32'hb5164456),
	.w2(32'h369815eb),
	.w3(32'h35a75c85),
	.w4(32'h34016b74),
	.w5(32'hb640ca11),
	.w6(32'hb6338653),
	.w7(32'h3642f876),
	.w8(32'hb644cc02),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a18bd),
	.w1(32'h395274ca),
	.w2(32'h3935a5c4),
	.w3(32'h395257fb),
	.w4(32'h38c5a95f),
	.w5(32'h37a90081),
	.w6(32'h397e8a78),
	.w7(32'h39290897),
	.w8(32'h389c61e4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6736180),
	.w1(32'h36cfb06b),
	.w2(32'h35e3e88a),
	.w3(32'hb675b6e7),
	.w4(32'h37165549),
	.w5(32'h37064c67),
	.w6(32'hb694bfbc),
	.w7(32'h3754fee8),
	.w8(32'h36ba57c0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6606f98),
	.w1(32'h37205989),
	.w2(32'h37964aca),
	.w3(32'hb7620c0e),
	.w4(32'hb79b0fb3),
	.w5(32'hb715391b),
	.w6(32'hb7908474),
	.w7(32'hb6d41355),
	.w8(32'h369285cf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab12100),
	.w1(32'h39ab1e1b),
	.w2(32'hb8fe9460),
	.w3(32'h3a8d1b02),
	.w4(32'hb6321595),
	.w5(32'hb9b005f3),
	.w6(32'h3a1e8104),
	.w7(32'hb9e91080),
	.w8(32'hba916d6d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e758b0),
	.w1(32'hb9904e15),
	.w2(32'hb974c226),
	.w3(32'hb81634e5),
	.w4(32'hb996f53a),
	.w5(32'hb9712b3c),
	.w6(32'hb837b628),
	.w7(32'hb97cffbc),
	.w8(32'hb93e79e6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368ddf6f),
	.w1(32'hb819141d),
	.w2(32'hb80cadce),
	.w3(32'hb76669cd),
	.w4(32'hb82bdfc3),
	.w5(32'hb84bd91f),
	.w6(32'h372ddc03),
	.w7(32'hb6f406d9),
	.w8(32'h3741e04c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39298479),
	.w1(32'hb8a587f5),
	.w2(32'hb81aadb6),
	.w3(32'hb794a338),
	.w4(32'hb98fd8c6),
	.w5(32'hb9ac0fbe),
	.w6(32'h37dab4ac),
	.w7(32'hb92d0646),
	.w8(32'hb9a139fe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e7ae51),
	.w1(32'hb95059b0),
	.w2(32'h3916e2bd),
	.w3(32'hb82f7bc3),
	.w4(32'hb9a4745d),
	.w5(32'hb99889d9),
	.w6(32'hb8c90917),
	.w7(32'hb9b613bf),
	.w8(32'hba079518),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e62fb),
	.w1(32'hb972c5e1),
	.w2(32'hb8c19d3b),
	.w3(32'h37f95d8c),
	.w4(32'hb9a8e950),
	.w5(32'hb9489847),
	.w6(32'hb880e4d7),
	.w7(32'hb9ae1205),
	.w8(32'hb9921a97),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69df137),
	.w1(32'hb6065cb9),
	.w2(32'hb60a1f01),
	.w3(32'hb6403f7d),
	.w4(32'h330aa9b4),
	.w5(32'hb4c43fdf),
	.w6(32'hb63f69f4),
	.w7(32'hb369a309),
	.w8(32'hb4ba8966),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9938f64),
	.w1(32'hb9ab03bf),
	.w2(32'hb9318f27),
	.w3(32'hb95415f7),
	.w4(32'hba048f1e),
	.w5(32'hb9f604eb),
	.w6(32'hb9bb1822),
	.w7(32'hba054eb4),
	.w8(32'hb9f515d6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39458349),
	.w1(32'h38ea3f53),
	.w2(32'h38de7e03),
	.w3(32'h391e7de9),
	.w4(32'h387cbf92),
	.w5(32'h37a4d0b7),
	.w6(32'h39682154),
	.w7(32'h38a597c1),
	.w8(32'hb67765b8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a099c8),
	.w1(32'h38f4269d),
	.w2(32'h3929e068),
	.w3(32'h39464e30),
	.w4(32'h37b64a2a),
	.w5(32'h37a6a1ac),
	.w6(32'h398dbc26),
	.w7(32'h3886ca4f),
	.w8(32'hb894d495),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39290356),
	.w1(32'hb9b1bfb0),
	.w2(32'hb99f0b6b),
	.w3(32'hb88b08ef),
	.w4(32'hba2eeb47),
	.w5(32'hba19cd1e),
	.w6(32'hb917ddce),
	.w7(32'hb9f6c32c),
	.w8(32'hb973a2aa),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388122af),
	.w1(32'hba1fb6e7),
	.w2(32'hb9acf0cd),
	.w3(32'hb9ead655),
	.w4(32'hba94958d),
	.w5(32'hba799ac1),
	.w6(32'h3899be6a),
	.w7(32'hba70e2f3),
	.w8(32'hba894e9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388d0484),
	.w1(32'hb871d21d),
	.w2(32'h38e059f6),
	.w3(32'hb76e3514),
	.w4(32'hb912d2f1),
	.w5(32'hb97537d6),
	.w6(32'h381a58d6),
	.w7(32'hb90b5369),
	.w8(32'hb9a88117),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f9fab),
	.w1(32'h3908a3f7),
	.w2(32'h391ba74d),
	.w3(32'h3a037cfd),
	.w4(32'h39f10df3),
	.w5(32'h39d128ae),
	.w6(32'hb75ead34),
	.w7(32'h388b33d2),
	.w8(32'hb98d505d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77bc755),
	.w1(32'hb6d98eb7),
	.w2(32'hb7242785),
	.w3(32'hb717c68c),
	.w4(32'h3582a2ab),
	.w5(32'hb58244ad),
	.w6(32'hb73f7a4b),
	.w7(32'h35d39105),
	.w8(32'hb6801a65),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6bcbb15),
	.w1(32'hb996b03d),
	.w2(32'hb8769b9f),
	.w3(32'h3a195929),
	.w4(32'hb89d7b2b),
	.w5(32'hb9653273),
	.w6(32'hb9eaccce),
	.w7(32'hb9a9d9c0),
	.w8(32'hba4258cd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ee7b18),
	.w1(32'hb85bf788),
	.w2(32'hb83951ed),
	.w3(32'hb74d70f8),
	.w4(32'hb9778e1d),
	.w5(32'hb907b41f),
	.w6(32'hb99e9ab5),
	.w7(32'hb9ac14bc),
	.w8(32'hb988d9f3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393791e8),
	.w1(32'hb948961f),
	.w2(32'hb90fa88f),
	.w3(32'h372b0e21),
	.w4(32'hb9b5fc21),
	.w5(32'hb99c1081),
	.w6(32'h399e5d9d),
	.w7(32'hb8a04361),
	.w8(32'hb895d594),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cf1ee1),
	.w1(32'hb9288f06),
	.w2(32'hb8f9c893),
	.w3(32'h38141c45),
	.w4(32'hb92850b6),
	.w5(32'hb93fa5aa),
	.w6(32'h384a29da),
	.w7(32'hb80b514c),
	.w8(32'hb8c4bd26),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f773f),
	.w1(32'h38022f98),
	.w2(32'hb84732cc),
	.w3(32'h395b9e76),
	.w4(32'hb5d064e3),
	.w5(32'hb920f8f5),
	.w6(32'h37d87e0e),
	.w7(32'hb948f33e),
	.w8(32'hb9e1432e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb776f9af),
	.w1(32'hb7477462),
	.w2(32'hb673ae14),
	.w3(32'hb6cd16e0),
	.w4(32'hb6c65822),
	.w5(32'hb690c390),
	.w6(32'hb6ecc873),
	.w7(32'hb6655aeb),
	.w8(32'hb638761f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7affecf),
	.w1(32'hb4ea3eee),
	.w2(32'h36cbf53f),
	.w3(32'hb7ffac5a),
	.w4(32'hb75ac7aa),
	.w5(32'h375f5817),
	.w6(32'hb80b79be),
	.w7(32'hb73fdcb3),
	.w8(32'h377b7c6d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce8d4d),
	.w1(32'h3733df19),
	.w2(32'hb8cc844b),
	.w3(32'h3a229326),
	.w4(32'h38d6468c),
	.w5(32'hb8163de9),
	.w6(32'h38579f3c),
	.w7(32'hb9cd2000),
	.w8(32'hba3b4860),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2dc94),
	.w1(32'h39248c92),
	.w2(32'h3980f395),
	.w3(32'h39bc2712),
	.w4(32'h391ac5dc),
	.w5(32'h3999e7fd),
	.w6(32'h3982d426),
	.w7(32'h3908a061),
	.w8(32'h3965fca9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c7e17),
	.w1(32'h390056c8),
	.w2(32'h3898bf60),
	.w3(32'h38bdd124),
	.w4(32'hb8528708),
	.w5(32'h38734c17),
	.w6(32'h386f72a7),
	.w7(32'hb6368bea),
	.w8(32'h38ee9010),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dd1770),
	.w1(32'hb90e9727),
	.w2(32'hb900b4ef),
	.w3(32'h38d0ae40),
	.w4(32'hb8936722),
	.w5(32'hb92d09c7),
	.w6(32'h3907941a),
	.w7(32'h3829b62e),
	.w8(32'hb7ee05ae),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f03482),
	.w1(32'h39bdc2fa),
	.w2(32'h398d84d7),
	.w3(32'h396272d2),
	.w4(32'h37f14e86),
	.w5(32'hb820fa8f),
	.w6(32'h39c308ac),
	.w7(32'h38a8f80c),
	.w8(32'hb87cbd7f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ea7ab8),
	.w1(32'hb98c6b36),
	.w2(32'hb9c0b82d),
	.w3(32'h393011cf),
	.w4(32'hb99f2970),
	.w5(32'hb9e39453),
	.w6(32'hb85ab220),
	.w7(32'hb9b5447f),
	.w8(32'hb9dd377e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3609446f),
	.w1(32'h35caa201),
	.w2(32'h36bbcdbd),
	.w3(32'hb560bfa5),
	.w4(32'hb6f959f8),
	.w5(32'hb6871277),
	.w6(32'hb583dd00),
	.w7(32'hb6bd58f1),
	.w8(32'hb6a4da29),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47c877),
	.w1(32'hb7dd95b0),
	.w2(32'h393c9e6e),
	.w3(32'h399668f5),
	.w4(32'hba0dfdee),
	.w5(32'hb9f758de),
	.w6(32'h39f247b3),
	.w7(32'hb8073a6f),
	.w8(32'hb8d58fc4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb503925d),
	.w1(32'hb41d37aa),
	.w2(32'h351bf2ec),
	.w3(32'hb6aced0d),
	.w4(32'hb68e04bf),
	.w5(32'hb6523aa5),
	.w6(32'hb6760971),
	.w7(32'hb61e85fd),
	.w8(32'hb5d86dfb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c973d),
	.w1(32'h382dd7b7),
	.w2(32'h389b6d2d),
	.w3(32'h38a1bd79),
	.w4(32'hb8ae0535),
	.w5(32'hb8bfd229),
	.w6(32'h39138c60),
	.w7(32'hb840ce0e),
	.w8(32'hb8f963b5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69a8119),
	.w1(32'h36ef950e),
	.w2(32'h36d896d7),
	.w3(32'hb63d57e2),
	.w4(32'h372927fd),
	.w5(32'h379d286f),
	.w6(32'h3707aede),
	.w7(32'h374a3169),
	.w8(32'h37f17d9d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393c80d5),
	.w1(32'h389cfade),
	.w2(32'h38d7de11),
	.w3(32'h39e9a6b4),
	.w4(32'h3982c698),
	.w5(32'h3990b5e5),
	.w6(32'h3819e3f7),
	.w7(32'h386e5013),
	.w8(32'h37ae65fa),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb630dc6e),
	.w1(32'hb5d9017f),
	.w2(32'hb557624c),
	.w3(32'hb5f63179),
	.w4(32'h3384cf3a),
	.w5(32'h353c70d3),
	.w6(32'hb63434a5),
	.w7(32'hb4b4f53b),
	.w8(32'h3483a9c0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3933bde6),
	.w1(32'h38578861),
	.w2(32'hb738d9b6),
	.w3(32'hb879024f),
	.w4(32'hb916d46a),
	.w5(32'hb960790b),
	.w6(32'h385df73b),
	.w7(32'hb850fc13),
	.w8(32'hb9544d6c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a705ca),
	.w1(32'hb5f4eeb3),
	.w2(32'hb5d3dbc2),
	.w3(32'hb65f094e),
	.w4(32'hb5b62961),
	.w5(32'hb4be9d21),
	.w6(32'hb6816914),
	.w7(32'hb651f9be),
	.w8(32'hb49f9f5c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399247d1),
	.w1(32'hb981f227),
	.w2(32'hb9381377),
	.w3(32'h392b8303),
	.w4(32'hb9990378),
	.w5(32'hba18a5ff),
	.w6(32'h39675f6d),
	.w7(32'hb933bc8b),
	.w8(32'hb9f20e99),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a29b2b),
	.w1(32'hb9ab67c8),
	.w2(32'hb988e929),
	.w3(32'h394fb635),
	.w4(32'hb8cc2de2),
	.w5(32'hb8b23292),
	.w6(32'hb99e7960),
	.w7(32'hb9815cdc),
	.w8(32'hb9b7a039),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b4ab00),
	.w1(32'h35e33362),
	.w2(32'h359e7628),
	.w3(32'hb6fbfe99),
	.w4(32'hb616f581),
	.w5(32'hb6a6b709),
	.w6(32'hb58958f5),
	.w7(32'hb5f67f38),
	.w8(32'hb6acce2f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7148a14),
	.w1(32'hb66b71f4),
	.w2(32'hb68ccf8a),
	.w3(32'hb6ee86b2),
	.w4(32'hb586c675),
	.w5(32'hb64368d0),
	.w6(32'hb6bf4806),
	.w7(32'hb602203b),
	.w8(32'hb6a0ae0d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6512c),
	.w1(32'h3994f3a5),
	.w2(32'h39815ba0),
	.w3(32'h3930bf2d),
	.w4(32'hb84bb885),
	.w5(32'hb86eb598),
	.w6(32'h39b22268),
	.w7(32'h3886e240),
	.w8(32'hb9846ef8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e90cb),
	.w1(32'hb91e3faf),
	.w2(32'hb8daf420),
	.w3(32'h3945e916),
	.w4(32'hb9ab914a),
	.w5(32'hb9f32069),
	.w6(32'h392390ce),
	.w7(32'hb98c81c3),
	.w8(32'hba1dc771),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a876848),
	.w1(32'hb9242a4b),
	.w2(32'hb9bc72bb),
	.w3(32'h3a8e115f),
	.w4(32'h390c2539),
	.w5(32'hb8d7d47d),
	.w6(32'h3923f2a6),
	.w7(32'hba339ec4),
	.w8(32'hba799c10),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1755bb),
	.w1(32'hb96ad8b0),
	.w2(32'hb6668768),
	.w3(32'h39d1bd90),
	.w4(32'hb9ba3164),
	.w5(32'hba0fffa2),
	.w6(32'h39fdd7ec),
	.w7(32'hb9ddc1a2),
	.w8(32'hba7604fd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c570db),
	.w1(32'h391c122e),
	.w2(32'h39b914d3),
	.w3(32'h385bfb22),
	.w4(32'hb812d2b9),
	.w5(32'h38e315cf),
	.w6(32'h399f6879),
	.w7(32'h39239e4e),
	.w8(32'hb8b951e4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb832ff0f),
	.w1(32'hb73661a5),
	.w2(32'hb7021801),
	.w3(32'hb7deb2ac),
	.w4(32'h3706ac8d),
	.w5(32'h36e541e8),
	.w6(32'hb7f9238c),
	.w7(32'h3522ee18),
	.w8(32'h3644e878),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cff3f),
	.w1(32'hb690c779),
	.w2(32'hb6844126),
	.w3(32'hb6b5ad32),
	.w4(32'hb5989309),
	.w5(32'hb58357ab),
	.w6(32'hb6f13f3f),
	.w7(32'hb6570400),
	.w8(32'hb62ad70d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74e3a60),
	.w1(32'hb6262a0a),
	.w2(32'h36012150),
	.w3(32'hb73bc819),
	.w4(32'hb5983ef3),
	.w5(32'h35dde4be),
	.w6(32'hb7190afa),
	.w7(32'hb65f8f03),
	.w8(32'hb3459102),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cba5cb),
	.w1(32'h386847b1),
	.w2(32'h386cf0af),
	.w3(32'hb6ca48a6),
	.w4(32'h3901573b),
	.w5(32'h38eed249),
	.w6(32'h37ad3c6e),
	.w7(32'h38eefd40),
	.w8(32'h37d19f22),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de47cf),
	.w1(32'h388c9f5d),
	.w2(32'h388a7a3f),
	.w3(32'h39c43ac6),
	.w4(32'h37927937),
	.w5(32'h3879873f),
	.w6(32'h38bf9eb9),
	.w7(32'hb940fa38),
	.w8(32'hb988e7f0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37697831),
	.w1(32'h37061241),
	.w2(32'h36f05d4f),
	.w3(32'h36a1fc70),
	.w4(32'hb4833d39),
	.w5(32'h36cca783),
	.w6(32'h377f9a01),
	.w7(32'h3682e3c4),
	.w8(32'h36ab0383),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d31ba3),
	.w1(32'h38d40989),
	.w2(32'h390a8007),
	.w3(32'h3907ecd6),
	.w4(32'hb92accdc),
	.w5(32'hb872acc6),
	.w6(32'h39b30249),
	.w7(32'hb817b713),
	.w8(32'hb8d18c47),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39874189),
	.w1(32'h389bd30c),
	.w2(32'h391e39bd),
	.w3(32'h3943b5f0),
	.w4(32'h386ab194),
	.w5(32'h37ac62c7),
	.w6(32'h39330d28),
	.w7(32'hb83e056b),
	.w8(32'hb8cb60c3),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886cd1c),
	.w1(32'hb6187732),
	.w2(32'hb876350f),
	.w3(32'h3960ff22),
	.w4(32'h389b5eb4),
	.w5(32'h38584251),
	.w6(32'h387b9295),
	.w7(32'hb83e4cde),
	.w8(32'hb8a6e569),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916bd19),
	.w1(32'hb993b408),
	.w2(32'hb9719611),
	.w3(32'h38a5315f),
	.w4(32'hb9722329),
	.w5(32'hb9cebfad),
	.w6(32'hb88e54a0),
	.w7(32'hb9a0f996),
	.w8(32'hb9e5ba27),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bc1fd),
	.w1(32'h38182400),
	.w2(32'h38a6cdac),
	.w3(32'h39cccd16),
	.w4(32'hb94dacf6),
	.w5(32'hb9bd98f9),
	.w6(32'h39c90eb9),
	.w7(32'hb99da68c),
	.w8(32'hba029284),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70b9b9d),
	.w1(32'hb52743b3),
	.w2(32'hb5252b20),
	.w3(32'hb6864361),
	.w4(32'h362413dc),
	.w5(32'h3689cdfe),
	.w6(32'hb6fb9782),
	.w7(32'hb61d3391),
	.w8(32'h354c3c8f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb802629e),
	.w1(32'hb6c2c4fb),
	.w2(32'hb7129f10),
	.w3(32'hb7ac4d19),
	.w4(32'h3683f17a),
	.w5(32'h36710213),
	.w6(32'hb7d5b74f),
	.w7(32'hb5b512f2),
	.w8(32'hb3ee1fb5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79096aa),
	.w1(32'hb70986b5),
	.w2(32'hb720fd17),
	.w3(32'hb7486828),
	.w4(32'hb5cd9a86),
	.w5(32'hb66ab899),
	.w6(32'hb76fd7e1),
	.w7(32'hb66379be),
	.w8(32'hb6abb7d6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e52201),
	.w1(32'h3684f6a7),
	.w2(32'h3739ac2d),
	.w3(32'h371f7f8f),
	.w4(32'hb415e309),
	.w5(32'h3713e229),
	.w6(32'h36c08bbf),
	.w7(32'h3469c608),
	.w8(32'h3618e496),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397799eb),
	.w1(32'h396bbbe2),
	.w2(32'h3978e409),
	.w3(32'h3919d2f6),
	.w4(32'h38f12e50),
	.w5(32'h38d018d3),
	.w6(32'h3905c450),
	.w7(32'h38d2ba06),
	.w8(32'h389db799),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bf4e8c),
	.w1(32'h3796afed),
	.w2(32'h36b120c1),
	.w3(32'h36cca61c),
	.w4(32'hb5033d45),
	.w5(32'hb679bfb2),
	.w6(32'h37a8813d),
	.w7(32'h378739f6),
	.w8(32'h368f082c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a018bc7),
	.w1(32'h39ba2cec),
	.w2(32'h39b0a485),
	.w3(32'h3928b383),
	.w4(32'hb805a1bc),
	.w5(32'h382c1241),
	.w6(32'h3981ea12),
	.w7(32'hb809928f),
	.w8(32'hb9224371),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3908c6c0),
	.w1(32'h3930fd23),
	.w2(32'h3961b7a4),
	.w3(32'h381c28f1),
	.w4(32'h3841a932),
	.w5(32'h390b7e9a),
	.w6(32'h38c89f17),
	.w7(32'h38f25877),
	.w8(32'hba545d83),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918ad40),
	.w1(32'hb92264c9),
	.w2(32'hba2371c5),
	.w3(32'h388e14f4),
	.w4(32'hba2e7874),
	.w5(32'hba3f5cbb),
	.w6(32'h39221325),
	.w7(32'h39127e87),
	.w8(32'hb957b5ef),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00bc8f),
	.w1(32'hbad419f0),
	.w2(32'hba82d122),
	.w3(32'hbb657591),
	.w4(32'hbb1838e3),
	.w5(32'hb9c6791e),
	.w6(32'h3a32c84b),
	.w7(32'hb9941e7a),
	.w8(32'hba3878dd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1157ee),
	.w1(32'h39a905ca),
	.w2(32'hb8ef86e3),
	.w3(32'h3a1ba01b),
	.w4(32'hba093d35),
	.w5(32'hb99ba9ed),
	.w6(32'h38ae4983),
	.w7(32'h38dd3fa6),
	.w8(32'h3905bfca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a897151),
	.w1(32'h3a3bcdb3),
	.w2(32'h3a06825f),
	.w3(32'h3a49a4bf),
	.w4(32'hb992ca3f),
	.w5(32'hb7b3ee52),
	.w6(32'h39c31ae3),
	.w7(32'h3a0354d4),
	.w8(32'hba49a095),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7bc50),
	.w1(32'hba265259),
	.w2(32'hb9988418),
	.w3(32'hb97e623f),
	.w4(32'hb981245e),
	.w5(32'hba364af6),
	.w6(32'h390505c8),
	.w7(32'hb9dacc58),
	.w8(32'h39c459d4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a909ba9),
	.w1(32'h3995c436),
	.w2(32'h3a6daf21),
	.w3(32'hbaf251fd),
	.w4(32'hb91b08cc),
	.w5(32'h3b909c03),
	.w6(32'hba021265),
	.w7(32'hbad7df30),
	.w8(32'hb9ee0b40),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a662099),
	.w1(32'hb95fb36d),
	.w2(32'hb8fc33f9),
	.w3(32'h394935f3),
	.w4(32'hbabce5e9),
	.w5(32'hba3f26e6),
	.w6(32'h3a203e7d),
	.w7(32'hba001ea9),
	.w8(32'h3b1752cf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad45824),
	.w1(32'h3a2e7579),
	.w2(32'h3ac2d599),
	.w3(32'h3aa10e88),
	.w4(32'h3a7bfb8f),
	.w5(32'h3a9e0e99),
	.w6(32'h3a4086d2),
	.w7(32'h3ac26895),
	.w8(32'h38cb4532),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19848e),
	.w1(32'h3a02cf1a),
	.w2(32'h392dd190),
	.w3(32'h3a486da1),
	.w4(32'h377f7c3e),
	.w5(32'hb9cf60f9),
	.w6(32'h395e671c),
	.w7(32'h393c920b),
	.w8(32'hba398ad8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ea1ee),
	.w1(32'hb9125c42),
	.w2(32'hb986817f),
	.w3(32'h39294bd4),
	.w4(32'hb94d229a),
	.w5(32'hb9956a50),
	.w6(32'hb8eb6f60),
	.w7(32'hb9862a14),
	.w8(32'hbacb01e5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93387d2),
	.w1(32'hb7f8728d),
	.w2(32'hba125b68),
	.w3(32'h39361b5c),
	.w4(32'hba06263e),
	.w5(32'hba029ff4),
	.w6(32'hb9bb6a04),
	.w7(32'hb99269ca),
	.w8(32'hbae5da27),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34588d),
	.w1(32'hba6435ae),
	.w2(32'hbb69f0c7),
	.w3(32'hbb2c5253),
	.w4(32'h39a760d1),
	.w5(32'hbb2c5804),
	.w6(32'h3aa82443),
	.w7(32'hbb896dfa),
	.w8(32'hb89eb53e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd6032),
	.w1(32'hba5cfc91),
	.w2(32'h388d6219),
	.w3(32'h3a6d4703),
	.w4(32'hb97ecdea),
	.w5(32'hb8b872a6),
	.w6(32'hb9e09018),
	.w7(32'h38edc5dd),
	.w8(32'h3b1fc3fe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfdb91),
	.w1(32'hbb1219d3),
	.w2(32'hbad7807d),
	.w3(32'hb99a4cd3),
	.w4(32'hba445c84),
	.w5(32'hb8de2b17),
	.w6(32'hbb217438),
	.w7(32'hbb04c92d),
	.w8(32'h394cf5d0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f7f59),
	.w1(32'hba0b87bf),
	.w2(32'hbb2ae17d),
	.w3(32'h397b3f19),
	.w4(32'hba063b3e),
	.w5(32'hba812da6),
	.w6(32'hbaf836c0),
	.w7(32'hba9b4ed7),
	.w8(32'h39fd5593),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b10ee),
	.w1(32'h3a49a906),
	.w2(32'h39acb7ff),
	.w3(32'h388cb587),
	.w4(32'hba1c2999),
	.w5(32'hba51cfd3),
	.w6(32'hbacecec5),
	.w7(32'hbabc65a7),
	.w8(32'h3aa7190b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80c72c),
	.w1(32'hba402333),
	.w2(32'hb91e1674),
	.w3(32'hba758988),
	.w4(32'h3a057675),
	.w5(32'hb9996b23),
	.w6(32'h3a4346d8),
	.w7(32'h3a5c99d3),
	.w8(32'h3a39ee89),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30f4d7),
	.w1(32'hb8c2d762),
	.w2(32'h3a427524),
	.w3(32'h3a4d6e85),
	.w4(32'hb9353695),
	.w5(32'h3a876f54),
	.w6(32'hb911c973),
	.w7(32'h3a7156a2),
	.w8(32'hba649fcb),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e073b),
	.w1(32'h38a774e3),
	.w2(32'hbabc7b8a),
	.w3(32'hbb02c19d),
	.w4(32'hba538d4d),
	.w5(32'hb9dcbe1d),
	.w6(32'hba5f23bc),
	.w7(32'hba505f97),
	.w8(32'h3a813506),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0c1c9),
	.w1(32'h3b0d2871),
	.w2(32'hbb8e275e),
	.w3(32'hbad68102),
	.w4(32'hbb14b5a1),
	.w5(32'h3a9b89e4),
	.w6(32'h3b4eb497),
	.w7(32'hba2b6860),
	.w8(32'hbaacf72e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad89a3a),
	.w1(32'hb967c31b),
	.w2(32'hb81120b4),
	.w3(32'hba634cf7),
	.w4(32'hba184bc7),
	.w5(32'hbabd338a),
	.w6(32'hba688e8b),
	.w7(32'hba648180),
	.w8(32'hb9ad1b18),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a397c35),
	.w1(32'h3a0ccb66),
	.w2(32'h39345ffe),
	.w3(32'h3a74eb26),
	.w4(32'hb8954d22),
	.w5(32'hb92692d6),
	.w6(32'h391b7cfd),
	.w7(32'h39d0ed58),
	.w8(32'hba9e7a0e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d6ab0),
	.w1(32'hbb6da3ed),
	.w2(32'h3a27bf47),
	.w3(32'hbab3d07a),
	.w4(32'hbafb7abd),
	.w5(32'hba8ed19b),
	.w6(32'hba82de40),
	.w7(32'hba8e8ea5),
	.w8(32'hba534a07),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule