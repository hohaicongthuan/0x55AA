module layer_10_featuremap_121(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8470e),
	.w1(32'h3a288142),
	.w2(32'h3aab15a6),
	.w3(32'h383bb1bf),
	.w4(32'h3a749811),
	.w5(32'h3ab59c78),
	.w6(32'hbaac8aef),
	.w7(32'hbabbdfe4),
	.w8(32'hba3460d7),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964359d),
	.w1(32'h39eb0827),
	.w2(32'h390ff1e7),
	.w3(32'h3a241f4c),
	.w4(32'h3a0adb75),
	.w5(32'h39d1071a),
	.w6(32'h38a3e59d),
	.w7(32'h39b197f7),
	.w8(32'h3979f2cb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a338f7c),
	.w1(32'hb9396684),
	.w2(32'hb910cdbe),
	.w3(32'h3a3b714d),
	.w4(32'hb9b245cb),
	.w5(32'hb9ba513a),
	.w6(32'h39592631),
	.w7(32'h39c7eb73),
	.w8(32'h3a29dc0f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4ed41),
	.w1(32'hb9854cc5),
	.w2(32'h3a95dd21),
	.w3(32'h38e6efc7),
	.w4(32'hba22c753),
	.w5(32'hba1445eb),
	.w6(32'h3a260060),
	.w7(32'h3a128929),
	.w8(32'h3a8fe404),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3304f4),
	.w1(32'hba1fdf93),
	.w2(32'hb9ee8d28),
	.w3(32'hb9cb7781),
	.w4(32'hba1327cb),
	.w5(32'hba7eec24),
	.w6(32'hba6be1c9),
	.w7(32'hba228634),
	.w8(32'hb7b6eec9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39022c39),
	.w1(32'h3a562e20),
	.w2(32'h39e7ddfb),
	.w3(32'hb9a7b114),
	.w4(32'h39f52009),
	.w5(32'h39c2b6d9),
	.w6(32'h3a5e3d15),
	.w7(32'h39811ab6),
	.w8(32'h3868d40b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e31dff),
	.w1(32'hb9938a8d),
	.w2(32'h3806a044),
	.w3(32'h3999b85f),
	.w4(32'hb9b845a3),
	.w5(32'hb9295f7c),
	.w6(32'hb934c54d),
	.w7(32'h38dd8fc1),
	.w8(32'h399a6340),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265502),
	.w1(32'h392085c7),
	.w2(32'hb8d307f8),
	.w3(32'h39fa5afa),
	.w4(32'h39497e6c),
	.w5(32'h386d2082),
	.w6(32'h38851924),
	.w7(32'hb89cacb9),
	.w8(32'hb87f4890),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b427fc),
	.w1(32'h3a213922),
	.w2(32'hb9557e43),
	.w3(32'hb8fb3432),
	.w4(32'h39fef628),
	.w5(32'h3818d94d),
	.w6(32'h3990e6f0),
	.w7(32'hb93b627b),
	.w8(32'hb915bd6c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42feee),
	.w1(32'h3a86d1d4),
	.w2(32'hb984106c),
	.w3(32'h3b0a1d5e),
	.w4(32'h39cd30e0),
	.w5(32'hb965c6f4),
	.w6(32'h3a20a8b5),
	.w7(32'hb967359b),
	.w8(32'h3800b7c2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a72d8e),
	.w1(32'h3970c993),
	.w2(32'h3a2ccabe),
	.w3(32'h39830a9f),
	.w4(32'h3949e146),
	.w5(32'h39b33d43),
	.w6(32'h3a929002),
	.w7(32'h3ae9ba49),
	.w8(32'h3acf0659),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00511c),
	.w1(32'hba0bf56e),
	.w2(32'h3a091269),
	.w3(32'h3a02eefc),
	.w4(32'hba3863d2),
	.w5(32'hba676bcd),
	.w6(32'hba3ad157),
	.w7(32'hb980b90e),
	.w8(32'hba0e8034),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae55752),
	.w1(32'h39e9e115),
	.w2(32'hba131b72),
	.w3(32'h3a92173b),
	.w4(32'h3a0ebb9d),
	.w5(32'hb9199af3),
	.w6(32'h3a3ec640),
	.w7(32'h38f85e43),
	.w8(32'h3990eb20),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c3f43),
	.w1(32'hb99bfec2),
	.w2(32'hba3b14c0),
	.w3(32'h3a908600),
	.w4(32'hb9cc8a25),
	.w5(32'hba49e976),
	.w6(32'h3a8476db),
	.w7(32'h3916ffaf),
	.w8(32'hb999af55),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39249102),
	.w1(32'hba008098),
	.w2(32'h3ae91743),
	.w3(32'hb9deadba),
	.w4(32'hba38af28),
	.w5(32'hba2da10e),
	.w6(32'hba64980e),
	.w7(32'hbaaa18b9),
	.w8(32'h399ab820),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9857fe),
	.w1(32'h3a4d472d),
	.w2(32'h3897d076),
	.w3(32'h3a227999),
	.w4(32'h3a0caec4),
	.w5(32'h39e2f166),
	.w6(32'h3a2b7ab1),
	.w7(32'hb9578cc9),
	.w8(32'h39bda544),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f395ea),
	.w1(32'h3a3e8038),
	.w2(32'h3945579d),
	.w3(32'h3a3418ef),
	.w4(32'h3993d69e),
	.w5(32'hb8720c12),
	.w6(32'h3a0a785a),
	.w7(32'hb8a79a2b),
	.w8(32'h396f5ac2),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a720bcd),
	.w1(32'hb9d3b976),
	.w2(32'hb992fb05),
	.w3(32'h3a1fe97e),
	.w4(32'hb95ceec2),
	.w5(32'h389121a2),
	.w6(32'hb9ba8b43),
	.w7(32'hb9a2710b),
	.w8(32'h3986ce64),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71a7a1),
	.w1(32'hb8c996b1),
	.w2(32'h380cd7e3),
	.w3(32'h39fa1b72),
	.w4(32'hb9914fe3),
	.w5(32'hb893ffd1),
	.w6(32'hb8b90fd6),
	.w7(32'hb7027d3c),
	.w8(32'h3a36dc00),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab277d),
	.w1(32'h3a307035),
	.w2(32'h3975c5b8),
	.w3(32'h39636cb2),
	.w4(32'h3a28f59c),
	.w5(32'h39f3a846),
	.w6(32'h39ef51a0),
	.w7(32'h39b4467f),
	.w8(32'h39a5c4bd),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b04f35),
	.w1(32'h3a23db0e),
	.w2(32'h39939aaa),
	.w3(32'h39a75377),
	.w4(32'h3a922de7),
	.w5(32'h3a4bcd59),
	.w6(32'h3a82c6b7),
	.w7(32'h3a17f22e),
	.w8(32'h3a19ab07),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3563d),
	.w1(32'hba7c8f88),
	.w2(32'h3a162228),
	.w3(32'h388a8767),
	.w4(32'hbaca456a),
	.w5(32'hba8e412c),
	.w6(32'hb99325bc),
	.w7(32'h3a669a96),
	.w8(32'h39924516),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bd696),
	.w1(32'h3af1c994),
	.w2(32'hb8fc4a83),
	.w3(32'h3ab66ad4),
	.w4(32'h3a884a61),
	.w5(32'hba767329),
	.w6(32'h3b09910c),
	.w7(32'hba1a8176),
	.w8(32'hb962aa44),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a8e3),
	.w1(32'h39c151f0),
	.w2(32'hba061d90),
	.w3(32'h3aaa2333),
	.w4(32'hb882b27f),
	.w5(32'hb9e5e929),
	.w6(32'h3a1a8533),
	.w7(32'hba1eea9a),
	.w8(32'hb9b4d79c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f591b),
	.w1(32'h3a2344d9),
	.w2(32'h37cd310a),
	.w3(32'h3a14ba51),
	.w4(32'h390326c4),
	.w5(32'hb9e109c7),
	.w6(32'h3a3c7467),
	.w7(32'hba12fdd4),
	.w8(32'hb8c8c17b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84bbd6),
	.w1(32'hb9996c92),
	.w2(32'hb9cca43e),
	.w3(32'h3a2c7d16),
	.w4(32'hb9c8209d),
	.w5(32'hba370ab1),
	.w6(32'hb7a3d9de),
	.w7(32'hba18d710),
	.w8(32'hb9c66499),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980ea45),
	.w1(32'h395c2ce8),
	.w2(32'h3872e751),
	.w3(32'hb9e3e01e),
	.w4(32'h39995d12),
	.w5(32'h39291ff9),
	.w6(32'h3947e2fc),
	.w7(32'h399a1344),
	.w8(32'h394e1b4e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9289783),
	.w1(32'hba37e2f9),
	.w2(32'hba4131fe),
	.w3(32'hb97242bc),
	.w4(32'hba870308),
	.w5(32'hba96cef9),
	.w6(32'hba5b0d5e),
	.w7(32'hba8bb9d3),
	.w8(32'hba378725),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72cfad),
	.w1(32'h3a962dbb),
	.w2(32'h38882743),
	.w3(32'hba77744b),
	.w4(32'h3a49400e),
	.w5(32'hb8ead1f7),
	.w6(32'h3ab7f57d),
	.w7(32'h3a0c2ebe),
	.w8(32'h3a2f45fa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b164328),
	.w1(32'h3b2a056c),
	.w2(32'h3a42d1bb),
	.w3(32'h3aa5a55e),
	.w4(32'h3af675ac),
	.w5(32'h3a07ba67),
	.w6(32'h3b137552),
	.w7(32'h3a085c4e),
	.w8(32'h3a6019c9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9110a3),
	.w1(32'h3a0de2eb),
	.w2(32'h3970c5bc),
	.w3(32'h3a435213),
	.w4(32'h3a543cb4),
	.w5(32'h3a2c55bb),
	.w6(32'h3a2f8f3a),
	.w7(32'h3a072526),
	.w8(32'h39f136db),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923fa05),
	.w1(32'h38c85f6d),
	.w2(32'h38d8c6a5),
	.w3(32'h39cb2ebf),
	.w4(32'h39551e8c),
	.w5(32'h39896c39),
	.w6(32'h395d47e9),
	.w7(32'h3948d7cb),
	.w8(32'h3982ee32),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4bed4c),
	.w1(32'h38510278),
	.w2(32'hb987a872),
	.w3(32'h3a39b0ff),
	.w4(32'hb95b3489),
	.w5(32'hba18b8f1),
	.w6(32'h39a82601),
	.w7(32'h38fdd32f),
	.w8(32'hb9a70549),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39015b19),
	.w1(32'hb91c94b6),
	.w2(32'h39c19761),
	.w3(32'hb98b2435),
	.w4(32'hba6768d7),
	.w5(32'hb9ae9aab),
	.w6(32'hb9b31516),
	.w7(32'h3a766cc7),
	.w8(32'hb9ead975),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90c4049),
	.w1(32'hb9021cb3),
	.w2(32'h39314b48),
	.w3(32'hba366197),
	.w4(32'hb54b69d1),
	.w5(32'h3753d2d6),
	.w6(32'hb9f58acb),
	.w7(32'h398f4f6a),
	.w8(32'h398c2df9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0831a),
	.w1(32'h395e0df9),
	.w2(32'h397f72c2),
	.w3(32'h38b57e3e),
	.w4(32'h39b13d3b),
	.w5(32'h39ad3489),
	.w6(32'h39cfc4ad),
	.w7(32'h395e8c36),
	.w8(32'h3952c1bc),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdbcff),
	.w1(32'h3ab6369a),
	.w2(32'h3a62aa87),
	.w3(32'h3ac472fd),
	.w4(32'h3a59846f),
	.w5(32'h3a37db4d),
	.w6(32'h3a86e920),
	.w7(32'h3a1cc3ff),
	.w8(32'h3a1d2534),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc8a31),
	.w1(32'h39ad6b32),
	.w2(32'hb901d3cc),
	.w3(32'h3a9e35db),
	.w4(32'h39290a39),
	.w5(32'hba308f5b),
	.w6(32'h396b48b6),
	.w7(32'h38d8311b),
	.w8(32'hba1c6190),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710992b),
	.w1(32'hb9ae0602),
	.w2(32'hba8426d7),
	.w3(32'h3920602f),
	.w4(32'hb9ef5860),
	.w5(32'hba8d3a98),
	.w6(32'hba6f2ecc),
	.w7(32'hba5765a6),
	.w8(32'hbaa153af),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39285e6f),
	.w1(32'h38fb888c),
	.w2(32'h3a1615b4),
	.w3(32'h39b81090),
	.w4(32'hb9714243),
	.w5(32'hb813de71),
	.w6(32'h391bcd63),
	.w7(32'h3a2b72c1),
	.w8(32'h3a244740),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02ddb2),
	.w1(32'h3aee859f),
	.w2(32'h3a5acac6),
	.w3(32'h390a7456),
	.w4(32'h3ab43f5c),
	.w5(32'h3a1f01a4),
	.w6(32'h3ac5dd1c),
	.w7(32'h3a75e4c8),
	.w8(32'h3a8e066c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d125a),
	.w1(32'h39c03ab5),
	.w2(32'h3a4485d6),
	.w3(32'h3a17e9a0),
	.w4(32'h39bb6576),
	.w5(32'h3a102ca3),
	.w6(32'h3a14ccc9),
	.w7(32'h3a4b2a50),
	.w8(32'h3a42f467),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dd0ad),
	.w1(32'h39f9ffba),
	.w2(32'hba16052e),
	.w3(32'h3a3a6119),
	.w4(32'h3a0a7433),
	.w5(32'hb93b188b),
	.w6(32'h3931c62e),
	.w7(32'hb8e4c5eb),
	.w8(32'hb900c277),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb4a42),
	.w1(32'h3954d931),
	.w2(32'hb9961de9),
	.w3(32'h3a23a1a3),
	.w4(32'h39cd701e),
	.w5(32'h38f59cde),
	.w6(32'hb9907ac1),
	.w7(32'hba8435f7),
	.w8(32'hb943e8d1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adddb41),
	.w1(32'hb8553eda),
	.w2(32'h37239538),
	.w3(32'h3a9f6938),
	.w4(32'hb992b120),
	.w5(32'hba5fcecf),
	.w6(32'h39b16932),
	.w7(32'hb9e11ec0),
	.w8(32'hba23e390),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefb628),
	.w1(32'hb9f43623),
	.w2(32'hba68136f),
	.w3(32'h3a8c2a1c),
	.w4(32'hba4788f7),
	.w5(32'hba78b272),
	.w6(32'h388ac213),
	.w7(32'hba4d2cc3),
	.w8(32'hb95b9096),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0718d),
	.w1(32'hba370757),
	.w2(32'h3ade0071),
	.w3(32'hb845b18c),
	.w4(32'hba6f2f21),
	.w5(32'hba9ca7c6),
	.w6(32'hba2d8cf5),
	.w7(32'hba7f8743),
	.w8(32'hb94ffc98),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc5328),
	.w1(32'h3a94bf87),
	.w2(32'h38cea981),
	.w3(32'hba11310c),
	.w4(32'h39f443f0),
	.w5(32'h399a452d),
	.w6(32'h3ac780db),
	.w7(32'h3942a0ca),
	.w8(32'h3aae72f5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41d823),
	.w1(32'h38adb9a6),
	.w2(32'hb908b740),
	.w3(32'h39ed1c15),
	.w4(32'h3819b006),
	.w5(32'h36079894),
	.w6(32'h36bfa8ae),
	.w7(32'h38df7d0b),
	.w8(32'h38bf9318),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394cf354),
	.w1(32'h3813b79a),
	.w2(32'hb93d6278),
	.w3(32'hb8c69a7d),
	.w4(32'hb8263c12),
	.w5(32'h387ce1da),
	.w6(32'hb900ca5e),
	.w7(32'hb9ee4574),
	.w8(32'hb9a34aab),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8067086),
	.w1(32'hb9d8f485),
	.w2(32'hb98698ae),
	.w3(32'h39238c11),
	.w4(32'hb9d95b4e),
	.w5(32'hb9ade979),
	.w6(32'hba5a2250),
	.w7(32'hba5d5c11),
	.w8(32'hb90ae9bd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50f2f5),
	.w1(32'h3a5e14ff),
	.w2(32'hba094dd8),
	.w3(32'h3a01e221),
	.w4(32'hb8907583),
	.w5(32'hb9a0423d),
	.w6(32'h3a008ca2),
	.w7(32'hba62eddd),
	.w8(32'hb9322ccf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866ea17),
	.w1(32'h3b0083e8),
	.w2(32'h3a6e86f6),
	.w3(32'h3936a020),
	.w4(32'h3b00b0ac),
	.w5(32'h3acdc0e8),
	.w6(32'h3ad495da),
	.w7(32'h3a2df60d),
	.w8(32'h3a5024c3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b618b93),
	.w1(32'h3a21b1c8),
	.w2(32'hb7590157),
	.w3(32'h3b2fe240),
	.w4(32'hb9b53216),
	.w5(32'hb9f476d3),
	.w6(32'h39b310e0),
	.w7(32'hb6ab09f7),
	.w8(32'hba08160e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390df428),
	.w1(32'hb918882b),
	.w2(32'hba49c5f3),
	.w3(32'hb8e6adf7),
	.w4(32'hb9033082),
	.w5(32'hba0a9657),
	.w6(32'hb95cde32),
	.w7(32'hb9dc492a),
	.w8(32'hb91b4ac6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b04fbb),
	.w1(32'h3ae7138b),
	.w2(32'h3a0564b6),
	.w3(32'h381c0cca),
	.w4(32'h3ac554b0),
	.w5(32'h3979a8c9),
	.w6(32'h3b0719b5),
	.w7(32'h3a93d4b3),
	.w8(32'h3aaad845),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a71b1),
	.w1(32'h3a2c5d46),
	.w2(32'h3a00fe25),
	.w3(32'h3a2019a9),
	.w4(32'h39d141f4),
	.w5(32'h3a064701),
	.w6(32'h3a01f255),
	.w7(32'h39a90f0e),
	.w8(32'h398032b7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05daa9),
	.w1(32'hba59fb9a),
	.w2(32'hba172c09),
	.w3(32'h39ff6f73),
	.w4(32'hbace7747),
	.w5(32'hbaa421b0),
	.w6(32'hba6cfc27),
	.w7(32'hba9fd7b1),
	.w8(32'hba1d9ecf),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e9802b),
	.w1(32'hb934b056),
	.w2(32'hb98b7691),
	.w3(32'hb99e6cec),
	.w4(32'hb9a997a6),
	.w5(32'hb9e9428b),
	.w6(32'hb8275903),
	.w7(32'hb8cacdb4),
	.w8(32'h373c5136),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18b416),
	.w1(32'h37a92eb6),
	.w2(32'hb90fe6ee),
	.w3(32'h39972e42),
	.w4(32'h38dee99f),
	.w5(32'h38ed43e5),
	.w6(32'h38fa0ec6),
	.w7(32'hb96bda1f),
	.w8(32'hb844c3a4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b1a417),
	.w1(32'hb91c0174),
	.w2(32'hb9baebf2),
	.w3(32'h39b743ff),
	.w4(32'hb932f1c2),
	.w5(32'hb9d9c552),
	.w6(32'hb9d30ad2),
	.w7(32'h3931ebf3),
	.w8(32'h399e4530),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a313aa7),
	.w1(32'h3a07aae1),
	.w2(32'h39f76695),
	.w3(32'h39ba799b),
	.w4(32'h39a43b50),
	.w5(32'h3a1a79aa),
	.w6(32'h39f16e2d),
	.w7(32'h39aba120),
	.w8(32'h3a05da4e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b810f),
	.w1(32'hb916c894),
	.w2(32'h382b98c5),
	.w3(32'h3926dc00),
	.w4(32'h3a18dfe3),
	.w5(32'hb7aa7b74),
	.w6(32'hba270a58),
	.w7(32'h3a283b3a),
	.w8(32'hb9b188c4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f427f),
	.w1(32'hb75f5377),
	.w2(32'h385f63fc),
	.w3(32'h381b57f3),
	.w4(32'hb7ddbd8c),
	.w5(32'hb8e8845b),
	.w6(32'hba17f946),
	.w7(32'hb9fbf18e),
	.w8(32'hb9c3a399),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ba055),
	.w1(32'hba16eda6),
	.w2(32'hb9c3847d),
	.w3(32'hb76ae255),
	.w4(32'hb9ee6107),
	.w5(32'hba3a3986),
	.w6(32'hba04ada3),
	.w7(32'hb9647777),
	.w8(32'hb8f5efa2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391122a5),
	.w1(32'hba6eb5ba),
	.w2(32'hba95d871),
	.w3(32'hb97c0e84),
	.w4(32'hba8e7b11),
	.w5(32'hba561b12),
	.w6(32'hba1d69f7),
	.w7(32'hba352c89),
	.w8(32'hb9925583),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97138f8),
	.w1(32'h3aa0f80b),
	.w2(32'h3a6b4c9f),
	.w3(32'hb9882f15),
	.w4(32'h3a8bded1),
	.w5(32'h3a90df6d),
	.w6(32'h3aa0c768),
	.w7(32'h3aa44116),
	.w8(32'h3a986321),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac361b9),
	.w1(32'h3b00a04c),
	.w2(32'h39ec7f08),
	.w3(32'h3aba22a5),
	.w4(32'h3a9835f7),
	.w5(32'hb974a1a2),
	.w6(32'h3ad6ee0b),
	.w7(32'hb83626cb),
	.w8(32'h3a18a09a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae10fa5),
	.w1(32'h3a67d26d),
	.w2(32'h398e2194),
	.w3(32'h3a6950dc),
	.w4(32'h3a7897be),
	.w5(32'h37cccc2c),
	.w6(32'h3a105a43),
	.w7(32'hb988e652),
	.w8(32'hba27e89a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2a7d1),
	.w1(32'hba3abf24),
	.w2(32'hba6217ff),
	.w3(32'h3ac22431),
	.w4(32'hbac2a127),
	.w5(32'hbaae35ef),
	.w6(32'hba8fff0a),
	.w7(32'hbac6c04b),
	.w8(32'hbab48924),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6bd883),
	.w1(32'h391ffd1d),
	.w2(32'h39edb239),
	.w3(32'hba728ad3),
	.w4(32'h398c6d7e),
	.w5(32'h39c085af),
	.w6(32'h374940f9),
	.w7(32'h39a4982a),
	.w8(32'h39fd3e5c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c626b),
	.w1(32'hb912c0fd),
	.w2(32'hb9223b57),
	.w3(32'h3a19248d),
	.w4(32'h382a1f14),
	.w5(32'h38526a82),
	.w6(32'hb8d25706),
	.w7(32'hb96cb1ba),
	.w8(32'hb8a13a49),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ef1a0),
	.w1(32'hb4f17b2e),
	.w2(32'hb8c712ac),
	.w3(32'h39705b32),
	.w4(32'h38fe2261),
	.w5(32'h38f7b346),
	.w6(32'h38775562),
	.w7(32'hb958fd1b),
	.w8(32'h370307cf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ab742),
	.w1(32'h39ac63ab),
	.w2(32'h390e71ca),
	.w3(32'h39aceb31),
	.w4(32'h3a1c217f),
	.w5(32'h39ebaf8c),
	.w6(32'h3a083688),
	.w7(32'h391c59d0),
	.w8(32'h3986f5e2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398846b3),
	.w1(32'hb8c31cd9),
	.w2(32'hb98b0d4a),
	.w3(32'h39ed992f),
	.w4(32'hb96e8fc6),
	.w5(32'hb9ae3d18),
	.w6(32'hb99b2315),
	.w7(32'hb9d252d8),
	.w8(32'hb8d195ff),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930d964),
	.w1(32'hb9929272),
	.w2(32'h3a6f4514),
	.w3(32'hb74c18ef),
	.w4(32'h3a6b070b),
	.w5(32'h3a51af39),
	.w6(32'h3876d4f4),
	.w7(32'hb98f62fc),
	.w8(32'hb9194cad),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a97cd),
	.w1(32'h39b04731),
	.w2(32'h39a0dbd7),
	.w3(32'h3ac5ca09),
	.w4(32'h3a485b13),
	.w5(32'h39d97b71),
	.w6(32'hb9a6fa17),
	.w7(32'hb929186f),
	.w8(32'hb90d3873),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6364d0),
	.w1(32'h3a33643b),
	.w2(32'h391cc0f9),
	.w3(32'h3a0abb64),
	.w4(32'h3a232ad9),
	.w5(32'h3810ff97),
	.w6(32'h3a6b852e),
	.w7(32'h39d3c627),
	.w8(32'h390bfa71),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9df474),
	.w1(32'h3a066c6c),
	.w2(32'hb884622f),
	.w3(32'h3a9232d0),
	.w4(32'h39204972),
	.w5(32'hba18c290),
	.w6(32'h38650ed6),
	.w7(32'hba297389),
	.w8(32'h38bc9353),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc6b34),
	.w1(32'h3a9c51f7),
	.w2(32'h3a6e35b6),
	.w3(32'h3821ccc7),
	.w4(32'h3aaed2c8),
	.w5(32'h3a8806d3),
	.w6(32'h3ab0b054),
	.w7(32'h3a626e50),
	.w8(32'h3a67a175),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd359),
	.w1(32'h3b17f036),
	.w2(32'h3a275a5d),
	.w3(32'h3ab0216d),
	.w4(32'h3adf4736),
	.w5(32'h3a256f6d),
	.w6(32'h3b23b739),
	.w7(32'h3a97cf65),
	.w8(32'h3ade5ac8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2a2a4),
	.w1(32'h3995db70),
	.w2(32'hb98af3c7),
	.w3(32'h3a679049),
	.w4(32'h38fe482c),
	.w5(32'hb8e94f66),
	.w6(32'h3a068fb0),
	.w7(32'hb88d598a),
	.w8(32'hb933860c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39821a2d),
	.w1(32'h3a7cd08c),
	.w2(32'h3a0c9bc9),
	.w3(32'h39bad075),
	.w4(32'h3a3b4ed9),
	.w5(32'h39fcb7b3),
	.w6(32'h3a82015b),
	.w7(32'h39d166bf),
	.w8(32'h3a399b32),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51ba02),
	.w1(32'h38cb300c),
	.w2(32'hb8238273),
	.w3(32'h3a3dff6c),
	.w4(32'h393a9a87),
	.w5(32'h39384473),
	.w6(32'hb932a3ff),
	.w7(32'hb8ac52e2),
	.w8(32'hb8daa09a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39038208),
	.w1(32'h3a30ed29),
	.w2(32'h3a6b9c8a),
	.w3(32'h399617d4),
	.w4(32'h384ff7e1),
	.w5(32'h3a05c6ed),
	.w6(32'h3a38afcc),
	.w7(32'h3a822c86),
	.w8(32'h3aab7dbf),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c8526),
	.w1(32'h3a9a777c),
	.w2(32'h3a65dd89),
	.w3(32'h39aeb32d),
	.w4(32'h3aab8467),
	.w5(32'h3aa792a9),
	.w6(32'h3aafb4c9),
	.w7(32'h3a94bb6d),
	.w8(32'h3a86dab3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcd30d),
	.w1(32'h39dd7f59),
	.w2(32'h3a1620da),
	.w3(32'h3abf4768),
	.w4(32'hb9e898de),
	.w5(32'h38f76686),
	.w6(32'h3a14d789),
	.w7(32'hb9a0fd85),
	.w8(32'hba00d2fb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f6708),
	.w1(32'h3a1d365a),
	.w2(32'h39a93aab),
	.w3(32'h39625dac),
	.w4(32'h3a6c01fd),
	.w5(32'h3a1b9859),
	.w6(32'h3a15a629),
	.w7(32'h39f13297),
	.w8(32'h39b09d12),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc0d07),
	.w1(32'h39fe0b9c),
	.w2(32'hba1a4b23),
	.w3(32'h3ab0db04),
	.w4(32'hb8f53535),
	.w5(32'hb9ee3539),
	.w6(32'h399c7b26),
	.w7(32'hb9f02749),
	.w8(32'hb96d10da),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391667c3),
	.w1(32'h3a39a60e),
	.w2(32'h39c1b850),
	.w3(32'h39c7cc8f),
	.w4(32'h3a85ae35),
	.w5(32'h3a14852a),
	.w6(32'h3a880838),
	.w7(32'h39f4de1a),
	.w8(32'h3a019a6f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f95fe4),
	.w1(32'h394dd716),
	.w2(32'hb97f2e09),
	.w3(32'h39db94bd),
	.w4(32'h39b370cc),
	.w5(32'h391fd280),
	.w6(32'h39c25fd4),
	.w7(32'h3912274e),
	.w8(32'h374a8121),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafa315),
	.w1(32'h3ab3d7d5),
	.w2(32'h391b2717),
	.w3(32'h3a86e5f9),
	.w4(32'h3ab58865),
	.w5(32'h39cf197c),
	.w6(32'h3aaf538f),
	.w7(32'h3a557ecf),
	.w8(32'h39ec17c1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8beef),
	.w1(32'h3ac0dc21),
	.w2(32'h3a20b2df),
	.w3(32'h3ab75a08),
	.w4(32'h3aeba3d6),
	.w5(32'h3aa69c04),
	.w6(32'h3addda24),
	.w7(32'h3a6566b5),
	.w8(32'h3a3a1f91),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f3509),
	.w1(32'h3b56ef42),
	.w2(32'h3a5dbb7c),
	.w3(32'h3b40c26a),
	.w4(32'h3b187deb),
	.w5(32'h3a2668be),
	.w6(32'h3b52cb49),
	.w7(32'h3a58c202),
	.w8(32'h3abbf769),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac48a3c),
	.w1(32'hb8824e7a),
	.w2(32'hb9d3e2aa),
	.w3(32'h3a54de69),
	.w4(32'hb9952ddc),
	.w5(32'hb9cd33d8),
	.w6(32'h38bdd5e6),
	.w7(32'h366b33bf),
	.w8(32'h38649f20),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8819af),
	.w1(32'h39b44354),
	.w2(32'h39f8ced0),
	.w3(32'h3a8565a8),
	.w4(32'h39cd3062),
	.w5(32'h3a20e1f1),
	.w6(32'hb87881e1),
	.w7(32'hb9d321ea),
	.w8(32'hba67deda),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba101917),
	.w1(32'h39c0d5ac),
	.w2(32'hb913262c),
	.w3(32'h392ce832),
	.w4(32'h39a60aea),
	.w5(32'hb995023e),
	.w6(32'h37beb8de),
	.w7(32'hb902aff4),
	.w8(32'h39cbbd67),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b11f),
	.w1(32'h38e29cc8),
	.w2(32'hba60aa3a),
	.w3(32'h3a90e497),
	.w4(32'h39cfbf12),
	.w5(32'hba23bda3),
	.w6(32'h3918c154),
	.w7(32'hba5d0c83),
	.w8(32'h38dabfd0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f8c92),
	.w1(32'h39aa63b6),
	.w2(32'hb935c7e3),
	.w3(32'h3a3baef8),
	.w4(32'hb8485b67),
	.w5(32'hba1a6a73),
	.w6(32'h3811eb8b),
	.w7(32'h385d6399),
	.w8(32'h38b83163),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e99ab),
	.w1(32'h3ace32de),
	.w2(32'h39f8d70d),
	.w3(32'h3a2006e8),
	.w4(32'h3abe5494),
	.w5(32'h3a39544a),
	.w6(32'h3aaf6b11),
	.w7(32'h39c6c7af),
	.w8(32'h39ea0f00),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25d9e6),
	.w1(32'hb924ad45),
	.w2(32'hbada46f1),
	.w3(32'h3b478798),
	.w4(32'hba6bc424),
	.w5(32'hbb1b7cfa),
	.w6(32'hba04637a),
	.w7(32'hbab9b4ef),
	.w8(32'hbaa888f9),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ecf46),
	.w1(32'hba97f115),
	.w2(32'hbb299931),
	.w3(32'h3b1365b5),
	.w4(32'hbabb3659),
	.w5(32'hbabfb174),
	.w6(32'hba910519),
	.w7(32'hbb1219b6),
	.w8(32'hbaa64cc8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aa9f3),
	.w1(32'h3a97dff8),
	.w2(32'h39e9f313),
	.w3(32'h3a6ccb94),
	.w4(32'h39ecb79f),
	.w5(32'h390808e1),
	.w6(32'h3a7bf50e),
	.w7(32'h38a1e496),
	.w8(32'h38ef19ff),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879d56c),
	.w1(32'hb8cc78de),
	.w2(32'h373222ac),
	.w3(32'hb906978a),
	.w4(32'hb3b214b1),
	.w5(32'h3902774c),
	.w6(32'h39232fbc),
	.w7(32'hb82a8efb),
	.w8(32'h3903c0d3),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25c861),
	.w1(32'h39dd2108),
	.w2(32'h39e59b60),
	.w3(32'h3a478855),
	.w4(32'h39dae1f0),
	.w5(32'h38e35792),
	.w6(32'h3a123580),
	.w7(32'hb84eab90),
	.w8(32'h374959f5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb781c8da),
	.w1(32'h3a152099),
	.w2(32'h39aa76ac),
	.w3(32'hb97eb6df),
	.w4(32'h3996f74e),
	.w5(32'h39abd77e),
	.w6(32'h39d66a94),
	.w7(32'h39b75062),
	.w8(32'h39c10386),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393adb72),
	.w1(32'hb9916608),
	.w2(32'hb9aa95fa),
	.w3(32'h3907cde2),
	.w4(32'h3875f0a6),
	.w5(32'hb98293e1),
	.w6(32'h38a54013),
	.w7(32'h39bf9d0d),
	.w8(32'h39c2d3d1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e41d95),
	.w1(32'h3a0b3d1f),
	.w2(32'h362ca3d5),
	.w3(32'hb6322dfa),
	.w4(32'h3a7dc450),
	.w5(32'h3a35990f),
	.w6(32'h3a4867de),
	.w7(32'h39f38739),
	.w8(32'h39d20bbf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2ead5),
	.w1(32'h39bca445),
	.w2(32'hb9f3e499),
	.w3(32'h3a59d2a4),
	.w4(32'h37637c07),
	.w5(32'hb968e206),
	.w6(32'h3a4a7d71),
	.w7(32'hb9e84a32),
	.w8(32'h3875e048),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ab9e9),
	.w1(32'hba9261d8),
	.w2(32'hbabd56f3),
	.w3(32'h39e0a138),
	.w4(32'hba847a6e),
	.w5(32'hbaad802e),
	.w6(32'hba520ed9),
	.w7(32'hbad031c2),
	.w8(32'hbab1cc3d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8589ad0),
	.w1(32'hb709ee8f),
	.w2(32'hb8819802),
	.w3(32'hb9800c99),
	.w4(32'hb8d60cb2),
	.w5(32'hb9312bf1),
	.w6(32'h39ababde),
	.w7(32'hb99da7ba),
	.w8(32'hba22c09c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a441c61),
	.w1(32'h39cd1ea2),
	.w2(32'h392918c4),
	.w3(32'h3a810401),
	.w4(32'h3923efc7),
	.w5(32'hba236882),
	.w6(32'h386b08ff),
	.w7(32'hb94e9678),
	.w8(32'hba3b1ad4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a01424),
	.w1(32'h3955cb92),
	.w2(32'hb954b6b2),
	.w3(32'hb9aad8a4),
	.w4(32'h38bc5aec),
	.w5(32'hb899a500),
	.w6(32'h397e94b9),
	.w7(32'hb9f2ee4c),
	.w8(32'hb9a71f07),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93ef0a),
	.w1(32'h39880ef6),
	.w2(32'hb9737e93),
	.w3(32'h3a5a0bc0),
	.w4(32'hb9af3936),
	.w5(32'hb9fe4e3d),
	.w6(32'h39afaa16),
	.w7(32'hb820f65e),
	.w8(32'h390b4d30),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a913662),
	.w1(32'h3975b81c),
	.w2(32'hba1008bd),
	.w3(32'h3a5ac345),
	.w4(32'h39580068),
	.w5(32'h36826aeb),
	.w6(32'h3a1225f5),
	.w7(32'hba24258f),
	.w8(32'hba0d3b2a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efd26e),
	.w1(32'h39d11d18),
	.w2(32'h3917a89e),
	.w3(32'hb8177363),
	.w4(32'h39aaba13),
	.w5(32'h38f0f6b0),
	.w6(32'h3a038af6),
	.w7(32'h38fb9309),
	.w8(32'h39076c5b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb756b7b1),
	.w1(32'h39a1baed),
	.w2(32'h39392dd1),
	.w3(32'hb88282a4),
	.w4(32'h395b9b96),
	.w5(32'h3892aff2),
	.w6(32'h39deff85),
	.w7(32'h39756b1e),
	.w8(32'h3919c15c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390478a5),
	.w1(32'h39bafb5e),
	.w2(32'h38f836e8),
	.w3(32'h38a3a107),
	.w4(32'h39a18b8f),
	.w5(32'h38e07ad7),
	.w6(32'h39e1a2bc),
	.w7(32'h38e9753b),
	.w8(32'h385eaaba),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cd39d),
	.w1(32'hba904707),
	.w2(32'h39060d19),
	.w3(32'hb7412061),
	.w4(32'hbaa89988),
	.w5(32'hba9a6f2f),
	.w6(32'hba656ff9),
	.w7(32'hb98f4297),
	.w8(32'hba3a1844),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d68bd),
	.w1(32'hb8a351c6),
	.w2(32'hb95df3db),
	.w3(32'h3989588d),
	.w4(32'hba3e097a),
	.w5(32'hb9c08431),
	.w6(32'hb8c7adc2),
	.w7(32'hb931ac2d),
	.w8(32'h3a6d5762),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a628f68),
	.w1(32'h3983a5cf),
	.w2(32'h38bf2698),
	.w3(32'h3a6668e0),
	.w4(32'h3a02e142),
	.w5(32'h3a4b7545),
	.w6(32'h39bda139),
	.w7(32'h3a065ba6),
	.w8(32'h39ad0e14),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17eb6e),
	.w1(32'h3a609e22),
	.w2(32'h37f1505e),
	.w3(32'h3a45dbf6),
	.w4(32'h3a816f9f),
	.w5(32'h3a7dcaed),
	.w6(32'h39ea4195),
	.w7(32'hb85542a9),
	.w8(32'h38a2e64e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f7ad38),
	.w1(32'h394b50ba),
	.w2(32'h38ad2ca6),
	.w3(32'h3a6d17aa),
	.w4(32'h39792a46),
	.w5(32'h38dd710b),
	.w6(32'h3940fc1a),
	.w7(32'hb87cd6bf),
	.w8(32'hb6719f72),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6c2a2),
	.w1(32'hbaf935e2),
	.w2(32'hb93e3e50),
	.w3(32'h38fa06c5),
	.w4(32'hbae8103d),
	.w5(32'hba781eb6),
	.w6(32'hbaeb6983),
	.w7(32'hbaaa93ed),
	.w8(32'hbad0443b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbfc64),
	.w1(32'h3af4c36f),
	.w2(32'h3a7f49a9),
	.w3(32'hba8833ee),
	.w4(32'h3b1aca4b),
	.w5(32'h3b08bcb1),
	.w6(32'h3abf0a9f),
	.w7(32'h39e6912c),
	.w8(32'h3a19bc0f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accea6d),
	.w1(32'h3a85e5fc),
	.w2(32'h3a1fad14),
	.w3(32'h3b112ee4),
	.w4(32'h3ac516f3),
	.w5(32'h3aa4b535),
	.w6(32'h3a8ae41f),
	.w7(32'h3a434cac),
	.w8(32'h3a3ef4e4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a538ebd),
	.w1(32'h39056c44),
	.w2(32'hb8d48c67),
	.w3(32'h3a849839),
	.w4(32'h37c044a6),
	.w5(32'hb93dc0d9),
	.w6(32'h378c2972),
	.w7(32'hb8bda71d),
	.w8(32'hb982ef1f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29fc2f),
	.w1(32'h39df513a),
	.w2(32'h389d8807),
	.w3(32'h3a25a58a),
	.w4(32'h39774dd8),
	.w5(32'hb8812327),
	.w6(32'h39f3b888),
	.w7(32'h3916781f),
	.w8(32'h393bb476),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad76f1),
	.w1(32'h3a0cb00e),
	.w2(32'hba0f1bb8),
	.w3(32'h3a43ebec),
	.w4(32'h381eca43),
	.w5(32'hba11e587),
	.w6(32'h3a0c0c30),
	.w7(32'hb9823db1),
	.w8(32'hba2843aa),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5830ba3),
	.w1(32'h359e6e39),
	.w2(32'h3717cd6d),
	.w3(32'hb742d7a8),
	.w4(32'h362d427c),
	.w5(32'h3719e740),
	.w6(32'h373867cb),
	.w7(32'h371ecf7a),
	.w8(32'h376c12a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38adce3f),
	.w1(32'h390693a7),
	.w2(32'hb825b368),
	.w3(32'h388ac140),
	.w4(32'h3716bd7b),
	.w5(32'hb94fc8ac),
	.w6(32'h33743694),
	.w7(32'hb7b7619d),
	.w8(32'hb96dea47),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902821d),
	.w1(32'h38e02939),
	.w2(32'h37907ea9),
	.w3(32'h38b5b513),
	.w4(32'h373fd997),
	.w5(32'hb83c28fe),
	.w6(32'h3848333c),
	.w7(32'h37504d0d),
	.w8(32'hb869d744),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2d03),
	.w1(32'h393bb523),
	.w2(32'hb80c602e),
	.w3(32'h39c1caf3),
	.w4(32'h38c345bd),
	.w5(32'h38989ae7),
	.w6(32'h399d0bce),
	.w7(32'hb89b8d64),
	.w8(32'h38831ad3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a58c9),
	.w1(32'hb92b10c9),
	.w2(32'hba07cf15),
	.w3(32'h397a3fb6),
	.w4(32'hb9a7fdf8),
	.w5(32'hba11a62b),
	.w6(32'h38cbe280),
	.w7(32'hb9c6d141),
	.w8(32'hba0144e8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67dd80),
	.w1(32'h39ccc9e0),
	.w2(32'h39002efe),
	.w3(32'h3a179eec),
	.w4(32'hb86289d5),
	.w5(32'hb980761f),
	.w6(32'h3a0496fe),
	.w7(32'hb893c6bf),
	.w8(32'hb909bf51),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3afd14),
	.w1(32'h39a834ef),
	.w2(32'hb844c3a7),
	.w3(32'h3a0805d0),
	.w4(32'h3979d32b),
	.w5(32'hb796c2f4),
	.w6(32'h39ba2b4c),
	.w7(32'hb8860d97),
	.w8(32'h368e4c7f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5bd76),
	.w1(32'h3a01583a),
	.w2(32'hb7e6bf5e),
	.w3(32'h3a696563),
	.w4(32'h395e9461),
	.w5(32'hb9771bbe),
	.w6(32'h3a3f239d),
	.w7(32'hb92166c5),
	.w8(32'hb9774dff),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a715053),
	.w1(32'h39fa264b),
	.w2(32'h395b1764),
	.w3(32'h3a589f27),
	.w4(32'h39b19600),
	.w5(32'h3920fc18),
	.w6(32'h3a1d39c2),
	.w7(32'h391a5290),
	.w8(32'h38fb20d2),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eda36a),
	.w1(32'h39460979),
	.w2(32'h397640cc),
	.w3(32'h39aca3bd),
	.w4(32'h397bcdb3),
	.w5(32'h38b549cb),
	.w6(32'h393dd9ed),
	.w7(32'h392a054f),
	.w8(32'h3889ffd0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaedfdc),
	.w1(32'h3a27e7a4),
	.w2(32'h380273a7),
	.w3(32'h3a534526),
	.w4(32'h38eda575),
	.w5(32'hb8d84628),
	.w6(32'h3a2c365b),
	.w7(32'hb90927fb),
	.w8(32'h389d43c3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8d88a),
	.w1(32'h392867c4),
	.w2(32'hb8a5f85f),
	.w3(32'h39bcd8c2),
	.w4(32'h390098de),
	.w5(32'hb7b756c4),
	.w6(32'h396e2115),
	.w7(32'hb783cf45),
	.w8(32'h380c109b),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac67480),
	.w1(32'h3a3fe9f0),
	.w2(32'h39d5b7a8),
	.w3(32'h3a8e01da),
	.w4(32'h39a500c2),
	.w5(32'h38c982d2),
	.w6(32'h3a1a8da4),
	.w7(32'h38c6f21c),
	.w8(32'h398f4949),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1d2bd),
	.w1(32'h3a05ffb4),
	.w2(32'h3a2852d2),
	.w3(32'h39888beb),
	.w4(32'h3992f870),
	.w5(32'h39dd2d78),
	.w6(32'h397b75db),
	.w7(32'hb5786f1a),
	.w8(32'h3968855f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb58fe279),
	.w1(32'h36db339d),
	.w2(32'h35b04ed5),
	.w3(32'h3781b235),
	.w4(32'h36fbbe29),
	.w5(32'hb56585fe),
	.w6(32'h35a4969d),
	.w7(32'h36df1bee),
	.w8(32'h36af6ebc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35734ae5),
	.w1(32'hb683b216),
	.w2(32'hb77ad267),
	.w3(32'h359a9920),
	.w4(32'h36bb23cf),
	.w5(32'hb6a15096),
	.w6(32'h370d2ecb),
	.w7(32'hb6820337),
	.w8(32'h36e67cc1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37172c75),
	.w1(32'h376f52b9),
	.w2(32'h370da849),
	.w3(32'hb5c742a8),
	.w4(32'h370baf47),
	.w5(32'h377ae908),
	.w6(32'hb680297c),
	.w7(32'h361e5cfb),
	.w8(32'h37535df7),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27717b),
	.w1(32'h39b8f440),
	.w2(32'h3a391262),
	.w3(32'h39ad9104),
	.w4(32'hb8dacc99),
	.w5(32'h3932c27c),
	.w6(32'h394afe7b),
	.w7(32'hb94b4351),
	.w8(32'hb8fa9ab3),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab16a86),
	.w1(32'h3a68e393),
	.w2(32'hb8eb7976),
	.w3(32'h3a7c62b2),
	.w4(32'h3a78c41b),
	.w5(32'h39d0babd),
	.w6(32'h39b00a00),
	.w7(32'h3a068c14),
	.w8(32'h39e844c3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fd56a5),
	.w1(32'h373f5571),
	.w2(32'h3635268a),
	.w3(32'hb75afb52),
	.w4(32'h36e24476),
	.w5(32'hb5c48316),
	.w6(32'hb62ce9b7),
	.w7(32'hb6c310cd),
	.w8(32'h363dcc9e),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa15c81),
	.w1(32'h39ac401e),
	.w2(32'hb9713f15),
	.w3(32'h3a44cc5f),
	.w4(32'h38cb02ad),
	.w5(32'hb95cf25d),
	.w6(32'h39b0beb5),
	.w7(32'hb96135d3),
	.w8(32'h386224a9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c30bc),
	.w1(32'h399d3831),
	.w2(32'hb9442b52),
	.w3(32'h3a37fa40),
	.w4(32'hb8a97888),
	.w5(32'hb9bc27c1),
	.w6(32'h39ce9386),
	.w7(32'hb9e235a9),
	.w8(32'hb9e86a14),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84b89c),
	.w1(32'h39ef2594),
	.w2(32'hb8cf0384),
	.w3(32'h3a4964bf),
	.w4(32'h3755de89),
	.w5(32'hb9de3969),
	.w6(32'h3a0d4e21),
	.w7(32'hb9228c03),
	.w8(32'hb9e3ee3e),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe6c0a),
	.w1(32'h3969bb35),
	.w2(32'h36cd4468),
	.w3(32'h397021f2),
	.w4(32'hb7c1fbf7),
	.w5(32'hb953c254),
	.w6(32'h385f23bb),
	.w7(32'hb94ff31a),
	.w8(32'hb99808ca),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c21ab3),
	.w1(32'h38c483df),
	.w2(32'h399b5b48),
	.w3(32'hb834c80a),
	.w4(32'hb8ba03da),
	.w5(32'h38365b58),
	.w6(32'hb8d81f8a),
	.w7(32'hb825634e),
	.w8(32'hb8af3abf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a05f3),
	.w1(32'hb760e79b),
	.w2(32'h3638422a),
	.w3(32'hb9319347),
	.w4(32'hb9109492),
	.w5(32'hb840946b),
	.w6(32'hb99ea305),
	.w7(32'h384f1201),
	.w8(32'h3902aa0c),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0148d4),
	.w1(32'h395c5b0a),
	.w2(32'hb89c7b26),
	.w3(32'h3947c694),
	.w4(32'h3872a6c2),
	.w5(32'hb8899f09),
	.w6(32'h37cc3893),
	.w7(32'hb8fb972f),
	.w8(32'h38b1ad29),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393bb59e),
	.w1(32'hb8b0741b),
	.w2(32'h35e9289f),
	.w3(32'h39b52db4),
	.w4(32'h39b93bf8),
	.w5(32'hb9cab142),
	.w6(32'hb7805c2f),
	.w7(32'h381314a1),
	.w8(32'hb91f8324),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cb4c1),
	.w1(32'hb946ae41),
	.w2(32'hb989c692),
	.w3(32'hb9b92370),
	.w4(32'hb98f1098),
	.w5(32'hb9b03103),
	.w6(32'hb9a5f03f),
	.w7(32'hb93983e6),
	.w8(32'hb992b1ff),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76e8cfc),
	.w1(32'hb7073707),
	.w2(32'h36cabe64),
	.w3(32'h36cd2f15),
	.w4(32'hb6218e02),
	.w5(32'h36859a41),
	.w6(32'h378a5092),
	.w7(32'h35cddca5),
	.w8(32'h37638abf),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6467caf),
	.w1(32'h368c508a),
	.w2(32'h3682922a),
	.w3(32'hb682a137),
	.w4(32'h36b51c16),
	.w5(32'h36965ed5),
	.w6(32'h3728d0a9),
	.w7(32'h37152c21),
	.w8(32'h37308717),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e5950),
	.w1(32'h39bd5a14),
	.w2(32'hb752fbb7),
	.w3(32'h39b572a4),
	.w4(32'h37b8532b),
	.w5(32'hb921011b),
	.w6(32'h3904294b),
	.w7(32'hb9298e7a),
	.w8(32'hb96b8843),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62b7789),
	.w1(32'h3803b71a),
	.w2(32'hb6b22829),
	.w3(32'h36bac5b5),
	.w4(32'h38084e49),
	.w5(32'h361624ca),
	.w6(32'h381a9128),
	.w7(32'h37b4858a),
	.w8(32'hb782a83e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c5b77),
	.w1(32'h3a1a3d26),
	.w2(32'h38531396),
	.w3(32'h3a3b3502),
	.w4(32'h39a9fef0),
	.w5(32'h3924e8ac),
	.w6(32'h3a2df826),
	.w7(32'hb8d64fc2),
	.w8(32'h390a7368),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70ab434),
	.w1(32'hb850a581),
	.w2(32'hb8a0e239),
	.w3(32'h38760828),
	.w4(32'hb70a82c7),
	.w5(32'hb8e542d8),
	.w6(32'h37abd5c6),
	.w7(32'h38be4acc),
	.w8(32'hb7e667f0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba234242),
	.w1(32'hba06b0d9),
	.w2(32'hba10eb80),
	.w3(32'hba1c188d),
	.w4(32'hba05d375),
	.w5(32'hb9f06f29),
	.w6(32'hba4c0cb4),
	.w7(32'hb9e8c513),
	.w8(32'hb9bca4ac),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8607547),
	.w1(32'hb788cda1),
	.w2(32'hb7a0e790),
	.w3(32'hb84c22b1),
	.w4(32'hb7d2448b),
	.w5(32'hb7a2eded),
	.w6(32'hb83a8dd0),
	.w7(32'hb811e50f),
	.w8(32'hb803bff4),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b31116),
	.w1(32'h3752392f),
	.w2(32'hb8a90b06),
	.w3(32'hb7c2eb73),
	.w4(32'hb84cf916),
	.w5(32'hb8d4d12c),
	.w6(32'hb8c5c97e),
	.w7(32'hb7fd5fbc),
	.w8(32'h37c13407),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a787df3),
	.w1(32'h3a1ffcda),
	.w2(32'h38e15956),
	.w3(32'h3a28bb23),
	.w4(32'h394e8ef6),
	.w5(32'hb91f7735),
	.w6(32'h3a0ad9e5),
	.w7(32'hb7eb7d7b),
	.w8(32'hb98d58df),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9feff),
	.w1(32'h3a30b9ad),
	.w2(32'hb8e26e87),
	.w3(32'h3a8c07aa),
	.w4(32'hb8a43943),
	.w5(32'hb9d98378),
	.w6(32'h396543b2),
	.w7(32'hb9a501fa),
	.w8(32'hb7aa69ec),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9431190),
	.w1(32'hb5e189ff),
	.w2(32'hb94613cc),
	.w3(32'hb980968c),
	.w4(32'hb93c541c),
	.w5(32'hb94d7d80),
	.w6(32'hb8853c46),
	.w7(32'hb8b66aac),
	.w8(32'hb8dbcbc1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace2739),
	.w1(32'h3a09b3fe),
	.w2(32'hb8983b84),
	.w3(32'h3a9d9193),
	.w4(32'h38879f8c),
	.w5(32'hb998a535),
	.w6(32'h3a4b7461),
	.w7(32'hb9e3f1d1),
	.w8(32'hb9aeb38d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39197088),
	.w1(32'h38172cd8),
	.w2(32'h37356803),
	.w3(32'h38ac53f8),
	.w4(32'hb838e739),
	.w5(32'hb8341544),
	.w6(32'h378a689d),
	.w7(32'hb8a5cea2),
	.w8(32'hb8956200),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafcb22),
	.w1(32'h3a91a037),
	.w2(32'h398ed89f),
	.w3(32'h3a6a9762),
	.w4(32'h3a89719b),
	.w5(32'h38aef81b),
	.w6(32'hb9346e8b),
	.w7(32'h3a0b744c),
	.w8(32'h38d723c5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39903167),
	.w1(32'h398166a8),
	.w2(32'h3797fc57),
	.w3(32'h399b7815),
	.w4(32'h3916b6bd),
	.w5(32'hb91d3e56),
	.w6(32'hb8455801),
	.w7(32'hb87a100a),
	.w8(32'hb991f03c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeae1e2),
	.w1(32'h39f029b9),
	.w2(32'hb990d47e),
	.w3(32'h3a8c83c6),
	.w4(32'h37f56690),
	.w5(32'hb975f04b),
	.w6(32'h3a32f629),
	.w7(32'hb9bbe508),
	.w8(32'hb91ecfcd),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38826b6f),
	.w1(32'h3880d225),
	.w2(32'h378fb1df),
	.w3(32'h388d8255),
	.w4(32'h38e6097f),
	.w5(32'h38b1c1a9),
	.w6(32'h38edcbc5),
	.w7(32'h383622ed),
	.w8(32'h3832fd60),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d28ab),
	.w1(32'h3a039abf),
	.w2(32'h39b240de),
	.w3(32'h3951a16d),
	.w4(32'h38d94cad),
	.w5(32'h3928fc52),
	.w6(32'h380ae900),
	.w7(32'hb91e5636),
	.w8(32'h39197775),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37237777),
	.w1(32'hb4875d23),
	.w2(32'h35b4e107),
	.w3(32'h361b3c71),
	.w4(32'hb5f02a3d),
	.w5(32'h35e29b12),
	.w6(32'hb69285b6),
	.w7(32'hb59b4b85),
	.w8(32'h3616cf6b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39194a5a),
	.w1(32'h38a2fe7c),
	.w2(32'hb6abec8d),
	.w3(32'h3908b07a),
	.w4(32'h38cc46ad),
	.w5(32'hb7e2d06b),
	.w6(32'hb7fd36bf),
	.w7(32'h37bf0d7e),
	.w8(32'hb7ef600f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381fba0d),
	.w1(32'h38412861),
	.w2(32'h378ab72f),
	.w3(32'h3825e0a8),
	.w4(32'h384d9475),
	.w5(32'h37b75881),
	.w6(32'h37d34a91),
	.w7(32'h36c6bbc9),
	.w8(32'h37ac0015),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3987c3e7),
	.w1(32'h398f13b0),
	.w2(32'h38a6b946),
	.w3(32'hb7ae520c),
	.w4(32'h3909ace5),
	.w5(32'hb878370d),
	.w6(32'hb933e1f9),
	.w7(32'h37d044e3),
	.w8(32'hb8d13b98),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3518697d),
	.w1(32'hb7628f95),
	.w2(32'h36b98439),
	.w3(32'hb609b1f8),
	.w4(32'hb747fa3c),
	.w5(32'h3709c2a2),
	.w6(32'hb743102a),
	.w7(32'h3565d9ed),
	.w8(32'h35947002),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84ce865),
	.w1(32'hb759b73b),
	.w2(32'hb7a51ac4),
	.w3(32'hb7cb1cc5),
	.w4(32'h36313f1c),
	.w5(32'h36c2a269),
	.w6(32'hb78ebdd2),
	.w7(32'hb7239ff0),
	.w8(32'hb70f2f5a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ad1c49),
	.w1(32'h3802bf85),
	.w2(32'h37736534),
	.w3(32'h368f954b),
	.w4(32'h37b7647c),
	.w5(32'h373af6c5),
	.w6(32'h37991edf),
	.w7(32'h371ba20c),
	.w8(32'h377b34f4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15a269),
	.w1(32'h39bad53a),
	.w2(32'hb92fa764),
	.w3(32'h3a00b69c),
	.w4(32'h3834069f),
	.w5(32'hb9813546),
	.w6(32'h39917fe4),
	.w7(32'hb90f32a3),
	.w8(32'hb9e2aafa),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383caf16),
	.w1(32'hb7c64e47),
	.w2(32'h374fb943),
	.w3(32'h380e556a),
	.w4(32'hb8226056),
	.w5(32'hb84647ff),
	.w6(32'h37fd4994),
	.w7(32'h37829fc4),
	.w8(32'hb6b24773),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ac4bf),
	.w1(32'hb8e52488),
	.w2(32'hb8dd7b1a),
	.w3(32'hb7d60434),
	.w4(32'hb7109b16),
	.w5(32'hb8e53a2e),
	.w6(32'hb957e36d),
	.w7(32'hb6fadda6),
	.w8(32'hb865ca6c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af78d17),
	.w1(32'h3987b833),
	.w2(32'hba377da5),
	.w3(32'h3a88ecf0),
	.w4(32'h39986728),
	.w5(32'hb957dd28),
	.w6(32'h398f3b70),
	.w7(32'h37d4ff82),
	.w8(32'h39ea6acd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dfb6bb),
	.w1(32'h38c90134),
	.w2(32'h38a1b391),
	.w3(32'h39c78d5a),
	.w4(32'hb92b7c6f),
	.w5(32'hb900f771),
	.w6(32'hb94880b1),
	.w7(32'hba05255a),
	.w8(32'hba150ccf),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8506bc3),
	.w1(32'h369bed58),
	.w2(32'hb7b2848a),
	.w3(32'hb875c792),
	.w4(32'hb7472e9b),
	.w5(32'hb7a62cb5),
	.w6(32'hb88d39d1),
	.w7(32'h3696e8b3),
	.w8(32'hb50fd421),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3607ca35),
	.w1(32'h37a69022),
	.w2(32'hb7f0f1dc),
	.w3(32'h34cb008b),
	.w4(32'h38089a94),
	.w5(32'hb74664f5),
	.w6(32'h3765c622),
	.w7(32'hb71b3d53),
	.w8(32'h35af814a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4e36ac2),
	.w1(32'hb660dfb7),
	.w2(32'h37990417),
	.w3(32'h3851f0d2),
	.w4(32'hb5e7638f),
	.w5(32'h38779124),
	.w6(32'h3714a086),
	.w7(32'hb5857660),
	.w8(32'h3834c689),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36df8311),
	.w1(32'hb303fe13),
	.w2(32'h35f9c6d1),
	.w3(32'h37244982),
	.w4(32'hb58d0ca6),
	.w5(32'hb51e3109),
	.w6(32'h368269c0),
	.w7(32'hb61c2dc9),
	.w8(32'h36df45cf),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a1ed4),
	.w1(32'h393ca068),
	.w2(32'h38c77f0e),
	.w3(32'h389635b0),
	.w4(32'h38227b9e),
	.w5(32'hb7a47cb9),
	.w6(32'h38b910c4),
	.w7(32'hb7dcb9db),
	.w8(32'hb906ba7d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd7850),
	.w1(32'h3a359b58),
	.w2(32'h39fa39c7),
	.w3(32'h3ac224e2),
	.w4(32'h3a43d1a5),
	.w5(32'h39dac844),
	.w6(32'h3a1a02b2),
	.w7(32'h390b0564),
	.w8(32'hb970a012),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a603869),
	.w1(32'hb76f5007),
	.w2(32'hb9159aba),
	.w3(32'h3a252153),
	.w4(32'hb419d973),
	.w5(32'h38b15954),
	.w6(32'h39d18d25),
	.w7(32'hb9a3171b),
	.w8(32'hb8f1aeb0),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adf940),
	.w1(32'h3981aa5b),
	.w2(32'hb81eb192),
	.w3(32'h3942bc9b),
	.w4(32'h38ba935f),
	.w5(32'h36c92978),
	.w6(32'h38f188b0),
	.w7(32'hb94193a5),
	.w8(32'hb82586fc),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6881f6),
	.w1(32'h39216555),
	.w2(32'hb9d71c74),
	.w3(32'h3a52c305),
	.w4(32'hb92e8d66),
	.w5(32'hba0fcb50),
	.w6(32'h3a0542c9),
	.w7(32'hb9c587b3),
	.w8(32'hb9de2e06),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d24d9),
	.w1(32'h3831680e),
	.w2(32'hb7da6eda),
	.w3(32'h38f7edb3),
	.w4(32'h384e8e67),
	.w5(32'h37a78819),
	.w6(32'h385655c1),
	.w7(32'hb66134ea),
	.w8(32'hb7b4f7bd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6028cfc),
	.w1(32'hb68200bc),
	.w2(32'h35989727),
	.w3(32'h3651d97d),
	.w4(32'hb66bd7ef),
	.w5(32'hb629675d),
	.w6(32'hb5c5b07f),
	.w7(32'h35abdb67),
	.w8(32'h369c36c0),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ff3acc),
	.w1(32'h378513fe),
	.w2(32'h375b20be),
	.w3(32'hb6a8038a),
	.w4(32'h379b6950),
	.w5(32'h37998dc4),
	.w6(32'h374dcf57),
	.w7(32'h37d43e86),
	.w8(32'h3821f6fa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d7861f),
	.w1(32'h36a8dec6),
	.w2(32'h373080a6),
	.w3(32'hb7bfca91),
	.w4(32'h37130733),
	.w5(32'h3764d53e),
	.w6(32'h361af551),
	.w7(32'h37aa2d1c),
	.w8(32'h37e6e407),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c5260),
	.w1(32'h3980c6ae),
	.w2(32'h385568a4),
	.w3(32'h39fc92ee),
	.w4(32'h39105dff),
	.w5(32'h377232cb),
	.w6(32'h399880f4),
	.w7(32'hb900ac09),
	.w8(32'hb92dc0a3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80c9ad9),
	.w1(32'h37366aea),
	.w2(32'h393ae8f1),
	.w3(32'h38c5d11b),
	.w4(32'h387a6320),
	.w5(32'hb98df26f),
	.w6(32'hb9560e05),
	.w7(32'hb86e2efd),
	.w8(32'hb9867cfb),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30573a),
	.w1(32'h3956b8e2),
	.w2(32'hb8f35c4d),
	.w3(32'h39f75fce),
	.w4(32'h37aff98e),
	.w5(32'hb99e4303),
	.w6(32'h3960b99f),
	.w7(32'hb9702b95),
	.w8(32'hb9f7eb5c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90159dc),
	.w1(32'hb8c10fc1),
	.w2(32'hb918623b),
	.w3(32'hb94ff70f),
	.w4(32'hb911da21),
	.w5(32'hb904613d),
	.w6(32'hb93de5ed),
	.w7(32'hb8f462cc),
	.w8(32'hb95d35ba),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a643d40),
	.w1(32'h38dbd513),
	.w2(32'hb99d9d5c),
	.w3(32'h3a2d853b),
	.w4(32'hb86fadbb),
	.w5(32'hb9f75805),
	.w6(32'h39c4608d),
	.w7(32'hb9871954),
	.w8(32'hba118076),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a79ce6d),
	.w1(32'h39fc3ac7),
	.w2(32'hb92c691f),
	.w3(32'h3a220652),
	.w4(32'h3929a1a1),
	.w5(32'hb9120e1b),
	.w6(32'h3a09f208),
	.w7(32'h3623b113),
	.w8(32'h37d149ff),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c0993),
	.w1(32'h39161b8e),
	.w2(32'hb94fd5ad),
	.w3(32'h3a6c9b9e),
	.w4(32'h391e1ec5),
	.w5(32'hb8adc274),
	.w6(32'h398b7c38),
	.w7(32'h3856846e),
	.w8(32'h39323486),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7909ea2),
	.w1(32'hb68d00ee),
	.w2(32'h36457b3e),
	.w3(32'hb79410e9),
	.w4(32'h351f865b),
	.w5(32'h3729afc6),
	.w6(32'hb4c0eb77),
	.w7(32'h373e60ae),
	.w8(32'h378c586f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b19f58),
	.w1(32'h371b60af),
	.w2(32'hb6881d8e),
	.w3(32'hb668b9b2),
	.w4(32'h372a5c82),
	.w5(32'hb61edd51),
	.w6(32'h36d06e8a),
	.w7(32'h34a10186),
	.w8(32'h36945e85),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08e4e7),
	.w1(32'h39b02073),
	.w2(32'h3978937f),
	.w3(32'h39f51996),
	.w4(32'h394d2597),
	.w5(32'hb8203541),
	.w6(32'h394ead78),
	.w7(32'h3764fef3),
	.w8(32'hb95ff3c3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae19091),
	.w1(32'h3a510282),
	.w2(32'hb887f473),
	.w3(32'h3a864c61),
	.w4(32'hb8b6371f),
	.w5(32'hba028686),
	.w6(32'h3a37609a),
	.w7(32'hb9ffd530),
	.w8(32'hba1b7d0c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a710335),
	.w1(32'h3997b3be),
	.w2(32'hb85b6460),
	.w3(32'h3a2a9006),
	.w4(32'h38dfa1b6),
	.w5(32'hb80b3994),
	.w6(32'h39913ceb),
	.w7(32'hb954bb88),
	.w8(32'hb8e38d30),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38676db7),
	.w1(32'h386d8136),
	.w2(32'h358398eb),
	.w3(32'h372a63e2),
	.w4(32'h36acaea7),
	.w5(32'h36767dfa),
	.w6(32'h37428c2b),
	.w7(32'h3754fb05),
	.w8(32'h37d53e14),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f0291f),
	.w1(32'h36ebb91e),
	.w2(32'h378ab051),
	.w3(32'hb6b2fa73),
	.w4(32'h36778ce3),
	.w5(32'h37aeeca0),
	.w6(32'hb76ccc2d),
	.w7(32'hb68b889c),
	.w8(32'h37772482),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377dc3ce),
	.w1(32'h37cb12bc),
	.w2(32'h376276a8),
	.w3(32'h373bad02),
	.w4(32'hb6d7455e),
	.w5(32'h37bb17ce),
	.w6(32'h374db055),
	.w7(32'h3756c479),
	.w8(32'h375d5009),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8bbce),
	.w1(32'hb96b0295),
	.w2(32'hb936dd64),
	.w3(32'hb8b377ac),
	.w4(32'hb97d85bd),
	.w5(32'hb952dfa0),
	.w6(32'hb880764d),
	.w7(32'hb926587c),
	.w8(32'hb954943f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6c446),
	.w1(32'h39d3cc50),
	.w2(32'hb79ba580),
	.w3(32'h3a658ed2),
	.w4(32'h3950ee37),
	.w5(32'h387923d2),
	.w6(32'h3a024fd5),
	.w7(32'h398cbd3a),
	.w8(32'h399a0dfe),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3843fd8d),
	.w1(32'hb8b6cb69),
	.w2(32'h37a9342c),
	.w3(32'hb877745d),
	.w4(32'hb91d51d7),
	.w5(32'hb8a9a9d8),
	.w6(32'h37a46831),
	.w7(32'hb8a121e9),
	.w8(32'h36a0cc62),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39350c4b),
	.w1(32'h389073a2),
	.w2(32'h37411c68),
	.w3(32'h397586f5),
	.w4(32'h38aacc3b),
	.w5(32'hb9405616),
	.w6(32'h38ac1125),
	.w7(32'h38ce3d0f),
	.w8(32'hb99aafbc),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a445332),
	.w1(32'h39a3e965),
	.w2(32'h38f744c6),
	.w3(32'h3a2a83ba),
	.w4(32'h39055277),
	.w5(32'h38cc2022),
	.w6(32'h39c69731),
	.w7(32'hb8e19d79),
	.w8(32'hb88ec3ca),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7926511),
	.w1(32'hb64ea37f),
	.w2(32'h35772e15),
	.w3(32'hb780d923),
	.w4(32'hb481ee22),
	.w5(32'h360426a0),
	.w6(32'hb5bba93f),
	.w7(32'h343cf879),
	.w8(32'h360d737c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b159cc),
	.w1(32'hb724afbd),
	.w2(32'hb680901c),
	.w3(32'hb63a73b4),
	.w4(32'hb6ccdbc9),
	.w5(32'hb66aaeb3),
	.w6(32'hb741520a),
	.w7(32'hb6835d65),
	.w8(32'hb33b0783),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862ada1),
	.w1(32'h37ddbfdb),
	.w2(32'hb772f3d2),
	.w3(32'h3743b9a3),
	.w4(32'hb622f2d9),
	.w5(32'hb843807b),
	.w6(32'h38106c1d),
	.w7(32'hb85f04e3),
	.w8(32'hb7b05963),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb785d502),
	.w1(32'h37b34fe1),
	.w2(32'h34ab5ed7),
	.w3(32'hb782af40),
	.w4(32'h37ac0f76),
	.w5(32'hb4bf4688),
	.w6(32'h37bc2073),
	.w7(32'h34b18a68),
	.w8(32'hb6807f4e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f40334),
	.w1(32'h370eacc7),
	.w2(32'hb921a1d2),
	.w3(32'hb881e380),
	.w4(32'hb8aaf87a),
	.w5(32'hb915498e),
	.w6(32'hb880a0de),
	.w7(32'hb900240b),
	.w8(32'hb8abbf5f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a655c62),
	.w1(32'h3a536d6f),
	.w2(32'hb810ce29),
	.w3(32'h3a2ce9ae),
	.w4(32'h39555cc6),
	.w5(32'hb9b16804),
	.w6(32'h39e3978c),
	.w7(32'hb9a05a16),
	.w8(32'hb9699d8e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a126cb8),
	.w1(32'h37ee24ba),
	.w2(32'hb8fbdf88),
	.w3(32'h39e3d4d2),
	.w4(32'hb8b36b2d),
	.w5(32'hb97fa321),
	.w6(32'h3955890e),
	.w7(32'hb98263b5),
	.w8(32'hb9875f48),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70a60ff),
	.w1(32'hb760c332),
	.w2(32'h372db430),
	.w3(32'hb64dcd6a),
	.w4(32'hb605084f),
	.w5(32'h3737883c),
	.w6(32'hb7aa182a),
	.w7(32'h36622c4b),
	.w8(32'h372d1cea),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a054ae7),
	.w1(32'h39be942c),
	.w2(32'hb874edab),
	.w3(32'h39c758d6),
	.w4(32'h38df3268),
	.w5(32'hb9326534),
	.w6(32'h396e72a6),
	.w7(32'hb7262af9),
	.w8(32'hb9a479e3),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0817d),
	.w1(32'h38289a7d),
	.w2(32'h38f2e9ae),
	.w3(32'h398b9cb3),
	.w4(32'h388c43ad),
	.w5(32'h393218a8),
	.w6(32'h38f634e5),
	.w7(32'hb8015477),
	.w8(32'h391024fe),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39740747),
	.w1(32'h390dd852),
	.w2(32'hb9248e07),
	.w3(32'h39853a2d),
	.w4(32'h391144b9),
	.w5(32'hb95486f6),
	.w6(32'h391b4480),
	.w7(32'hb79f1b66),
	.w8(32'hb9aa396c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b611d9),
	.w1(32'h39449b68),
	.w2(32'hb9397e2d),
	.w3(32'h39a2b4f6),
	.w4(32'h391fa5ed),
	.w5(32'hb90b5196),
	.w6(32'h3988e676),
	.w7(32'hb707e950),
	.w8(32'hb89e501a),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3831acc8),
	.w1(32'hb6c484e8),
	.w2(32'hb5d2582b),
	.w3(32'h3832ffbc),
	.w4(32'h36940a84),
	.w5(32'h37893313),
	.w6(32'h36901375),
	.w7(32'hb726a23a),
	.w8(32'h3786fcbf),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a11723),
	.w1(32'h37445555),
	.w2(32'hb8a0cc51),
	.w3(32'h3823d14d),
	.w4(32'hb69ebd24),
	.w5(32'hb9005ec0),
	.w6(32'hb7b1e51c),
	.w7(32'hb8136ecc),
	.w8(32'hb89fdd8d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ff9c48),
	.w1(32'h35ab7c41),
	.w2(32'hb70ae035),
	.w3(32'h370f05de),
	.w4(32'h339c067f),
	.w5(32'hb669917d),
	.w6(32'h3562e13d),
	.w7(32'h35372cae),
	.w8(32'h377da3ee),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37083dd7),
	.w1(32'hb71c1547),
	.w2(32'hb73170c8),
	.w3(32'h369e80d3),
	.w4(32'hb6d066a0),
	.w5(32'hb75f5b29),
	.w6(32'hb71d3f14),
	.w7(32'hb79d19bd),
	.w8(32'hb6c11f35),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7a018),
	.w1(32'hb9746a21),
	.w2(32'hb95f6c35),
	.w3(32'hb8f58010),
	.w4(32'hb9afb395),
	.w5(32'hb9d73e1a),
	.w6(32'hb9d5d1bb),
	.w7(32'hb9a9d9e6),
	.w8(32'hb9c0016e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad409e2),
	.w1(32'h3a3492e1),
	.w2(32'hb889db28),
	.w3(32'h3a859f04),
	.w4(32'h39555180),
	.w5(32'hb96af946),
	.w6(32'h3a35907c),
	.w7(32'hb909ce69),
	.w8(32'h38ed4289),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9345ab),
	.w1(32'h3a37bfee),
	.w2(32'h3846e326),
	.w3(32'h3a3ffe8f),
	.w4(32'h39e17a69),
	.w5(32'h38be0170),
	.w6(32'h39e229c9),
	.w7(32'h37aec333),
	.w8(32'h391209f9),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62f32f),
	.w1(32'h38b003dc),
	.w2(32'hb997c490),
	.w3(32'h39f94c50),
	.w4(32'hb95bc320),
	.w5(32'hb9a853be),
	.w6(32'h391082c3),
	.w7(32'hb987967e),
	.w8(32'hb899de07),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3873197f),
	.w1(32'h36fa0272),
	.w2(32'hb80ec663),
	.w3(32'h385e5e26),
	.w4(32'h3820499a),
	.w5(32'hb79fc256),
	.w6(32'h388f1c9c),
	.w7(32'h36b11c9e),
	.w8(32'hb7d696aa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cd59bb),
	.w1(32'h36b5639d),
	.w2(32'h36a9216a),
	.w3(32'h36827f6e),
	.w4(32'hb5b2c470),
	.w5(32'hb5e66de6),
	.w6(32'hb64bd3e9),
	.w7(32'hb620300a),
	.w8(32'h36d57111),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b26454),
	.w1(32'hb4bb80c8),
	.w2(32'h369b3329),
	.w3(32'hb7020d53),
	.w4(32'hb61dbb9e),
	.w5(32'hb63c6da3),
	.w6(32'hb703a1cd),
	.w7(32'h36ca72b5),
	.w8(32'h375944f4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379a9ca6),
	.w1(32'h3784f641),
	.w2(32'h358e2c6b),
	.w3(32'h3648d990),
	.w4(32'h3658c474),
	.w5(32'hb732a332),
	.w6(32'h369e7bab),
	.w7(32'h3784aead),
	.w8(32'h3753d3b6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a720bd),
	.w1(32'h39807c66),
	.w2(32'h39e9eae6),
	.w3(32'h392ad7a8),
	.w4(32'h394733e2),
	.w5(32'h3985ed50),
	.w6(32'hb8d807cb),
	.w7(32'h390cfde1),
	.w8(32'h394b8fd8),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d8853),
	.w1(32'hb67b1408),
	.w2(32'hb7db95bd),
	.w3(32'hb8aa3826),
	.w4(32'hb73aec23),
	.w5(32'hb6e6cd69),
	.w6(32'hb83886ba),
	.w7(32'h36f60d49),
	.w8(32'hb7aedd3d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c5bf08),
	.w1(32'h36302856),
	.w2(32'hb9451e2c),
	.w3(32'hb96b68ad),
	.w4(32'hb8ed8b92),
	.w5(32'hb960c731),
	.w6(32'hb95dbabe),
	.w7(32'hb915f008),
	.w8(32'hb92192e0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83e292c),
	.w1(32'hb7d43149),
	.w2(32'hb884117f),
	.w3(32'hb895b744),
	.w4(32'hb7c8bb17),
	.w5(32'hb899c8d4),
	.w6(32'hb7da3dbc),
	.w7(32'h38308bab),
	.w8(32'h32de7804),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371a6db4),
	.w1(32'h379eaa15),
	.w2(32'h34ed2916),
	.w3(32'h37092406),
	.w4(32'h378fc889),
	.w5(32'hb6b6a3d2),
	.w6(32'h3765bce8),
	.w7(32'h3726c611),
	.w8(32'hb768aa24),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80cae2a),
	.w1(32'hb5c48589),
	.w2(32'h36b86e80),
	.w3(32'hb841f50d),
	.w4(32'hb7742cde),
	.w5(32'h37b13847),
	.w6(32'hb8178909),
	.w7(32'hb6ea6836),
	.w8(32'h38197b16),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378aebe6),
	.w1(32'h3697f076),
	.w2(32'hb619bdeb),
	.w3(32'hb60cbd11),
	.w4(32'h3779bab5),
	.w5(32'hb6b4086c),
	.w6(32'h37b17208),
	.w7(32'h37617917),
	.w8(32'h35d151c2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09296b),
	.w1(32'h3962883a),
	.w2(32'h38fc9d3c),
	.w3(32'h3a00e935),
	.w4(32'h3914301a),
	.w5(32'h3880dede),
	.w6(32'h3987bc92),
	.w7(32'hb8a7c973),
	.w8(32'hb7745904),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3823f145),
	.w1(32'h3757b168),
	.w2(32'hb5694672),
	.w3(32'h372a17e6),
	.w4(32'hb785a641),
	.w5(32'hb6f1b0fd),
	.w6(32'hb7865cf1),
	.w7(32'hb725d793),
	.w8(32'hb3c53258),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e8648),
	.w1(32'h3ad038e8),
	.w2(32'h3abb2c35),
	.w3(32'h3ad544e7),
	.w4(32'h3a6c3a81),
	.w5(32'h3aaf852b),
	.w6(32'hb9e4ddb7),
	.w7(32'hb9f17b31),
	.w8(32'hb993ea34),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule