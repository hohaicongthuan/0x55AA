module layer_10_featuremap_69(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3cb98c),
	.w1(32'h3c161254),
	.w2(32'h3b3d75b4),
	.w3(32'h3c2b2e9e),
	.w4(32'h3ba30444),
	.w5(32'h3be25c39),
	.w6(32'hbc8b5612),
	.w7(32'hbbb67a99),
	.w8(32'hbc15c46d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d479),
	.w1(32'hbc7a8eb6),
	.w2(32'hbbfc79a1),
	.w3(32'h3bc72343),
	.w4(32'hbb26ccd6),
	.w5(32'hba1a3e5f),
	.w6(32'hbc5a7422),
	.w7(32'hbc340a7c),
	.w8(32'h3cb4be53),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1119a4),
	.w1(32'hbb55914a),
	.w2(32'h3c3342c1),
	.w3(32'hbac1d1be),
	.w4(32'hbb9fcaf5),
	.w5(32'h3afe9f8d),
	.w6(32'h3c8252ad),
	.w7(32'h3af406fe),
	.w8(32'hbc0d6e39),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb7e60),
	.w1(32'h3c03d636),
	.w2(32'hbc195acb),
	.w3(32'hbbf968b7),
	.w4(32'hbb8cfab5),
	.w5(32'hbc0d7c85),
	.w6(32'hbcde6029),
	.w7(32'hbcb0f008),
	.w8(32'h3bbd69c3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8414dd),
	.w1(32'hbb74a7fa),
	.w2(32'hbc1cb568),
	.w3(32'hbaa8aa5a),
	.w4(32'hbb71e595),
	.w5(32'hbcb7dabd),
	.w6(32'h3c651fe1),
	.w7(32'h3bf2c8d3),
	.w8(32'hbcd7232f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4d09),
	.w1(32'h3c36a6d8),
	.w2(32'h3c05e509),
	.w3(32'hbb1f1214),
	.w4(32'h3c91ff20),
	.w5(32'h3c1ddfcb),
	.w6(32'h3ab13a75),
	.w7(32'h3c5e50bc),
	.w8(32'h3b7946cd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4bda7),
	.w1(32'h3b132f8a),
	.w2(32'hbbbe2621),
	.w3(32'h3b3ad963),
	.w4(32'hbb29ecb3),
	.w5(32'h3b8f806f),
	.w6(32'hbaa48f7c),
	.w7(32'hbb510f7f),
	.w8(32'h3bd4dd6f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2511a3),
	.w1(32'hbbb1fc69),
	.w2(32'hba57987d),
	.w3(32'h3be031cf),
	.w4(32'h3b385e54),
	.w5(32'hba66c51d),
	.w6(32'h3bf92013),
	.w7(32'h3bb52045),
	.w8(32'h3b0d9d68),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b320982),
	.w1(32'h3bab5468),
	.w2(32'h3bc141f1),
	.w3(32'h38957b3f),
	.w4(32'h3add40a6),
	.w5(32'h3b444ff5),
	.w6(32'h39c6a7a9),
	.w7(32'hbb8e8908),
	.w8(32'h3c150c82),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2539a0),
	.w1(32'hbb9d1f7e),
	.w2(32'h3a32b9eb),
	.w3(32'hba05d11a),
	.w4(32'hbb5cc4d4),
	.w5(32'hbb44b96f),
	.w6(32'h3bfe6c8d),
	.w7(32'hbac32dcf),
	.w8(32'hbb5a4e7b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97202c),
	.w1(32'h39093c7f),
	.w2(32'h3c25c2fa),
	.w3(32'hbafd0d81),
	.w4(32'hbb2b11c8),
	.w5(32'h3c3337ef),
	.w6(32'hbac8087b),
	.w7(32'hbb6f4d20),
	.w8(32'hbb866bc5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c277120),
	.w1(32'h3c190bd4),
	.w2(32'hb9ead0ba),
	.w3(32'hbb43be0b),
	.w4(32'hbc300e23),
	.w5(32'hbb125b77),
	.w6(32'hbcab6561),
	.w7(32'hbc8d5f53),
	.w8(32'hbaf3787a),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba961d6b),
	.w1(32'hbafe0203),
	.w2(32'hba9864ba),
	.w3(32'h399ed953),
	.w4(32'hbafd37f0),
	.w5(32'h3c099b0e),
	.w6(32'hbad22d1d),
	.w7(32'hbb4fc78e),
	.w8(32'h3968f220),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba0bd),
	.w1(32'h3b7e81d0),
	.w2(32'hbb761543),
	.w3(32'h3c031315),
	.w4(32'h3bdc48f1),
	.w5(32'h3bd8f381),
	.w6(32'h3b146fd6),
	.w7(32'h3c016f4a),
	.w8(32'h3c7cf9f8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c6ed1),
	.w1(32'hbc1e0a0b),
	.w2(32'h3b1ec80d),
	.w3(32'h3c21f057),
	.w4(32'h3b7f5ba1),
	.w5(32'h3bd45ca1),
	.w6(32'h3c4b6d71),
	.w7(32'h3beaa365),
	.w8(32'h3c0e520b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39786062),
	.w1(32'hbbcbf7b8),
	.w2(32'h3b29dffb),
	.w3(32'h3b1d95d1),
	.w4(32'hbbbcf206),
	.w5(32'hb9bdfcf8),
	.w6(32'h3c1868ae),
	.w7(32'h3ad55372),
	.w8(32'h39192ce3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5402),
	.w1(32'h3a1c7ad1),
	.w2(32'h3b53ba9c),
	.w3(32'hb9e20a0d),
	.w4(32'hbb100a24),
	.w5(32'h3c29a104),
	.w6(32'h394ff2b4),
	.w7(32'hbabe8cf1),
	.w8(32'h3c79fc97),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08788e),
	.w1(32'hbab035ba),
	.w2(32'hba41c353),
	.w3(32'h3ba51fc8),
	.w4(32'hb92b2948),
	.w5(32'h3afd6a40),
	.w6(32'h3c7eb36f),
	.w7(32'h3c35ef00),
	.w8(32'h3b970123),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e5f2d),
	.w1(32'h3bc56eea),
	.w2(32'h3af7167c),
	.w3(32'h3b1af93d),
	.w4(32'h3b30679a),
	.w5(32'hbad42a93),
	.w6(32'hbb7cc51c),
	.w7(32'hbb5bdeb1),
	.w8(32'hbb906487),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399690a7),
	.w1(32'hba8137ca),
	.w2(32'h39dedb41),
	.w3(32'hbc6f2dd1),
	.w4(32'hbc5829aa),
	.w5(32'hbae96ddc),
	.w6(32'hbc8e276f),
	.w7(32'hbcbfcf5c),
	.w8(32'h3a56ad44),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388dc64a),
	.w1(32'h3ab4d9b6),
	.w2(32'h3c0b59c1),
	.w3(32'hba642b0e),
	.w4(32'hba3d90cb),
	.w5(32'hbb5c66f8),
	.w6(32'h3b43baf7),
	.w7(32'h3af6ad5f),
	.w8(32'hbb365216),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22a975),
	.w1(32'h3b786a46),
	.w2(32'h3b847b08),
	.w3(32'hbb9fa918),
	.w4(32'h3ba018c1),
	.w5(32'hba3a3fca),
	.w6(32'hbc4f1f7a),
	.w7(32'hbc31572b),
	.w8(32'hbca0e6f8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb721bd),
	.w1(32'h3b24803d),
	.w2(32'hbbb8e99a),
	.w3(32'hbba73fc6),
	.w4(32'h39e0f7ba),
	.w5(32'hbbcf71a7),
	.w6(32'hbc858387),
	.w7(32'hbba20215),
	.w8(32'hbb25ae3b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8240),
	.w1(32'hbae9048b),
	.w2(32'h3bb1f482),
	.w3(32'hbaf42086),
	.w4(32'h39fae2ae),
	.w5(32'h3b4f8c69),
	.w6(32'hbb075bb9),
	.w7(32'h3a1740e6),
	.w8(32'h3a4a1f62),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3985c),
	.w1(32'h3c0dfa84),
	.w2(32'h3c496d91),
	.w3(32'h3bd07aa4),
	.w4(32'h3b768ccf),
	.w5(32'h3c375500),
	.w6(32'hbb2858af),
	.w7(32'hbaa11e42),
	.w8(32'h3a9b091c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b98372),
	.w1(32'hbb1d70df),
	.w2(32'h3ac8fa68),
	.w3(32'hbc38f77e),
	.w4(32'hbc7d28c5),
	.w5(32'hbb82eaa8),
	.w6(32'hbbf686a2),
	.w7(32'hbc57369f),
	.w8(32'hbb602b9b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48904c),
	.w1(32'hbb4bd7e3),
	.w2(32'hb9869fa8),
	.w3(32'h3c1b9387),
	.w4(32'h3ad7c904),
	.w5(32'hbafebe85),
	.w6(32'hba413677),
	.w7(32'hbb6a61c5),
	.w8(32'hb98841ab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460a94),
	.w1(32'hba58026d),
	.w2(32'h3bba4880),
	.w3(32'h3b15b547),
	.w4(32'hbab9e02b),
	.w5(32'h3b07e5ce),
	.w6(32'hbb2e3b01),
	.w7(32'hbab62085),
	.w8(32'hbba82056),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35f0df),
	.w1(32'hbc1fcffb),
	.w2(32'hbadecb24),
	.w3(32'h3c695764),
	.w4(32'hbb445fe9),
	.w5(32'h3b1cbec1),
	.w6(32'h3b4391f4),
	.w7(32'hbc66e43c),
	.w8(32'h3b2ef6fa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7379eb),
	.w1(32'hbbd1c42d),
	.w2(32'hb9663769),
	.w3(32'h3b74fa91),
	.w4(32'hbb2f1a6e),
	.w5(32'h39936511),
	.w6(32'h3bc212fe),
	.w7(32'h39f19d11),
	.w8(32'hb9c81793),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5ffa9),
	.w1(32'h3ac61ee2),
	.w2(32'h3b001336),
	.w3(32'h3b37fe0b),
	.w4(32'h3ba1a599),
	.w5(32'h3919dd54),
	.w6(32'h3b2fb3ac),
	.w7(32'h3b9942b6),
	.w8(32'h3c27e43c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba207214),
	.w1(32'h3bab90df),
	.w2(32'hbc07c9a6),
	.w3(32'h39b04dac),
	.w4(32'h3c0a3309),
	.w5(32'hbc00becb),
	.w6(32'h3bb34d9e),
	.w7(32'h3c510207),
	.w8(32'hba946532),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c3e92),
	.w1(32'hbb94cc71),
	.w2(32'hbb405d7b),
	.w3(32'hbbce046a),
	.w4(32'h3a36c7a6),
	.w5(32'hbbc92c83),
	.w6(32'hba48163b),
	.w7(32'h3baffe6e),
	.w8(32'hbb7eda80),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba57c15),
	.w1(32'hbb9bb94a),
	.w2(32'hbb4d02ce),
	.w3(32'hbbc26bd1),
	.w4(32'hbb9851f9),
	.w5(32'h3ab3d9f4),
	.w6(32'hbb67b4f1),
	.w7(32'hbb360e1e),
	.w8(32'hbb759a5f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5976ed),
	.w1(32'h3bcee6ca),
	.w2(32'hbb6ea1a9),
	.w3(32'hbb10562d),
	.w4(32'h3bce3970),
	.w5(32'hbb6abdc1),
	.w6(32'h3b4cfe4b),
	.w7(32'h3c5e14eb),
	.w8(32'hbb19da90),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f45a),
	.w1(32'hbb8125d5),
	.w2(32'h3c0417a3),
	.w3(32'hba200e7a),
	.w4(32'hbb0929fd),
	.w5(32'h3b7c357e),
	.w6(32'h3a13c471),
	.w7(32'hbaeaac47),
	.w8(32'h3be9ebae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1dda7),
	.w1(32'h3bdc2080),
	.w2(32'h3b14e6e1),
	.w3(32'h39bf8f64),
	.w4(32'h3b8ae53e),
	.w5(32'hbb28c1f8),
	.w6(32'h3b70a0e8),
	.w7(32'h3cb20ddf),
	.w8(32'hbbb4b05f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5649d),
	.w1(32'hba3ba6f2),
	.w2(32'hba0bd3d2),
	.w3(32'h3bc44d35),
	.w4(32'h3bb1f560),
	.w5(32'hbb194848),
	.w6(32'h3b270bad),
	.w7(32'h3b34660a),
	.w8(32'hbb642f7a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9520d6),
	.w1(32'hbbd4df5b),
	.w2(32'h3b0780ec),
	.w3(32'h3b4a9b57),
	.w4(32'h39bba863),
	.w5(32'hbbd47ab4),
	.w6(32'hba29142e),
	.w7(32'hbbe26dd0),
	.w8(32'hbb5e6574),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc31974),
	.w1(32'hbbb763c0),
	.w2(32'hbb797040),
	.w3(32'hbc00eddd),
	.w4(32'hbb51a4cc),
	.w5(32'hba92eb56),
	.w6(32'hbbd7c3ec),
	.w7(32'hbbbd1c7d),
	.w8(32'h3ad0ff38),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe9cd),
	.w1(32'h3b088226),
	.w2(32'hbb7453ac),
	.w3(32'h3c711521),
	.w4(32'h3c787652),
	.w5(32'hbbf8d66f),
	.w6(32'h3cd1408b),
	.w7(32'h3cb6236e),
	.w8(32'hbbc5aec2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae78222),
	.w1(32'h39d954b5),
	.w2(32'hbb0fe785),
	.w3(32'hbb061ddd),
	.w4(32'h3adab3e0),
	.w5(32'h3b01d9a9),
	.w6(32'hba30d95e),
	.w7(32'h3b0eeb09),
	.w8(32'h3c0c52af),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb5080),
	.w1(32'h3b190ba0),
	.w2(32'h3b3fd7d8),
	.w3(32'h3a2e2953),
	.w4(32'h3bc83542),
	.w5(32'h39d02dba),
	.w6(32'h3b0c036d),
	.w7(32'h3b1a52b0),
	.w8(32'h3a858b2f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39762934),
	.w1(32'hb9713868),
	.w2(32'hb9d27fdb),
	.w3(32'h3b58a581),
	.w4(32'h3b0f576f),
	.w5(32'hbafb3309),
	.w6(32'h3b8229b8),
	.w7(32'h3b94641b),
	.w8(32'h3bab9e8c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc99659),
	.w1(32'hbc4077b5),
	.w2(32'hbc05f196),
	.w3(32'h3bc79cea),
	.w4(32'hbba29ed0),
	.w5(32'hbbe3ab75),
	.w6(32'h3c0f5373),
	.w7(32'hbbea7c0a),
	.w8(32'hbbae943d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85446c),
	.w1(32'hbbb6697d),
	.w2(32'hbb99b811),
	.w3(32'hbbb4f194),
	.w4(32'hbbdbeef7),
	.w5(32'hb9542dbf),
	.w6(32'hbb9b2dee),
	.w7(32'hbbe8ba90),
	.w8(32'h3ad50c62),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a34f0),
	.w1(32'hbc0aed9a),
	.w2(32'hbb58a5b4),
	.w3(32'h3b480166),
	.w4(32'hbb02ee23),
	.w5(32'hba39c652),
	.w6(32'h3b77d804),
	.w7(32'hbb999338),
	.w8(32'hbb9fa529),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16b445),
	.w1(32'hbb041d84),
	.w2(32'hbb70f979),
	.w3(32'hbb36f5ad),
	.w4(32'h3b9f19a3),
	.w5(32'hbb107443),
	.w6(32'h38d7eb24),
	.w7(32'h3bd8f30c),
	.w8(32'hbab6acc7),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa29de6),
	.w1(32'hbaa07326),
	.w2(32'h3b9e9350),
	.w3(32'hbab718f7),
	.w4(32'hba071388),
	.w5(32'h3b3306d0),
	.w6(32'hbab90058),
	.w7(32'h38660ed0),
	.w8(32'h3b68ff85),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa4756),
	.w1(32'h3b8a549d),
	.w2(32'h3acde959),
	.w3(32'h3b9c9b96),
	.w4(32'h3be4bb88),
	.w5(32'hbc2b9e15),
	.w6(32'h39ba1ea4),
	.w7(32'h3b8140e1),
	.w8(32'hbb6e48e1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe43753),
	.w1(32'hbbbec4b9),
	.w2(32'hbb8a58a8),
	.w3(32'hbba4e72c),
	.w4(32'hbc02aee9),
	.w5(32'hb8e2c2ae),
	.w6(32'hbbfa05b0),
	.w7(32'h3b2ad316),
	.w8(32'hbaf3aa3b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae99057),
	.w1(32'hbc0263e3),
	.w2(32'h3abc0b8d),
	.w3(32'h399c5052),
	.w4(32'hbb93ba3d),
	.w5(32'hbb50c932),
	.w6(32'h3b99e3ba),
	.w7(32'hbb6da809),
	.w8(32'hbba70392),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd7468),
	.w1(32'hbbbdb59d),
	.w2(32'hbb4d0da5),
	.w3(32'hbb7f3a6c),
	.w4(32'hbc39054d),
	.w5(32'hbb7ce792),
	.w6(32'hbc11bd1c),
	.w7(32'hbafd9676),
	.w8(32'hbc591cad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf67d59),
	.w1(32'hbbf856cf),
	.w2(32'h396b5ef4),
	.w3(32'hbbfef3db),
	.w4(32'hbb6dd767),
	.w5(32'h3ac0117c),
	.w6(32'hbc8e8ab6),
	.w7(32'hbc63077e),
	.w8(32'h3b875a65),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96806a9),
	.w1(32'hbb3bdb5b),
	.w2(32'h38d92673),
	.w3(32'h3aff106b),
	.w4(32'hbb90fd58),
	.w5(32'hbb2a5d64),
	.w6(32'h3abf413a),
	.w7(32'h3c11c934),
	.w8(32'h3c106753),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c3bb5),
	.w1(32'h3a83f424),
	.w2(32'h3b831784),
	.w3(32'h3b4079ef),
	.w4(32'h3b04373f),
	.w5(32'h3b3d201b),
	.w6(32'h3c55703d),
	.w7(32'h3c4fc563),
	.w8(32'h3bc14bee),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a1217c),
	.w1(32'hb9f4c7e4),
	.w2(32'hbb3e8d92),
	.w3(32'hbb4422d8),
	.w4(32'hbb0a7c49),
	.w5(32'hbba46d78),
	.w6(32'h39fea119),
	.w7(32'hbb9b3120),
	.w8(32'hbb9376b4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f8a92),
	.w1(32'h3bf08d4c),
	.w2(32'h391d3bff),
	.w3(32'hb9ab0d76),
	.w4(32'h3c068fb8),
	.w5(32'h3a5a92dd),
	.w6(32'h3b037b02),
	.w7(32'h3c109df6),
	.w8(32'hbbd60bb4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0e0fe),
	.w1(32'hbb914721),
	.w2(32'h3a0edc19),
	.w3(32'h3b2ee1dc),
	.w4(32'h3bd030cf),
	.w5(32'hbb3f3294),
	.w6(32'hbb213c92),
	.w7(32'h3c17c202),
	.w8(32'h3b16d9d2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87758a),
	.w1(32'hbb05f557),
	.w2(32'h3c1197b3),
	.w3(32'hbb3acb9d),
	.w4(32'h3aa4a906),
	.w5(32'h3b9b9342),
	.w6(32'h3a49f085),
	.w7(32'h3b7e16f8),
	.w8(32'hbaf749df),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba056246),
	.w1(32'hbac3fd98),
	.w2(32'hbaa39e24),
	.w3(32'h3c16027c),
	.w4(32'h3b938dcd),
	.w5(32'h3a01f1fd),
	.w6(32'h3b62356a),
	.w7(32'h3a662d36),
	.w8(32'h39f72ba8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b605e),
	.w1(32'h3b206100),
	.w2(32'h3b2cbed8),
	.w3(32'h3be16e43),
	.w4(32'h3b56097b),
	.w5(32'h3b6e1531),
	.w6(32'h3c4b6182),
	.w7(32'hb991cb3e),
	.w8(32'h3ba32f79),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dfe67),
	.w1(32'hbaeacf2b),
	.w2(32'h3b58d25f),
	.w3(32'h3b95806c),
	.w4(32'hba6bfd32),
	.w5(32'h3b35794f),
	.w6(32'h3b82a7a6),
	.w7(32'hbb06443a),
	.w8(32'h3bb9d8dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a630da9),
	.w1(32'h3a673e84),
	.w2(32'hbb8ef8f0),
	.w3(32'h3b141b66),
	.w4(32'h3b1b7fa6),
	.w5(32'hbc3c80ac),
	.w6(32'h3bbe92b5),
	.w7(32'h3c1d7e34),
	.w8(32'h3c88e272),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94c3d9),
	.w1(32'hbba5740f),
	.w2(32'h3a2c765c),
	.w3(32'hbc227bab),
	.w4(32'hbbe9d317),
	.w5(32'h3a73b4b6),
	.w6(32'h3c4ea5df),
	.w7(32'h3c4df983),
	.w8(32'h3b5ae678),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4523a6),
	.w1(32'h3b3885dc),
	.w2(32'h3b75855f),
	.w3(32'h3b8fad99),
	.w4(32'h3b9a0bbb),
	.w5(32'hbb0c58cf),
	.w6(32'h3bde077f),
	.w7(32'h3ba359bf),
	.w8(32'hbab49955),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5e900),
	.w1(32'hbb8fa665),
	.w2(32'hbc142c30),
	.w3(32'h3b26ba77),
	.w4(32'hbb198f52),
	.w5(32'hbc1f1e9e),
	.w6(32'h3b0a5870),
	.w7(32'hbaf5122c),
	.w8(32'hbc0b2970),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9933068),
	.w1(32'hbbd8fec5),
	.w2(32'hb8a0032e),
	.w3(32'h3b15903d),
	.w4(32'hbb904f1f),
	.w5(32'hbb1984d8),
	.w6(32'h3ba7d2d6),
	.w7(32'hbaba6451),
	.w8(32'hbb859241),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf559eb),
	.w1(32'hbb073fe7),
	.w2(32'hbb48e55a),
	.w3(32'h3af1a5d0),
	.w4(32'hbb5073b3),
	.w5(32'hbb1a37d7),
	.w6(32'hbb2af105),
	.w7(32'hbb84037a),
	.w8(32'hbb6d9aca),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c04f5),
	.w1(32'hbb9e1516),
	.w2(32'h3bb3d105),
	.w3(32'hbb964d0f),
	.w4(32'hbb16aa2b),
	.w5(32'h3af7c282),
	.w6(32'hbb810721),
	.w7(32'hbbb36c86),
	.w8(32'h39e4b77c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fec20),
	.w1(32'hbc01f033),
	.w2(32'hbbac25d0),
	.w3(32'h3b928f29),
	.w4(32'hbb8b6e90),
	.w5(32'hbc0e970c),
	.w6(32'h3bdad9a1),
	.w7(32'hbbd5171b),
	.w8(32'hbc31edb8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a96ca),
	.w1(32'hb9a84408),
	.w2(32'hbc4401b9),
	.w3(32'hbbdac432),
	.w4(32'hbba1093f),
	.w5(32'hbbd624e6),
	.w6(32'hbc1bee80),
	.w7(32'hbc1441a8),
	.w8(32'hbb80bb9e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda7dd3),
	.w1(32'hbc1857aa),
	.w2(32'h3bfd8c0a),
	.w3(32'h3bd39f96),
	.w4(32'hba8e46ac),
	.w5(32'h3ba5ca9d),
	.w6(32'h3c0c1b73),
	.w7(32'hbb64e40c),
	.w8(32'h3c3d7c0d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9ac5f),
	.w1(32'h3bca93aa),
	.w2(32'hbba50d84),
	.w3(32'h3bd8e57f),
	.w4(32'h3c55a6ee),
	.w5(32'hbb50edac),
	.w6(32'h3c581a0a),
	.w7(32'h3caf1f26),
	.w8(32'hbb0530f0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a5418),
	.w1(32'hbb9a1ba4),
	.w2(32'hbbd13d0c),
	.w3(32'h398f0807),
	.w4(32'hbab21b06),
	.w5(32'hbc0b58f3),
	.w6(32'h3a601da8),
	.w7(32'hb9c5c5c4),
	.w8(32'hbb07447b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba81b52),
	.w1(32'hbb9a95fc),
	.w2(32'h3b2e7dbc),
	.w3(32'hbba34f33),
	.w4(32'hbb815618),
	.w5(32'h3ba4af2f),
	.w6(32'h3ac2fe05),
	.w7(32'h3aacb859),
	.w8(32'hbb71b87e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccf617),
	.w1(32'hbbb5b958),
	.w2(32'h3b905869),
	.w3(32'h398aa8e6),
	.w4(32'hbae32a1a),
	.w5(32'h3ae87912),
	.w6(32'hbc0db287),
	.w7(32'hba4ee021),
	.w8(32'hbba9842c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af859),
	.w1(32'hbbbf0b84),
	.w2(32'hbad60933),
	.w3(32'h393fd488),
	.w4(32'hbb50bbe9),
	.w5(32'h3989b70b),
	.w6(32'hbbd74213),
	.w7(32'h3b6b1915),
	.w8(32'h3ad4e48b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89790cb),
	.w1(32'h3c0491a8),
	.w2(32'hba050701),
	.w3(32'h3b4751d5),
	.w4(32'h3bd9a4b2),
	.w5(32'hba1a480e),
	.w6(32'h3b7c97a5),
	.w7(32'h3b2cd562),
	.w8(32'h3a45736c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44fcb4),
	.w1(32'hb9be695a),
	.w2(32'hbb2d8b85),
	.w3(32'h3d02db6d),
	.w4(32'h3bd526fb),
	.w5(32'hbb163359),
	.w6(32'h3cac0252),
	.w7(32'hba72bf42),
	.w8(32'hbbd062d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea8bc2),
	.w1(32'hbbfde090),
	.w2(32'hba9e7dac),
	.w3(32'hbbdf51bb),
	.w4(32'hbbf5ebfc),
	.w5(32'hbb853161),
	.w6(32'hbbf1319b),
	.w7(32'hbbcb1c1d),
	.w8(32'hbad5d535),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe47e09),
	.w1(32'hbb3fd4d1),
	.w2(32'h3b0cabae),
	.w3(32'hbaed6d5b),
	.w4(32'hba1e3b75),
	.w5(32'h3b708d25),
	.w6(32'hba9112c1),
	.w7(32'hb8b7c57f),
	.w8(32'hbb81333a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74a7c),
	.w1(32'h3baca5be),
	.w2(32'hbbe852fd),
	.w3(32'h3afcd3f6),
	.w4(32'h3c0c55c6),
	.w5(32'hbba76b05),
	.w6(32'hbbeacbb2),
	.w7(32'h3c158256),
	.w8(32'hbba083b4),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a740a74),
	.w1(32'h3b292ffa),
	.w2(32'hbbc1c5e0),
	.w3(32'h3b505202),
	.w4(32'h3bcf10e9),
	.w5(32'hbaeab812),
	.w6(32'h3b8537af),
	.w7(32'h3c22e202),
	.w8(32'hbb64520b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5af63a),
	.w1(32'hbb06db1b),
	.w2(32'h3b91a85d),
	.w3(32'hb9ea6507),
	.w4(32'hbbb6e05a),
	.w5(32'hbaa85356),
	.w6(32'h3ae12c02),
	.w7(32'hbbc399fa),
	.w8(32'h3c09363b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb931ba6),
	.w1(32'h3b0aad8a),
	.w2(32'hba8cedbc),
	.w3(32'h386130ec),
	.w4(32'h3b7e6e5d),
	.w5(32'hbb019633),
	.w6(32'h3bc08751),
	.w7(32'h3bc99a5f),
	.w8(32'hbb0c5945),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0add9c),
	.w1(32'hba918983),
	.w2(32'h3961534f),
	.w3(32'hbb1b17d6),
	.w4(32'hba789917),
	.w5(32'h3b148d2f),
	.w6(32'h3a566f1f),
	.w7(32'h3b0334c9),
	.w8(32'h3b70fcf7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0be9e0),
	.w1(32'h3b827056),
	.w2(32'hb9fb7cdf),
	.w3(32'h3b9443d7),
	.w4(32'h3bde7688),
	.w5(32'hbbcb2a3e),
	.w6(32'h3bf605cd),
	.w7(32'h3c144ae5),
	.w8(32'hbbeb03fb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb046515),
	.w1(32'hbb272014),
	.w2(32'hbb902432),
	.w3(32'h3aad6893),
	.w4(32'hbbadbee0),
	.w5(32'hbba10514),
	.w6(32'hbc27a898),
	.w7(32'hbb443493),
	.w8(32'hbc354582),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd5a0),
	.w1(32'h3af53e21),
	.w2(32'hbabdd260),
	.w3(32'hbabf5a5f),
	.w4(32'hb8c69028),
	.w5(32'hbb64199d),
	.w6(32'hbb9ff206),
	.w7(32'h3a38316f),
	.w8(32'h3b98fdb6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7d2c1),
	.w1(32'hbb288baa),
	.w2(32'h3b7fc0e4),
	.w3(32'h393311a1),
	.w4(32'h3a69f1a7),
	.w5(32'h3a5b0d4c),
	.w6(32'h3ae1ead2),
	.w7(32'h3b94b11d),
	.w8(32'hbb8f0755),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08a812),
	.w1(32'hbb976d30),
	.w2(32'hbace77ac),
	.w3(32'h3a9a1203),
	.w4(32'h3ae7a018),
	.w5(32'h3b99a835),
	.w6(32'hbac3e4a2),
	.w7(32'hbaef79e5),
	.w8(32'h3bce9fda),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7bfd2),
	.w1(32'h3b993f87),
	.w2(32'h3ad72341),
	.w3(32'h3c79f930),
	.w4(32'h3c89462e),
	.w5(32'h3b0deec9),
	.w6(32'h3c9c5c1c),
	.w7(32'h3c9a68d6),
	.w8(32'h3b6d82b1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34b385),
	.w1(32'hb9915fda),
	.w2(32'h3b6d2bda),
	.w3(32'h3b9d603b),
	.w4(32'h3b8309c6),
	.w5(32'hbb669ce3),
	.w6(32'h3bf2a232),
	.w7(32'h3bef0286),
	.w8(32'hbabfb879),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d47771),
	.w1(32'hbbbf4b7c),
	.w2(32'h3ba86aa2),
	.w3(32'hb7ced7ba),
	.w4(32'hbbae72e5),
	.w5(32'h3a97aded),
	.w6(32'h3a389dc2),
	.w7(32'hbba103e4),
	.w8(32'hbb806886),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc7d0b),
	.w1(32'h3bb34b67),
	.w2(32'h3bafacc7),
	.w3(32'h3b3a2bfc),
	.w4(32'h3bad8184),
	.w5(32'h3abf4578),
	.w6(32'hbbd4c862),
	.w7(32'hbbb30d38),
	.w8(32'h3bedbc2c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00ba6a),
	.w1(32'h3a5a9adb),
	.w2(32'hbb6d7a3e),
	.w3(32'h3b0081ba),
	.w4(32'h3ba0a189),
	.w5(32'hbb63666f),
	.w6(32'h3c3b370e),
	.w7(32'h3c513065),
	.w8(32'hbb556cf4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1b7d8),
	.w1(32'hbbeee108),
	.w2(32'h3a1cf4ae),
	.w3(32'hbc02ec48),
	.w4(32'hbc0bceac),
	.w5(32'hbb0c67a4),
	.w6(32'hbbb6902f),
	.w7(32'hbbfe3412),
	.w8(32'hbb2f060f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc98ac),
	.w1(32'hba087b83),
	.w2(32'h3b172c70),
	.w3(32'hbbab8228),
	.w4(32'hb8a3f1f3),
	.w5(32'h3b3b4e85),
	.w6(32'hbc2f6a32),
	.w7(32'h3a3d9589),
	.w8(32'hbbc8ca75),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045770),
	.w1(32'h39feb41e),
	.w2(32'hbc27d5c9),
	.w3(32'hbb093b26),
	.w4(32'h3c02c940),
	.w5(32'h3ba667d7),
	.w6(32'hbbe6719d),
	.w7(32'h3bb851d7),
	.w8(32'h3b4c62bc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f4600),
	.w1(32'hbbb473ba),
	.w2(32'h380b39e7),
	.w3(32'h3bf72057),
	.w4(32'h3c7e3470),
	.w5(32'h3c383560),
	.w6(32'hbaa5c555),
	.w7(32'h39e0e91f),
	.w8(32'h3c2af772),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82eff0),
	.w1(32'hbbce0f17),
	.w2(32'hbb845707),
	.w3(32'h3bdecf4e),
	.w4(32'h3c2fe77b),
	.w5(32'h3ac2c9f7),
	.w6(32'h3c45ba7f),
	.w7(32'h3c465426),
	.w8(32'h3ad7523c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460c53),
	.w1(32'h3ab44732),
	.w2(32'hbbbf3146),
	.w3(32'hbb376c76),
	.w4(32'h3b68a2cc),
	.w5(32'h3b63950b),
	.w6(32'hbaaf9815),
	.w7(32'h3bc8d5fe),
	.w8(32'h3bc304f2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9699ff),
	.w1(32'h3b27368c),
	.w2(32'hba9d1cfe),
	.w3(32'h3b31b40f),
	.w4(32'h3bfc5d31),
	.w5(32'h3ab31327),
	.w6(32'h3b894c8e),
	.w7(32'h3c2d6272),
	.w8(32'h3b00e6e4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f493),
	.w1(32'hbbb5b124),
	.w2(32'hbbcda63d),
	.w3(32'hbad258d6),
	.w4(32'hb9ea44a4),
	.w5(32'hbc26df4d),
	.w6(32'h3a838fa4),
	.w7(32'hb9b3526b),
	.w8(32'hbc2da5c3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3286),
	.w1(32'hbaa8660d),
	.w2(32'hbad41130),
	.w3(32'hbc2bad77),
	.w4(32'hbb9cc5f3),
	.w5(32'hbb87ed36),
	.w6(32'hbbb40e90),
	.w7(32'hba420f4a),
	.w8(32'hbb0bce62),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108734),
	.w1(32'hba187498),
	.w2(32'hbc083591),
	.w3(32'h3ad8927e),
	.w4(32'hbb261732),
	.w5(32'h3b394d2d),
	.w6(32'h3b25df5d),
	.w7(32'hbb3b9cc8),
	.w8(32'hb9a46593),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59c81f),
	.w1(32'h3b9d530e),
	.w2(32'hbc1c14dc),
	.w3(32'h3b310358),
	.w4(32'h3c2f9d40),
	.w5(32'hbbc554ca),
	.w6(32'hbb4ed6e8),
	.w7(32'h3b674c06),
	.w8(32'hb9f067d7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b34e11),
	.w1(32'hbc4700fb),
	.w2(32'hbb39766b),
	.w3(32'h3ba807f4),
	.w4(32'hbc5292f8),
	.w5(32'hb72da14a),
	.w6(32'h3c130549),
	.w7(32'hbc786d59),
	.w8(32'hba027c4f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb966594d),
	.w1(32'h3b5b7f50),
	.w2(32'hbbe6bbef),
	.w3(32'h3b8a358c),
	.w4(32'h3c16a048),
	.w5(32'hbb962db2),
	.w6(32'h3a550017),
	.w7(32'h3b369871),
	.w8(32'hbba174c2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef381c),
	.w1(32'hbbe565d6),
	.w2(32'hba448b41),
	.w3(32'hbba93305),
	.w4(32'hbbc8414b),
	.w5(32'hbaeb1bfb),
	.w6(32'hbbe306f1),
	.w7(32'hbbf3686c),
	.w8(32'h3a639c34),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78167b),
	.w1(32'h3b8efcb4),
	.w2(32'hb90b29c5),
	.w3(32'hbb875355),
	.w4(32'h3bf05424),
	.w5(32'hba983fd0),
	.w6(32'hbb02eed5),
	.w7(32'h3c2aebe1),
	.w8(32'hbb53c9ec),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f49a),
	.w1(32'h3c0c09dc),
	.w2(32'hbb85c469),
	.w3(32'hbae9e5fe),
	.w4(32'h3b459c58),
	.w5(32'hbb257f0b),
	.w6(32'hbb4e0d78),
	.w7(32'h3c1e6a24),
	.w8(32'h3bdcbfdb),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a7df3),
	.w1(32'h3b1181e9),
	.w2(32'h3acc2f75),
	.w3(32'h3b0ce91d),
	.w4(32'h3a94b5e4),
	.w5(32'h3b09ec55),
	.w6(32'h3a8974fb),
	.w7(32'h3ab16837),
	.w8(32'h3b0a76a3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5b6e4),
	.w1(32'h3872da0b),
	.w2(32'hbac1062a),
	.w3(32'h3a6d4c1f),
	.w4(32'hbacbd408),
	.w5(32'hbad557b3),
	.w6(32'h3b16a74a),
	.w7(32'h3b3b77c1),
	.w8(32'hbb6b9ae6),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74bc9e),
	.w1(32'hbb53a8b8),
	.w2(32'hbb024b76),
	.w3(32'h3a24a71c),
	.w4(32'h3a236132),
	.w5(32'hb9ae99dd),
	.w6(32'hbad981fc),
	.w7(32'hbb369bb5),
	.w8(32'hbb1d45c9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5ebee),
	.w1(32'hbb8c0d62),
	.w2(32'hbb155697),
	.w3(32'h3b0e7919),
	.w4(32'h3bb33154),
	.w5(32'h3a42c5ff),
	.w6(32'hbaae750f),
	.w7(32'hb9dac023),
	.w8(32'hbb72333b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f7b71),
	.w1(32'hbb91b737),
	.w2(32'h3b87d38c),
	.w3(32'h3b933410),
	.w4(32'h3b856f55),
	.w5(32'hba84cd77),
	.w6(32'h3aa24532),
	.w7(32'h3a8e7f6c),
	.w8(32'h3bce0ca8),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb805cf1),
	.w1(32'hba6b9b1a),
	.w2(32'hbc1cb873),
	.w3(32'hbb0351f2),
	.w4(32'h3b90cbea),
	.w5(32'h3c11e0e8),
	.w6(32'h3b1239d1),
	.w7(32'h3c13fe99),
	.w8(32'hbbbb1ebd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21f048),
	.w1(32'hbb541c9a),
	.w2(32'hbb0cc6c9),
	.w3(32'h3b1148ce),
	.w4(32'h3ba26c5e),
	.w5(32'hbb864601),
	.w6(32'hbbcb3969),
	.w7(32'h3bc8afb0),
	.w8(32'h3a254b07),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d50c3),
	.w1(32'hbb11d22d),
	.w2(32'hbb7b6b27),
	.w3(32'h3b8410ec),
	.w4(32'hbab50077),
	.w5(32'hba82129c),
	.w6(32'h3bc07470),
	.w7(32'hbb89af75),
	.w8(32'h381dc713),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb334c43),
	.w1(32'hbaa3ac22),
	.w2(32'hbb9401ea),
	.w3(32'hba24e8b1),
	.w4(32'h3a693402),
	.w5(32'hbb602726),
	.w6(32'h3a40cb23),
	.w7(32'h3b8d76a2),
	.w8(32'hbb45d616),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb5a3),
	.w1(32'hbb0ad742),
	.w2(32'hbb4b3103),
	.w3(32'hbb0b24d2),
	.w4(32'hba93e4d6),
	.w5(32'hbb5b1e4f),
	.w6(32'hbaf3ffbe),
	.w7(32'hbb01c37b),
	.w8(32'hbbde92d6),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81a76a),
	.w1(32'h39a6e743),
	.w2(32'h3b04acf5),
	.w3(32'hbb87f747),
	.w4(32'h3ba8730b),
	.w5(32'h3b3ebafb),
	.w6(32'hbbd886bb),
	.w7(32'h3b697707),
	.w8(32'hba733a4c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d7fd),
	.w1(32'h3af143da),
	.w2(32'h3b1c12c6),
	.w3(32'h3be21d1a),
	.w4(32'h3b4f8644),
	.w5(32'hbbc7e31f),
	.w6(32'h3b486ea0),
	.w7(32'hbafb6bc7),
	.w8(32'hbada4dcc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ab951),
	.w1(32'hbb19dfc7),
	.w2(32'hbbe229a8),
	.w3(32'hbc0d90dd),
	.w4(32'hbc0bfff9),
	.w5(32'hbba21f5a),
	.w6(32'h3a87506e),
	.w7(32'h3a1f5429),
	.w8(32'hba86e1c1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c468f35),
	.w1(32'h3b5bf04b),
	.w2(32'hbba3532b),
	.w3(32'h3c811c74),
	.w4(32'h3b06bac7),
	.w5(32'hbbaa7639),
	.w6(32'h3c72648b),
	.w7(32'h3baf0660),
	.w8(32'hbb5dd9ba),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a6a78),
	.w1(32'hbbc64e39),
	.w2(32'hbbbdf126),
	.w3(32'h3b97b4eb),
	.w4(32'hbbc48c99),
	.w5(32'h3b650f62),
	.w6(32'h3b889c77),
	.w7(32'hbaec3ed8),
	.w8(32'h3b4e1a37),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae55a5f),
	.w1(32'hba6e774d),
	.w2(32'hbbd2f996),
	.w3(32'hbaea12ed),
	.w4(32'h3c2ea6d3),
	.w5(32'hbbf999d0),
	.w6(32'hba9c935c),
	.w7(32'hba837770),
	.w8(32'hba16cff1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bb736),
	.w1(32'h3c5ad0b1),
	.w2(32'h3b10ac76),
	.w3(32'hbaf38b80),
	.w4(32'h3bc3eb1a),
	.w5(32'h3bf98988),
	.w6(32'h3ae546cc),
	.w7(32'h3c2a2f6f),
	.w8(32'h3b8f6306),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd66aa),
	.w1(32'h3b7d49ef),
	.w2(32'hbb1cc21e),
	.w3(32'h3be6d574),
	.w4(32'h3c6b2fe7),
	.w5(32'hba64aea5),
	.w6(32'h3bf8a13c),
	.w7(32'h3c225be2),
	.w8(32'h3a182071),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc096ea8),
	.w1(32'hbb744dae),
	.w2(32'h3badbb30),
	.w3(32'h3aa39dcf),
	.w4(32'hbbfd6918),
	.w5(32'hbb46cef4),
	.w6(32'hbbbbd928),
	.w7(32'hbc100fb3),
	.w8(32'hbbea4142),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99647c),
	.w1(32'hbb022860),
	.w2(32'hbb3a59ea),
	.w3(32'hb98f2bbe),
	.w4(32'h3b8b179d),
	.w5(32'h3ad2b4c4),
	.w6(32'hbbafbb82),
	.w7(32'hb95e409c),
	.w8(32'h3b13a309),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2113fb),
	.w1(32'hbc27e48b),
	.w2(32'hbb278ce8),
	.w3(32'h3c3c6d87),
	.w4(32'hbc0e2fef),
	.w5(32'hbae86f20),
	.w6(32'h3c9a6fe9),
	.w7(32'hbc300bdd),
	.w8(32'hbab042fb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec299),
	.w1(32'hbb8e301b),
	.w2(32'hbb0ecfda),
	.w3(32'h3b777f3a),
	.w4(32'h39dcae8f),
	.w5(32'h3a0a9dd2),
	.w6(32'h3b9f3927),
	.w7(32'h3a113bf0),
	.w8(32'hbbad0aaa),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3aaac),
	.w1(32'hbb9e9167),
	.w2(32'hbbd07389),
	.w3(32'h3b9c6911),
	.w4(32'h3ae4c933),
	.w5(32'h3ac9ce39),
	.w6(32'hbab23d99),
	.w7(32'hbb52a2cd),
	.w8(32'h3b12dc60),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3a3b7),
	.w1(32'h3917d5b5),
	.w2(32'h3b5aac23),
	.w3(32'h3bbcc3e7),
	.w4(32'h3a94b641),
	.w5(32'h3ac4a717),
	.w6(32'h3b018512),
	.w7(32'hba308f92),
	.w8(32'h3b878ed7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad14623),
	.w1(32'hbb28748e),
	.w2(32'hbb0d3d3c),
	.w3(32'h3be90567),
	.w4(32'h3b2aaa8a),
	.w5(32'hbb4d6b78),
	.w6(32'h3bb7c8ee),
	.w7(32'h3b3cc4ae),
	.w8(32'hbb156184),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba297a5),
	.w1(32'hbb7d65bd),
	.w2(32'hbb0ff23e),
	.w3(32'hbb38d5ed),
	.w4(32'hbb3947d3),
	.w5(32'hbc0b53a9),
	.w6(32'hbb2075b4),
	.w7(32'hbb35d932),
	.w8(32'hbb45b3e0),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc11658),
	.w1(32'hbbbdddff),
	.w2(32'hba1bb959),
	.w3(32'hbbd7656a),
	.w4(32'hbb47d8a2),
	.w5(32'h3a9f2c79),
	.w6(32'h391d9f44),
	.w7(32'hbb7d7bc5),
	.w8(32'h3ab51ca4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acce297),
	.w1(32'h3a2fa110),
	.w2(32'hbbf2aaa0),
	.w3(32'h3b876daa),
	.w4(32'h3b76fe64),
	.w5(32'hbc4dfe2d),
	.w6(32'h3b8b71e8),
	.w7(32'h3b7ce058),
	.w8(32'hbc819998),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc223c1c),
	.w1(32'hbc354c1e),
	.w2(32'h3b887aa6),
	.w3(32'hbb1fe191),
	.w4(32'hbc8ee90e),
	.w5(32'h3c13732a),
	.w6(32'hbbdf7eec),
	.w7(32'hbc679884),
	.w8(32'h3c097943),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f6b38),
	.w1(32'hbb3306a7),
	.w2(32'hbacab595),
	.w3(32'h3bca9d2f),
	.w4(32'h3c3592c3),
	.w5(32'hba196971),
	.w6(32'h3af3e1d1),
	.w7(32'h3bdf8e37),
	.w8(32'hba09cfa4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e2c74),
	.w1(32'hbbf2a340),
	.w2(32'hbb6d223d),
	.w3(32'hb9f2f675),
	.w4(32'hbba977a4),
	.w5(32'hbb9c7823),
	.w6(32'hb936a1a5),
	.w7(32'hbc0ee971),
	.w8(32'hbb86a267),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79fb3),
	.w1(32'hbb9333ae),
	.w2(32'hb9344d5a),
	.w3(32'hbb8ecad0),
	.w4(32'hbb81b16b),
	.w5(32'h39ed7675),
	.w6(32'hbb6eddea),
	.w7(32'hbb72a54c),
	.w8(32'h3a39b9e4),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241b86),
	.w1(32'h39b99541),
	.w2(32'hbbaaa7a7),
	.w3(32'h3b94635f),
	.w4(32'h3b0016dc),
	.w5(32'hbbbc91ef),
	.w6(32'h3b4cb64b),
	.w7(32'h3aa75b26),
	.w8(32'hbbbeb441),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb303a84),
	.w1(32'hbba2be73),
	.w2(32'hbaff9216),
	.w3(32'h3a89eb72),
	.w4(32'hbb112769),
	.w5(32'h3a951c5c),
	.w6(32'hb931f415),
	.w7(32'hbb92bbff),
	.w8(32'h3b240fd2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07036a),
	.w1(32'hba6b17ee),
	.w2(32'hbb5d8305),
	.w3(32'h3c0067db),
	.w4(32'h3bc26224),
	.w5(32'hba764dfa),
	.w6(32'h3ab519ff),
	.w7(32'hbb864474),
	.w8(32'hbb86dedd),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5602ba),
	.w1(32'hbb45800d),
	.w2(32'hbaadaadf),
	.w3(32'hbb2eecf1),
	.w4(32'h39d7864f),
	.w5(32'hbb23b286),
	.w6(32'hbb6e3d0e),
	.w7(32'hba54eeb6),
	.w8(32'hba3daa65),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc324550),
	.w1(32'hbc2acfb9),
	.w2(32'h3b04bb48),
	.w3(32'hbbc9c875),
	.w4(32'hbb8ff3e3),
	.w5(32'h3bf1daa4),
	.w6(32'hbc12d3e7),
	.w7(32'hbc554c84),
	.w8(32'h3c0ef412),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a190652),
	.w1(32'hbb22b0ac),
	.w2(32'hbab7af7c),
	.w3(32'h3c094d85),
	.w4(32'h3b68954d),
	.w5(32'hb8a8a2a7),
	.w6(32'h3c21b829),
	.w7(32'h3b50f694),
	.w8(32'hbaa9a486),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a754434),
	.w1(32'h3a57a4d4),
	.w2(32'hbc0a314c),
	.w3(32'h3b5ec79e),
	.w4(32'h3b6d47c5),
	.w5(32'hbc4b26a2),
	.w6(32'h3b177769),
	.w7(32'h3b19e8ce),
	.w8(32'hbc115c24),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb977fcd),
	.w1(32'hbc2d074f),
	.w2(32'hbbcdf944),
	.w3(32'hba615183),
	.w4(32'hbc1ccb0f),
	.w5(32'hbb4235b4),
	.w6(32'hbb2fe3e7),
	.w7(32'hbc0a1ec1),
	.w8(32'hbc3af6b4),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b9712),
	.w1(32'h3b5ffc81),
	.w2(32'h3ba1fc4a),
	.w3(32'hbb5ce7c0),
	.w4(32'h3b17b44a),
	.w5(32'hb9f002bb),
	.w6(32'hbc0157d7),
	.w7(32'hbbbcff28),
	.w8(32'hbb106081),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da0bb),
	.w1(32'hbb94c51b),
	.w2(32'h3aea543d),
	.w3(32'hbb1340e7),
	.w4(32'hbb8f1338),
	.w5(32'h3b2e1cb6),
	.w6(32'hbc0272bd),
	.w7(32'hbb84f942),
	.w8(32'h3ab5d4aa),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864986),
	.w1(32'h3a774445),
	.w2(32'hbb14de81),
	.w3(32'h3a9d3dc1),
	.w4(32'h3a6f66ae),
	.w5(32'hbb51ddce),
	.w6(32'h394a6652),
	.w7(32'h3a91da90),
	.w8(32'hbbb03be1),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32dbb0),
	.w1(32'h3b02c29d),
	.w2(32'h37d0f2bc),
	.w3(32'h3c4855cd),
	.w4(32'h3b6ce7a1),
	.w5(32'hbb056dee),
	.w6(32'h3b82d4e0),
	.w7(32'hbaeda11c),
	.w8(32'hbb54de3a),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0c85a),
	.w1(32'hbab45f85),
	.w2(32'hbb2dee82),
	.w3(32'hbb12b238),
	.w4(32'hbabdaeb3),
	.w5(32'hbb0853fb),
	.w6(32'hbb5b8c2b),
	.w7(32'hbbe1243f),
	.w8(32'hbbc35594),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba292e45),
	.w1(32'hbb1b355c),
	.w2(32'hbc0f5911),
	.w3(32'h3ad00d25),
	.w4(32'h3b03484b),
	.w5(32'hbc64ebfb),
	.w6(32'hbb0511e6),
	.w7(32'hba084f37),
	.w8(32'hbc38def9),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90ab2),
	.w1(32'h39a4842b),
	.w2(32'hbc28f68c),
	.w3(32'hbc7c3d01),
	.w4(32'h3ca6cfc8),
	.w5(32'hbc9f09e9),
	.w6(32'hbc92485a),
	.w7(32'h3c7b29b3),
	.w8(32'hbca29744),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dc714),
	.w1(32'h3bc6f1b0),
	.w2(32'hbb765aa4),
	.w3(32'hbb92460a),
	.w4(32'h3c68ac28),
	.w5(32'hbb844864),
	.w6(32'hbc953b09),
	.w7(32'h3cd9740a),
	.w8(32'hbae4b0d7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f154ee),
	.w1(32'hbbb8ebb9),
	.w2(32'hbb47874b),
	.w3(32'h3a836138),
	.w4(32'hbb1d4740),
	.w5(32'hbc1d8d52),
	.w6(32'h3a012bd7),
	.w7(32'hbb487f41),
	.w8(32'hbc31f8ef),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb166502),
	.w1(32'h3c729440),
	.w2(32'hbaa3f7bd),
	.w3(32'hbc558345),
	.w4(32'h3cb52609),
	.w5(32'hba5e153f),
	.w6(32'hbc5897b6),
	.w7(32'hbad7b238),
	.w8(32'h3aabd782),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4850),
	.w1(32'h3abff6b1),
	.w2(32'h3bbf04c5),
	.w3(32'hbb32c596),
	.w4(32'hbb3ecc85),
	.w5(32'hbb77e34e),
	.w6(32'hbb0659f7),
	.w7(32'hbb1225ed),
	.w8(32'hbbce4b07),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca15da),
	.w1(32'h3c47f5ac),
	.w2(32'hbabc76ba),
	.w3(32'h3b049b5e),
	.w4(32'h3c85bf0c),
	.w5(32'hbb2198b6),
	.w6(32'hbbb7e85b),
	.w7(32'h3c84a78b),
	.w8(32'hbb6ec3fd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d941),
	.w1(32'hba30121c),
	.w2(32'hbc4b4878),
	.w3(32'h3ba9bc5e),
	.w4(32'h3abc3764),
	.w5(32'hbc2a3a01),
	.w6(32'h3b12024c),
	.w7(32'h3b11bfa0),
	.w8(32'hbafb944c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ac8ee),
	.w1(32'h3b9b8a49),
	.w2(32'h3b628eac),
	.w3(32'hbc650da1),
	.w4(32'h3ab41a79),
	.w5(32'hb9d20280),
	.w6(32'hbc1c5eb2),
	.w7(32'h3bd2df07),
	.w8(32'hbc46383f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c136432),
	.w1(32'h3c22470b),
	.w2(32'h3ad7b004),
	.w3(32'h3bdbb2fd),
	.w4(32'h3b902bfb),
	.w5(32'h3b37f7f2),
	.w6(32'hbb689741),
	.w7(32'hbaf7df38),
	.w8(32'hbb3e3f2f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aec27),
	.w1(32'h3b94dc39),
	.w2(32'hb93de99d),
	.w3(32'h3bdef249),
	.w4(32'h3c2c2adb),
	.w5(32'hba4f46b8),
	.w6(32'h3b937d76),
	.w7(32'h3c82b1e6),
	.w8(32'hbb814dc0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0589ac),
	.w1(32'h3c766e0f),
	.w2(32'hbc37e82a),
	.w3(32'hbb62212d),
	.w4(32'h3c129eae),
	.w5(32'hbc64966b),
	.w6(32'hbbf26055),
	.w7(32'h3c23a7fd),
	.w8(32'hbb89470a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4a17),
	.w1(32'h3baeed24),
	.w2(32'h3ac3402c),
	.w3(32'hbbd26ff0),
	.w4(32'h3c716403),
	.w5(32'h3b0afd28),
	.w6(32'hbc0e54b6),
	.w7(32'h3c28982a),
	.w8(32'h3b70be82),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f1deb),
	.w1(32'h3b070028),
	.w2(32'hbbb66f9a),
	.w3(32'hba997ab6),
	.w4(32'hbacf2775),
	.w5(32'h3aa65a9a),
	.w6(32'h393767e4),
	.w7(32'h3952ea0b),
	.w8(32'h3b36fb81),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00148b),
	.w1(32'hbc5fc4c9),
	.w2(32'h3979834f),
	.w3(32'h3c0f1944),
	.w4(32'hbcc5601c),
	.w5(32'h3ba93b07),
	.w6(32'h3c4655f6),
	.w7(32'hbc35c291),
	.w8(32'h3b9834ce),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e8184),
	.w1(32'h39af43a1),
	.w2(32'hbb8de5a3),
	.w3(32'h3b9ac687),
	.w4(32'h3a3fdba2),
	.w5(32'hbb9340fe),
	.w6(32'h3ba6d69e),
	.w7(32'h3bdb4fc8),
	.w8(32'hbc0ef48c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be342),
	.w1(32'hbbd413ab),
	.w2(32'h3c460c08),
	.w3(32'hbb422c69),
	.w4(32'h3bd70552),
	.w5(32'h3c52db13),
	.w6(32'hbb63afc1),
	.w7(32'h3c064f5b),
	.w8(32'h3c4684ff),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ca1a0),
	.w1(32'hbb1211f0),
	.w2(32'hb930a373),
	.w3(32'hbb09d90e),
	.w4(32'hbb5f3c11),
	.w5(32'hb9893a8c),
	.w6(32'h3c22f421),
	.w7(32'hbad5cd72),
	.w8(32'h396ba2bb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20e8c4),
	.w1(32'h3a465e8a),
	.w2(32'h3b320792),
	.w3(32'hbb41102e),
	.w4(32'hbb455a6c),
	.w5(32'hbb4dd5a4),
	.w6(32'h3a28461a),
	.w7(32'hbac548dc),
	.w8(32'h3b3a5cef),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee9551),
	.w1(32'h3be9f42d),
	.w2(32'hbabe0edb),
	.w3(32'h3b429982),
	.w4(32'h3b0e1a3a),
	.w5(32'hbb67680e),
	.w6(32'h3b70ee53),
	.w7(32'hbb7fb015),
	.w8(32'hbb16e910),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54a7e9),
	.w1(32'h3b6449fc),
	.w2(32'hbc15d7c7),
	.w3(32'hbc3fda0a),
	.w4(32'h3c393e9d),
	.w5(32'hbc1e1aa1),
	.w6(32'hbc11c8a3),
	.w7(32'h3b05d7e8),
	.w8(32'hbb617e15),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69e483),
	.w1(32'h3bc465b7),
	.w2(32'h39978d17),
	.w3(32'hbc0a37b1),
	.w4(32'h3ba3b9c2),
	.w5(32'hbb46c4ff),
	.w6(32'hbb0afa13),
	.w7(32'h3b0b7e25),
	.w8(32'h39f265b3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ca862),
	.w1(32'h3c595f01),
	.w2(32'hbc0d768f),
	.w3(32'hbbd013f2),
	.w4(32'h3c67f109),
	.w5(32'hbc059830),
	.w6(32'hbb8eb315),
	.w7(32'hbb498dea),
	.w8(32'hbb8f4a3b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f270),
	.w1(32'h3bbeb256),
	.w2(32'h3b168398),
	.w3(32'hbbb08d26),
	.w4(32'h3c8674b0),
	.w5(32'h3b82d996),
	.w6(32'hb9676ed1),
	.w7(32'h3c96d3ab),
	.w8(32'hbb059da3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c8f94),
	.w1(32'h3bb8526f),
	.w2(32'hbb0c0f28),
	.w3(32'h3c3d9123),
	.w4(32'h3ba170ff),
	.w5(32'hbc41d359),
	.w6(32'h3a1999f9),
	.w7(32'h3b8e3189),
	.w8(32'hbc27767e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eec58),
	.w1(32'h3bdf4f0e),
	.w2(32'hbc649662),
	.w3(32'hbc45e30e),
	.w4(32'h3c36a63b),
	.w5(32'hbc5dd3df),
	.w6(32'hbbf01f5d),
	.w7(32'h3b8d8a8f),
	.w8(32'hbb84df23),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbf49),
	.w1(32'hbbec9940),
	.w2(32'hba994a76),
	.w3(32'h3c7ecb77),
	.w4(32'h3bbf559f),
	.w5(32'h3b051caf),
	.w6(32'h3c418d9d),
	.w7(32'h3c4b969a),
	.w8(32'h3af98ed1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f9dfa),
	.w1(32'hbbbd4893),
	.w2(32'hba7cc5cc),
	.w3(32'hbabcbd08),
	.w4(32'h3ac80dfe),
	.w5(32'hb9ba8fc2),
	.w6(32'hbbc56bd1),
	.w7(32'hbc035362),
	.w8(32'h3ba5e9ad),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe0f50),
	.w1(32'hbc260f20),
	.w2(32'hbbc2628c),
	.w3(32'hbb3d1cc8),
	.w4(32'hbbd2da95),
	.w5(32'hbbb984c6),
	.w6(32'h3c29e644),
	.w7(32'h3c0169b0),
	.w8(32'hbbdd2589),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2d451),
	.w1(32'h3bb4bcd5),
	.w2(32'hba8ad691),
	.w3(32'hbae7eedd),
	.w4(32'h3c1dbb38),
	.w5(32'h3ae24990),
	.w6(32'hbbd2aaf5),
	.w7(32'hba93df92),
	.w8(32'h3b49362b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b824905),
	.w1(32'hbb7a344d),
	.w2(32'hbbeef104),
	.w3(32'hbb52286a),
	.w4(32'hbc338143),
	.w5(32'hbbad4525),
	.w6(32'h3acd32e1),
	.w7(32'hbbccfee3),
	.w8(32'hba8f9ff0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6983cb),
	.w1(32'hb91411d8),
	.w2(32'hbae038a3),
	.w3(32'h3a932eb5),
	.w4(32'h3c110194),
	.w5(32'hb98cc763),
	.w6(32'h3b3b2f16),
	.w7(32'h3c80ca65),
	.w8(32'hbad60641),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6b4f),
	.w1(32'hbb00ea5e),
	.w2(32'hbba01875),
	.w3(32'hbac835af),
	.w4(32'hbb83ecef),
	.w5(32'hba862fdb),
	.w6(32'hbab6fc6d),
	.w7(32'hbaa6cd2e),
	.w8(32'hbbcf17da),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebd941),
	.w1(32'hbaf28922),
	.w2(32'h3c1986ec),
	.w3(32'hbb835bd8),
	.w4(32'h3b2fd54e),
	.w5(32'h3b8c3de0),
	.w6(32'hbc0a2dda),
	.w7(32'hbacd5cdc),
	.w8(32'h3bf35ac4),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37121b01),
	.w1(32'hbbc2926d),
	.w2(32'hbacdd529),
	.w3(32'h3a8927c3),
	.w4(32'hbab0906e),
	.w5(32'h3a7a00c4),
	.w6(32'h39b806eb),
	.w7(32'hbc003ef9),
	.w8(32'hbad65fa5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57233c),
	.w1(32'hbbd613aa),
	.w2(32'hb9f67303),
	.w3(32'h3bb660fe),
	.w4(32'h3a44874a),
	.w5(32'h399b4986),
	.w6(32'h3be33cc5),
	.w7(32'h3b834cb0),
	.w8(32'hb9a9ce7d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0977cc),
	.w1(32'hb9981948),
	.w2(32'h3b91c642),
	.w3(32'h3b244087),
	.w4(32'hba91159c),
	.w5(32'hba8f2c2a),
	.w6(32'hb998c622),
	.w7(32'h39ba9cd8),
	.w8(32'hba7a85bd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0273a7),
	.w1(32'h3be8ef5a),
	.w2(32'hbba54e0c),
	.w3(32'hbbb7bfc9),
	.w4(32'h3c004f17),
	.w5(32'hbbce9063),
	.w6(32'h3a608d41),
	.w7(32'hbc33242e),
	.w8(32'hbb2a02f7),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc168370),
	.w1(32'hba04900b),
	.w2(32'h3aefe03d),
	.w3(32'hbc1abc21),
	.w4(32'hbbb25da2),
	.w5(32'h3b7279b1),
	.w6(32'hbbb376ff),
	.w7(32'hbbf9ada9),
	.w8(32'h3b6c6be2),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9448d8),
	.w1(32'hbb5740bc),
	.w2(32'h3adf6b17),
	.w3(32'h3b97f1fc),
	.w4(32'hbae82785),
	.w5(32'hbb27fc54),
	.w6(32'h3bd5dad7),
	.w7(32'h3a545482),
	.w8(32'hbae752e2),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87e531),
	.w1(32'h3b0d96ad),
	.w2(32'h3afc221e),
	.w3(32'h3c06c31c),
	.w4(32'hbb2467f7),
	.w5(32'h3aaed303),
	.w6(32'h3ba1641c),
	.w7(32'h3ba15ea3),
	.w8(32'hbb0c5209),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a4440),
	.w1(32'hba8d90b1),
	.w2(32'h38a046dd),
	.w3(32'h3c0b3250),
	.w4(32'h3bc671ab),
	.w5(32'hba849233),
	.w6(32'h3be14b62),
	.w7(32'h3b959e1d),
	.w8(32'h3b04879e),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dc520),
	.w1(32'hbb35ae4a),
	.w2(32'h3a1f26e0),
	.w3(32'h3b67921b),
	.w4(32'h3bd388c4),
	.w5(32'h3c201a9f),
	.w6(32'hba8a0183),
	.w7(32'hba817381),
	.w8(32'h3c149da8),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11cee8),
	.w1(32'hbbbd6cad),
	.w2(32'hbb332890),
	.w3(32'hbb757073),
	.w4(32'hbb550a6c),
	.w5(32'hbbba9726),
	.w6(32'hbae03c0f),
	.w7(32'h3b1b7ad3),
	.w8(32'hbb8c0de3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb809d50),
	.w1(32'h3ae0244e),
	.w2(32'hbafbeca1),
	.w3(32'hbba96c6e),
	.w4(32'hbae72131),
	.w5(32'hbb3cc2d2),
	.w6(32'hbb2c0680),
	.w7(32'h3ada4493),
	.w8(32'h3ae3d086),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ff921),
	.w1(32'hbc13a1b6),
	.w2(32'hbabd4160),
	.w3(32'hbc5e8eef),
	.w4(32'hbc206978),
	.w5(32'h3b0c6671),
	.w6(32'hbbfe4153),
	.w7(32'hbc285568),
	.w8(32'h3b279f77),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb070cf1),
	.w1(32'h3ba38b4d),
	.w2(32'hbbd1689c),
	.w3(32'h3bc42076),
	.w4(32'h3ac88d42),
	.w5(32'hbadaf976),
	.w6(32'hbb5db520),
	.w7(32'hbb28a7ab),
	.w8(32'hbbd56579),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14fc82),
	.w1(32'h3c17b47d),
	.w2(32'hbbba5574),
	.w3(32'hbb98b1a8),
	.w4(32'h3c5dd6be),
	.w5(32'h3bd3951b),
	.w6(32'hbc2a9cab),
	.w7(32'h3a4f8953),
	.w8(32'h3b59306a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53d4fe),
	.w1(32'hbba0c8c4),
	.w2(32'h392041e4),
	.w3(32'hba3a95c2),
	.w4(32'h3b892826),
	.w5(32'hba3712c5),
	.w6(32'h3b837005),
	.w7(32'h3c4629e9),
	.w8(32'h39cb7ed7),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e1e9),
	.w1(32'h3a013bf7),
	.w2(32'h3c33f05f),
	.w3(32'hb90a0702),
	.w4(32'hb90ba3c9),
	.w5(32'h3bcde4f0),
	.w6(32'h3813e582),
	.w7(32'h3a568ca2),
	.w8(32'h3c12ef01),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27fc92),
	.w1(32'hbbfb8215),
	.w2(32'hba179a47),
	.w3(32'hbb7cc007),
	.w4(32'hbc828dad),
	.w5(32'h3a75228c),
	.w6(32'hb80b8c51),
	.w7(32'hbc261f1f),
	.w8(32'hba81f1c3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8e7ae),
	.w1(32'hbb9ff5dd),
	.w2(32'h3bdf7580),
	.w3(32'h3b151581),
	.w4(32'hbb26c744),
	.w5(32'h3b1715da),
	.w6(32'h397a7730),
	.w7(32'hbb8920c5),
	.w8(32'hba95f12c),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9ba0b),
	.w1(32'h3ca9cc49),
	.w2(32'h39bf9685),
	.w3(32'h3cbe5e97),
	.w4(32'h3c8040aa),
	.w5(32'h3b8b5f97),
	.w6(32'h3c44c0e8),
	.w7(32'h3c88a2b6),
	.w8(32'h3b38f24f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf10156),
	.w1(32'hbcc12c75),
	.w2(32'hb8a2c594),
	.w3(32'hbc3bec5d),
	.w4(32'hbbad0b64),
	.w5(32'hbbf40fa4),
	.w6(32'hbb9ca432),
	.w7(32'hbba9500b),
	.w8(32'hbbbd4892),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb844b9b),
	.w1(32'hbc05bd1d),
	.w2(32'h3b3ef5d9),
	.w3(32'hbbc20e20),
	.w4(32'h3bc5a126),
	.w5(32'hbb6e1d16),
	.w6(32'hbbfa97dc),
	.w7(32'h3b9e51c0),
	.w8(32'hbc9b4d6b),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8da749),
	.w1(32'h3c80f028),
	.w2(32'h3bf6fab7),
	.w3(32'h3cf573c1),
	.w4(32'h3ccbb8ea),
	.w5(32'h3bbca30f),
	.w6(32'h3a3dd92b),
	.w7(32'h3bf874a9),
	.w8(32'h3b4795c0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba49497),
	.w1(32'hb9f6476a),
	.w2(32'hbb81a6d9),
	.w3(32'h3c20e34b),
	.w4(32'h3ba529ce),
	.w5(32'hbb96ceee),
	.w6(32'h3c3954e6),
	.w7(32'h3c0d7a0b),
	.w8(32'hbb5d032c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb749820),
	.w1(32'hbb13a63d),
	.w2(32'hbc48164a),
	.w3(32'hbb8e4836),
	.w4(32'hbaf96d48),
	.w5(32'hbb92e220),
	.w6(32'hbb9c9514),
	.w7(32'hbb34e210),
	.w8(32'hbc172f5b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13a6c3),
	.w1(32'h39eed6ff),
	.w2(32'hbc15b7cc),
	.w3(32'hbc03aaef),
	.w4(32'h3bdef659),
	.w5(32'hbc1cd6a3),
	.w6(32'hbb99403a),
	.w7(32'hbbb29796),
	.w8(32'hbbd673fd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f520),
	.w1(32'h3bfc13dd),
	.w2(32'hb73f0013),
	.w3(32'hbbe248a6),
	.w4(32'h3c1aa4b2),
	.w5(32'hbb059e8c),
	.w6(32'hbb572ad1),
	.w7(32'h3b537388),
	.w8(32'hbaa226e7),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55d15b),
	.w1(32'hbc018b32),
	.w2(32'hbad5b5ea),
	.w3(32'hbb54d101),
	.w4(32'h3b4e8a1e),
	.w5(32'h3aa97b9e),
	.w6(32'h3bbba357),
	.w7(32'h3c861057),
	.w8(32'h39e18a50),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afee269),
	.w1(32'hbbde0a6e),
	.w2(32'hbb03eda4),
	.w3(32'h3ba2e747),
	.w4(32'hbbd5e808),
	.w5(32'hba808b69),
	.w6(32'h3b9a79af),
	.w7(32'h39ac9019),
	.w8(32'h3abeabd7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb947b6d3),
	.w1(32'h3b969447),
	.w2(32'h3b9a310c),
	.w3(32'h3aee92ea),
	.w4(32'h3bc2b1d3),
	.w5(32'h3b458c61),
	.w6(32'h37d6c94f),
	.w7(32'h3b94d359),
	.w8(32'h3ad3dcc7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedb0bf),
	.w1(32'h3b414d17),
	.w2(32'hbbc3ff91),
	.w3(32'hb99ab7e2),
	.w4(32'h3b03a46d),
	.w5(32'hb9bb78a2),
	.w6(32'hba7dd15d),
	.w7(32'hbaf2b9f9),
	.w8(32'hbace751d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90cf01),
	.w1(32'hbba58d4b),
	.w2(32'hbb69ed50),
	.w3(32'hbb21775a),
	.w4(32'hbb445f06),
	.w5(32'hbb9ffc92),
	.w6(32'hbbda58f0),
	.w7(32'hbc0ccf9b),
	.w8(32'hb97ddc3f),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fa006),
	.w1(32'hb9f31961),
	.w2(32'h3ac77c9b),
	.w3(32'hbb61d662),
	.w4(32'hbbd711a1),
	.w5(32'h3b4c1b79),
	.w6(32'hbb1c8f5f),
	.w7(32'hbc11f60f),
	.w8(32'hba4f9c35),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8669a2),
	.w1(32'hbab6600d),
	.w2(32'hbb3fb0fa),
	.w3(32'hbc2bb2e4),
	.w4(32'hbc20b8c0),
	.w5(32'hbb968793),
	.w6(32'hbbe629ef),
	.w7(32'hbc0d11bc),
	.w8(32'hbc1449e8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc581e77),
	.w1(32'hba68052b),
	.w2(32'hbc8f2f38),
	.w3(32'hbb4d1db9),
	.w4(32'h3c113ebb),
	.w5(32'hbc8a4863),
	.w6(32'hbc1b3198),
	.w7(32'h3c66925d),
	.w8(32'hbc272674),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62f57f),
	.w1(32'h3c220c0d),
	.w2(32'h3c333f66),
	.w3(32'hbc51a1c4),
	.w4(32'h3cb7c66d),
	.w5(32'h3c1b748b),
	.w6(32'hbc601c3c),
	.w7(32'h3b4dd8b8),
	.w8(32'h3c67b8f1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2a446),
	.w1(32'hbc10a0e7),
	.w2(32'hbb405f0d),
	.w3(32'hbc2805bc),
	.w4(32'hbcbdc8af),
	.w5(32'hbae0ffc9),
	.w6(32'hbb51f558),
	.w7(32'hbc801b0f),
	.w8(32'h3bae427c),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1142d),
	.w1(32'h3ba89156),
	.w2(32'h3a4b5732),
	.w3(32'hbb5520c9),
	.w4(32'h3bb8c9ae),
	.w5(32'hbc18bca5),
	.w6(32'hbbca7c24),
	.w7(32'h3b2686fe),
	.w8(32'hbc049698),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5670ba),
	.w1(32'h3bd01351),
	.w2(32'hb83d778e),
	.w3(32'hbb8008a5),
	.w4(32'h3c01582e),
	.w5(32'h3b8f4e7a),
	.w6(32'hbbc44177),
	.w7(32'hbbc686dd),
	.w8(32'h3b8e71a8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc116b02),
	.w1(32'hba27f6ff),
	.w2(32'hba121e50),
	.w3(32'h3b1e7bbe),
	.w4(32'h3b5f7c2a),
	.w5(32'hbba71955),
	.w6(32'h3b8ee6d2),
	.w7(32'h3a63d99c),
	.w8(32'hbaee39e6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc5899),
	.w1(32'hbadcc749),
	.w2(32'hbad3da3b),
	.w3(32'hbc54027d),
	.w4(32'hbbfc63bf),
	.w5(32'hbc4517e4),
	.w6(32'hbc27508e),
	.w7(32'hbba3f00f),
	.w8(32'hbc34f88f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b778d69),
	.w1(32'h3c681134),
	.w2(32'h39c39f41),
	.w3(32'h3b4ff22d),
	.w4(32'h3c9d3198),
	.w5(32'hbb14c059),
	.w6(32'hbbd2b11d),
	.w7(32'h3ba39dd0),
	.w8(32'hb9ae88bc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53ecea),
	.w1(32'h3bec4dde),
	.w2(32'hbaae2660),
	.w3(32'h3bbcede5),
	.w4(32'h3be14e5f),
	.w5(32'hbb75e4bd),
	.w6(32'hba3bce05),
	.w7(32'h3989846e),
	.w8(32'hbb90e325),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd57db),
	.w1(32'h3bc62fa5),
	.w2(32'hbc148aaf),
	.w3(32'h3c5d00e0),
	.w4(32'h3c069393),
	.w5(32'hbbd6aa04),
	.w6(32'h3c08a931),
	.w7(32'h3b8458d0),
	.w8(32'h3b2ad420),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc881540),
	.w1(32'hbc7b7ae4),
	.w2(32'hba45722d),
	.w3(32'hbc45ac6e),
	.w4(32'hbc45f853),
	.w5(32'hbbd1f024),
	.w6(32'hbbd03766),
	.w7(32'hbb585ef8),
	.w8(32'hbc3523cb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09833f),
	.w1(32'hbbc5f445),
	.w2(32'hbb19d6e7),
	.w3(32'hbae1a90d),
	.w4(32'h3b73b102),
	.w5(32'hbb8a852f),
	.w6(32'hbb51a4bf),
	.w7(32'h38a79b88),
	.w8(32'hbbbb2857),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3010a),
	.w1(32'h3b630e7e),
	.w2(32'hba5c5ec4),
	.w3(32'hbb84c29c),
	.w4(32'h3b938d3b),
	.w5(32'hbbb4284c),
	.w6(32'hbc17ff07),
	.w7(32'h3b884d65),
	.w8(32'hbb91aa21),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a2801),
	.w1(32'h3bc4e23e),
	.w2(32'hbbc85895),
	.w3(32'h397b0af2),
	.w4(32'h3c01bfbb),
	.w5(32'hbc1638c9),
	.w6(32'hbc497061),
	.w7(32'hba7a0daf),
	.w8(32'hbc43d867),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2119f4),
	.w1(32'h38d2e286),
	.w2(32'h3c10dd8f),
	.w3(32'h3bcac853),
	.w4(32'h3c1711f3),
	.w5(32'h3ba752a0),
	.w6(32'hbac28dd3),
	.w7(32'h3a858033),
	.w8(32'hbb234564),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60e98e),
	.w1(32'h3b0ddcb6),
	.w2(32'hbc829ac7),
	.w3(32'hba5eea75),
	.w4(32'h3c00dd82),
	.w5(32'hbc73106a),
	.w6(32'hbbfc3c78),
	.w7(32'hbc036781),
	.w8(32'hbc50ab6b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912ed14),
	.w1(32'h3bece067),
	.w2(32'hbbe153d8),
	.w3(32'hbc1edd13),
	.w4(32'h3c943b39),
	.w5(32'hbc2b5a34),
	.w6(32'hbc4dde84),
	.w7(32'h3c52721e),
	.w8(32'hb7cf8517),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e97be),
	.w1(32'hbb67ddb6),
	.w2(32'h3b1d1259),
	.w3(32'hbc1436d7),
	.w4(32'hbb0eee97),
	.w5(32'h3b532f19),
	.w6(32'hbafebf72),
	.w7(32'hbbb992a7),
	.w8(32'h3b8e8525),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2daa4d),
	.w1(32'h3c3d70f2),
	.w2(32'hbb903db6),
	.w3(32'hbb1f337d),
	.w4(32'hbacfe554),
	.w5(32'hbc046b99),
	.w6(32'hbb025249),
	.w7(32'hbbf4bf0d),
	.w8(32'hbc2217a0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66d5fa),
	.w1(32'hbbea6ad4),
	.w2(32'hbb84b4fe),
	.w3(32'hbb9ced6e),
	.w4(32'h395e70b2),
	.w5(32'hba8452dd),
	.w6(32'hba1690fe),
	.w7(32'h3c25f1ed),
	.w8(32'hbad3c129),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f99267),
	.w1(32'h3c08defb),
	.w2(32'hbc7347b9),
	.w3(32'hbb564295),
	.w4(32'h3b354bf2),
	.w5(32'hbc6a3e84),
	.w6(32'hbb2d4e96),
	.w7(32'h3b00b08d),
	.w8(32'hbc91cc13),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8f60a),
	.w1(32'h3cd5fc27),
	.w2(32'hbb85b6b7),
	.w3(32'hbc4df64b),
	.w4(32'h3cb6dda8),
	.w5(32'h3b4e4ce3),
	.w6(32'hbc75d055),
	.w7(32'h3bfa25ea),
	.w8(32'h3c0d5881),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11bab5),
	.w1(32'hba954d34),
	.w2(32'h3ad387db),
	.w3(32'hbbdccbb9),
	.w4(32'hba8b1012),
	.w5(32'hbb2b1478),
	.w6(32'hbb3058a3),
	.w7(32'hbb8da60c),
	.w8(32'hbb793dfa),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa61951),
	.w1(32'hbb9d3c90),
	.w2(32'hb9ed68a8),
	.w3(32'hbbc2d10a),
	.w4(32'hbc3115ce),
	.w5(32'hb8d48001),
	.w6(32'hbb8fc301),
	.w7(32'hba90a317),
	.w8(32'hbad16f1c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eac265),
	.w1(32'hbb2df92d),
	.w2(32'hb8bd41b2),
	.w3(32'h3a1a21f8),
	.w4(32'hbb4f94bb),
	.w5(32'hbb360152),
	.w6(32'hbad4d1d7),
	.w7(32'hbba50904),
	.w8(32'hbb59966e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f20be),
	.w1(32'hbb28ba47),
	.w2(32'hba4b3e38),
	.w3(32'hbb8b43aa),
	.w4(32'hba6aa1af),
	.w5(32'hbb531e56),
	.w6(32'hbb9fc9cd),
	.w7(32'hbb1323d1),
	.w8(32'h3b156014),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe47841),
	.w1(32'hbbb60b05),
	.w2(32'hba1d6f88),
	.w3(32'hbc96b377),
	.w4(32'hbb25b273),
	.w5(32'hbaffd315),
	.w6(32'hbc28baba),
	.w7(32'hbbc1db4c),
	.w8(32'hbb8da3ba),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0efcc6),
	.w1(32'h3bca3bf7),
	.w2(32'hbbe80223),
	.w3(32'h3bef8fe6),
	.w4(32'h3bd6a945),
	.w5(32'h3a222e20),
	.w6(32'hb90a44bf),
	.w7(32'h3b88271e),
	.w8(32'hbbeea75d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dc4fe),
	.w1(32'h3bb44ebf),
	.w2(32'hbb28952e),
	.w3(32'hbb55d5e7),
	.w4(32'hbbb4a541),
	.w5(32'hbbda0a34),
	.w6(32'hbc60ebb6),
	.w7(32'hbc93499e),
	.w8(32'h3a5f2030),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa68d3f),
	.w1(32'h3b1491b9),
	.w2(32'h3b431695),
	.w3(32'hbb8e4c25),
	.w4(32'h3a7f8273),
	.w5(32'hb8a7da5c),
	.w6(32'hbaeb30da),
	.w7(32'h3a8cb6cb),
	.w8(32'h3acda9ea),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b677a62),
	.w1(32'h3a0d03e0),
	.w2(32'hbbb20ff1),
	.w3(32'h3bdb71ae),
	.w4(32'h3ae68f1b),
	.w5(32'hbb9de088),
	.w6(32'h3a3c1dd4),
	.w7(32'hbb4e81f9),
	.w8(32'hbb0e3af3),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule