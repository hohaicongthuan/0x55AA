module LineBuffer(data_in, data_out, Clk, valid_in, Rst);
    parameter DATA_WIDTH = 8;
    parameter BUFFER_DEPTH = 97;

    input  Clk, valid_in, Rst;
    input  [DATA_WIDTH - 1:0] data_in;

    output reg [DATA_WIDTH - 1:0] data_out;

	reg [DATA_WIDTH - 1:0] Buffer [BUFFER_DEPTH - 1:0];
	 
    always @ (posedge Clk or negedge Rst) begin
        if (!Rst) begin
            Buffer[0] <= 0;
            Buffer[1] <= 0;
            Buffer[2] <= 0;
            Buffer[3] <= 0;
            Buffer[4] <= 0;
            Buffer[5] <= 0;
            Buffer[6] <= 0;
            Buffer[7] <= 0;
            Buffer[8] <= 0;
            Buffer[9] <= 0;
            Buffer[10] <= 0;
            Buffer[11] <= 0;
            Buffer[12] <= 0;
            Buffer[13] <= 0;
            Buffer[14] <= 0;
            Buffer[15] <= 0;
            Buffer[16] <= 0;
            Buffer[17] <= 0;
            Buffer[18] <= 0;
            Buffer[19] <= 0;
            Buffer[20] <= 0;
            Buffer[21] <= 0;
            Buffer[22] <= 0;
            Buffer[23] <= 0;
            Buffer[24] <= 0;
            Buffer[25] <= 0;
            Buffer[26] <= 0;
            Buffer[27] <= 0;
            Buffer[28] <= 0;
            Buffer[29] <= 0;
            Buffer[30] <= 0;
            Buffer[31] <= 0;
            Buffer[32] <= 0;
            Buffer[33] <= 0;
            Buffer[34] <= 0;
            Buffer[35] <= 0;
            Buffer[36] <= 0;
            Buffer[37] <= 0;
            Buffer[38] <= 0;
            Buffer[39] <= 0;
            Buffer[40] <= 0;
            Buffer[41] <= 0;
            Buffer[42] <= 0;
            Buffer[43] <= 0;
            Buffer[44] <= 0;
            Buffer[45] <= 0;
            Buffer[46] <= 0;
            Buffer[47] <= 0;
            Buffer[48] <= 0;
            Buffer[49] <= 0;
            Buffer[50] <= 0;
            Buffer[51] <= 0;
            Buffer[52] <= 0;
            Buffer[53] <= 0;
            Buffer[54] <= 0;
            Buffer[55] <= 0;
            Buffer[56] <= 0;
            Buffer[57] <= 0;
            Buffer[58] <= 0;
            Buffer[59] <= 0;
            Buffer[60] <= 0;
            Buffer[61] <= 0;
            Buffer[62] <= 0;
            Buffer[63] <= 0;
            Buffer[64] <= 0;
            Buffer[65] <= 0;
            Buffer[66] <= 0;
            Buffer[67] <= 0;
            Buffer[68] <= 0;
            Buffer[69] <= 0;
            Buffer[70] <= 0;
            Buffer[71] <= 0;
            Buffer[72] <= 0;
            Buffer[73] <= 0;
            Buffer[74] <= 0;
            Buffer[75] <= 0;
            Buffer[76] <= 0;
            Buffer[77] <= 0;
            Buffer[78] <= 0;
            Buffer[79] <= 0;
            Buffer[80] <= 0;
            Buffer[81] <= 0;
            Buffer[82] <= 0;
            Buffer[83] <= 0;
            Buffer[84] <= 0;
            Buffer[85] <= 0;
            Buffer[86] <= 0;
            Buffer[87] <= 0;
            Buffer[88] <= 0;
            Buffer[89] <= 0;
            Buffer[90] <= 0;
            Buffer[91] <= 0;
            Buffer[92] <= 0;
            Buffer[93] <= 0;
            Buffer[94] <= 0;
            Buffer[95] <= 0;
            Buffer[96] <= 0;
        end else
        if (valid_in) begin
            data_out <= Buffer[BUFFER_DEPTH - 1];
            
            Buffer[1] <= Buffer[0];
            Buffer[2] <= Buffer[1];
            Buffer[3] <= Buffer[2];
            Buffer[4] <= Buffer[3];
            Buffer[5] <= Buffer[4];
            Buffer[6] <= Buffer[5];
            Buffer[7] <= Buffer[6];
            Buffer[8] <= Buffer[7];
            Buffer[9] <= Buffer[8];
            Buffer[10] <= Buffer[9];
            Buffer[11] <= Buffer[10];
            Buffer[12] <= Buffer[11];
            Buffer[13] <= Buffer[12];
            Buffer[14] <= Buffer[13];
            Buffer[15] <= Buffer[14];
            Buffer[16] <= Buffer[15];
            Buffer[17] <= Buffer[16];
            Buffer[18] <= Buffer[17];
            Buffer[19] <= Buffer[18];
            Buffer[20] <= Buffer[19];
            Buffer[21] <= Buffer[20];
            Buffer[22] <= Buffer[21];
            Buffer[23] <= Buffer[22];
            Buffer[24] <= Buffer[23];
            Buffer[25] <= Buffer[24];
            Buffer[26] <= Buffer[25];
            Buffer[27] <= Buffer[26];
            Buffer[28] <= Buffer[27];
            Buffer[29] <= Buffer[28];
            Buffer[30] <= Buffer[29];
            Buffer[31] <= Buffer[30];
            Buffer[32] <= Buffer[31];
            Buffer[33] <= Buffer[32];
            Buffer[34] <= Buffer[33];
            Buffer[35] <= Buffer[34];
            Buffer[36] <= Buffer[35];
            Buffer[37] <= Buffer[36];
            Buffer[38] <= Buffer[37];
            Buffer[39] <= Buffer[38];
            Buffer[40] <= Buffer[39];
            Buffer[41] <= Buffer[40];
            Buffer[42] <= Buffer[41];
            Buffer[43] <= Buffer[42];
            Buffer[44] <= Buffer[43];
            Buffer[45] <= Buffer[44];
            Buffer[46] <= Buffer[45];
            Buffer[47] <= Buffer[46];
            Buffer[48] <= Buffer[47];
            Buffer[49] <= Buffer[48];
            Buffer[50] <= Buffer[49];
            Buffer[51] <= Buffer[50];
            Buffer[52] <= Buffer[51];
            Buffer[53] <= Buffer[52];
            Buffer[54] <= Buffer[53];
            Buffer[55] <= Buffer[54];
            Buffer[56] <= Buffer[55];
            Buffer[57] <= Buffer[56];
            Buffer[58] <= Buffer[57];
            Buffer[59] <= Buffer[58];
            Buffer[60] <= Buffer[59];
            Buffer[61] <= Buffer[60];
            Buffer[62] <= Buffer[61];
            Buffer[63] <= Buffer[62];
            Buffer[64] <= Buffer[63];
            Buffer[65] <= Buffer[64];
            Buffer[66] <= Buffer[65];
            Buffer[67] <= Buffer[66];
            Buffer[68] <= Buffer[67];
            Buffer[69] <= Buffer[68];
            Buffer[70] <= Buffer[69];
            Buffer[71] <= Buffer[70];
            Buffer[72] <= Buffer[71];
            Buffer[73] <= Buffer[72];
            Buffer[74] <= Buffer[73];
            Buffer[75] <= Buffer[74];
            Buffer[76] <= Buffer[75];
            Buffer[77] <= Buffer[76];
            Buffer[78] <= Buffer[77];
            Buffer[79] <= Buffer[78];
            Buffer[80] <= Buffer[79];
            Buffer[81] <= Buffer[80];
            Buffer[82] <= Buffer[81];
            Buffer[83] <= Buffer[82];
            Buffer[84] <= Buffer[83];
            Buffer[85] <= Buffer[84];
            Buffer[86] <= Buffer[85];
            Buffer[87] <= Buffer[86];
            Buffer[88] <= Buffer[87];
            Buffer[89] <= Buffer[88];
            Buffer[90] <= Buffer[89];
            Buffer[91] <= Buffer[90];
            Buffer[92] <= Buffer[91];
            Buffer[93] <= Buffer[92];
            Buffer[94] <= Buffer[93];
            Buffer[95] <= Buffer[94];
            Buffer[96] <= Buffer[95];
            
            Buffer[0] <= data_in;
        end else begin
            Buffer[0] <= Buffer[0];
            Buffer[1] <= Buffer[1];
            Buffer[2] <= Buffer[2];
            Buffer[3] <= Buffer[3];
            Buffer[4] <= Buffer[4];
            Buffer[5] <= Buffer[5];
            Buffer[6] <= Buffer[6];
            Buffer[7] <= Buffer[7];
            Buffer[8] <= Buffer[8];
            Buffer[9] <= Buffer[9];
            Buffer[10] <= Buffer[10];
            Buffer[11] <= Buffer[11];
            Buffer[12] <= Buffer[12];
            Buffer[13] <= Buffer[13];
            Buffer[14] <= Buffer[14];
            Buffer[15] <= Buffer[15];
            Buffer[16] <= Buffer[16];
            Buffer[17] <= Buffer[17];
            Buffer[18] <= Buffer[18];
            Buffer[19] <= Buffer[19];
            Buffer[20] <= Buffer[20];
            Buffer[21] <= Buffer[21];
            Buffer[22] <= Buffer[22];
            Buffer[23] <= Buffer[23];
            Buffer[24] <= Buffer[24];
            Buffer[25] <= Buffer[25];
            Buffer[26] <= Buffer[26];
            Buffer[27] <= Buffer[27];
            Buffer[28] <= Buffer[28];
            Buffer[29] <= Buffer[29];
            Buffer[30] <= Buffer[30];
            Buffer[31] <= Buffer[31];
            Buffer[32] <= Buffer[32];
            Buffer[33] <= Buffer[33];
            Buffer[34] <= Buffer[34];
            Buffer[35] <= Buffer[35];
            Buffer[36] <= Buffer[36];
            Buffer[37] <= Buffer[37];
            Buffer[38] <= Buffer[38];
            Buffer[39] <= Buffer[39];
            Buffer[40] <= Buffer[40];
            Buffer[41] <= Buffer[41];
            Buffer[42] <= Buffer[42];
            Buffer[43] <= Buffer[43];
            Buffer[44] <= Buffer[44];
            Buffer[45] <= Buffer[45];
            Buffer[46] <= Buffer[46];
            Buffer[47] <= Buffer[47];
            Buffer[48] <= Buffer[48];
            Buffer[49] <= Buffer[49];
            Buffer[50] <= Buffer[50];
            Buffer[51] <= Buffer[51];
            Buffer[52] <= Buffer[52];
            Buffer[53] <= Buffer[53];
            Buffer[54] <= Buffer[54];
            Buffer[55] <= Buffer[55];
            Buffer[56] <= Buffer[56];
            Buffer[57] <= Buffer[57];
            Buffer[58] <= Buffer[58];
            Buffer[59] <= Buffer[59];
            Buffer[60] <= Buffer[60];
            Buffer[61] <= Buffer[61];
            Buffer[62] <= Buffer[62];
            Buffer[63] <= Buffer[63];
            Buffer[64] <= Buffer[64];
            Buffer[65] <= Buffer[65];
            Buffer[66] <= Buffer[66];
            Buffer[67] <= Buffer[67];
            Buffer[68] <= Buffer[68];
            Buffer[69] <= Buffer[69];
            Buffer[70] <= Buffer[70];
            Buffer[71] <= Buffer[71];
            Buffer[72] <= Buffer[72];
            Buffer[73] <= Buffer[73];
            Buffer[74] <= Buffer[74];
            Buffer[75] <= Buffer[75];
            Buffer[76] <= Buffer[76];
            Buffer[77] <= Buffer[77];
            Buffer[78] <= Buffer[78];
            Buffer[79] <= Buffer[79];
            Buffer[80] <= Buffer[80];
            Buffer[81] <= Buffer[81];
            Buffer[82] <= Buffer[82];
            Buffer[83] <= Buffer[83];
            Buffer[84] <= Buffer[84];
            Buffer[85] <= Buffer[85];
            Buffer[86] <= Buffer[86];
            Buffer[87] <= Buffer[87];
            Buffer[88] <= Buffer[88];
            Buffer[89] <= Buffer[89];
            Buffer[90] <= Buffer[90];
            Buffer[91] <= Buffer[91];
            Buffer[92] <= Buffer[92];
            Buffer[93] <= Buffer[93];
            Buffer[94] <= Buffer[94];
            Buffer[95] <= Buffer[95];
            Buffer[96] <= Buffer[96];
        end
	end
endmodule