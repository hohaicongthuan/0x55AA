module layer_10_featuremap_175(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91e3951),
	.w1(32'hb8032629),
	.w2(32'hb823e6c5),
	.w3(32'hb917329d),
	.w4(32'hb50b316b),
	.w5(32'h370bc24d),
	.w6(32'hb911744d),
	.w7(32'h3751e880),
	.w8(32'hb790ab14),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e687c),
	.w1(32'h3b92d552),
	.w2(32'h3bb27502),
	.w3(32'h3c10a3df),
	.w4(32'hbaf8de87),
	.w5(32'h39b45ce4),
	.w6(32'h3bd6ca5d),
	.w7(32'hbb7e46f6),
	.w8(32'h39d21329),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a28c3f),
	.w1(32'hb76c3e27),
	.w2(32'hb80e6831),
	.w3(32'hb884bee5),
	.w4(32'hb637e833),
	.w5(32'hb7af1a05),
	.w6(32'hb8814d79),
	.w7(32'hb6f2b2d5),
	.w8(32'hb7f27b12),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bcdc48),
	.w1(32'hba49927b),
	.w2(32'hbaa20297),
	.w3(32'h3a0e6815),
	.w4(32'h3a367a56),
	.w5(32'h3924e314),
	.w6(32'hb9db21ac),
	.w7(32'hbaa2b988),
	.w8(32'hba9718b3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54836a),
	.w1(32'h38561001),
	.w2(32'h3a6498f1),
	.w3(32'hba6288a8),
	.w4(32'hba1c575b),
	.w5(32'h395ae670),
	.w6(32'hba5ab463),
	.w7(32'hba63e7d4),
	.w8(32'hba148613),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb931f54d),
	.w1(32'hb7b0bf3a),
	.w2(32'hb854c7c4),
	.w3(32'hb915aa13),
	.w4(32'hb7edca92),
	.w5(32'hb89bdb99),
	.w6(32'hb90fe920),
	.w7(32'hb73d7474),
	.w8(32'hb8acbdcf),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e018a),
	.w1(32'h3b8145a5),
	.w2(32'h3c11ca0d),
	.w3(32'hba90802f),
	.w4(32'h3be26d55),
	.w5(32'h3c2a0e5d),
	.w6(32'hbb978bac),
	.w7(32'h3b81dc4c),
	.w8(32'h3c1e28fc),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f5d23),
	.w1(32'h3c313df7),
	.w2(32'h3bf3154f),
	.w3(32'h3c89a6e5),
	.w4(32'h3c8b9b9e),
	.w5(32'h3c371de6),
	.w6(32'h3c4052ae),
	.w7(32'h3b86d18a),
	.w8(32'h3bd5e25d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f3c52),
	.w1(32'hba47b386),
	.w2(32'h3a508c5b),
	.w3(32'h3a29d98f),
	.w4(32'hbacdccfd),
	.w5(32'h3a76b2d1),
	.w6(32'h3a0fc668),
	.w7(32'hba2695b0),
	.w8(32'h399ad9a1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c958ba6),
	.w1(32'h3b59b492),
	.w2(32'h3c88010d),
	.w3(32'h3c89fcfb),
	.w4(32'hb960452e),
	.w5(32'h3bf84092),
	.w6(32'h3c4b6a28),
	.w7(32'hb90f9303),
	.w8(32'h3bd1ef4f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff9971),
	.w1(32'h3afef539),
	.w2(32'h3b1b293b),
	.w3(32'h3ac9ad39),
	.w4(32'h3a0c55c1),
	.w5(32'h3ac7c52f),
	.w6(32'h3ace199c),
	.w7(32'h39b20e56),
	.w8(32'h3a7eb479),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88eebe),
	.w1(32'hbbbfde4d),
	.w2(32'h3b8081c6),
	.w3(32'h3ba23fb0),
	.w4(32'hba4d095f),
	.w5(32'h3bf0f42b),
	.w6(32'hba638412),
	.w7(32'hbbc6ca71),
	.w8(32'h3c192dc5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c03bd),
	.w1(32'h3bb436fd),
	.w2(32'h3ca3dba8),
	.w3(32'h3c28924b),
	.w4(32'h3b806cc4),
	.w5(32'h3c569f34),
	.w6(32'h3be30f98),
	.w7(32'h3b8b77f0),
	.w8(32'h3c3eaf9e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fbb7),
	.w1(32'h3c159c97),
	.w2(32'h3c4eec7b),
	.w3(32'h3b41edb5),
	.w4(32'h3bd8ba06),
	.w5(32'h3c0658c3),
	.w6(32'h3b9fb37f),
	.w7(32'h3bd14c1b),
	.w8(32'h3bc68e9f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c151c2d),
	.w1(32'hbad9bd44),
	.w2(32'h3b09baa9),
	.w3(32'h3bc9701f),
	.w4(32'hbbe2c2f1),
	.w5(32'hbb790b3e),
	.w6(32'h3c044a89),
	.w7(32'hbbaf1de5),
	.w8(32'hbb2ed6c6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72566f),
	.w1(32'h3b232a27),
	.w2(32'h3c3caa2f),
	.w3(32'h3c5390e2),
	.w4(32'hba9a4587),
	.w5(32'h3b0b608f),
	.w6(32'h3c608598),
	.w7(32'h3b5430f2),
	.w8(32'h3b67b5c4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d8b078),
	.w1(32'hb9d970fa),
	.w2(32'hb9bbf58a),
	.w3(32'hb8b80cdd),
	.w4(32'hb9cefb8f),
	.w5(32'hb9ae9474),
	.w6(32'hb9d4b166),
	.w7(32'hba9a4ee3),
	.w8(32'hba7c94fa),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c823376),
	.w1(32'h3c1e45bd),
	.w2(32'h3c779534),
	.w3(32'h3c6d2261),
	.w4(32'h3bd2e5ce),
	.w5(32'h3c87f2c0),
	.w6(32'h3c21fbc9),
	.w7(32'h3a189202),
	.w8(32'h3c02b9d4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd97b5b),
	.w1(32'h3b9c4501),
	.w2(32'h3c38c219),
	.w3(32'h3b9c4681),
	.w4(32'h3b7f1ea8),
	.w5(32'h3c224811),
	.w6(32'h3af2107b),
	.w7(32'h3a5bdd8b),
	.w8(32'h3bbc0d7e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901f065),
	.w1(32'hb8f7ad42),
	.w2(32'hb8cd7138),
	.w3(32'hb99516b7),
	.w4(32'hb9aee6f2),
	.w5(32'hb942239a),
	.w6(32'hb9a10e3f),
	.w7(32'hb9823177),
	.w8(32'hb827111d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4a86e),
	.w1(32'hb88e0b76),
	.w2(32'hb929e040),
	.w3(32'hb9d73066),
	.w4(32'h367e36d7),
	.w5(32'hb909a8f3),
	.w6(32'hb9ebb9fe),
	.w7(32'hb87f89d0),
	.w8(32'hb98e2f89),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c15b),
	.w1(32'hbb994470),
	.w2(32'h3b205b6d),
	.w3(32'hbb16dc71),
	.w4(32'hbbef7bb9),
	.w5(32'h36f47c84),
	.w6(32'hbaae3bdd),
	.w7(32'hbbe9e19b),
	.w8(32'h38922466),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1be62e),
	.w1(32'h3ad27474),
	.w2(32'h3c3add30),
	.w3(32'h3cd9b788),
	.w4(32'h3aeda5c5),
	.w5(32'h3c3428d0),
	.w6(32'h3ca098b4),
	.w7(32'hbb395b37),
	.w8(32'h3c5bd33f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f3a4f),
	.w1(32'h398d5732),
	.w2(32'h3c3f7800),
	.w3(32'h3c60dfc5),
	.w4(32'hbc06bc57),
	.w5(32'h3ac7896c),
	.w6(32'h3c48c467),
	.w7(32'hbc0ac61a),
	.w8(32'h3addc86a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceac77c),
	.w1(32'h3ad7be9c),
	.w2(32'h3c4ba4ae),
	.w3(32'h3cc1f7d4),
	.w4(32'hbbbca803),
	.w5(32'h3b4bf228),
	.w6(32'h3cb2d75f),
	.w7(32'hbc2e9846),
	.w8(32'h39b0637a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8482ffc),
	.w1(32'hb904f471),
	.w2(32'h3a1230d3),
	.w3(32'h3875ad0a),
	.w4(32'hb95c5a5d),
	.w5(32'h3a04e2e7),
	.w6(32'h37d7ce24),
	.w7(32'hb94a8615),
	.w8(32'hb8e28863),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55ab8b),
	.w1(32'hb9c33e60),
	.w2(32'hba0c3204),
	.w3(32'hba31c6a4),
	.w4(32'hb97c05c8),
	.w5(32'hb9ea793e),
	.w6(32'hba2457d2),
	.w7(32'hb9ba96ca),
	.w8(32'hba21681e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a345f0d),
	.w1(32'hbb70da47),
	.w2(32'h3c0d539a),
	.w3(32'h3a0ee549),
	.w4(32'hbbcb82b8),
	.w5(32'hbbc122b7),
	.w6(32'h3a58773a),
	.w7(32'hbba51700),
	.w8(32'hbb244b4d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae18550),
	.w1(32'hbb5d06bb),
	.w2(32'h3a809d83),
	.w3(32'h3a2880fd),
	.w4(32'hbb8a6c9b),
	.w5(32'h3a0fcffb),
	.w6(32'h3b7647fd),
	.w7(32'hbb5994d7),
	.w8(32'h3a41591c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05bad0),
	.w1(32'hbba67c39),
	.w2(32'h3c01b1e2),
	.w3(32'h3c011976),
	.w4(32'hbc0854c9),
	.w5(32'hba5d0be5),
	.w6(32'h3c109e3a),
	.w7(32'hbc094e2d),
	.w8(32'hba6af897),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9169615),
	.w1(32'hb8d893b8),
	.w2(32'hb8b73111),
	.w3(32'hb9109376),
	.w4(32'hb8d75ba8),
	.w5(32'hb8d0260d),
	.w6(32'hb9254ecb),
	.w7(32'hb9144704),
	.w8(32'hb8e8cc30),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38591255),
	.w1(32'hb70285ec),
	.w2(32'hb8f39984),
	.w3(32'hb856a4e8),
	.w4(32'hb91c9fd7),
	.w5(32'hb9a1fbe0),
	.w6(32'hb97ebc41),
	.w7(32'hb987e9e1),
	.w8(32'hb9c07958),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb4322),
	.w1(32'hba4809b6),
	.w2(32'h3b982dbd),
	.w3(32'h3b6ce738),
	.w4(32'hbb8d56d6),
	.w5(32'h37c6c413),
	.w6(32'h3b52abc0),
	.w7(32'hbb6bd6b6),
	.w8(32'hb853fade),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c14a9),
	.w1(32'hb9432cdd),
	.w2(32'h3a82e35e),
	.w3(32'h3c043b05),
	.w4(32'hba7a1ff1),
	.w5(32'hb926227c),
	.w6(32'h3bea72a2),
	.w7(32'hba9bb143),
	.w8(32'hb8021ab7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d0316),
	.w1(32'h3a4c4453),
	.w2(32'h3a1bb33c),
	.w3(32'h3949c4d2),
	.w4(32'h39de8f4d),
	.w5(32'hb90804f2),
	.w6(32'h39f0c691),
	.w7(32'h3a86e885),
	.w8(32'h3ab2ad63),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed8c0f),
	.w1(32'h3b1d81a3),
	.w2(32'h3b953f0e),
	.w3(32'h3abdec29),
	.w4(32'h3b8be55a),
	.w5(32'h3bc8f60c),
	.w6(32'hbb03edc0),
	.w7(32'h395be107),
	.w8(32'h3b2e6bb1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9db0a1),
	.w1(32'hbaad5da1),
	.w2(32'h3ba041f9),
	.w3(32'h3c0fe119),
	.w4(32'hbbdad787),
	.w5(32'hbadfde7a),
	.w6(32'hbb1a4ac0),
	.w7(32'hbc76759a),
	.w8(32'hba9e910d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1de92d),
	.w1(32'hbb876f96),
	.w2(32'h3c1f5638),
	.w3(32'h3ce4a058),
	.w4(32'hbc998d5a),
	.w5(32'hbb91ca74),
	.w6(32'h3cd13213),
	.w7(32'hbc9c2138),
	.w8(32'hbaa66683),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb538a5),
	.w1(32'hbc1431bd),
	.w2(32'h3bcfb53d),
	.w3(32'h3ca15391),
	.w4(32'hbc8c924b),
	.w5(32'hba4ddb32),
	.w6(32'h3cbe0bfd),
	.w7(32'hbc7e1af8),
	.w8(32'h3bb5ac25),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb3d79),
	.w1(32'h39e5c7e1),
	.w2(32'h3a4fd0b3),
	.w3(32'h3b9c2a41),
	.w4(32'hbb117aa8),
	.w5(32'hbad71dcc),
	.w6(32'h3b8258a7),
	.w7(32'hbb2909c1),
	.w8(32'hba340cfd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907f59e),
	.w1(32'h3900bbdc),
	.w2(32'hb90f5a37),
	.w3(32'hb879ed32),
	.w4(32'h3998e9e7),
	.w5(32'hb65929c3),
	.w6(32'hb99df1d5),
	.w7(32'h396adb9c),
	.w8(32'hb8ee3533),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d9ed2),
	.w1(32'hb9d0e292),
	.w2(32'hba121f5b),
	.w3(32'hba85dc65),
	.w4(32'hb98992df),
	.w5(32'hb9c81921),
	.w6(32'hba63c9fe),
	.w7(32'hb9abe2e0),
	.w8(32'hb9cbc47f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d794),
	.w1(32'hbb6301bd),
	.w2(32'hba262bf8),
	.w3(32'h3b19b73d),
	.w4(32'hbb850a2a),
	.w5(32'hba188185),
	.w6(32'h3b1a4c8d),
	.w7(32'hbac9adea),
	.w8(32'h3ab0aa59),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca63067),
	.w1(32'h3b013fae),
	.w2(32'h3c6eb699),
	.w3(32'h3c92cb5b),
	.w4(32'h3b3c78de),
	.w5(32'h3bf96b32),
	.w6(32'h3c9d25cb),
	.w7(32'h3c0fb458),
	.w8(32'h3c1ce91e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94556e),
	.w1(32'hbb4cdb7f),
	.w2(32'h3c174e18),
	.w3(32'h3c4cecf8),
	.w4(32'hbc316a37),
	.w5(32'hbaab2583),
	.w6(32'h3c42b518),
	.w7(32'hbc3f0d48),
	.w8(32'hbb2ca360),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbddfdc),
	.w1(32'h39a88b39),
	.w2(32'h3c3bf735),
	.w3(32'h3c85d94a),
	.w4(32'hbc063c10),
	.w5(32'h3979e1cd),
	.w6(32'h3c5175f8),
	.w7(32'hbc180152),
	.w8(32'hb99aa647),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8d7f1),
	.w1(32'h39a31770),
	.w2(32'h3bab297b),
	.w3(32'h3c91349a),
	.w4(32'hbb055ea3),
	.w5(32'h3913edef),
	.w6(32'h3c462857),
	.w7(32'hbbb899b4),
	.w8(32'hba15b959),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c204bca),
	.w1(32'h3c5bbabc),
	.w2(32'h3cb66b1b),
	.w3(32'h3c3e35c1),
	.w4(32'h3c6328b9),
	.w5(32'h3ca11ca4),
	.w6(32'hbb2f077d),
	.w7(32'h39f2c282),
	.w8(32'h3bc13686),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90cc70b),
	.w1(32'hb8f8efcb),
	.w2(32'h3939e87e),
	.w3(32'hba3959d2),
	.w4(32'hb96a0679),
	.w5(32'h3984dd31),
	.w6(32'hb9bb943e),
	.w7(32'hb8bf32a1),
	.w8(32'h3981daca),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8d424),
	.w1(32'hb93131be),
	.w2(32'hbb02b6cf),
	.w3(32'h3aaa2f16),
	.w4(32'h3a8aa8b9),
	.w5(32'h39a2b22e),
	.w6(32'h3ae2322e),
	.w7(32'h3af1b66e),
	.w8(32'h3b0b55c6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9badbcb),
	.w1(32'h39cc6dfa),
	.w2(32'h3a5b79a8),
	.w3(32'hba3040d9),
	.w4(32'h39a736d2),
	.w5(32'h3a88d149),
	.w6(32'hba04dc80),
	.w7(32'h39a845c0),
	.w8(32'h3a85c3c5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46f4f6),
	.w1(32'h3b27decc),
	.w2(32'h3c1adbda),
	.w3(32'h3c2326e5),
	.w4(32'h37fcdc75),
	.w5(32'h3b90a94a),
	.w6(32'h3bc040a4),
	.w7(32'hbb1bc2ce),
	.w8(32'h3afa18ad),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5971cf),
	.w1(32'h3a6a52c7),
	.w2(32'h3b18a250),
	.w3(32'h3b44f57f),
	.w4(32'h3a5dfea1),
	.w5(32'h3b2209a6),
	.w6(32'h3b03bbc1),
	.w7(32'hb9a52752),
	.w8(32'h3a8df81d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c883ee2),
	.w1(32'h3bb8d55b),
	.w2(32'h3c6342ea),
	.w3(32'h3c605d33),
	.w4(32'h3b80cd4f),
	.w5(32'h3c0d220f),
	.w6(32'h3bd70a13),
	.w7(32'hbab07251),
	.w8(32'h3b4e849f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0ec1),
	.w1(32'hba4cd9c7),
	.w2(32'h39fabbfa),
	.w3(32'h3b552e02),
	.w4(32'h3a9d618c),
	.w5(32'h3aea1dc0),
	.w6(32'h3b1836c5),
	.w7(32'hba7c79d3),
	.w8(32'hb97974c1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe1cd8),
	.w1(32'h39bc86df),
	.w2(32'h39d3f2a6),
	.w3(32'h395e6f43),
	.w4(32'hb6e23b81),
	.w5(32'hb80a7234),
	.w6(32'h390b371d),
	.w7(32'hb9865f83),
	.w8(32'hb99e698a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8643499),
	.w1(32'hb78ff30a),
	.w2(32'hb7d45397),
	.w3(32'hb85c630a),
	.w4(32'hb5ab2177),
	.w5(32'hb7b72a29),
	.w6(32'hb89812bd),
	.w7(32'hb858c2a8),
	.w8(32'hb81bdc4f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921e931),
	.w1(32'hb9d61955),
	.w2(32'h3a310683),
	.w3(32'h37e874a9),
	.w4(32'hb9f33bf4),
	.w5(32'h39a2d98e),
	.w6(32'h38e1abfa),
	.w7(32'hba12227f),
	.w8(32'h39d2d411),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f3570),
	.w1(32'hbb3de863),
	.w2(32'hb9240d81),
	.w3(32'hb8f1610c),
	.w4(32'hbb5b8044),
	.w5(32'hba0421c0),
	.w6(32'h3ad6160e),
	.w7(32'hbb03536e),
	.w8(32'h38caa128),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac59a2f),
	.w1(32'hb8833c03),
	.w2(32'h3a723649),
	.w3(32'h37f57c28),
	.w4(32'hba9ba37d),
	.w5(32'hb98d9f14),
	.w6(32'h3a676caa),
	.w7(32'hb9f056a1),
	.w8(32'h3a61a97c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4532be),
	.w1(32'h3b9146e4),
	.w2(32'h3bda3ad0),
	.w3(32'h3c2e612b),
	.w4(32'h3ba57c43),
	.w5(32'h3bb0c6e4),
	.w6(32'h3bed4403),
	.w7(32'h3b290c83),
	.w8(32'h3b1c1e56),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25d580),
	.w1(32'h3b27db0c),
	.w2(32'h3b94af0d),
	.w3(32'h3c2360c3),
	.w4(32'h3bbc02a8),
	.w5(32'h3b1002cb),
	.w6(32'h3c07998a),
	.w7(32'h3ba70ad4),
	.w8(32'h3ba7a2ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb946ec19),
	.w1(32'hb7b57436),
	.w2(32'hb9267dbb),
	.w3(32'hb91eac63),
	.w4(32'h383f099e),
	.w5(32'hb8b169bc),
	.w6(32'hb9678b0c),
	.w7(32'h373069cb),
	.w8(32'hb8f7360d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954a36a),
	.w1(32'hb82df84e),
	.w2(32'hb9071a3c),
	.w3(32'hb9171e18),
	.w4(32'h380d0327),
	.w5(32'hb887a31d),
	.w6(32'hb943c0c0),
	.w7(32'hb7bf648c),
	.w8(32'hb909d71c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983127f),
	.w1(32'hb852d293),
	.w2(32'h386a0eca),
	.w3(32'hb9eff71f),
	.w4(32'hb9e55a99),
	.w5(32'hb9db44bf),
	.w6(32'hb9dd9f8e),
	.w7(32'hb9e3f543),
	.w8(32'hb9e22457),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f258a9),
	.w1(32'hb93c7003),
	.w2(32'hb988da77),
	.w3(32'hb9cad1a8),
	.w4(32'hb8b5ff3d),
	.w5(32'hb92e1bcb),
	.w6(32'hb9ceeb48),
	.w7(32'hb8fdf7f6),
	.w8(32'hb97d40c6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cf00b),
	.w1(32'h3c2b2e04),
	.w2(32'h3c6f0cf0),
	.w3(32'h3c697c32),
	.w4(32'h3c2a37bd),
	.w5(32'h3aabfdd0),
	.w6(32'h3c0a1ba9),
	.w7(32'h3bbc60a7),
	.w8(32'h3bcd8f64),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1dd7e),
	.w1(32'h3b068d60),
	.w2(32'h3c60af4a),
	.w3(32'h3c8dc4fa),
	.w4(32'hbaf6322c),
	.w5(32'h3c2325e3),
	.w6(32'h3c607474),
	.w7(32'hbbe1663c),
	.w8(32'h3bb7f32e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caebb9a),
	.w1(32'hba9f0ee4),
	.w2(32'h3c24f98b),
	.w3(32'h3ca14ea2),
	.w4(32'hbb43d1a6),
	.w5(32'h3bff9d5d),
	.w6(32'h3c90eba8),
	.w7(32'hbb7967a0),
	.w8(32'h3c02e277),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d043187),
	.w1(32'hbc0af031),
	.w2(32'h3c828b31),
	.w3(32'h3cce2ce2),
	.w4(32'hbc97662c),
	.w5(32'h3a831fa2),
	.w6(32'h3cd9fdcc),
	.w7(32'hbcb98a49),
	.w8(32'h3ac66b5c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa32b7),
	.w1(32'hb82d5f24),
	.w2(32'hb9664bf0),
	.w3(32'hb9d25150),
	.w4(32'h38641500),
	.w5(32'hb8c6ee4b),
	.w6(32'hb9e6b4d2),
	.w7(32'hb78d9913),
	.w8(32'hb94f8c97),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba478fad),
	.w1(32'hb91f7fc0),
	.w2(32'hb9ef023c),
	.w3(32'hba247f10),
	.w4(32'hb76c7d18),
	.w5(32'hb9aa9ea7),
	.w6(32'hba349e19),
	.w7(32'hb91b1684),
	.w8(32'hb9f6a9ad),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fc57e),
	.w1(32'hb6c9ff1c),
	.w2(32'hb93e9a02),
	.w3(32'hba3c1f79),
	.w4(32'h38e3c74b),
	.w5(32'hb90a3027),
	.w6(32'hba3fd86c),
	.w7(32'h38397bd2),
	.w8(32'hb98452b4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b451eb4),
	.w1(32'h39787277),
	.w2(32'h3ae0a896),
	.w3(32'h3b4f83a0),
	.w4(32'h3aae095d),
	.w5(32'h3b1d562c),
	.w6(32'h3adbace2),
	.w7(32'h39e15fa5),
	.w8(32'h3a9ff95f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22a77d),
	.w1(32'hb8b68ad2),
	.w2(32'hb95ffef4),
	.w3(32'hba0b696e),
	.w4(32'hb785600b),
	.w5(32'hb9109856),
	.w6(32'hba1cb539),
	.w7(32'hb892a1ca),
	.w8(32'hb92a8cb0),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd31ade),
	.w1(32'h3b8d9dbe),
	.w2(32'h3b1d1a31),
	.w3(32'h3bdd6bcc),
	.w4(32'h3c0194f1),
	.w5(32'h3b5c1467),
	.w6(32'hb9380b0c),
	.w7(32'h3a1af8d9),
	.w8(32'hb9b703f9),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c652e43),
	.w1(32'h3b4b8305),
	.w2(32'h3c0400fa),
	.w3(32'h3c30f3f0),
	.w4(32'h3b5e9ff4),
	.w5(32'h3be151ef),
	.w6(32'h3c071dce),
	.w7(32'h3b2ec98f),
	.w8(32'h3b1a9730),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c821241),
	.w1(32'h3b98aad5),
	.w2(32'h3c3f9ce2),
	.w3(32'h3c57efcd),
	.w4(32'hbb07aad6),
	.w5(32'h3b208917),
	.w6(32'h3bce2004),
	.w7(32'hbbf06ab7),
	.w8(32'hba8f46fa),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c094b77),
	.w1(32'h3b17da76),
	.w2(32'h3c02a9de),
	.w3(32'h3be215e4),
	.w4(32'h399b355f),
	.w5(32'h3b87efda),
	.w6(32'h3be073b1),
	.w7(32'hba143bf8),
	.w8(32'h3b65865d),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1a507),
	.w1(32'h3a7e747c),
	.w2(32'h3bd2917b),
	.w3(32'h3ae2f4b6),
	.w4(32'h3a1e4889),
	.w5(32'h3ad96e43),
	.w6(32'hba802160),
	.w7(32'hbaaae750),
	.w8(32'h3b54dc8c),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d8bf),
	.w1(32'h397bf2a9),
	.w2(32'h3b797a46),
	.w3(32'h3bd1753e),
	.w4(32'hbab6fb38),
	.w5(32'hb6b0769d),
	.w6(32'h3bd43eef),
	.w7(32'hba9ab806),
	.w8(32'hb9de13bf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b819476),
	.w1(32'h3b237c7f),
	.w2(32'h3bdde620),
	.w3(32'h3b6d3ed8),
	.w4(32'h3b39ce6b),
	.w5(32'h3be8bc8a),
	.w6(32'hba333c00),
	.w7(32'hbb001efc),
	.w8(32'h3b17babb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fbae9),
	.w1(32'h3677db44),
	.w2(32'hb7a647d0),
	.w3(32'hb87def30),
	.w4(32'h36a60106),
	.w5(32'hb814deea),
	.w6(32'hb8a16fce),
	.w7(32'hb6c24a80),
	.w8(32'hb886a6d3),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85c9010),
	.w1(32'hb8367707),
	.w2(32'hb8b8d54c),
	.w3(32'hb8539778),
	.w4(32'hb83c77a9),
	.w5(32'hb8c599ac),
	.w6(32'hb6a12643),
	.w7(32'h37d1a652),
	.w8(32'hb81e1862),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95bbd30),
	.w1(32'hb991459f),
	.w2(32'hb9d85be8),
	.w3(32'h3986bd74),
	.w4(32'hb73420bc),
	.w5(32'hb944baab),
	.w6(32'hb8f4f865),
	.w7(32'hb904f9bd),
	.w8(32'hb6aea38a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c795f),
	.w1(32'hb8cd015a),
	.w2(32'h375330a0),
	.w3(32'h388c2489),
	.w4(32'hb9df72ab),
	.w5(32'hb9df78d5),
	.w6(32'hb930c6af),
	.w7(32'hba3d2a0f),
	.w8(32'hb9b14c52),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91a6d3),
	.w1(32'hbb003287),
	.w2(32'hbb7f30b3),
	.w3(32'h3c81e8f6),
	.w4(32'hbb8fe7e5),
	.w5(32'hbbd521bb),
	.w6(32'h3c4273ec),
	.w7(32'hbc369edc),
	.w8(32'hbbe988d0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01bd16),
	.w1(32'hba91a354),
	.w2(32'hba4998b8),
	.w3(32'hba9d9ae6),
	.w4(32'hbb0fbc0f),
	.w5(32'hbab90c36),
	.w6(32'h3a05d403),
	.w7(32'hbaa8d97e),
	.w8(32'hba4fd679),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dfb23),
	.w1(32'h3b10eaea),
	.w2(32'h3bada9d0),
	.w3(32'h3bdbc294),
	.w4(32'hbb3f1222),
	.w5(32'h3a60d262),
	.w6(32'h3b9c9f4f),
	.w7(32'hbb29b9ed),
	.w8(32'hb894a129),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b28bf),
	.w1(32'h3b391563),
	.w2(32'h3c03e7ec),
	.w3(32'h3c906804),
	.w4(32'h3bec53f1),
	.w5(32'h3c2963fa),
	.w6(32'h3c39d11a),
	.w7(32'h3b291082),
	.w8(32'h3bb4b9ad),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07f182),
	.w1(32'hbb7e83b9),
	.w2(32'h3b7ee2ae),
	.w3(32'h3c012db0),
	.w4(32'hbbc7048c),
	.w5(32'hbae8cc75),
	.w6(32'h3b77a940),
	.w7(32'hbc1652ca),
	.w8(32'hbae4d4ff),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a94bc),
	.w1(32'h3c08cf3d),
	.w2(32'h3c406231),
	.w3(32'h3c1dceeb),
	.w4(32'h3a81aa7b),
	.w5(32'h3b95d96c),
	.w6(32'h3a89d69c),
	.w7(32'hba1308a9),
	.w8(32'h3b7b9a04),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc27920),
	.w1(32'hbb8ee196),
	.w2(32'h3acc17ad),
	.w3(32'h3b91b44a),
	.w4(32'hbbdf1a18),
	.w5(32'hbb2a00ac),
	.w6(32'h3b01ce89),
	.w7(32'hbc160781),
	.w8(32'hbb873e0b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2fe5e),
	.w1(32'h3bdb9585),
	.w2(32'h3c39f3ee),
	.w3(32'h3ca9fbbc),
	.w4(32'h3bb1b001),
	.w5(32'h3bb45841),
	.w6(32'h3c9cf750),
	.w7(32'h3b0083b6),
	.w8(32'h3b92679b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c619b52),
	.w1(32'h3ac4e298),
	.w2(32'h3b3ea5f5),
	.w3(32'h3c4350ad),
	.w4(32'hbae04221),
	.w5(32'hbb82b62a),
	.w6(32'h3be6ab10),
	.w7(32'hbb74b9fe),
	.w8(32'hbb2cdc0a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b15f8),
	.w1(32'h38e64cc4),
	.w2(32'h3be6d422),
	.w3(32'h3c67fe6a),
	.w4(32'hbbe1cf6a),
	.w5(32'hbad9b459),
	.w6(32'h3c1c0f43),
	.w7(32'hbc241039),
	.w8(32'hbb55cf14),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8971c28),
	.w1(32'hb99bc074),
	.w2(32'hba249636),
	.w3(32'hba673b34),
	.w4(32'hba1b7347),
	.w5(32'hb901a9a5),
	.w6(32'hba75000a),
	.w7(32'hba3b6aeb),
	.w8(32'hba66b567),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7cde4d),
	.w1(32'h3aee43bf),
	.w2(32'h3c3a2d8f),
	.w3(32'h3c3df4df),
	.w4(32'hbaac27fc),
	.w5(32'h3bab0691),
	.w6(32'h3c44678b),
	.w7(32'hb9207a5a),
	.w8(32'h3bb439a7),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c64ef29),
	.w1(32'h3aabb975),
	.w2(32'h3bdbfeae),
	.w3(32'h3c599dc0),
	.w4(32'h3ac294f0),
	.w5(32'h3bb1f640),
	.w6(32'h3bc5bf02),
	.w7(32'h3a38c7c1),
	.w8(32'h3c1ea3c3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93dc26),
	.w1(32'h3adc2ce4),
	.w2(32'h3c04b065),
	.w3(32'h3c1a3ae4),
	.w4(32'hbb0241da),
	.w5(32'h3bbd7029),
	.w6(32'hbae54049),
	.w7(32'hbc30e506),
	.w8(32'h3a8f3e86),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1076b3),
	.w1(32'hbbbe8e18),
	.w2(32'hbba5556b),
	.w3(32'h3cddf0a5),
	.w4(32'hbc8d8c9b),
	.w5(32'hbc18cbed),
	.w6(32'h3c940b57),
	.w7(32'hbc679d60),
	.w8(32'hbbb4fda2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c709969),
	.w1(32'hb9c140dc),
	.w2(32'h3c5971be),
	.w3(32'h3c4165a6),
	.w4(32'hbbb25528),
	.w5(32'h3bb9ef10),
	.w6(32'h3c2d588d),
	.w7(32'hbbe06666),
	.w8(32'h3acd71d8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c693de6),
	.w1(32'h3c211fdc),
	.w2(32'h3c398b2a),
	.w3(32'h3c16e4b1),
	.w4(32'h3c119e1a),
	.w5(32'h3bc9005f),
	.w6(32'hbba190e2),
	.w7(32'hbbb15812),
	.w8(32'h3b95af3b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981df41),
	.w1(32'hba5063f6),
	.w2(32'hba9dea3e),
	.w3(32'hbab06c46),
	.w4(32'hbac1790b),
	.w5(32'h38e98305),
	.w6(32'hba89064e),
	.w7(32'hbb3781c4),
	.w8(32'hbb3351ce),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8be19),
	.w1(32'h3c4d7a28),
	.w2(32'h3ba4fa0c),
	.w3(32'h3c7ee082),
	.w4(32'h3bb5067e),
	.w5(32'h3ad865d3),
	.w6(32'hbbba343c),
	.w7(32'hbc7f2a23),
	.w8(32'hbc102722),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d039e),
	.w1(32'hbb9d3ec5),
	.w2(32'hba1920b1),
	.w3(32'h3b8ab5b0),
	.w4(32'hba8aa2a9),
	.w5(32'h3b0b6f1c),
	.w6(32'h3b140fc9),
	.w7(32'hba600db8),
	.w8(32'h3b66e69e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cf8d9),
	.w1(32'hb95c4707),
	.w2(32'h3a4a2e59),
	.w3(32'h37818419),
	.w4(32'hba275187),
	.w5(32'h3a09f9fb),
	.w6(32'hb9969547),
	.w7(32'hba82f11a),
	.w8(32'h398af568),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76c6c),
	.w1(32'h3b11d1ac),
	.w2(32'h3b49cab4),
	.w3(32'h3b33d287),
	.w4(32'hb998a186),
	.w5(32'hb9447100),
	.w6(32'h3b386cc3),
	.w7(32'hba436e71),
	.w8(32'hb82369a4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf0005),
	.w1(32'h3b3b0e5a),
	.w2(32'h3c3f399e),
	.w3(32'h3ba314ff),
	.w4(32'h3b4e08bd),
	.w5(32'h3c0e3bd4),
	.w6(32'h3b93bb84),
	.w7(32'h3b6ba59f),
	.w8(32'h3c07d758),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6c7f0),
	.w1(32'hbaf3c7e0),
	.w2(32'h3bf7bbd5),
	.w3(32'h3bf9c95d),
	.w4(32'hbb901047),
	.w5(32'h3b1004b7),
	.w6(32'h3be2da00),
	.w7(32'hbbdc4425),
	.w8(32'hb97a960d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbaf26),
	.w1(32'hba631099),
	.w2(32'h3a81a1e2),
	.w3(32'h3c0c5067),
	.w4(32'hbb4b5395),
	.w5(32'hba8479ca),
	.w6(32'h3bf04ed8),
	.w7(32'hbb8acf47),
	.w8(32'hbac8224a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38f7c8),
	.w1(32'h3b300d05),
	.w2(32'h3b935fe6),
	.w3(32'h3bfa8c5e),
	.w4(32'hba8f31f1),
	.w5(32'h3abea2c6),
	.w6(32'h3bcd505c),
	.w7(32'hbb2a369e),
	.w8(32'h3acc5d8f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3c926),
	.w1(32'hbb473070),
	.w2(32'h3ad4bbf8),
	.w3(32'h3be49053),
	.w4(32'hbb3e217b),
	.w5(32'h3b34b1b9),
	.w6(32'h3b885abf),
	.w7(32'hbbed30fb),
	.w8(32'hba20724c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c316209),
	.w1(32'h3b2b8884),
	.w2(32'h3c00f5c1),
	.w3(32'h3be33102),
	.w4(32'hbace4df4),
	.w5(32'hb95c5cad),
	.w6(32'h3bbcf88b),
	.w7(32'hb8b9e669),
	.w8(32'h3b1d7c94),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0293e3),
	.w1(32'hb925fc37),
	.w2(32'h3b68af50),
	.w3(32'h3bef6f61),
	.w4(32'hbacda9b0),
	.w5(32'h3aed5579),
	.w6(32'h3bd650fc),
	.w7(32'hbb23fa97),
	.w8(32'h3a99b77a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399447af),
	.w1(32'h39862a7b),
	.w2(32'h3902042b),
	.w3(32'h3984ebfc),
	.w4(32'h39867e78),
	.w5(32'h38a1023b),
	.w6(32'h39328ee6),
	.w7(32'h38a97430),
	.w8(32'hb8fa1261),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac498f3),
	.w1(32'h3a6b1538),
	.w2(32'h398fb139),
	.w3(32'h3a87f10b),
	.w4(32'h3934f48b),
	.w5(32'hb9f75e94),
	.w6(32'h3a47ab9c),
	.w7(32'hb94a6ce0),
	.w8(32'hb983d349),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37066005),
	.w1(32'hb996c083),
	.w2(32'hb9850518),
	.w3(32'h397ae584),
	.w4(32'hb95a3228),
	.w5(32'hb974d627),
	.w6(32'h38f7b590),
	.w7(32'hb932f765),
	.w8(32'hb9470812),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f53e65),
	.w1(32'hba549526),
	.w2(32'h3909701e),
	.w3(32'h3905132b),
	.w4(32'hbaa3e105),
	.w5(32'hba3446a9),
	.w6(32'h395f80f6),
	.w7(32'hba8b52d4),
	.w8(32'hbaa922e7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155c1c),
	.w1(32'hbb938f40),
	.w2(32'h3ae51f1b),
	.w3(32'h3bda25b2),
	.w4(32'hbbf65052),
	.w5(32'hbb07cd83),
	.w6(32'h3be77f8d),
	.w7(32'hbbced5dd),
	.w8(32'hbaf5622b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0309ef),
	.w1(32'h3ad5a6f8),
	.w2(32'h3b43fa17),
	.w3(32'h3a48a13c),
	.w4(32'hba24b3cb),
	.w5(32'h3a99bad7),
	.w6(32'h39308237),
	.w7(32'hbab66358),
	.w8(32'h3980b3dd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19de8c),
	.w1(32'h3a9b684e),
	.w2(32'h3b9c6dd1),
	.w3(32'h3b226266),
	.w4(32'h3b62f2f0),
	.w5(32'h3b72dadc),
	.w6(32'hbb7850ca),
	.w7(32'hbb10bcd0),
	.w8(32'hb818f2b5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8673e),
	.w1(32'h3b4ff18f),
	.w2(32'h3c171046),
	.w3(32'h3c6d8275),
	.w4(32'hbb7897c0),
	.w5(32'h3b0db26d),
	.w6(32'h3c2ee392),
	.w7(32'hbbb576b1),
	.w8(32'h3b4846dd),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f2e035),
	.w1(32'hb96cfe0d),
	.w2(32'hb8d2fe73),
	.w3(32'hba0350ae),
	.w4(32'hb9a9dbb0),
	.w5(32'hb9751703),
	.w6(32'hba1dff1f),
	.w7(32'hb9e019cd),
	.w8(32'hb9afd4f2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0467a1),
	.w1(32'h383c4a29),
	.w2(32'h3a5f2d97),
	.w3(32'hba2d8124),
	.w4(32'hb9eaf5ec),
	.w5(32'h39c0c90b),
	.w6(32'hb90c8969),
	.w7(32'h37aeac0c),
	.w8(32'h3a2f9d69),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d6ee5),
	.w1(32'hb9025a69),
	.w2(32'hb84cd0ed),
	.w3(32'hb91deaaf),
	.w4(32'hb915077e),
	.w5(32'hb8a15716),
	.w6(32'hb93cf3cc),
	.w7(32'hb9146231),
	.w8(32'hb85fb39b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0e49f),
	.w1(32'h39a56f8f),
	.w2(32'h3a79beb3),
	.w3(32'h3af45bea),
	.w4(32'hb93982be),
	.w5(32'h38ff155a),
	.w6(32'h3afd00aa),
	.w7(32'h3a4241f3),
	.w8(32'h3aa6282c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e00ee),
	.w1(32'h3ba90d56),
	.w2(32'h3c0882af),
	.w3(32'h3b85b6cd),
	.w4(32'h3bdf63a4),
	.w5(32'h3c4de9a3),
	.w6(32'h3a6752ad),
	.w7(32'h3adcc571),
	.w8(32'h3bebc8ee),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01b98f),
	.w1(32'hb9c4af7f),
	.w2(32'h3bff7fb3),
	.w3(32'h3bbe9913),
	.w4(32'hbb5f19eb),
	.w5(32'h3b291307),
	.w6(32'h3bae70e1),
	.w7(32'hba9acf5d),
	.w8(32'h3b8b60cf),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adad61c),
	.w1(32'h3afba0fd),
	.w2(32'h3a9165e8),
	.w3(32'h3a4bb36c),
	.w4(32'h3abfa951),
	.w5(32'h39aa52db),
	.w6(32'hba7bb3e0),
	.w7(32'hb98a0d92),
	.w8(32'h38ecd1d6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68a45a),
	.w1(32'h3a814788),
	.w2(32'h3afb6a2a),
	.w3(32'h3b9b1d6d),
	.w4(32'h3ae05127),
	.w5(32'h3b2b679c),
	.w6(32'h3b989caa),
	.w7(32'h3a02352c),
	.w8(32'h3b09d984),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5a6e),
	.w1(32'h3a40864d),
	.w2(32'h3b2d6be7),
	.w3(32'h3ba530d4),
	.w4(32'hba992418),
	.w5(32'h3a1f144d),
	.w6(32'h3b1e4fc1),
	.w7(32'hbb40327e),
	.w8(32'hb92124f1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2d099),
	.w1(32'h3a65d98e),
	.w2(32'h3b81dd8d),
	.w3(32'h3b991d0a),
	.w4(32'h39cb575f),
	.w5(32'h3aedc603),
	.w6(32'h3bbc2624),
	.w7(32'h39fff28c),
	.w8(32'h3a8f2c60),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c716591),
	.w1(32'h3b3300fc),
	.w2(32'h3bbfe4bf),
	.w3(32'h3c287732),
	.w4(32'hbb70cfc2),
	.w5(32'hbb539a1b),
	.w6(32'h3bf3ec64),
	.w7(32'hbb99e6e8),
	.w8(32'hbb6bfdcb),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3aa548),
	.w1(32'h3bc92024),
	.w2(32'h3c2f1771),
	.w3(32'h3c1bb507),
	.w4(32'h3b696e85),
	.w5(32'h3bfc5a70),
	.w6(32'h3b584201),
	.w7(32'h3a7b8b18),
	.w8(32'h3b948e79),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cbf91),
	.w1(32'hba5b0754),
	.w2(32'h3b7d7a5a),
	.w3(32'h3c171a15),
	.w4(32'hbb6df2a0),
	.w5(32'hba839964),
	.w6(32'h3bfc7863),
	.w7(32'hbbaf463e),
	.w8(32'h399cd5c8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a1793),
	.w1(32'h3b311fa5),
	.w2(32'h3b815f34),
	.w3(32'h3c0202c3),
	.w4(32'hba87a2be),
	.w5(32'hb90d71d9),
	.w6(32'h3bad4799),
	.w7(32'h38844743),
	.w8(32'h3b034416),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c516fec),
	.w1(32'h3b302d01),
	.w2(32'h3c1c5ada),
	.w3(32'h3c20c277),
	.w4(32'h3b9c7397),
	.w5(32'h3c0eb5e5),
	.w6(32'h3b005c22),
	.w7(32'hbb94a73e),
	.w8(32'h3a111c61),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46eaf3),
	.w1(32'h3b19b012),
	.w2(32'h3b0fc9cb),
	.w3(32'h3c0cd455),
	.w4(32'hbaf38e5f),
	.w5(32'hbb161d32),
	.w6(32'h3c03da07),
	.w7(32'hbb8ad467),
	.w8(32'hbb075116),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bded2ab),
	.w1(32'h3aafa8fe),
	.w2(32'h3bb093e1),
	.w3(32'h3b96f6b0),
	.w4(32'hba3e156f),
	.w5(32'h3aecd9fe),
	.w6(32'h3b9e0080),
	.w7(32'h3b078893),
	.w8(32'h3b812861),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69458b),
	.w1(32'h39caf178),
	.w2(32'h3b115f69),
	.w3(32'h3b1a1676),
	.w4(32'hba9ca571),
	.w5(32'h38c48b8c),
	.w6(32'h3b141f4f),
	.w7(32'hbab8dbbf),
	.w8(32'hb8130cb8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c593584),
	.w1(32'hbbd4a51a),
	.w2(32'h3bb5cc52),
	.w3(32'h3c7e6e47),
	.w4(32'hbbce2108),
	.w5(32'h3b78e541),
	.w6(32'h3c20b0c2),
	.w7(32'hbc4297c5),
	.w8(32'h3a955e33),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e4693),
	.w1(32'hba903cc7),
	.w2(32'hbb9c7b8f),
	.w3(32'h3c04c2a1),
	.w4(32'hbb318f2a),
	.w5(32'hbbac2311),
	.w6(32'h3be92cc0),
	.w7(32'hbba025bc),
	.w8(32'hbba2ba1b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35954daf),
	.w1(32'hb7a4fcba),
	.w2(32'hb7b510a8),
	.w3(32'h392ef453),
	.w4(32'h3975ba17),
	.w5(32'h3953df45),
	.w6(32'h38915a29),
	.w7(32'h39095f5b),
	.w8(32'h390ccc46),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7998943),
	.w1(32'h375c106a),
	.w2(32'h38a236be),
	.w3(32'h37d5dc58),
	.w4(32'h383f733c),
	.w5(32'h385c8d3f),
	.w6(32'hb893461a),
	.w7(32'hb907dfac),
	.w8(32'hb8f54f2f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b32f),
	.w1(32'h3818d7c5),
	.w2(32'h392c9d1a),
	.w3(32'h3b9b2658),
	.w4(32'hb9db06a4),
	.w5(32'hbb05bef8),
	.w6(32'h3b36224d),
	.w7(32'hbaa8e7c8),
	.w8(32'hb92c2cc4),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79b0a8),
	.w1(32'hb9875bbb),
	.w2(32'hba833501),
	.w3(32'h3c13fccd),
	.w4(32'hbbd80123),
	.w5(32'hbb9745ce),
	.w6(32'h3bddea67),
	.w7(32'hbc1365fc),
	.w8(32'hbb7aa66c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c421b),
	.w1(32'h3b5723f1),
	.w2(32'h3c5b35fe),
	.w3(32'h3c82828c),
	.w4(32'h3b50f677),
	.w5(32'h3c07f9f4),
	.w6(32'h3c1f2d72),
	.w7(32'h3a488644),
	.w8(32'h3bd76788),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88807e3),
	.w1(32'hb792998f),
	.w2(32'hb80a761e),
	.w3(32'hb83ab1f0),
	.w4(32'hb7808119),
	.w5(32'hb787d6a8),
	.w6(32'h37894cd8),
	.w7(32'h38888afe),
	.w8(32'hb81e3047),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e7348),
	.w1(32'h3ae7e804),
	.w2(32'h3c1bd760),
	.w3(32'h3c227b87),
	.w4(32'hba18880e),
	.w5(32'h3b830c9f),
	.w6(32'h3c20293e),
	.w7(32'hb81d6ddd),
	.w8(32'h3b5ff267),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c015c6b),
	.w1(32'h39c03a6e),
	.w2(32'h3b906526),
	.w3(32'h3bbe1a71),
	.w4(32'hbafab6f4),
	.w5(32'h393bc278),
	.w6(32'h3bb23e45),
	.w7(32'hba1fa110),
	.w8(32'h3b122632),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc25927),
	.w1(32'h3be2d34c),
	.w2(32'h3c589ffa),
	.w3(32'h3bc3f10c),
	.w4(32'h3b8a6ebd),
	.w5(32'h3be86ac2),
	.w6(32'hbbd3ef29),
	.w7(32'hbb1f66e3),
	.w8(32'h3b8cdc66),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d888c),
	.w1(32'hbb988934),
	.w2(32'h3bbb8db1),
	.w3(32'h3be77836),
	.w4(32'hbc21b478),
	.w5(32'hbab443c3),
	.w6(32'h3ba05298),
	.w7(32'hbc74016a),
	.w8(32'hbbe8fb01),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfb621),
	.w1(32'h3a7b40b8),
	.w2(32'h38d57321),
	.w3(32'h3bad7cc2),
	.w4(32'hb91a6809),
	.w5(32'hb9afc9c6),
	.w6(32'h3ba2f1c5),
	.w7(32'hbaf50442),
	.w8(32'h3a7f2651),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94e665),
	.w1(32'hbab9fa14),
	.w2(32'hba1d20c9),
	.w3(32'hbab38459),
	.w4(32'hbaa169ba),
	.w5(32'hb98dcf0c),
	.w6(32'hbaa6d352),
	.w7(32'hbb1e9441),
	.w8(32'hbac747c2),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beea5fd),
	.w1(32'hbb7e0236),
	.w2(32'h380d55fc),
	.w3(32'h3b95fbac),
	.w4(32'hbbba296f),
	.w5(32'hbaebd21f),
	.w6(32'h3bc7bdbd),
	.w7(32'hbbc6913d),
	.w8(32'hbaaf48f8),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7662ea),
	.w1(32'hba774afd),
	.w2(32'hb87de39f),
	.w3(32'h3c33681b),
	.w4(32'hbbff5220),
	.w5(32'hbb50556c),
	.w6(32'h3c068e4d),
	.w7(32'hbc062dc3),
	.w8(32'hbaa6228f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bd23c),
	.w1(32'hbbc54256),
	.w2(32'h399237c0),
	.w3(32'h3b90477c),
	.w4(32'hbbf45dd7),
	.w5(32'hbad801ad),
	.w6(32'h3ba5e261),
	.w7(32'hbc0a369e),
	.w8(32'hbacb9ede),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae06eb7),
	.w1(32'h3aa485e7),
	.w2(32'h3a9b81f8),
	.w3(32'h3afe9f41),
	.w4(32'h3adfa917),
	.w5(32'h3aac1489),
	.w6(32'hb9ef08e2),
	.w7(32'h387faf8f),
	.w8(32'h3a2b81c2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a096b50),
	.w1(32'h39990376),
	.w2(32'h39e00265),
	.w3(32'h392162ea),
	.w4(32'h372d38cd),
	.w5(32'hb87f0cfd),
	.w6(32'h3a09b694),
	.w7(32'h3a1d39b3),
	.w8(32'h3a0ce279),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53ac48),
	.w1(32'h3b4cc319),
	.w2(32'h3ba872ca),
	.w3(32'h3c012b1e),
	.w4(32'h3a7dc5b4),
	.w5(32'h3b21e350),
	.w6(32'h3bb6ec13),
	.w7(32'h3a198d38),
	.w8(32'h3b392e8b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25e29c),
	.w1(32'hb94ebdf4),
	.w2(32'h3a982a20),
	.w3(32'hba4b99b0),
	.w4(32'hba24797f),
	.w5(32'h3a425ba1),
	.w6(32'hbafa4696),
	.w7(32'hbab08f61),
	.w8(32'h3996337c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914253),
	.w1(32'hbb31c483),
	.w2(32'h3ae4c082),
	.w3(32'h3b739592),
	.w4(32'hbb569f0f),
	.w5(32'hba87c907),
	.w6(32'h3ba4d959),
	.w7(32'hbb705cdb),
	.w8(32'hbafcff47),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cb3ca),
	.w1(32'hb92d9fd8),
	.w2(32'h3a49722f),
	.w3(32'hba02395d),
	.w4(32'hba5e41ce),
	.w5(32'h393a6b6f),
	.w6(32'hb9b35ed2),
	.w7(32'hba928bc7),
	.w8(32'h3944e904),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201af6),
	.w1(32'hbaccd0e4),
	.w2(32'h3bd04fcd),
	.w3(32'h3b963111),
	.w4(32'h3a6b932b),
	.w5(32'h3c17b2f9),
	.w6(32'h3b86d6b9),
	.w7(32'hb993f442),
	.w8(32'h3c1265ec),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386cc2bf),
	.w1(32'hb960163d),
	.w2(32'hb90f3406),
	.w3(32'hb90693e6),
	.w4(32'hb959de7a),
	.w5(32'hb8b40d36),
	.w6(32'hb83d1f50),
	.w7(32'hb910f03a),
	.w8(32'hb8f9f213),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6b18),
	.w1(32'h3a25e35b),
	.w2(32'h3aa6f4e9),
	.w3(32'h3a1cf63b),
	.w4(32'h3a33a37b),
	.w5(32'h3a87c7a3),
	.w6(32'h39ded31e),
	.w7(32'h39c62af3),
	.w8(32'h3a7b1276),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdf08d),
	.w1(32'hb76c6c60),
	.w2(32'h3b2c31d6),
	.w3(32'h3bb4e707),
	.w4(32'hbb853501),
	.w5(32'hba91b4f6),
	.w6(32'h3bc4a83a),
	.w7(32'hbb970289),
	.w8(32'hbb1758a8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c40b4),
	.w1(32'hba9825bc),
	.w2(32'h3babdd19),
	.w3(32'h3c855cb7),
	.w4(32'hbab50309),
	.w5(32'h3c1cbdba),
	.w6(32'h3c4d0310),
	.w7(32'hbb3ddc21),
	.w8(32'h3b92e8ef),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff2f90),
	.w1(32'hbb7f298a),
	.w2(32'h3aa5f5cb),
	.w3(32'h3a727432),
	.w4(32'hbb93d23a),
	.w5(32'h3a1fea4d),
	.w6(32'h3b71ba35),
	.w7(32'hbb4b93c5),
	.w8(32'h3aeb8c09),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c3799),
	.w1(32'h3b258320),
	.w2(32'h3c2bb777),
	.w3(32'h3c1cdc6c),
	.w4(32'h3a4a754b),
	.w5(32'h3beb61a8),
	.w6(32'h3bf4b268),
	.w7(32'hbaeea5b6),
	.w8(32'h3bb5f584),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af718d4),
	.w1(32'hb918ffe4),
	.w2(32'h3b20e0f7),
	.w3(32'h3b0c9201),
	.w4(32'hba78af14),
	.w5(32'h386b5336),
	.w6(32'h39288778),
	.w7(32'hbb0e79fe),
	.w8(32'hba8f218f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c941c77),
	.w1(32'h3b035e21),
	.w2(32'h3c935584),
	.w3(32'h3c6baf87),
	.w4(32'hbba31af6),
	.w5(32'h3b8292dc),
	.w6(32'h3c5bb96b),
	.w7(32'h3ab7f770),
	.w8(32'h3bdd66ff),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7ef8d8),
	.w1(32'h3b07ffea),
	.w2(32'h3c1880d1),
	.w3(32'h3c398706),
	.w4(32'hbb3e3af8),
	.w5(32'h3b0bd00e),
	.w6(32'h3c13a3fd),
	.w7(32'hbb9d9bc1),
	.w8(32'h3b14a25c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24b6f2),
	.w1(32'hba378987),
	.w2(32'h3baf7181),
	.w3(32'h3be03c53),
	.w4(32'hbaccd04e),
	.w5(32'h3b0711ed),
	.w6(32'h3bba1b9c),
	.w7(32'hbac798a9),
	.w8(32'h3a98719c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91aaba1),
	.w1(32'hba318ba1),
	.w2(32'hba6754d5),
	.w3(32'hb9fefcfd),
	.w4(32'hba4e7d75),
	.w5(32'hbaa3bc1c),
	.w6(32'hb9fe4731),
	.w7(32'hba8d2abe),
	.w8(32'hba9c1e95),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be53771),
	.w1(32'h3a8ebc88),
	.w2(32'h3b5900ba),
	.w3(32'h3bc30398),
	.w4(32'hba1735c0),
	.w5(32'hb98749f6),
	.w6(32'h3b4062a5),
	.w7(32'hbb290386),
	.w8(32'hbb0f6a0b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7a9e3),
	.w1(32'hb85fddc1),
	.w2(32'hb8d2c18e),
	.w3(32'hb98aafc6),
	.w4(32'h37c6ffc9),
	.w5(32'hb81cabab),
	.w6(32'hb9912cc2),
	.w7(32'hb685fa68),
	.w8(32'hb8e1b726),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8546ec),
	.w1(32'hba6ad3c4),
	.w2(32'h3b1f3f21),
	.w3(32'hb819e4e0),
	.w4(32'hbb0564f1),
	.w5(32'h3a0295c2),
	.w6(32'h3a0fba64),
	.w7(32'hbaa2eb29),
	.w8(32'h3ad90d6d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b518a44),
	.w1(32'h3a41bd02),
	.w2(32'h3a94797e),
	.w3(32'h3b55b031),
	.w4(32'h3a1bbbc4),
	.w5(32'h3a32b9ae),
	.w6(32'h3b2c5656),
	.w7(32'hba014f4a),
	.w8(32'h3a3581dc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3757d0),
	.w1(32'h3aea4872),
	.w2(32'h3c18a9d2),
	.w3(32'h3c162f13),
	.w4(32'hb9b6db1c),
	.w5(32'h3b2f829d),
	.w6(32'h3c070c61),
	.w7(32'h39f33421),
	.w8(32'h3b85e805),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900028f),
	.w1(32'hb5cdef68),
	.w2(32'hb816168f),
	.w3(32'hb8c08bc7),
	.w4(32'h379d39ec),
	.w5(32'hb780383d),
	.w6(32'hb8df64e0),
	.w7(32'hb7c2822e),
	.w8(32'hb884a0f6),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac7380),
	.w1(32'h375e037e),
	.w2(32'h3920a0d0),
	.w3(32'h390b81a8),
	.w4(32'h39552ffd),
	.w5(32'h394992b8),
	.w6(32'hb89f0697),
	.w7(32'hb84fffe2),
	.w8(32'h376981b7),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4274b),
	.w1(32'h3a8161d3),
	.w2(32'h3ac60399),
	.w3(32'h3b9977cf),
	.w4(32'hba43ce34),
	.w5(32'hba067159),
	.w6(32'h3ab7a923),
	.w7(32'hbb6bd705),
	.w8(32'hbb1247ed),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ded04),
	.w1(32'hb9a8b721),
	.w2(32'h3bd7ffa0),
	.w3(32'h3c20d599),
	.w4(32'hbb354d8c),
	.w5(32'h3a93e9f0),
	.w6(32'h3be6dd75),
	.w7(32'hbb3f7166),
	.w8(32'h3ad8ffe2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b898219),
	.w1(32'hba09de98),
	.w2(32'h39196912),
	.w3(32'h3b9e4f8a),
	.w4(32'hb9fb66b0),
	.w5(32'h3afd9836),
	.w6(32'hba970709),
	.w7(32'hbbcbf632),
	.w8(32'h39eeb419),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f2393),
	.w1(32'h3987b3c3),
	.w2(32'h3ab035dc),
	.w3(32'h3ac5ebd5),
	.w4(32'h39be2cf2),
	.w5(32'h3ad97b33),
	.w6(32'h3af0668c),
	.w7(32'h38ddf8bb),
	.w8(32'h3b148db0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f1b84),
	.w1(32'h3c2105f9),
	.w2(32'h3cea702c),
	.w3(32'h3c8ed7ca),
	.w4(32'h3c259e53),
	.w5(32'h3cb7bbf0),
	.w6(32'h3be3ac84),
	.w7(32'h3c0acdf7),
	.w8(32'h3c4bde18),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03a39b),
	.w1(32'h3ab492eb),
	.w2(32'h3c5156cd),
	.w3(32'h3cc9a8cb),
	.w4(32'hbc2507e9),
	.w5(32'hbba61762),
	.w6(32'h3c912a56),
	.w7(32'hbca5021e),
	.w8(32'hbc018f8f),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb866478c),
	.w1(32'h3ac52670),
	.w2(32'h3ab6a972),
	.w3(32'h379b9b88),
	.w4(32'h3ae885d5),
	.w5(32'h3b1459f0),
	.w6(32'hba87b171),
	.w7(32'h3a422990),
	.w8(32'h3b139929),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8846e44),
	.w1(32'h38717d33),
	.w2(32'h382b910c),
	.w3(32'hb8040ed5),
	.w4(32'h392b7cef),
	.w5(32'h391a6517),
	.w6(32'hb8d6f053),
	.w7(32'h38b9b2ce),
	.w8(32'h38cfed43),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962b857),
	.w1(32'h3937f720),
	.w2(32'h39d1d650),
	.w3(32'hb903dbd3),
	.w4(32'h387b5058),
	.w5(32'h39e84f1c),
	.w6(32'hb84e66b4),
	.w7(32'h384b09b2),
	.w8(32'h39cf745c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d467d),
	.w1(32'hb8139f94),
	.w2(32'hb8a14db8),
	.w3(32'hb94d06eb),
	.w4(32'h37a15044),
	.w5(32'hb7d73e28),
	.w6(32'hb963fa94),
	.w7(32'hb7a8687b),
	.w8(32'hb8a7362e),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a965e0e),
	.w1(32'h3b385eeb),
	.w2(32'h3b92f65a),
	.w3(32'h3ae11ac7),
	.w4(32'h3b93b65c),
	.w5(32'h3b9a1650),
	.w6(32'hba1b0fd3),
	.w7(32'h3b1c45be),
	.w8(32'h3b8e500d),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fc5d4),
	.w1(32'h3af97733),
	.w2(32'h3b1d4f84),
	.w3(32'h3bdd5163),
	.w4(32'hbba06234),
	.w5(32'hbb0ee7ef),
	.w6(32'h3beca7c1),
	.w7(32'hba8f69ea),
	.w8(32'h3b80dc16),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8dcd6b),
	.w1(32'h3b8ee6ff),
	.w2(32'h3c4a73e3),
	.w3(32'h3c778411),
	.w4(32'hbb7bf639),
	.w5(32'h3b32934c),
	.w6(32'h3c30aa25),
	.w7(32'hbbef6b13),
	.w8(32'hbab8be45),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d39a),
	.w1(32'hbb2afa07),
	.w2(32'hba2a13e6),
	.w3(32'h3b33c7f8),
	.w4(32'hbb1659f1),
	.w5(32'hb95822a4),
	.w6(32'h3b292bb8),
	.w7(32'hba8644a2),
	.w8(32'h3ad1f58c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27e047),
	.w1(32'h3be6d3a6),
	.w2(32'h3c85edb9),
	.w3(32'h3befd766),
	.w4(32'h3accf0fe),
	.w5(32'h3c21365d),
	.w6(32'h3bd80e8f),
	.w7(32'h3af816c0),
	.w8(32'h3c04df25),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2291f4),
	.w1(32'h3938c760),
	.w2(32'h3a8d8659),
	.w3(32'h3b1273e7),
	.w4(32'h3a4198d9),
	.w5(32'h3ad4625c),
	.w6(32'h3a94423e),
	.w7(32'h36cb3d2a),
	.w8(32'h39a9df18),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3f426),
	.w1(32'hb9245663),
	.w2(32'hb9a74bc9),
	.w3(32'hb9a329b0),
	.w4(32'hb8a7c9de),
	.w5(32'hb9731582),
	.w6(32'hb9adb907),
	.w7(32'hb8faa1ab),
	.w8(32'hb9911185),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42f196),
	.w1(32'h3af0cd24),
	.w2(32'hb9e0aca5),
	.w3(32'h3b1c2e19),
	.w4(32'h3b123ffe),
	.w5(32'h3998828c),
	.w6(32'h39dbf593),
	.w7(32'hba99de7f),
	.w8(32'hbb324098),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ad710),
	.w1(32'hb95e3c3c),
	.w2(32'hba14b7d9),
	.w3(32'hba3444f7),
	.w4(32'hb8172c0c),
	.w5(32'hb9ab4916),
	.w6(32'hba45ce21),
	.w7(32'hb92e2e26),
	.w8(32'hb9fdb069),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50eb8f),
	.w1(32'h3ab25bf6),
	.w2(32'h3bcbea36),
	.w3(32'h3c2b416b),
	.w4(32'hbb05af0e),
	.w5(32'h38aa990f),
	.w6(32'h3c1299ed),
	.w7(32'hbb343bc7),
	.w8(32'h3a21c5ce),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a1dfc),
	.w1(32'hbb6d8e1b),
	.w2(32'h3a20ff0a),
	.w3(32'h3c476ebc),
	.w4(32'hbc102db8),
	.w5(32'hbb5be775),
	.w6(32'h3c740eaa),
	.w7(32'hbc1e72ff),
	.w8(32'hb9bb6727),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c605ea2),
	.w1(32'h3a908c1d),
	.w2(32'h3bec4a34),
	.w3(32'h3c252666),
	.w4(32'hbb8ddb21),
	.w5(32'h3a43377a),
	.w6(32'h3c182cd0),
	.w7(32'hbba3912d),
	.w8(32'h3acfd6e2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0222f8),
	.w1(32'h38777074),
	.w2(32'h3a2be671),
	.w3(32'h3ac16789),
	.w4(32'hb9d8e732),
	.w5(32'h3a64e8f8),
	.w6(32'h3b303f08),
	.w7(32'hb886a670),
	.w8(32'h3af3009f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c845b81),
	.w1(32'h3910d90a),
	.w2(32'h3bfab66d),
	.w3(32'h3c4ca1b6),
	.w4(32'hbbb9eaa5),
	.w5(32'hb8f6dc3d),
	.w6(32'h3c1ec721),
	.w7(32'hbc01bb3f),
	.w8(32'hbac79935),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaca7f),
	.w1(32'h3acf10c0),
	.w2(32'h3bce4594),
	.w3(32'h3bc7a749),
	.w4(32'h3a81cc83),
	.w5(32'h3b6640dc),
	.w6(32'h3bd0cb40),
	.w7(32'h3b3a75f0),
	.w8(32'h3b43cbe7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca5cd77),
	.w1(32'hba3c4dd5),
	.w2(32'h3c3f9f1f),
	.w3(32'h3c95d98b),
	.w4(32'hbb541844),
	.w5(32'h3bdd2bde),
	.w6(32'h3c2c664e),
	.w7(32'hbb5ebd71),
	.w8(32'h3bdab726),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d50700),
	.w1(32'h388c3760),
	.w2(32'hb85e2dbe),
	.w3(32'hb8664cff),
	.w4(32'h386e6342),
	.w5(32'hb774d2af),
	.w6(32'hb95cd43a),
	.w7(32'hb7c617d3),
	.w8(32'hb908708f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3d7d3),
	.w1(32'hb9d1f302),
	.w2(32'hb9306bc8),
	.w3(32'hb681090f),
	.w4(32'hb865537b),
	.w5(32'h3996a95c),
	.w6(32'h3863db7c),
	.w7(32'hb9b59653),
	.w8(32'hb80790ce),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c791377),
	.w1(32'h3a5f1af4),
	.w2(32'h3bf4ee71),
	.w3(32'h3c328119),
	.w4(32'hbaf732cd),
	.w5(32'h3b947ac6),
	.w6(32'h3bedb8fc),
	.w7(32'hbb7d28f7),
	.w8(32'h3b797bbd),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bcc23),
	.w1(32'hbb53ddbf),
	.w2(32'h3ba4ea26),
	.w3(32'h3c891be9),
	.w4(32'hbb0ad97e),
	.w5(32'h3baff4b6),
	.w6(32'h3c4598fc),
	.w7(32'hbb90c9f3),
	.w8(32'h3949d566),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a90ff),
	.w1(32'h3b0fe68e),
	.w2(32'h3bef43d2),
	.w3(32'h3c4d3c77),
	.w4(32'hbb9ef9ff),
	.w5(32'hba801501),
	.w6(32'h3c2f584a),
	.w7(32'hbbf2f4a2),
	.w8(32'hbb37d181),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab126b1),
	.w1(32'h3b3d9f1f),
	.w2(32'h3b7be45c),
	.w3(32'h3bba47ef),
	.w4(32'h3c0f2782),
	.w5(32'h3bb469fa),
	.w6(32'hbba06883),
	.w7(32'h39217614),
	.w8(32'h3b8d77d7),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39477cc5),
	.w1(32'h399db376),
	.w2(32'h3a22e171),
	.w3(32'h39abfa6b),
	.w4(32'h3a44033c),
	.w5(32'h3a0e01db),
	.w6(32'h39b7fe33),
	.w7(32'h3a4a9360),
	.w8(32'h3a2a93a0),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addcb51),
	.w1(32'h3a714ea5),
	.w2(32'hb998e62f),
	.w3(32'h3abf9a1d),
	.w4(32'h3a4155bc),
	.w5(32'hb8fbf4ce),
	.w6(32'h3abb8cec),
	.w7(32'h3a30829e),
	.w8(32'hb7b0e000),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f12fcb),
	.w1(32'hbae3a5ec),
	.w2(32'h3bcf8d1a),
	.w3(32'hba2edc81),
	.w4(32'h3b9cd6a3),
	.w5(32'h3c305b23),
	.w6(32'hbbd87fb7),
	.w7(32'hbb7e583a),
	.w8(32'h3ba5ed72),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51afd8),
	.w1(32'h3baf3b14),
	.w2(32'h3c6fe933),
	.w3(32'h3c4d0c63),
	.w4(32'h3bb07bcb),
	.w5(32'h3c68a742),
	.w6(32'h3bd02560),
	.w7(32'h3b89269d),
	.w8(32'h3c255a3f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8617b2),
	.w1(32'h3ba9ce94),
	.w2(32'h3ba26e70),
	.w3(32'h3b8961e2),
	.w4(32'h3bcdef10),
	.w5(32'h3bab1379),
	.w6(32'hbbad5929),
	.w7(32'hbb0e437b),
	.w8(32'hb955e9c8),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c260ad1),
	.w1(32'hbbb654cb),
	.w2(32'h395ad092),
	.w3(32'h3c19372e),
	.w4(32'hbbf2aac8),
	.w5(32'hbb02eae9),
	.w6(32'h3c0ff969),
	.w7(32'hbc00401d),
	.w8(32'hba71648f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c805e35),
	.w1(32'h3a1355a1),
	.w2(32'h3bf6547b),
	.w3(32'h3c641b41),
	.w4(32'hbbaa1317),
	.w5(32'h3a8764fc),
	.w6(32'h3c3b56fb),
	.w7(32'hbc0094b5),
	.w8(32'hb98bfd31),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93850dc),
	.w1(32'hb8b297d9),
	.w2(32'hb8c90804),
	.w3(32'hb913677f),
	.w4(32'hb880bbb0),
	.w5(32'hb8ad7ad5),
	.w6(32'hb9298326),
	.w7(32'hb8bf6d1a),
	.w8(32'hb8e7c64a),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c27d1),
	.w1(32'hb8ba47a7),
	.w2(32'hb90fa275),
	.w3(32'hb952c82c),
	.w4(32'hb819edf4),
	.w5(32'hb8b7211d),
	.w6(32'hb9504375),
	.w7(32'hb83936f8),
	.w8(32'hb8d95ab4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba879e4d),
	.w1(32'hb9ca9c08),
	.w2(32'hb946cbb7),
	.w3(32'hba854400),
	.w4(32'h39420a57),
	.w5(32'h39841e89),
	.w6(32'hba8c6296),
	.w7(32'h3990ebdc),
	.w8(32'h39b1de4a),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996b3b4),
	.w1(32'hb84899ea),
	.w2(32'hb8c89e96),
	.w3(32'hb98352ad),
	.w4(32'h36b3750f),
	.w5(32'hb851480c),
	.w6(32'hb9924df7),
	.w7(32'hb690e85f),
	.w8(32'hb8988e51),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74a0b0),
	.w1(32'h3b3e772c),
	.w2(32'h3b819795),
	.w3(32'h39dcda9c),
	.w4(32'h3b424541),
	.w5(32'h3b81b38c),
	.w6(32'hba0c04d9),
	.w7(32'h3ab2f4fc),
	.w8(32'h3b5a015b),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c83ea),
	.w1(32'hb8e40e5f),
	.w2(32'h3b9d6f34),
	.w3(32'h3c01d038),
	.w4(32'hbac5f5c2),
	.w5(32'h3b691c0f),
	.w6(32'h3be08b16),
	.w7(32'hbace7eab),
	.w8(32'h3b02d5bb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c200585),
	.w1(32'hba0c9d61),
	.w2(32'h3b233ef8),
	.w3(32'h3c1bc882),
	.w4(32'hba55fb7c),
	.w5(32'h3ad345d6),
	.w6(32'h3bba0aee),
	.w7(32'hba9c0aac),
	.w8(32'h38fa9da3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944abb5),
	.w1(32'hb8cc72d5),
	.w2(32'hb90cacac),
	.w3(32'hb96eea67),
	.w4(32'hb9109f3c),
	.w5(32'hb91f8464),
	.w6(32'hb9740986),
	.w7(32'hb94ced0f),
	.w8(32'hb9530237),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd16914),
	.w1(32'h3b8351eb),
	.w2(32'h3c370d3d),
	.w3(32'h3ba9c1af),
	.w4(32'h3bb0c479),
	.w5(32'h3c47605b),
	.w6(32'hbbd4c806),
	.w7(32'hbbcdd449),
	.w8(32'h3b9ea601),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71487a),
	.w1(32'h39acfbce),
	.w2(32'h3ac7b291),
	.w3(32'h3aff0770),
	.w4(32'hb99e49d8),
	.w5(32'h3a9ab309),
	.w6(32'h3a258aad),
	.w7(32'hba5b287a),
	.w8(32'h3a0d9d3a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39816e88),
	.w1(32'hb90c5ef4),
	.w2(32'hba4cea19),
	.w3(32'h39dab5b4),
	.w4(32'hb8bfbfb5),
	.w5(32'hb9fb36cc),
	.w6(32'h398ab857),
	.w7(32'hb8fea3b9),
	.w8(32'hb9c43911),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7326e6),
	.w1(32'h3b60406e),
	.w2(32'h3bd0bca5),
	.w3(32'h3b2bc31b),
	.w4(32'h3b5442c2),
	.w5(32'h3badb3e6),
	.w6(32'h3a919cc3),
	.w7(32'h3add4851),
	.w8(32'h3b814e30),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbf7b6),
	.w1(32'hb9c4b515),
	.w2(32'hb9943bda),
	.w3(32'hb9d74df9),
	.w4(32'hb9becee1),
	.w5(32'hb9acc1cf),
	.w6(32'hb9000df8),
	.w7(32'hb92dd6b2),
	.w8(32'hb9372e66),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1fe36),
	.w1(32'hba91194c),
	.w2(32'hbad11d77),
	.w3(32'h38d68ca9),
	.w4(32'hba93b2ed),
	.w5(32'hbac801b7),
	.w6(32'h3ac066b6),
	.w7(32'h3a1a8491),
	.w8(32'h39455a85),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a359c),
	.w1(32'hb913f95c),
	.w2(32'hb95e53b8),
	.w3(32'hb8bb9c35),
	.w4(32'hb89225a7),
	.w5(32'hb93cbf08),
	.w6(32'hb8ebd620),
	.w7(32'hb887142c),
	.w8(32'hb8f685d8),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979f0de),
	.w1(32'hb91964d9),
	.w2(32'hb90b8c3e),
	.w3(32'hb9410692),
	.w4(32'hb8c4ed95),
	.w5(32'hb8af7f3d),
	.w6(32'hb93c6537),
	.w7(32'hb8bf6227),
	.w8(32'hb8994121),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97fbd3),
	.w1(32'h396f6fd1),
	.w2(32'h3a874f2e),
	.w3(32'h3bb0d920),
	.w4(32'h3a9cfadf),
	.w5(32'h3a1e89ee),
	.w6(32'h3bc64e75),
	.w7(32'hba3546f4),
	.w8(32'hba826732),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b832a),
	.w1(32'h3a8c8db5),
	.w2(32'h3c469c6f),
	.w3(32'h3c1bafc6),
	.w4(32'hba9b1281),
	.w5(32'h3af7c056),
	.w6(32'h3c03a7d7),
	.w7(32'hb9320317),
	.w8(32'h3b445bad),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09796c),
	.w1(32'h3b66bd93),
	.w2(32'h3be446ee),
	.w3(32'h3ba4f5ab),
	.w4(32'h3b30c72d),
	.w5(32'h3bbda3e3),
	.w6(32'h3b2ce756),
	.w7(32'hba2ebd92),
	.w8(32'h3b3c8c7a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c230c8a),
	.w1(32'h3b7d9570),
	.w2(32'h3c3bcb17),
	.w3(32'h3c188394),
	.w4(32'h3b82c912),
	.w5(32'h3bd0ab99),
	.w6(32'h3b940741),
	.w7(32'h3baec814),
	.w8(32'h3bea842d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8905ad9),
	.w1(32'hb90e5c60),
	.w2(32'h3939ae9e),
	.w3(32'hb90bd572),
	.w4(32'hba02e919),
	.w5(32'hb907b6ba),
	.w6(32'h3851d806),
	.w7(32'hba1590bf),
	.w8(32'hb90a20bc),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dcd096),
	.w1(32'h3a509682),
	.w2(32'h39f42e9b),
	.w3(32'h392c7a5d),
	.w4(32'h39ff19eb),
	.w5(32'hb8a1dc28),
	.w6(32'h3879662c),
	.w7(32'h39c38448),
	.w8(32'hb833ea8a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848d941),
	.w1(32'h38244210),
	.w2(32'hb7aa0b3b),
	.w3(32'hb8631a58),
	.w4(32'h3870e8ae),
	.w5(32'hb6ea800f),
	.w6(32'hb8ac3a23),
	.w7(32'h38698dd8),
	.w8(32'hb6e30104),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91abb71),
	.w1(32'hb903699f),
	.w2(32'hb91beaeb),
	.w3(32'hb93e363f),
	.w4(32'hb8943087),
	.w5(32'hb8820b70),
	.w6(32'hb91836f0),
	.w7(32'h38a6217b),
	.w8(32'h38238182),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ca703),
	.w1(32'h3b207264),
	.w2(32'h3baf80bc),
	.w3(32'h3c0eab0b),
	.w4(32'hb9e79403),
	.w5(32'h3aa4779f),
	.w6(32'h3be7eaac),
	.w7(32'hbad00d15),
	.w8(32'hba56e193),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a265d38),
	.w1(32'h3a492688),
	.w2(32'h3a034afe),
	.w3(32'h3a030466),
	.w4(32'h3a4a39b6),
	.w5(32'h3a379f65),
	.w6(32'h39949723),
	.w7(32'h3a224bef),
	.w8(32'h3a34ae81),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d21b08),
	.w1(32'hbb713d70),
	.w2(32'h3b1233c2),
	.w3(32'h3a220d98),
	.w4(32'hbb8292b6),
	.w5(32'h3abeecd8),
	.w6(32'h3b3a72af),
	.w7(32'hbb248fb7),
	.w8(32'h3b47ee1e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6df204),
	.w1(32'h39845162),
	.w2(32'h3aaa9f6b),
	.w3(32'h3b60c37a),
	.w4(32'h399d7b58),
	.w5(32'h3a628c2e),
	.w6(32'h3b42a50b),
	.w7(32'hba72068f),
	.w8(32'hb8bf5a10),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d0b29f),
	.w1(32'hb8512313),
	.w2(32'h37841272),
	.w3(32'hb95f4432),
	.w4(32'hb8d1e9e2),
	.w5(32'hb781b64d),
	.w6(32'hb96f9413),
	.w7(32'hb8675a66),
	.w8(32'h385271fb),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b404379),
	.w1(32'h3a85598c),
	.w2(32'h3b11a8d1),
	.w3(32'h3b2a81be),
	.w4(32'h3a0fbb67),
	.w5(32'h3aad8cb8),
	.w6(32'h39da759c),
	.w7(32'h399cda06),
	.w8(32'h3a85e1c0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b07f75),
	.w1(32'h38af2fe4),
	.w2(32'h38b6bb0a),
	.w3(32'h378a6394),
	.w4(32'hb9016410),
	.w5(32'hb8c25aa0),
	.w6(32'h36e5cbdc),
	.w7(32'h35ac7239),
	.w8(32'h3988af71),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94665e),
	.w1(32'h3c1ec2c2),
	.w2(32'h3c9040f2),
	.w3(32'h3c4ce93a),
	.w4(32'h3bdeecc1),
	.w5(32'h3b98cd6a),
	.w6(32'h3c4ada76),
	.w7(32'h3b42490f),
	.w8(32'h3baa20db),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f130cc),
	.w1(32'h38c1412d),
	.w2(32'hb96721ac),
	.w3(32'hb90a0c04),
	.w4(32'h39e99a4e),
	.w5(32'h36a77b48),
	.w6(32'h38312f29),
	.w7(32'hb8808647),
	.w8(32'h38aa4a99),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1baf4d),
	.w1(32'hbb775b37),
	.w2(32'hbb34d1a1),
	.w3(32'h3c5c4580),
	.w4(32'h3b128566),
	.w5(32'h3aed88ee),
	.w6(32'h3c5546f7),
	.w7(32'hbb10ae55),
	.w8(32'hbb90b42c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule