module layer_10_featuremap_485(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa25bc),
	.w1(32'h3b46c7d9),
	.w2(32'h3ad34084),
	.w3(32'hbafd93ca),
	.w4(32'hba9c9017),
	.w5(32'h3b1168ef),
	.w6(32'hbb642d05),
	.w7(32'h3b9c1491),
	.w8(32'h3b619390),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828b13),
	.w1(32'hbae2fd50),
	.w2(32'h3bf8a508),
	.w3(32'h3b41e199),
	.w4(32'hbbb80e40),
	.w5(32'hbc196f6e),
	.w6(32'hba2cffa5),
	.w7(32'hbba517c9),
	.w8(32'hbb8b51e9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c095398),
	.w1(32'hbb3c7929),
	.w2(32'h3b7d1ec7),
	.w3(32'h3c46c107),
	.w4(32'hbbabf018),
	.w5(32'hbb6080e5),
	.w6(32'h3bcc0225),
	.w7(32'hbc0c697f),
	.w8(32'hbc23db86),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919cb88),
	.w1(32'h3b8d47f3),
	.w2(32'h3b6943f1),
	.w3(32'h3bd522a9),
	.w4(32'h3b60a963),
	.w5(32'hbb8bd368),
	.w6(32'h3b687b87),
	.w7(32'h3b856c08),
	.w8(32'h3bf2e77b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b017),
	.w1(32'hbb40e11a),
	.w2(32'h3b42920e),
	.w3(32'hb9950e81),
	.w4(32'hbbc6866b),
	.w5(32'hbb1f3060),
	.w6(32'h3bda275b),
	.w7(32'hbad133f0),
	.w8(32'hbb8eae43),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e7d1),
	.w1(32'hbba3df6b),
	.w2(32'h3b29f599),
	.w3(32'h3c89c6a6),
	.w4(32'hba3409f8),
	.w5(32'hbb56fa33),
	.w6(32'h392e71e1),
	.w7(32'hbc2bf005),
	.w8(32'hbbb39232),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f25e5),
	.w1(32'hbb82b2a6),
	.w2(32'h3ad5b3b1),
	.w3(32'h3a96df00),
	.w4(32'h3ab87ea8),
	.w5(32'hbbed6095),
	.w6(32'hbb783cde),
	.w7(32'h3b47a23e),
	.w8(32'h3be09456),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90a34a),
	.w1(32'h3b021738),
	.w2(32'hbaf153cb),
	.w3(32'hbbf09af5),
	.w4(32'h3b231dea),
	.w5(32'h3bf510dc),
	.w6(32'h3b8059ff),
	.w7(32'h3b959b2d),
	.w8(32'h3a5c0604),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa10cc),
	.w1(32'h3a02e297),
	.w2(32'hbad1752c),
	.w3(32'hbbf9077c),
	.w4(32'hbbf1aa74),
	.w5(32'hbc2d96e3),
	.w6(32'h38c0d1b7),
	.w7(32'hbbdb1243),
	.w8(32'h3a34966c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ce304),
	.w1(32'h3abf9d59),
	.w2(32'h3c009745),
	.w3(32'hbab2b7a6),
	.w4(32'hbadee7db),
	.w5(32'hbb8975bc),
	.w6(32'h3ae70ce3),
	.w7(32'h3951062f),
	.w8(32'h3b2183f3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be3cc),
	.w1(32'h3b9aff57),
	.w2(32'h3c2d3349),
	.w3(32'h3b580ca4),
	.w4(32'h3b9c4112),
	.w5(32'hbb963396),
	.w6(32'h3b08b800),
	.w7(32'hbae5fee4),
	.w8(32'h391a50e2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb489c),
	.w1(32'hbb02198e),
	.w2(32'h393a6cdc),
	.w3(32'hbb08fefa),
	.w4(32'hbb5dbc36),
	.w5(32'h3ad5a5a1),
	.w6(32'hbb0e067f),
	.w7(32'hbab307ac),
	.w8(32'hbad7908f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02ca0d),
	.w1(32'hbb9da7f7),
	.w2(32'h3ad5d558),
	.w3(32'hbb96e77c),
	.w4(32'h39294c3e),
	.w5(32'hbc33b8f8),
	.w6(32'hbab2643f),
	.w7(32'h39d4aec4),
	.w8(32'h3ace1247),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a9088),
	.w1(32'hba7efe89),
	.w2(32'h3c1abddb),
	.w3(32'h3b7d5870),
	.w4(32'hbbe22106),
	.w5(32'hbb4f5e79),
	.w6(32'h3b575520),
	.w7(32'hbb9d61a9),
	.w8(32'hbb6b599a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dc24e),
	.w1(32'h3ae6cd97),
	.w2(32'h3c00cb80),
	.w3(32'h3bbf716a),
	.w4(32'h3b5d2e98),
	.w5(32'hbafc8e3f),
	.w6(32'hbb1c4751),
	.w7(32'h3ae4799d),
	.w8(32'h3bd66e1d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd718c),
	.w1(32'h3c2fe520),
	.w2(32'h3b2b3878),
	.w3(32'h3c15a16a),
	.w4(32'h3bf4aee7),
	.w5(32'h3b8d34b8),
	.w6(32'h3bab724f),
	.w7(32'h3b7ad09f),
	.w8(32'h3b9ba8e5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc206740),
	.w1(32'hbb9cad00),
	.w2(32'hbb3a1213),
	.w3(32'hbb911449),
	.w4(32'hbbec844f),
	.w5(32'hbb9d9d9c),
	.w6(32'hbbba7722),
	.w7(32'hbb96b963),
	.w8(32'hbbf4963d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eb42c),
	.w1(32'hbad03e12),
	.w2(32'hbb80627c),
	.w3(32'hbb8f3959),
	.w4(32'hbc15e490),
	.w5(32'h3b299603),
	.w6(32'hbb93b357),
	.w7(32'hbae87dd1),
	.w8(32'h3ada9025),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdf375),
	.w1(32'hbb8bcdce),
	.w2(32'h3a2da0ba),
	.w3(32'hb7f48986),
	.w4(32'h3a62effc),
	.w5(32'hbc2d9bf3),
	.w6(32'hbb8e3c1e),
	.w7(32'h3b6f1071),
	.w8(32'hbb08de4d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b608e91),
	.w1(32'hbb5ceafc),
	.w2(32'h3b0945d7),
	.w3(32'h3a40cc5a),
	.w4(32'hbbaab310),
	.w5(32'hbab131ea),
	.w6(32'h3bcd5065),
	.w7(32'hbbf7b888),
	.w8(32'hba105e41),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbe705),
	.w1(32'h3b00374f),
	.w2(32'h3ac67156),
	.w3(32'h3bcd03d9),
	.w4(32'h3c139764),
	.w5(32'h3b938129),
	.w6(32'hbb9939b7),
	.w7(32'h3bc67f18),
	.w8(32'h3baa2aad),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb77424),
	.w1(32'hbb06b8b2),
	.w2(32'hbc046345),
	.w3(32'h3ad67b8f),
	.w4(32'hbc01c86b),
	.w5(32'hbb0816ae),
	.w6(32'h3c07ee9c),
	.w7(32'hbb3e0c2e),
	.w8(32'h3b99b4d9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01744d),
	.w1(32'hbb09820f),
	.w2(32'h3b84a6b7),
	.w3(32'h3cd51153),
	.w4(32'hbb4393c1),
	.w5(32'hbb90c63f),
	.w6(32'hba61bed3),
	.w7(32'hbb8635e7),
	.w8(32'hba2a61db),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520c01),
	.w1(32'h3afebdef),
	.w2(32'h3b2be34a),
	.w3(32'hbc75d9b5),
	.w4(32'h3b8721d5),
	.w5(32'h3b6643f1),
	.w6(32'hbbda02c5),
	.w7(32'h3a9ed28a),
	.w8(32'hbaf35b46),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6118e),
	.w1(32'h3b06c0f9),
	.w2(32'hbba48d37),
	.w3(32'h3b94cb92),
	.w4(32'h3ad7d6f4),
	.w5(32'hbc1ca281),
	.w6(32'h3b13bd93),
	.w7(32'h3b1c63af),
	.w8(32'h3c0d2ebf),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea9d23),
	.w1(32'hbba2ac51),
	.w2(32'hba990284),
	.w3(32'hbbabe24c),
	.w4(32'hbb882096),
	.w5(32'h3c9600ad),
	.w6(32'h3b999ae4),
	.w7(32'hbb9fbfb1),
	.w8(32'hbc269076),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb956c16),
	.w1(32'hbb153dcb),
	.w2(32'hbba0ce85),
	.w3(32'hb97388f5),
	.w4(32'h39ae63f3),
	.w5(32'hb9a017c3),
	.w6(32'hbbeafd95),
	.w7(32'h3a2813e1),
	.w8(32'h3b9bd738),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbada5a6),
	.w1(32'hbb342ecd),
	.w2(32'hbb12181b),
	.w3(32'h3b234d4a),
	.w4(32'hbb2594b9),
	.w5(32'hbbb912c8),
	.w6(32'h3b37a8c1),
	.w7(32'hbb68d374),
	.w8(32'hb9c047db),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7eb7c1),
	.w1(32'hb91d6d03),
	.w2(32'hbb8f9c3a),
	.w3(32'hbb2e06bd),
	.w4(32'hbb1fe00c),
	.w5(32'hbbd9ea57),
	.w6(32'h39d67941),
	.w7(32'h3a4e85e7),
	.w8(32'h3baf617e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a38da),
	.w1(32'h3b510c79),
	.w2(32'h3b3b25f6),
	.w3(32'h3c1a0a7d),
	.w4(32'h3943eedc),
	.w5(32'h3c0200a3),
	.w6(32'hbb579deb),
	.w7(32'h37bcc7cf),
	.w8(32'hbb5843af),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f956),
	.w1(32'h3b1d96d0),
	.w2(32'h3b8b9de5),
	.w3(32'h3a074824),
	.w4(32'h3b6f0d65),
	.w5(32'h3c5ea280),
	.w6(32'hbb41c773),
	.w7(32'h3b4f9976),
	.w8(32'h3bdd6889),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44d39b),
	.w1(32'hba4ffe67),
	.w2(32'hbab1f5e4),
	.w3(32'hb95afcf9),
	.w4(32'h399354e6),
	.w5(32'h3b0147bd),
	.w6(32'hba06a59a),
	.w7(32'h3acfb4cf),
	.w8(32'h3b551348),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab42eae),
	.w1(32'h3a92edbf),
	.w2(32'h3be8a7a9),
	.w3(32'h3bbbbd04),
	.w4(32'hbbc9be56),
	.w5(32'hbc0fb479),
	.w6(32'h3a4dea87),
	.w7(32'hbbacb3c4),
	.w8(32'hbb83a2d9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef9aae),
	.w1(32'hbaa4a4bf),
	.w2(32'hb9c2ed28),
	.w3(32'h3a9f2a17),
	.w4(32'hbbb8de50),
	.w5(32'hbbe2f2ca),
	.w6(32'hbb9aceaa),
	.w7(32'hbad7fd33),
	.w8(32'h37d08ec8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d1183),
	.w1(32'hbb347e59),
	.w2(32'hba9111b7),
	.w3(32'hbb829869),
	.w4(32'hbbfd0907),
	.w5(32'h3b0c31fd),
	.w6(32'h3815b853),
	.w7(32'h3a83faef),
	.w8(32'hbc2c0e74),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f2b1d),
	.w1(32'h3b84af46),
	.w2(32'hbbddd98e),
	.w3(32'hbbc0b66a),
	.w4(32'h3a5caa0d),
	.w5(32'hbbb43986),
	.w6(32'h3993c3a1),
	.w7(32'h3bad6443),
	.w8(32'hba7479ab),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc369920),
	.w1(32'hba0fc760),
	.w2(32'h3c1d15d3),
	.w3(32'hbc170e66),
	.w4(32'hbbdf6008),
	.w5(32'hbc2c53de),
	.w6(32'hbaff9728),
	.w7(32'hbb681aac),
	.w8(32'hbab513a5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c470070),
	.w1(32'hbb897351),
	.w2(32'hbb098fb4),
	.w3(32'h3c6afb31),
	.w4(32'hba87ae2e),
	.w5(32'hbabcfd70),
	.w6(32'h3c2d8e71),
	.w7(32'h3a6a373d),
	.w8(32'hba3f6c57),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b839ceb),
	.w1(32'h3ba09cf7),
	.w2(32'h3a072c60),
	.w3(32'h3c50d4f9),
	.w4(32'h3bbacaa0),
	.w5(32'hbabf1aaa),
	.w6(32'h3bd4509e),
	.w7(32'h39acc0e5),
	.w8(32'h3b568a2e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebc638),
	.w1(32'h3b7ecac0),
	.w2(32'hb9e471aa),
	.w3(32'hbb9dc729),
	.w4(32'h3b6213a0),
	.w5(32'h3c03fc2d),
	.w6(32'hbaa31547),
	.w7(32'hbb1c6215),
	.w8(32'h3b81f611),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984d9d3),
	.w1(32'hbb9a2f75),
	.w2(32'hbb259bfd),
	.w3(32'hbb1466d5),
	.w4(32'hbc32fe11),
	.w5(32'h3bf9e927),
	.w6(32'h3b1e38f3),
	.w7(32'hbc08833b),
	.w8(32'hbb106694),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943af2),
	.w1(32'hbafcc662),
	.w2(32'hbbd1ae44),
	.w3(32'hbbaad337),
	.w4(32'h3afc46a7),
	.w5(32'hbc3c7197),
	.w6(32'hbc1401c5),
	.w7(32'hbaf51ad6),
	.w8(32'h39bce56f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acebf13),
	.w1(32'hbbab8102),
	.w2(32'h3aad2a96),
	.w3(32'hba36e991),
	.w4(32'hbc3336f6),
	.w5(32'hbbde1944),
	.w6(32'h3b11de7e),
	.w7(32'hbc30fafd),
	.w8(32'hbbf592fc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2be5fb),
	.w1(32'h3be23ade),
	.w2(32'h3c463d16),
	.w3(32'h3c2d3b1f),
	.w4(32'h3b8614dd),
	.w5(32'h3c3895cf),
	.w6(32'h3bcdea9a),
	.w7(32'h3a9403f8),
	.w8(32'hbb58d89d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe14554),
	.w1(32'hb811f88a),
	.w2(32'hbb66ddad),
	.w3(32'hbc4e637c),
	.w4(32'hbaffcab5),
	.w5(32'hbc0bf38b),
	.w6(32'hbbf9aae8),
	.w7(32'h3aeef4b3),
	.w8(32'hbb6678f3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad850ac),
	.w1(32'h3bec6385),
	.w2(32'h3bca51dc),
	.w3(32'h3b833a84),
	.w4(32'hb91084c3),
	.w5(32'h3b02e5f7),
	.w6(32'h3b081d74),
	.w7(32'h3b8b1a31),
	.w8(32'h3bbd3d33),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87d7874),
	.w1(32'hbb7cfcc6),
	.w2(32'hbb63e9ba),
	.w3(32'hbb634185),
	.w4(32'h3bbf6ffe),
	.w5(32'hbae0665e),
	.w6(32'h3b21ac3c),
	.w7(32'hbbb964a7),
	.w8(32'h3b44f5c9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f374e),
	.w1(32'hb82c585b),
	.w2(32'hbb88c708),
	.w3(32'hbbd0ea8a),
	.w4(32'h3a8797eb),
	.w5(32'hbc36787e),
	.w6(32'h3b1ef8ea),
	.w7(32'hbb1d64a3),
	.w8(32'hbae2d134),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50f48f),
	.w1(32'h3b537be2),
	.w2(32'hbc19b319),
	.w3(32'hbaffbf25),
	.w4(32'h3b9a984d),
	.w5(32'h3c15dd65),
	.w6(32'h3aa80fd9),
	.w7(32'h3ac3e625),
	.w8(32'h3b5954f8),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50574f),
	.w1(32'h3ac04e23),
	.w2(32'hbc5f421b),
	.w3(32'hbb7f7bcf),
	.w4(32'h3b1ec5ba),
	.w5(32'h3c103cda),
	.w6(32'hbc1d2123),
	.w7(32'h3b78982c),
	.w8(32'hb9e0b074),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadbe15),
	.w1(32'hbb8b8f15),
	.w2(32'hb9a51b6a),
	.w3(32'hbc398802),
	.w4(32'h3a85bd87),
	.w5(32'hbb85ad40),
	.w6(32'hbc106137),
	.w7(32'hba4c3b66),
	.w8(32'hbbc9f447),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b1649),
	.w1(32'hba01ffe5),
	.w2(32'h3bd6fc7a),
	.w3(32'hbb5eb0ed),
	.w4(32'hbb6289ba),
	.w5(32'hbb2b5e6c),
	.w6(32'h3b975b9a),
	.w7(32'h3b147004),
	.w8(32'h3bf37c12),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bf629),
	.w1(32'h3a7ab80f),
	.w2(32'hbbf5c395),
	.w3(32'h3c303222),
	.w4(32'hbbc3bc82),
	.w5(32'hbb3467df),
	.w6(32'h3bce2897),
	.w7(32'hbb600f47),
	.w8(32'hbb8a7c94),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7b06),
	.w1(32'hbbc05a9a),
	.w2(32'hbbed5cb0),
	.w3(32'hbc0c48f3),
	.w4(32'hbbbe728d),
	.w5(32'hbac68baf),
	.w6(32'hbae46d0c),
	.w7(32'h3b8ae10c),
	.w8(32'h3ab1ceb7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6879e),
	.w1(32'hbbeccbdf),
	.w2(32'hbb13c9ef),
	.w3(32'hbba81dc0),
	.w4(32'hbbab3108),
	.w5(32'hbbf42169),
	.w6(32'h3bf0d6db),
	.w7(32'hbbc5b6c9),
	.w8(32'hbbadfe1b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926eb0),
	.w1(32'h3961ab18),
	.w2(32'h3c52aa73),
	.w3(32'h3c1f1686),
	.w4(32'hbc315779),
	.w5(32'hbc2e23db),
	.w6(32'h3b9a8aa2),
	.w7(32'hbbf2eb8c),
	.w8(32'hbc37ad90),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c9f14),
	.w1(32'hbb8183ac),
	.w2(32'h3b55762a),
	.w3(32'h3ca40384),
	.w4(32'hbb0a87fc),
	.w5(32'h3bc5553f),
	.w6(32'h3bc9b085),
	.w7(32'hbbbe7951),
	.w8(32'h3ac8fc18),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05143),
	.w1(32'h39970490),
	.w2(32'h3c40f2ea),
	.w3(32'hba48d3ec),
	.w4(32'hbb8c7c18),
	.w5(32'hbc5c6b87),
	.w6(32'hbac69804),
	.w7(32'hbb617194),
	.w8(32'hbb4e9b1b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc10057),
	.w1(32'hbbd244f9),
	.w2(32'hbafdfac2),
	.w3(32'h3c6a8bc5),
	.w4(32'hbc0753be),
	.w5(32'hbb7bb8ef),
	.w6(32'h3975af2a),
	.w7(32'hbbe897c9),
	.w8(32'hbbe63995),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a84dc),
	.w1(32'hbb56fe29),
	.w2(32'hbbac4f5e),
	.w3(32'hb6f9659d),
	.w4(32'h3adbc8a4),
	.w5(32'h3aee4dd5),
	.w6(32'hbbcabcfc),
	.w7(32'hbb8d6838),
	.w8(32'hbb2a629d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924e5a7),
	.w1(32'hbbfa4655),
	.w2(32'hbb8e4968),
	.w3(32'hbc19abf1),
	.w4(32'hbadeed76),
	.w5(32'h3bfc84cc),
	.w6(32'hbba3b4cb),
	.w7(32'hbbc367c5),
	.w8(32'hbb095bd4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d9aa8),
	.w1(32'hbb62fb17),
	.w2(32'hbb125a5d),
	.w3(32'hbb23cd82),
	.w4(32'hbba400d2),
	.w5(32'hbb602b8e),
	.w6(32'h3a203aa1),
	.w7(32'hbc18e814),
	.w8(32'hbc151baf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10775d),
	.w1(32'hba062df5),
	.w2(32'hbb2816dc),
	.w3(32'h3b3e5ea0),
	.w4(32'hbb9a9301),
	.w5(32'hbc1fdbf0),
	.w6(32'hba967796),
	.w7(32'h3a911652),
	.w8(32'h3a9e9fb9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94058a5),
	.w1(32'hbbcba806),
	.w2(32'h3b95e276),
	.w3(32'h3be2e1f3),
	.w4(32'hbbb28f01),
	.w5(32'h3b894b74),
	.w6(32'h3bd11c02),
	.w7(32'hbbc79d15),
	.w8(32'hb809125e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23b7ae),
	.w1(32'h3b9f87fb),
	.w2(32'hbadee49a),
	.w3(32'h3bb7bc72),
	.w4(32'h3c43271d),
	.w5(32'h3c2bf087),
	.w6(32'h38b15ac3),
	.w7(32'h3c43f75c),
	.w8(32'h3b9daeef),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc385851),
	.w1(32'hb9f39ff3),
	.w2(32'h3a1c3caa),
	.w3(32'hbb54dd25),
	.w4(32'hbb55bf4b),
	.w5(32'h3ad53271),
	.w6(32'hba970322),
	.w7(32'hbbbb86a0),
	.w8(32'hbb89c060),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dbfe22),
	.w1(32'hbbdd0653),
	.w2(32'hbbff732e),
	.w3(32'hbbbc332a),
	.w4(32'hbc2c2e43),
	.w5(32'hbb020c07),
	.w6(32'hbbc8adc2),
	.w7(32'hbc73a422),
	.w8(32'hbc506c50),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb815),
	.w1(32'hbc1b7646),
	.w2(32'h3996d26e),
	.w3(32'hbc04e73a),
	.w4(32'hbc056403),
	.w5(32'hbc167d22),
	.w6(32'hba9fefee),
	.w7(32'hbc62122f),
	.w8(32'hbc0393e0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd421c),
	.w1(32'h3b57f729),
	.w2(32'h3b2fed0f),
	.w3(32'h39af1fd7),
	.w4(32'h3bcc5912),
	.w5(32'hbc62575a),
	.w6(32'hb84f61dd),
	.w7(32'h3c100478),
	.w8(32'h3b85448f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07b328),
	.w1(32'h399973eb),
	.w2(32'h3a9647d9),
	.w3(32'h3c0a94a8),
	.w4(32'h39a1e90e),
	.w5(32'h3b0b7fed),
	.w6(32'h3b980694),
	.w7(32'h3a603d3d),
	.w8(32'h3b0c849f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34a6f2),
	.w1(32'h39bb82b0),
	.w2(32'hba830257),
	.w3(32'h3a99e4c1),
	.w4(32'h3a816940),
	.w5(32'h39ee1cb9),
	.w6(32'h3a7b2dd1),
	.w7(32'h3abcf29b),
	.w8(32'h3a7a72a7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381e64d2),
	.w1(32'h3b35da53),
	.w2(32'h3adc2295),
	.w3(32'h3ae13fe9),
	.w4(32'h3a131473),
	.w5(32'hba41c7ae),
	.w6(32'h3b216396),
	.w7(32'h38a12566),
	.w8(32'hba60fb80),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62a115),
	.w1(32'hba4b37f2),
	.w2(32'hbabddc2c),
	.w3(32'hba235717),
	.w4(32'hba643837),
	.w5(32'h378af3ea),
	.w6(32'hb9bb6717),
	.w7(32'hba87215e),
	.w8(32'hba2a363d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8517c7),
	.w1(32'h39d31c5d),
	.w2(32'h3a70b9f5),
	.w3(32'hbba655b1),
	.w4(32'h38b92f03),
	.w5(32'hba908ef0),
	.w6(32'hbb598488),
	.w7(32'hba9a3ec1),
	.w8(32'hba3b2224),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39836d77),
	.w1(32'hbb2e8519),
	.w2(32'h39325914),
	.w3(32'hba9592f0),
	.w4(32'h3a540bab),
	.w5(32'hb8f5d0e8),
	.w6(32'hba2cb7fb),
	.w7(32'h3a154d92),
	.w8(32'h3b2b4ca9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a24946),
	.w1(32'h39fad3d8),
	.w2(32'h3b0acd25),
	.w3(32'h39e7a27a),
	.w4(32'hb9b40758),
	.w5(32'hb89955d9),
	.w6(32'h3b0bf36b),
	.w7(32'hba3bfb75),
	.w8(32'hba81f7b8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f0a0a),
	.w1(32'h3b86d19b),
	.w2(32'h3aa15759),
	.w3(32'hb913136b),
	.w4(32'h3ac13093),
	.w5(32'hbb45d66b),
	.w6(32'hba90ef42),
	.w7(32'h3b10014b),
	.w8(32'hba2180af),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f68fc),
	.w1(32'h3a3581da),
	.w2(32'hba5d4dea),
	.w3(32'h3a460031),
	.w4(32'h391767ef),
	.w5(32'h3af34cac),
	.w6(32'h3af8866a),
	.w7(32'hb9d33669),
	.w8(32'h3b007474),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6df4c),
	.w1(32'h3aa7a8cc),
	.w2(32'h3ad5b7b1),
	.w3(32'hbac52507),
	.w4(32'h39b8de67),
	.w5(32'hba8ce2b9),
	.w6(32'hbafbc3d2),
	.w7(32'h3abcd73e),
	.w8(32'h3a5d2504),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae078b8),
	.w1(32'h3b138606),
	.w2(32'h3a03494f),
	.w3(32'h3ad267a4),
	.w4(32'h3b11b56e),
	.w5(32'hba2ba5e5),
	.w6(32'h39cf4c14),
	.w7(32'h3b05bbec),
	.w8(32'h37412712),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4eaee0),
	.w1(32'h3bb3e406),
	.w2(32'h3baf5030),
	.w3(32'h3aab0838),
	.w4(32'h3b970346),
	.w5(32'h3aac1177),
	.w6(32'h3b06891b),
	.w7(32'h3b33c0e3),
	.w8(32'h3b205f46),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf2b4b),
	.w1(32'h3a2f18f1),
	.w2(32'h3898df14),
	.w3(32'h3b8502d4),
	.w4(32'hb868c1a5),
	.w5(32'hb91369cf),
	.w6(32'h3b610ab4),
	.w7(32'hb949e1f0),
	.w8(32'h384210a6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6dfdc),
	.w1(32'h3ab35fce),
	.w2(32'h3a400ed3),
	.w3(32'h389ce0df),
	.w4(32'hb81aa42e),
	.w5(32'hba2f829a),
	.w6(32'h39738899),
	.w7(32'hba8f30c9),
	.w8(32'hba1472b7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b902e3),
	.w1(32'h3afdff1e),
	.w2(32'h3a6fa0ad),
	.w3(32'h36020bfb),
	.w4(32'h3b113fb2),
	.w5(32'hba296739),
	.w6(32'h38da8588),
	.w7(32'h3b3e8359),
	.w8(32'h3b0712b0),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2b191),
	.w1(32'hb9e7f2c9),
	.w2(32'h386bc7ba),
	.w3(32'hba783aa5),
	.w4(32'h3a4b8101),
	.w5(32'h3aa4351b),
	.w6(32'h39301f8f),
	.w7(32'hb938ebb3),
	.w8(32'hbaf88624),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d7926),
	.w1(32'h3b5f3b6c),
	.w2(32'h3a5aba4a),
	.w3(32'hba37cf90),
	.w4(32'h3b331087),
	.w5(32'h3be0ad30),
	.w6(32'hba2e90e7),
	.w7(32'hbab54121),
	.w8(32'h3b442514),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a031ae2),
	.w1(32'h3a10b16b),
	.w2(32'h3a2c7ea4),
	.w3(32'h3b20c7e4),
	.w4(32'h3b1c6374),
	.w5(32'h3b8447f2),
	.w6(32'h3959ca80),
	.w7(32'h3af6d132),
	.w8(32'h3b1372b4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67b150),
	.w1(32'h3a26ea0e),
	.w2(32'h3a9e530c),
	.w3(32'h3aaebdea),
	.w4(32'h3a99ac33),
	.w5(32'h3ad39b94),
	.w6(32'hb8e05f9e),
	.w7(32'hbaee5d21),
	.w8(32'hba2686b5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e00cb),
	.w1(32'hb9b327f8),
	.w2(32'hb945584e),
	.w3(32'h3a2aec48),
	.w4(32'hbaead3a1),
	.w5(32'hbb0ddb4e),
	.w6(32'hba8c87bf),
	.w7(32'h3a64eaf9),
	.w8(32'hb8b44f92),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395443f7),
	.w1(32'hbb90edb3),
	.w2(32'h3a09dcdf),
	.w3(32'hbb02ea67),
	.w4(32'hbb917498),
	.w5(32'h3ae72b30),
	.w6(32'hb9dff5aa),
	.w7(32'hbb54dcc8),
	.w8(32'hb9ec1541),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a670319),
	.w1(32'hba24da71),
	.w2(32'hba8217ae),
	.w3(32'h3b12ff51),
	.w4(32'hba5db0fc),
	.w5(32'h3a6be3fc),
	.w6(32'h3a71f042),
	.w7(32'hba6c96b2),
	.w8(32'hbb18aa1f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7c6ad),
	.w1(32'h3a2896e3),
	.w2(32'h3b138a06),
	.w3(32'h3a4f5c6d),
	.w4(32'h3af804a9),
	.w5(32'h3bb50cf3),
	.w6(32'h3a14dc67),
	.w7(32'h3a696a49),
	.w8(32'h3ac69006),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62958d),
	.w1(32'h39fe4da5),
	.w2(32'h3a69b89d),
	.w3(32'h3b53ea68),
	.w4(32'hbb0d67f1),
	.w5(32'hb7f02427),
	.w6(32'hbad6122d),
	.w7(32'hbb0dde67),
	.w8(32'hba8d0ea4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16bd14),
	.w1(32'h3b24aba4),
	.w2(32'h3b25d2f2),
	.w3(32'hb9bf27d4),
	.w4(32'h3860dd98),
	.w5(32'h3abe6df9),
	.w6(32'hba8254d2),
	.w7(32'h379adc70),
	.w8(32'h3918022d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6ddc3),
	.w1(32'h3ac678b6),
	.w2(32'h3acb012e),
	.w3(32'h3a473a1e),
	.w4(32'h3b1bcb52),
	.w5(32'h3a651ad0),
	.w6(32'hba85cabf),
	.w7(32'h3aabefa8),
	.w8(32'h3a4fa246),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6be84f),
	.w1(32'h3a2d2e34),
	.w2(32'hb92da49f),
	.w3(32'h3a1186b5),
	.w4(32'h39b5b496),
	.w5(32'hbb4ca17d),
	.w6(32'h3acb3948),
	.w7(32'h3a740ab8),
	.w8(32'hb999eab5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b6a43),
	.w1(32'h398d9396),
	.w2(32'hb9956ea6),
	.w3(32'hb9f1766f),
	.w4(32'h3a70b7a9),
	.w5(32'hb9bfcc8f),
	.w6(32'h3a694435),
	.w7(32'hba18b310),
	.w8(32'hbb11a9ef),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934a742),
	.w1(32'h399a43ce),
	.w2(32'h3a653691),
	.w3(32'hba092a18),
	.w4(32'hbad16dd9),
	.w5(32'h3a83eacf),
	.w6(32'hba885d20),
	.w7(32'hba08916a),
	.w8(32'hbb07b3d1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac60805),
	.w1(32'hb931cf6a),
	.w2(32'hbab7646d),
	.w3(32'h3a7d3a0d),
	.w4(32'hbae751a3),
	.w5(32'h3a9e591a),
	.w6(32'hba15ebf9),
	.w7(32'hbb568bfa),
	.w8(32'hbbaaaefb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0bce),
	.w1(32'hbb20e29f),
	.w2(32'hb9d5bb8a),
	.w3(32'hbb0d6dc2),
	.w4(32'hbafc834a),
	.w5(32'hb9523468),
	.w6(32'hbb7ffd80),
	.w7(32'h3ac48b60),
	.w8(32'hb9862515),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff864e),
	.w1(32'hb81d067a),
	.w2(32'h3aa18751),
	.w3(32'hbb205b86),
	.w4(32'hbb288a1b),
	.w5(32'hbaa279e5),
	.w6(32'h3918e5a7),
	.w7(32'hb9a1c485),
	.w8(32'h3954aa43),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac96949),
	.w1(32'hb9428a52),
	.w2(32'h3824b7bf),
	.w3(32'hba051162),
	.w4(32'hba49e3b1),
	.w5(32'h3a3a29ef),
	.w6(32'h3a351494),
	.w7(32'h3af60598),
	.w8(32'h3a4bb007),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8698066),
	.w1(32'h3b81da29),
	.w2(32'h3ae48637),
	.w3(32'h3a707588),
	.w4(32'h3b7073b7),
	.w5(32'hbabf2c9f),
	.w6(32'h3a1b6ca8),
	.w7(32'h3af513c9),
	.w8(32'hba349f92),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb06f7),
	.w1(32'hba6063ed),
	.w2(32'hbad7e59c),
	.w3(32'hbaf2cbb4),
	.w4(32'h3a98d757),
	.w5(32'h3a01eb8e),
	.w6(32'hba891ba9),
	.w7(32'hb9e797d6),
	.w8(32'hba2f801f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a931f0a),
	.w1(32'h3a3946b0),
	.w2(32'h3ad94488),
	.w3(32'h3add4c77),
	.w4(32'h3a334405),
	.w5(32'h39866d69),
	.w6(32'h37641c8d),
	.w7(32'h3ad00a79),
	.w8(32'h3abbae61),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbf0a0),
	.w1(32'h3b0eb265),
	.w2(32'h3b1cac33),
	.w3(32'h3a630083),
	.w4(32'h3a8d8165),
	.w5(32'h3b434f33),
	.w6(32'h3a79ab17),
	.w7(32'h3a14e1e2),
	.w8(32'h3a062eee),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aedbc),
	.w1(32'hba50cbee),
	.w2(32'hbb132708),
	.w3(32'h3a073cad),
	.w4(32'hba96540c),
	.w5(32'hba977468),
	.w6(32'hb83c02b6),
	.w7(32'h39f3bec2),
	.w8(32'h3ab881c0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba877d2f),
	.w1(32'hb907c2d2),
	.w2(32'h3a1f1109),
	.w3(32'h3a5091d3),
	.w4(32'h39e8fa22),
	.w5(32'h3b5fb9c1),
	.w6(32'h3a65e399),
	.w7(32'h3ab790cc),
	.w8(32'h3a4e58f5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a050889),
	.w1(32'h38ac6ec6),
	.w2(32'h3b070ad3),
	.w3(32'h3b094089),
	.w4(32'hb9c0666a),
	.w5(32'h3bb5c9c0),
	.w6(32'h39b38272),
	.w7(32'hb92ceab2),
	.w8(32'h39e1c141),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a842f78),
	.w1(32'h3b041dea),
	.w2(32'h3b454050),
	.w3(32'h3af4c197),
	.w4(32'h3a865eff),
	.w5(32'h3b8ab48a),
	.w6(32'h3a30ba75),
	.w7(32'h3b1d904c),
	.w8(32'h3ad95bd0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d70f3),
	.w1(32'hbb1fa4b6),
	.w2(32'hb9e18dac),
	.w3(32'h3b0db039),
	.w4(32'hbb3ba02a),
	.w5(32'h3a9a891e),
	.w6(32'h3ab9c7f4),
	.w7(32'h3a17704b),
	.w8(32'h3ac257a4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972194),
	.w1(32'h3ac80ea4),
	.w2(32'hb909b6fd),
	.w3(32'h3a933e83),
	.w4(32'h3b12630e),
	.w5(32'h3b951795),
	.w6(32'h39f65489),
	.w7(32'hb99d3095),
	.w8(32'h3afe1135),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71efda),
	.w1(32'h3a80d611),
	.w2(32'h39b60e81),
	.w3(32'hba5cede9),
	.w4(32'h3aafa555),
	.w5(32'hb9d52bfb),
	.w6(32'h3abd05b5),
	.w7(32'hba14e16d),
	.w8(32'hbad9cf4b),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84b576),
	.w1(32'hba49e116),
	.w2(32'h39c9a69d),
	.w3(32'hbae36918),
	.w4(32'hba622029),
	.w5(32'hbb3205a0),
	.w6(32'hbb147652),
	.w7(32'h39d74586),
	.w8(32'h3a6146e2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993d10c),
	.w1(32'h3a255342),
	.w2(32'hba647e9a),
	.w3(32'hba111f5d),
	.w4(32'h3afffe8c),
	.w5(32'h3b11a21a),
	.w6(32'hba3c594a),
	.w7(32'h380451be),
	.w8(32'hb9b04cdc),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb292ec9),
	.w1(32'h3ad04d1b),
	.w2(32'h3a2259be),
	.w3(32'hbaf93aa5),
	.w4(32'h397e768a),
	.w5(32'hb9e099bd),
	.w6(32'hbb2707b8),
	.w7(32'h3abcf793),
	.w8(32'h3a07f652),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13b457),
	.w1(32'h3a1e5fb1),
	.w2(32'hb9c2635b),
	.w3(32'hb8eebe7f),
	.w4(32'h3a9c0420),
	.w5(32'h3b624fdc),
	.w6(32'h3ad81666),
	.w7(32'h3abb5818),
	.w8(32'hb8dd4325),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0faa41),
	.w1(32'h3a5f2fe6),
	.w2(32'h3a2b5a17),
	.w3(32'h3a9063ee),
	.w4(32'hba859589),
	.w5(32'h3919170e),
	.w6(32'hb930b512),
	.w7(32'hba809c0a),
	.w8(32'hbb05cf20),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b2034),
	.w1(32'h3b190d67),
	.w2(32'h399b7476),
	.w3(32'hb93ba96b),
	.w4(32'h3a94132c),
	.w5(32'hba85cd35),
	.w6(32'hbade98c1),
	.w7(32'hba16b7ca),
	.w8(32'h3a0e97d0),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925ae46),
	.w1(32'h3b6441b2),
	.w2(32'h3a8b71f8),
	.w3(32'hbac930c9),
	.w4(32'h3b3bf47c),
	.w5(32'h3ab7b689),
	.w6(32'hb73ece5d),
	.w7(32'h3b275273),
	.w8(32'h39e8498a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c0de8),
	.w1(32'h3b521db0),
	.w2(32'h3a82fdfd),
	.w3(32'h39735de7),
	.w4(32'h38da1537),
	.w5(32'hbb34d320),
	.w6(32'h390584c0),
	.w7(32'h3a87d798),
	.w8(32'hb989231c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff70ca),
	.w1(32'h38a9f885),
	.w2(32'h3ab290be),
	.w3(32'hba787597),
	.w4(32'h3b3546a7),
	.w5(32'h3bb56421),
	.w6(32'h3ab7ceb7),
	.w7(32'h3ae01ecb),
	.w8(32'h3a995ce9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a1c12d),
	.w1(32'hb967ad3e),
	.w2(32'hbabd676a),
	.w3(32'h3b27dd93),
	.w4(32'h38e70258),
	.w5(32'hbb38d40e),
	.w6(32'hb983e33b),
	.w7(32'h3a409568),
	.w8(32'hba45bf21),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d04dfa),
	.w1(32'hbb03379a),
	.w2(32'hba324891),
	.w3(32'hb7afc601),
	.w4(32'hba6633d6),
	.w5(32'h39e53af9),
	.w6(32'h3a25ff5e),
	.w7(32'hba648a9c),
	.w8(32'h38ac0926),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc7eff),
	.w1(32'hba862724),
	.w2(32'h399ade73),
	.w3(32'hbaa0d6be),
	.w4(32'hbace93da),
	.w5(32'h3a9b1a70),
	.w6(32'hbabc3204),
	.w7(32'hb8c2865b),
	.w8(32'hba6826c7),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dc9a7),
	.w1(32'h39af8d90),
	.w2(32'hba3c9c99),
	.w3(32'hbaa91385),
	.w4(32'hb9cbc2de),
	.w5(32'hbadb6de0),
	.w6(32'h3981f602),
	.w7(32'h394678ae),
	.w8(32'h3a6d0bb8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9901a36),
	.w1(32'hbb2cb9c6),
	.w2(32'hbb26aa1c),
	.w3(32'hb8d69a89),
	.w4(32'h37074389),
	.w5(32'h3b804dbc),
	.w6(32'hb9801b6d),
	.w7(32'hbaddd3b7),
	.w8(32'h3ab2c343),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb365e48),
	.w1(32'h3adc4147),
	.w2(32'h3afa1c55),
	.w3(32'h3aa88ff3),
	.w4(32'h3a5ac101),
	.w5(32'h3968c0b8),
	.w6(32'hb957747d),
	.w7(32'h3a0abd12),
	.w8(32'h39d78fe0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bbf6b7),
	.w1(32'h3b3bede2),
	.w2(32'h3b0baf87),
	.w3(32'h3aac5d1b),
	.w4(32'h3abad5a5),
	.w5(32'hb94140b7),
	.w6(32'h3a841995),
	.w7(32'h3a43332f),
	.w8(32'h3b06a7ae),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a064c99),
	.w1(32'hba37ce49),
	.w2(32'hba47aec3),
	.w3(32'h3aa78831),
	.w4(32'h3a0b32a7),
	.w5(32'h3a95a773),
	.w6(32'h3ac7b84b),
	.w7(32'hb9e561e2),
	.w8(32'h3951f654),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84f6d2),
	.w1(32'h39e52c0c),
	.w2(32'h3a08c076),
	.w3(32'hb8a7c04e),
	.w4(32'h3a087703),
	.w5(32'h3a6765e6),
	.w6(32'hbaf599ba),
	.w7(32'h3ade6247),
	.w8(32'h3ae33657),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b062e21),
	.w1(32'hbaaa2266),
	.w2(32'h3b12641f),
	.w3(32'h3a5e110d),
	.w4(32'hba85d97f),
	.w5(32'hbac7a392),
	.w6(32'h3a551f8c),
	.w7(32'hb91fb013),
	.w8(32'hba599298),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c0445),
	.w1(32'hba099ec9),
	.w2(32'h39a58dd7),
	.w3(32'hbab2c8f8),
	.w4(32'h3880e752),
	.w5(32'h3ad8237b),
	.w6(32'hbae1ea23),
	.w7(32'hba56563e),
	.w8(32'hb8d4521a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1403c2),
	.w1(32'hba057dca),
	.w2(32'hb9e27899),
	.w3(32'h3a95924b),
	.w4(32'hb920484f),
	.w5(32'h3ac94cbf),
	.w6(32'h3a8b8b6a),
	.w7(32'hb81644e9),
	.w8(32'h3abf4149),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88a125),
	.w1(32'h3ae6390c),
	.w2(32'h3ad16ccb),
	.w3(32'h3accad8e),
	.w4(32'h3a94073d),
	.w5(32'hbacb869d),
	.w6(32'h3a1d96a3),
	.w7(32'hba8cf7bb),
	.w8(32'hba8f767c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0d3bb),
	.w1(32'h3a6b1818),
	.w2(32'h3a4f741c),
	.w3(32'hba10e51a),
	.w4(32'hbb11c220),
	.w5(32'hba559d25),
	.w6(32'h385ed7dc),
	.w7(32'hbb692344),
	.w8(32'hbb190147),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8350f3),
	.w1(32'h3ab01a4e),
	.w2(32'h3b299925),
	.w3(32'hba7418de),
	.w4(32'h3aae6b14),
	.w5(32'h3aa2304f),
	.w6(32'hbb2e1618),
	.w7(32'h39905b31),
	.w8(32'hba71a99f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a426f54),
	.w1(32'hbaf9de46),
	.w2(32'hba99be76),
	.w3(32'hb9f2eece),
	.w4(32'hba0bcf2a),
	.w5(32'h3addb5c8),
	.w6(32'hbadc57dc),
	.w7(32'hbaf78144),
	.w8(32'hba258756),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa165f6),
	.w1(32'h3a139bf2),
	.w2(32'h3a0e4102),
	.w3(32'hb9d0ea98),
	.w4(32'hba5966e5),
	.w5(32'h3aa1ac06),
	.w6(32'hbaba8ded),
	.w7(32'h3a84c1f9),
	.w8(32'hb98dcd70),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade9727),
	.w1(32'h3b84656c),
	.w2(32'h3b10aab7),
	.w3(32'h3a694739),
	.w4(32'h3b1d0deb),
	.w5(32'hbac58747),
	.w6(32'h39ef81e9),
	.w7(32'h3b2976b8),
	.w8(32'h39afa4f8),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90f69d),
	.w1(32'hba025a59),
	.w2(32'hbac76d63),
	.w3(32'hbb3967cc),
	.w4(32'hb8d177e2),
	.w5(32'hbb090c60),
	.w6(32'h3948af21),
	.w7(32'hba1886e0),
	.w8(32'h3a0a110a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0dd61),
	.w1(32'h390eb3ba),
	.w2(32'h3a9dccc4),
	.w3(32'hb9fbff72),
	.w4(32'h3a6dce87),
	.w5(32'h3acf24da),
	.w6(32'h3791c459),
	.w7(32'h3a826555),
	.w8(32'h3aada638),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad05495),
	.w1(32'hb9890b63),
	.w2(32'hb9919193),
	.w3(32'h396a9014),
	.w4(32'h3a67fdab),
	.w5(32'h3aac4117),
	.w6(32'hb992cf3d),
	.w7(32'h3abff37d),
	.w8(32'hba2ed1a5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd323d),
	.w1(32'h3a975815),
	.w2(32'h399d5772),
	.w3(32'h39dc8469),
	.w4(32'hb9a40722),
	.w5(32'hbb282a57),
	.w6(32'h3a8d1356),
	.w7(32'h3a99f95b),
	.w8(32'hba238bed),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbb605),
	.w1(32'h3ab5f461),
	.w2(32'hba1a488a),
	.w3(32'h39f3e746),
	.w4(32'h3a396a61),
	.w5(32'hb979f61a),
	.w6(32'h3b041a58),
	.w7(32'h3a9ebb0b),
	.w8(32'h390da6bb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04305f),
	.w1(32'h3a36f952),
	.w2(32'h39bc5827),
	.w3(32'hba8e5d65),
	.w4(32'hbaca2e6f),
	.w5(32'hbb53ef73),
	.w6(32'h3a728030),
	.w7(32'hb9b75c69),
	.w8(32'hbaa21c09),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada2ad7),
	.w1(32'h3a516827),
	.w2(32'hb9e84900),
	.w3(32'h3a2fd962),
	.w4(32'h3abdb919),
	.w5(32'hb8608a97),
	.w6(32'h3a3b2502),
	.w7(32'h3a9de3d8),
	.w8(32'hba702209),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c8be8),
	.w1(32'h3b41d9ee),
	.w2(32'h3ab4655c),
	.w3(32'hba835ff0),
	.w4(32'h3ab8927b),
	.w5(32'h3b22d4ee),
	.w6(32'hb97f1356),
	.w7(32'h3a529a83),
	.w8(32'h3b804fc2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfcb10),
	.w1(32'hba976ef2),
	.w2(32'hbb22dbe9),
	.w3(32'hbabcdc2f),
	.w4(32'hb9137783),
	.w5(32'h3a06c659),
	.w6(32'h3ab9873d),
	.w7(32'hb9f1be18),
	.w8(32'h3a1e6b6a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba386309),
	.w1(32'h3b5dc794),
	.w2(32'h3a6477b1),
	.w3(32'h3b003aac),
	.w4(32'h3b355564),
	.w5(32'h3b1e8c65),
	.w6(32'h3a5990ed),
	.w7(32'h3b0681f7),
	.w8(32'h3a4fc31c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397927dc),
	.w1(32'hb9f243eb),
	.w2(32'h3a52e023),
	.w3(32'h3b413382),
	.w4(32'hb9a00814),
	.w5(32'h397a9e91),
	.w6(32'h3aa034f8),
	.w7(32'h3a6c3e85),
	.w8(32'h3a3e7ea8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98487d),
	.w1(32'hba667f82),
	.w2(32'hbb3824fa),
	.w3(32'hbb0dcf63),
	.w4(32'hb9763ddc),
	.w5(32'hba611329),
	.w6(32'h3a82640d),
	.w7(32'h3abfe3d3),
	.w8(32'h3a3e8b51),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6696a8),
	.w1(32'h388c5511),
	.w2(32'h395cfdc2),
	.w3(32'hb98bb0a5),
	.w4(32'h3af25b03),
	.w5(32'h3be9c780),
	.w6(32'h3aaa3f37),
	.w7(32'h3b3095b4),
	.w8(32'h3b47b637),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eb013),
	.w1(32'hbb645f2c),
	.w2(32'hbac234f9),
	.w3(32'h3afe88d9),
	.w4(32'hb9273a57),
	.w5(32'h3bf51697),
	.w6(32'h3ab06fa0),
	.w7(32'hbb20181b),
	.w8(32'hb9a8415d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7e05c),
	.w1(32'hbae55f57),
	.w2(32'hbb68a85b),
	.w3(32'hbb2fee58),
	.w4(32'hbb03f06e),
	.w5(32'hbb4f2827),
	.w6(32'hbb99c58b),
	.w7(32'hbb0e70b0),
	.w8(32'hbb16f10a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5405),
	.w1(32'hb9f43d92),
	.w2(32'h3a53804e),
	.w3(32'hbae42916),
	.w4(32'hb9c0f7bc),
	.w5(32'h39b2917f),
	.w6(32'hbb567eea),
	.w7(32'hbaaaf4ff),
	.w8(32'hba913979),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00fefb),
	.w1(32'h3b123413),
	.w2(32'h3a952335),
	.w3(32'hbadddd06),
	.w4(32'h3ad26dff),
	.w5(32'h3a0ba14e),
	.w6(32'hbae62aa9),
	.w7(32'h3b15ca57),
	.w8(32'h3b65cc4b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435af8),
	.w1(32'hb90de80f),
	.w2(32'h39823c67),
	.w3(32'h3b4862a7),
	.w4(32'hbac776a3),
	.w5(32'h3aac59a9),
	.w6(32'h3adb0205),
	.w7(32'hba5f8d90),
	.w8(32'h3a9b845e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac729fe),
	.w1(32'h3b08341d),
	.w2(32'hb9200113),
	.w3(32'h3aac9909),
	.w4(32'h3ab90e2f),
	.w5(32'hba794ca9),
	.w6(32'h3a46f645),
	.w7(32'h3a807559),
	.w8(32'h3a315521),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a73a511),
	.w1(32'hba36b30a),
	.w2(32'hb97fa72c),
	.w3(32'h39bb39c8),
	.w4(32'h39beb61a),
	.w5(32'h3aa22b25),
	.w6(32'h3afb8c1f),
	.w7(32'h3a586023),
	.w8(32'h3a32dd65),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1d99a),
	.w1(32'h3a839ac3),
	.w2(32'h39b30280),
	.w3(32'h385be456),
	.w4(32'hb970c57d),
	.w5(32'h39ff9d82),
	.w6(32'h3a37c66a),
	.w7(32'hbab900d0),
	.w8(32'hb9b7d2a6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a956697),
	.w1(32'hba1145a9),
	.w2(32'h395fddf6),
	.w3(32'h39fbaeea),
	.w4(32'hbad6fc04),
	.w5(32'hb9890673),
	.w6(32'hbac92d1d),
	.w7(32'hbb3d650f),
	.w8(32'hbb2055c1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88b235),
	.w1(32'h3b2910e9),
	.w2(32'h3b0a5366),
	.w3(32'hbb1078ca),
	.w4(32'hb98cb79a),
	.w5(32'hb910afcb),
	.w6(32'hba8f76f2),
	.w7(32'hbb67d6a2),
	.w8(32'hbb522e73),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86ec6d),
	.w1(32'h3ae4577d),
	.w2(32'h3b04e338),
	.w3(32'hb97142af),
	.w4(32'h3991482a),
	.w5(32'hba205bd1),
	.w6(32'hbafdb10a),
	.w7(32'h3a43eb6b),
	.w8(32'h3990de7a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae63ba2),
	.w1(32'h3b08b6a5),
	.w2(32'h3b18f227),
	.w3(32'h3adaf039),
	.w4(32'h3b114c79),
	.w5(32'h3afdfb80),
	.w6(32'h398fc63f),
	.w7(32'h3b4a4a57),
	.w8(32'h3b0388f6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432caa),
	.w1(32'h3ae186ed),
	.w2(32'h3af8ec6c),
	.w3(32'h3adc2a89),
	.w4(32'h3aa1d0d1),
	.w5(32'h3a861e5f),
	.w6(32'h3b10d6e2),
	.w7(32'h3a822392),
	.w8(32'h3a1f7a29),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7df254),
	.w1(32'h3a912f97),
	.w2(32'h3a382b94),
	.w3(32'h3abb9e87),
	.w4(32'h3a486edf),
	.w5(32'h3ad26aff),
	.w6(32'hb83ef0de),
	.w7(32'h3a106f21),
	.w8(32'h39184f09),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70c851),
	.w1(32'hba9aff09),
	.w2(32'hb9501b37),
	.w3(32'h3ac195d7),
	.w4(32'h3ac7f7ff),
	.w5(32'h3b137686),
	.w6(32'h3977c150),
	.w7(32'h397d1713),
	.w8(32'h399662e9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a2892),
	.w1(32'h3b420528),
	.w2(32'h3ab77e4a),
	.w3(32'hbad2423f),
	.w4(32'h3b0c5e45),
	.w5(32'hba85c56f),
	.w6(32'hbac2e7f3),
	.w7(32'h3b6ae4d3),
	.w8(32'h3b38ff65),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa62238),
	.w1(32'h391b3291),
	.w2(32'hba6a002a),
	.w3(32'h3ad450fc),
	.w4(32'hba1efabe),
	.w5(32'hbb0bd7f1),
	.w6(32'h3a398cfb),
	.w7(32'hb9629f8d),
	.w8(32'hbb0b98aa),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961662a),
	.w1(32'hbad11f2b),
	.w2(32'h3aaad940),
	.w3(32'hba15432b),
	.w4(32'hbac9148c),
	.w5(32'hba8fde3c),
	.w6(32'hb82a02e3),
	.w7(32'hb9f550a1),
	.w8(32'h39acbaf5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5799e2),
	.w1(32'h3aca6b58),
	.w2(32'h3b245718),
	.w3(32'h3ad777d2),
	.w4(32'h3aac9113),
	.w5(32'h3ab7cdcf),
	.w6(32'h39f5a8b2),
	.w7(32'h3a91e200),
	.w8(32'h3afd1913),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6610d6),
	.w1(32'h3988f3f3),
	.w2(32'hbaa2a728),
	.w3(32'h39fbf859),
	.w4(32'h382d8031),
	.w5(32'hbb3327ae),
	.w6(32'h3a777549),
	.w7(32'hb9b8742a),
	.w8(32'hbaf65688),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fcddf4),
	.w1(32'h3b1d02e1),
	.w2(32'h3a9e12d0),
	.w3(32'hbb141286),
	.w4(32'hb8f94c34),
	.w5(32'hba36ca04),
	.w6(32'hba07478c),
	.w7(32'h3b1f1e06),
	.w8(32'h39b128ee),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b5f13),
	.w1(32'h3b3656b1),
	.w2(32'h3b373d66),
	.w3(32'h3a3d0dda),
	.w4(32'h3b094314),
	.w5(32'h3bbf3104),
	.w6(32'h3b319eb6),
	.w7(32'h3aedc6fd),
	.w8(32'h3b151765),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7e961),
	.w1(32'h3b029a89),
	.w2(32'h39bb85d6),
	.w3(32'h3afb6b36),
	.w4(32'hb9ff41c3),
	.w5(32'h39b61c80),
	.w6(32'h397b59cf),
	.w7(32'hba928d24),
	.w8(32'h39162f3a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41e313),
	.w1(32'hba778346),
	.w2(32'hb9c89b84),
	.w3(32'h39d8323a),
	.w4(32'hbab482fe),
	.w5(32'h3afbc269),
	.w6(32'hb8ee7723),
	.w7(32'hbabd7eff),
	.w8(32'h39bb9c81),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0951f2),
	.w1(32'h3ae01289),
	.w2(32'hbaa3ef97),
	.w3(32'h3a21987e),
	.w4(32'h3ac585f9),
	.w5(32'h3ab45363),
	.w6(32'hba0ed9ab),
	.w7(32'h3af6a181),
	.w8(32'h3afe7428),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f22ba),
	.w1(32'h3a7ecfda),
	.w2(32'hbb0d80ef),
	.w3(32'h399ada5f),
	.w4(32'h3acf3042),
	.w5(32'hbb2c9256),
	.w6(32'hb98de335),
	.w7(32'h3ad78fd0),
	.w8(32'hba2aec8e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926bb1),
	.w1(32'h3ab46248),
	.w2(32'h3a22342d),
	.w3(32'hbace3c91),
	.w4(32'h3a8ec67c),
	.w5(32'h39e52395),
	.w6(32'hba7ac673),
	.w7(32'h3a936464),
	.w8(32'hbb0ff7d3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b366c),
	.w1(32'h39da131e),
	.w2(32'h39be8228),
	.w3(32'h3b0578f4),
	.w4(32'hb98bba0d),
	.w5(32'hb8568dc4),
	.w6(32'hb9cd46c1),
	.w7(32'hbb682041),
	.w8(32'hbb007143),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd84e5),
	.w1(32'h39eb493a),
	.w2(32'h3a9041ed),
	.w3(32'hba9949ea),
	.w4(32'hb98e95ba),
	.w5(32'h3ab8af68),
	.w6(32'hbb0a4ed3),
	.w7(32'hbb29ff56),
	.w8(32'hbad47065),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a346261),
	.w1(32'hb9b93d33),
	.w2(32'h3922f4fb),
	.w3(32'h3aac83d2),
	.w4(32'hba396a45),
	.w5(32'h3b354e32),
	.w6(32'hbb0eb35b),
	.w7(32'hbab25698),
	.w8(32'hb903a0d3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb123f3f),
	.w1(32'hba169399),
	.w2(32'h3a33797f),
	.w3(32'hbb07be04),
	.w4(32'h3b40f20f),
	.w5(32'h3b122b26),
	.w6(32'hbaf35f17),
	.w7(32'h3ae18be6),
	.w8(32'h3afcef1e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cba4f6),
	.w1(32'hbaed4381),
	.w2(32'hbadd52a3),
	.w3(32'h3ae94c14),
	.w4(32'hba41d80d),
	.w5(32'hbb038b56),
	.w6(32'hb95afda4),
	.w7(32'hb8139678),
	.w8(32'h3a26d5dd),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9c4c4),
	.w1(32'hbaeff2f8),
	.w2(32'hb98db28d),
	.w3(32'h3922d2a7),
	.w4(32'hbab19030),
	.w5(32'h3b8c5d7f),
	.w6(32'hb9348d69),
	.w7(32'hba85da8e),
	.w8(32'h3ab24e7a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78398e6),
	.w1(32'hbb26ef42),
	.w2(32'hb86bdba3),
	.w3(32'hb8e89fc9),
	.w4(32'hba7ff1bf),
	.w5(32'hba871139),
	.w6(32'h3a079b49),
	.w7(32'hbb1fe810),
	.w8(32'h39f290bb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97a86a),
	.w1(32'h3a0581ca),
	.w2(32'h39589954),
	.w3(32'h37a2ca44),
	.w4(32'h3b064ee3),
	.w5(32'h3bf8fe1a),
	.w6(32'hb982cfd6),
	.w7(32'h3a9fe98a),
	.w8(32'h3a6e0acd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39036077),
	.w1(32'hbb3a1122),
	.w2(32'hbb8c673c),
	.w3(32'h3b2c12ce),
	.w4(32'h39577dce),
	.w5(32'h3b8104e3),
	.w6(32'h3a60a3d7),
	.w7(32'h385b98dd),
	.w8(32'h381fccb8),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb761cce),
	.w1(32'hb80f7a39),
	.w2(32'h3918e6d4),
	.w3(32'h396cf963),
	.w4(32'h39be5272),
	.w5(32'h3adee5c1),
	.w6(32'hbaef2908),
	.w7(32'h3a3a7dd6),
	.w8(32'hb9f5b104),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95cf9a6),
	.w1(32'hb90ffbd3),
	.w2(32'h38fae308),
	.w3(32'hba9b5307),
	.w4(32'hb80b1286),
	.w5(32'hbaa4afed),
	.w6(32'hba4a7c2d),
	.w7(32'h3aaaace5),
	.w8(32'h3875ad04),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1323f9),
	.w1(32'h3aa0990f),
	.w2(32'hba7090c7),
	.w3(32'h3a4329e4),
	.w4(32'h39a16ddb),
	.w5(32'hbb2d4050),
	.w6(32'hb9375ca1),
	.w7(32'h3a8ad273),
	.w8(32'h385c8176),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2af06d),
	.w1(32'h3b414d25),
	.w2(32'h3b661604),
	.w3(32'hbb357a16),
	.w4(32'h3b1ad80e),
	.w5(32'h39c73b2f),
	.w6(32'h3a1e97c4),
	.w7(32'h3b0b6188),
	.w8(32'h3af3abb2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b773831),
	.w1(32'h3ac16e38),
	.w2(32'h3ac6fed2),
	.w3(32'h3b30e1be),
	.w4(32'h3a92bf49),
	.w5(32'hb80fd3a5),
	.w6(32'h3b0f29de),
	.w7(32'h3a57d752),
	.w8(32'hbab1e76c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a69103),
	.w1(32'h3a87e5d1),
	.w2(32'h3a2524a7),
	.w3(32'h39f1b6da),
	.w4(32'h3aaa60ee),
	.w5(32'h3b80c94d),
	.w6(32'hb923334e),
	.w7(32'h392c1c4f),
	.w8(32'hba42f4cb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a6711),
	.w1(32'h39aef458),
	.w2(32'hba2725d6),
	.w3(32'h39fd16a0),
	.w4(32'hbb327918),
	.w5(32'h3a848c09),
	.w6(32'hbaee9ed6),
	.w7(32'hbaa3f1ea),
	.w8(32'hbb3d1081),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6982fb),
	.w1(32'h3add9177),
	.w2(32'h398d4df3),
	.w3(32'hbb0d394c),
	.w4(32'h3aef9780),
	.w5(32'h39e5eace),
	.w6(32'hbad5c6b1),
	.w7(32'hb92dd549),
	.w8(32'h3aba9613),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97ca40),
	.w1(32'hbb0f6cdd),
	.w2(32'hbb227883),
	.w3(32'h38ef5cb8),
	.w4(32'hbb4b8349),
	.w5(32'hbc034a5b),
	.w6(32'hba088299),
	.w7(32'h3b6fe43a),
	.w8(32'h3ba819c9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e5b1f),
	.w1(32'h38a8140c),
	.w2(32'h3acbcdbc),
	.w3(32'h3a44e38f),
	.w4(32'h3b86b24a),
	.w5(32'h3b47b4a8),
	.w6(32'h3b941db5),
	.w7(32'hbb857653),
	.w8(32'hbb6fd76f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb1683),
	.w1(32'h3c0f3392),
	.w2(32'h3c26b463),
	.w3(32'h3a92c049),
	.w4(32'hbbfa02ec),
	.w5(32'hbb9ff542),
	.w6(32'hbb70e3dd),
	.w7(32'hbb24c245),
	.w8(32'h3b3219ac),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba14a51),
	.w1(32'hbab43bc0),
	.w2(32'h3b5dadd9),
	.w3(32'h3993b6b7),
	.w4(32'hbb1a3673),
	.w5(32'h3a6e9e21),
	.w6(32'h3af5b877),
	.w7(32'h3b00f692),
	.w8(32'h3b2f1a7e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb9463),
	.w1(32'hbbf265ca),
	.w2(32'hbbcb26a8),
	.w3(32'h3b97500d),
	.w4(32'h3a5dd4ef),
	.w5(32'h3bcff1c8),
	.w6(32'h3bb11d14),
	.w7(32'h3b05d437),
	.w8(32'h3b3ec3ec),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e30f6),
	.w1(32'hbae58d6d),
	.w2(32'h3b832ff6),
	.w3(32'h3adf0b14),
	.w4(32'hbb69bcac),
	.w5(32'hbb676985),
	.w6(32'hba0c4c60),
	.w7(32'hbba17a4c),
	.w8(32'hbbf6c158),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad509fa),
	.w1(32'h3b098130),
	.w2(32'h3b192ac1),
	.w3(32'hbb97a388),
	.w4(32'hbb8cde63),
	.w5(32'hbb88c337),
	.w6(32'hbbf0a42f),
	.w7(32'h3a764c80),
	.w8(32'h3a9c5d87),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04ef4b),
	.w1(32'h3b8030e8),
	.w2(32'h3b6aeabc),
	.w3(32'hbb908ab6),
	.w4(32'hba3c5630),
	.w5(32'h3a24a1ec),
	.w6(32'hbaaa0751),
	.w7(32'h3b327379),
	.w8(32'h3bba9f54),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35fcd),
	.w1(32'hbc980485),
	.w2(32'hbc66bb1a),
	.w3(32'h3bcb8b92),
	.w4(32'h3c2d3e20),
	.w5(32'h3ca00503),
	.w6(32'h3c0a0860),
	.w7(32'hbb7a023e),
	.w8(32'hbb37df1d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff754b),
	.w1(32'hbb9cbffa),
	.w2(32'hbae7b51f),
	.w3(32'hbba3b9c9),
	.w4(32'h3b4daa8f),
	.w5(32'h38eab84e),
	.w6(32'h3bf83757),
	.w7(32'h3aac731d),
	.w8(32'hba375569),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc59e7b),
	.w1(32'hba0d8763),
	.w2(32'h3a8a9f5d),
	.w3(32'h3bbe0fba),
	.w4(32'h3b1139af),
	.w5(32'hbc14cb79),
	.w6(32'h3c094436),
	.w7(32'hb96d47e3),
	.w8(32'hb9b0fab4),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745526),
	.w1(32'h3bdda91a),
	.w2(32'h3a84ed2d),
	.w3(32'hbac15d63),
	.w4(32'h3c1ab3bf),
	.w5(32'h3c03f673),
	.w6(32'h3a6f9030),
	.w7(32'h3c48fb11),
	.w8(32'h3b98547c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41e450),
	.w1(32'hba821dff),
	.w2(32'h3a980d48),
	.w3(32'h3c4041e3),
	.w4(32'hb9bdb0d6),
	.w5(32'h3b229bc5),
	.w6(32'h3c05134f),
	.w7(32'h39022f65),
	.w8(32'h3b79351d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83d426),
	.w1(32'hba9d0200),
	.w2(32'hb9644f0f),
	.w3(32'h3ae8bd18),
	.w4(32'hbb6008c9),
	.w5(32'hbbd99fbd),
	.w6(32'h3b45cb16),
	.w7(32'h3a13e952),
	.w8(32'h3b26f0d9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e4a78),
	.w1(32'h3bd9d9cc),
	.w2(32'h3bf0f4bd),
	.w3(32'hbb2b3df2),
	.w4(32'hba24cc57),
	.w5(32'hba5bc6e9),
	.w6(32'hb9b9a078),
	.w7(32'h3b424470),
	.w8(32'h3b501fcf),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc89929),
	.w1(32'h3bed7020),
	.w2(32'h3bf8847c),
	.w3(32'h3b837bf1),
	.w4(32'hbb0825fd),
	.w5(32'hba9603a7),
	.w6(32'hbaaf2565),
	.w7(32'h3b3441b4),
	.w8(32'h3b8b0423),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0decf6),
	.w1(32'h3b2d2c92),
	.w2(32'h3bbc858b),
	.w3(32'h3a479c80),
	.w4(32'h3a346bc5),
	.w5(32'h3af39071),
	.w6(32'hbaad80c0),
	.w7(32'hbb3921f3),
	.w8(32'hbb6e1a50),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5737e8),
	.w1(32'hbc2ceae0),
	.w2(32'hbc4024b6),
	.w3(32'h3ba0b928),
	.w4(32'h3c4f416f),
	.w5(32'h3c6b5a7a),
	.w6(32'hb98d505c),
	.w7(32'hbbd3ae97),
	.w8(32'hbb1fad98),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42d927),
	.w1(32'hbc125e71),
	.w2(32'hbc251203),
	.w3(32'h3ba75de7),
	.w4(32'h3b87d614),
	.w5(32'h3c88c987),
	.w6(32'h3c559e2b),
	.w7(32'hbb98499b),
	.w8(32'hbbf35cfc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f6d8),
	.w1(32'hbb232ea5),
	.w2(32'hbb26dc2e),
	.w3(32'h3acf9400),
	.w4(32'hbc17e2f5),
	.w5(32'hbbe6e7a2),
	.w6(32'hbab31920),
	.w7(32'h3b92f1c7),
	.w8(32'h3bbe20fc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a405c2b),
	.w1(32'hbb01d075),
	.w2(32'hbae16814),
	.w3(32'hbbf42d31),
	.w4(32'h3b748b53),
	.w5(32'h3b5393b6),
	.w6(32'hba94cdd2),
	.w7(32'hb9cd2ade),
	.w8(32'h3b8accab),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c48d),
	.w1(32'hbb24b062),
	.w2(32'h3bacada5),
	.w3(32'hbb664075),
	.w4(32'hbbc16f7f),
	.w5(32'hbabe86fd),
	.w6(32'hb8e7766c),
	.w7(32'hbb01de94),
	.w8(32'h3b2106dc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0652c),
	.w1(32'hbbd9659c),
	.w2(32'hb7b9b933),
	.w3(32'h3b20bf82),
	.w4(32'h3b18b1cf),
	.w5(32'h3b13e0ac),
	.w6(32'h3940a95a),
	.w7(32'hbb3b1737),
	.w8(32'hbbcced48),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa370fa),
	.w1(32'h3bec9fdd),
	.w2(32'h3c4d2fe4),
	.w3(32'h3b7e6fbb),
	.w4(32'hbc2172cf),
	.w5(32'hbc5e591f),
	.w6(32'hbb2f769e),
	.w7(32'h3aef15bd),
	.w8(32'h39964273),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c575ec5),
	.w1(32'hbabe75d1),
	.w2(32'hbb82a626),
	.w3(32'hbbae21e6),
	.w4(32'h3ac701f8),
	.w5(32'hbaeb1fed),
	.w6(32'h39850954),
	.w7(32'h3b5e1747),
	.w8(32'h39454aff),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d97c7),
	.w1(32'hbb43818e),
	.w2(32'hbac3ab6c),
	.w3(32'h3b8a074f),
	.w4(32'h3ba51a16),
	.w5(32'hbb1f9e34),
	.w6(32'h3b519e79),
	.w7(32'h3ba7e504),
	.w8(32'h3b459467),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09e02d),
	.w1(32'hbbaa6e51),
	.w2(32'hbb2356a1),
	.w3(32'h3b5b9b0c),
	.w4(32'hbc042202),
	.w5(32'hbc2b970e),
	.w6(32'h3c03c8be),
	.w7(32'h3b671dfa),
	.w8(32'h3b91ee4d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc746b15),
	.w1(32'hbb770bae),
	.w2(32'hbb16c3cd),
	.w3(32'h3b1e2a72),
	.w4(32'hbb78f02a),
	.w5(32'hbb09c9a5),
	.w6(32'hbbcfd913),
	.w7(32'h3b9db92f),
	.w8(32'h3b816429),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79e91f),
	.w1(32'h3bacf3ab),
	.w2(32'h3b59f6c1),
	.w3(32'h3ada74cd),
	.w4(32'h3baba7ae),
	.w5(32'h3b98746e),
	.w6(32'hbb1fc016),
	.w7(32'h3c06644a),
	.w8(32'h3c1dce2f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8b333),
	.w1(32'h3b54ddca),
	.w2(32'h3bc9bae3),
	.w3(32'h3a9bf341),
	.w4(32'hb9066cad),
	.w5(32'hba571f7f),
	.w6(32'h3c04ab5e),
	.w7(32'h3c1f34a2),
	.w8(32'h3bd821ad),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb501a),
	.w1(32'h3b3a64be),
	.w2(32'h3bf7418e),
	.w3(32'h3a9cee03),
	.w4(32'hbba90169),
	.w5(32'hbb51439c),
	.w6(32'h3ba73bb2),
	.w7(32'h39da0c62),
	.w8(32'hbb0e166e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7454),
	.w1(32'hbbc82e53),
	.w2(32'hbbc33d01),
	.w3(32'hbc227144),
	.w4(32'h39fc7857),
	.w5(32'hbaeb6c15),
	.w6(32'h3b03ba91),
	.w7(32'h3c0bc325),
	.w8(32'h3c44d23d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef2e3b),
	.w1(32'h3a9ad92a),
	.w2(32'hba55d5fc),
	.w3(32'hba2be917),
	.w4(32'hbba85643),
	.w5(32'hbbc98586),
	.w6(32'h3bdb211b),
	.w7(32'h39bc3071),
	.w8(32'hba8a8f0e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb358752),
	.w1(32'h3ba2eede),
	.w2(32'h3af3743f),
	.w3(32'h3bbb6a7d),
	.w4(32'hbb3602fb),
	.w5(32'hbab85845),
	.w6(32'hbbf9dd83),
	.w7(32'h3b988618),
	.w8(32'h3bf08a30),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb376cca),
	.w1(32'h392ae423),
	.w2(32'h3b443ce9),
	.w3(32'h3a2b6c41),
	.w4(32'h3b585188),
	.w5(32'h3b4fe428),
	.w6(32'hba3f5af0),
	.w7(32'hbb314258),
	.w8(32'h392105e7),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d85a),
	.w1(32'hbae79f3f),
	.w2(32'hba2820fc),
	.w3(32'h3ace413d),
	.w4(32'hbc01d05d),
	.w5(32'hbc19473c),
	.w6(32'h3a7dfc8b),
	.w7(32'hbb8e744e),
	.w8(32'hba0a8d55),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92daa2),
	.w1(32'hbaeff8b6),
	.w2(32'hba32e70b),
	.w3(32'hbbf038bf),
	.w4(32'h3a5db4f0),
	.w5(32'h3ae691da),
	.w6(32'hbb68baf8),
	.w7(32'h3b185b97),
	.w8(32'h3b57697c),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c0e53),
	.w1(32'hbb235795),
	.w2(32'hbb61900b),
	.w3(32'h3810ca3e),
	.w4(32'hbb258d61),
	.w5(32'hbba7b55b),
	.w6(32'h3b06944e),
	.w7(32'hbac4a7cc),
	.w8(32'h3b1c44f7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03a160),
	.w1(32'hbbc5f1dc),
	.w2(32'hbb1e8f1f),
	.w3(32'hbba84b23),
	.w4(32'hbc0ca847),
	.w5(32'hbbb337f2),
	.w6(32'h3af8668b),
	.w7(32'hbb87c963),
	.w8(32'hbbbd03c1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e2fcf),
	.w1(32'h390733d6),
	.w2(32'h3b454f04),
	.w3(32'hbb298cea),
	.w4(32'hbb8bfd4e),
	.w5(32'hbb4f7a20),
	.w6(32'hbbdb4db2),
	.w7(32'hbb73ae57),
	.w8(32'hbb695ec9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5edcb),
	.w1(32'hbaa26869),
	.w2(32'h3be1ce78),
	.w3(32'hbb20bb02),
	.w4(32'hbc1836a4),
	.w5(32'hbbfc29c0),
	.w6(32'hbb8235cb),
	.w7(32'hbbed9cb6),
	.w8(32'hbbf1f8a1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c95d5),
	.w1(32'h3b3781c5),
	.w2(32'hbb0b98dc),
	.w3(32'h3a574de7),
	.w4(32'hbaeb95c2),
	.w5(32'h3b089ac6),
	.w6(32'hbb677eaf),
	.w7(32'hbbbaf1af),
	.w8(32'hbb0479ab),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09cdd2),
	.w1(32'h3c23425a),
	.w2(32'h3b868e51),
	.w3(32'hbb12b8b3),
	.w4(32'hbb3a94ba),
	.w5(32'hba48021c),
	.w6(32'hbb37ba59),
	.w7(32'h3bb0a7e2),
	.w8(32'h3b364002),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4931cc),
	.w1(32'hb9837123),
	.w2(32'hbb48440c),
	.w3(32'hbb63892e),
	.w4(32'h3b89b793),
	.w5(32'h3bae8b77),
	.w6(32'hbb425d80),
	.w7(32'h3be240ef),
	.w8(32'h3a0d5b6e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9624d),
	.w1(32'hbc41fd9e),
	.w2(32'hbbf135a1),
	.w3(32'h3c113ccb),
	.w4(32'hbb6d4aab),
	.w5(32'hbb808970),
	.w6(32'hba94b537),
	.w7(32'hbabc9d76),
	.w8(32'hbaca7790),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc024380),
	.w1(32'hbb6aeef7),
	.w2(32'hbab07d55),
	.w3(32'hbb0fd3fd),
	.w4(32'h39ec0c79),
	.w5(32'hbb3d0fca),
	.w6(32'h3a129cf1),
	.w7(32'hba06fc63),
	.w8(32'hbb29c4b1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86c744),
	.w1(32'h39d5d9eb),
	.w2(32'hba43d002),
	.w3(32'hb9e068a3),
	.w4(32'h3bb72460),
	.w5(32'h3b906e83),
	.w6(32'h3b161f9c),
	.w7(32'hb9be9d4f),
	.w8(32'h3ae8e4d1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9aabe),
	.w1(32'h3b8653c1),
	.w2(32'h3bd7f507),
	.w3(32'hba00b095),
	.w4(32'hbb658af8),
	.w5(32'hbbfe166d),
	.w6(32'h3ad80ce1),
	.w7(32'h3b03b213),
	.w8(32'h3ad47a31),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b7331),
	.w1(32'h3c1cc72b),
	.w2(32'h3b7cd5ed),
	.w3(32'h3ba9c275),
	.w4(32'hbb31701b),
	.w5(32'hbc2098ac),
	.w6(32'h3b70cd90),
	.w7(32'h3b87b2c7),
	.w8(32'h3a821ea1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa37ba),
	.w1(32'hbc27f6f2),
	.w2(32'hbc3857f0),
	.w3(32'hbbc74a94),
	.w4(32'h3bb2bc63),
	.w5(32'h3c9829f0),
	.w6(32'h3b1551cd),
	.w7(32'h3b03190a),
	.w8(32'h39fa4b7f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a6d8c),
	.w1(32'hbb909b56),
	.w2(32'hbba07580),
	.w3(32'h3b2224fa),
	.w4(32'hbb600c33),
	.w5(32'hb86ec534),
	.w6(32'h3a8bd232),
	.w7(32'h3a91a966),
	.w8(32'h3b5ed61d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2504ec),
	.w1(32'h3b3b1c46),
	.w2(32'hb9ccc56a),
	.w3(32'h3bc887a3),
	.w4(32'h3ac84dcc),
	.w5(32'h3a8d2b60),
	.w6(32'hbabaf2eb),
	.w7(32'h3b71a7af),
	.w8(32'h3bd28beb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88fca5),
	.w1(32'hbc32e7db),
	.w2(32'hbbd4c547),
	.w3(32'h3b1efc6e),
	.w4(32'hbbac9461),
	.w5(32'hbb89e2fd),
	.w6(32'h3b3be33e),
	.w7(32'h373f7e5c),
	.w8(32'h3b7b31df),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea674f),
	.w1(32'hbc135553),
	.w2(32'hbbd59783),
	.w3(32'hbb965e3d),
	.w4(32'hbb0e42f7),
	.w5(32'h399a4dc7),
	.w6(32'hba5bc1d4),
	.w7(32'hbb036b34),
	.w8(32'hbb083bd7),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4b5ae),
	.w1(32'h3b95f1a0),
	.w2(32'hb9d05766),
	.w3(32'h3b201b51),
	.w4(32'hb80a56fb),
	.w5(32'hbb98e76b),
	.w6(32'hbbd6d296),
	.w7(32'h3bbb6b3b),
	.w8(32'h3b4a2b96),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba53309),
	.w1(32'h3c00579c),
	.w2(32'h3c305e66),
	.w3(32'h3ab6e009),
	.w4(32'hbc70e890),
	.w5(32'hbc44554c),
	.w6(32'hbafe479e),
	.w7(32'hbbc5ee6f),
	.w8(32'hbb991ef3),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b924bb1),
	.w1(32'h3b79fcc1),
	.w2(32'hb9c5dfc6),
	.w3(32'hbc22c2af),
	.w4(32'hbb41bf47),
	.w5(32'hbadd2d77),
	.w6(32'hbbcbc50e),
	.w7(32'hbb998bf4),
	.w8(32'hbb8b4fb7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba516826),
	.w1(32'hbb9388f1),
	.w2(32'h38935a1a),
	.w3(32'h3a3245a4),
	.w4(32'hbbad889a),
	.w5(32'hbbdcf70b),
	.w6(32'hbaef30d8),
	.w7(32'hbbad28dc),
	.w8(32'hbb85d7da),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba876423),
	.w1(32'hbaa23fff),
	.w2(32'h399c1ae6),
	.w3(32'hbbdde97c),
	.w4(32'hbb09b407),
	.w5(32'hbbc0f7f1),
	.w6(32'hbbcb8a03),
	.w7(32'hbb3445ec),
	.w8(32'hbb055a33),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule