module layer_8_featuremap_145(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849584),
	.w1(32'hbb7dde62),
	.w2(32'hbc694879),
	.w3(32'hbb8a5049),
	.w4(32'hbaeab8d2),
	.w5(32'h3a4e0742),
	.w6(32'hba3ac94a),
	.w7(32'hbc3a9bf3),
	.w8(32'h3d170618),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb522943),
	.w1(32'hbc053fc5),
	.w2(32'hbaf292af),
	.w3(32'hbc5997c5),
	.w4(32'h3b7fc7fa),
	.w5(32'h3c51b1f3),
	.w6(32'h3a7c1dc4),
	.w7(32'hbb0c53db),
	.w8(32'h3cdb9445),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c757bc4),
	.w1(32'h3c03a926),
	.w2(32'hbb8c2e43),
	.w3(32'h3aa80412),
	.w4(32'hb9b1b83e),
	.w5(32'hbcaa9de1),
	.w6(32'h3bda3f15),
	.w7(32'h3cbf9fac),
	.w8(32'hbc80b0f9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbeb3c2),
	.w1(32'hbb7672a1),
	.w2(32'hbc02b890),
	.w3(32'h3b89ef7e),
	.w4(32'hbb85d2c9),
	.w5(32'h3bd2e281),
	.w6(32'h3be6fdd5),
	.w7(32'hba12182a),
	.w8(32'h3c7b231e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a99ef),
	.w1(32'hba5c75e7),
	.w2(32'h3b8cb5ee),
	.w3(32'h3ae469a2),
	.w4(32'h3ad8e98e),
	.w5(32'hbb0603c2),
	.w6(32'hba8d7ff2),
	.w7(32'h3b05075b),
	.w8(32'h3c9a8822),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f944b),
	.w1(32'h3c20b767),
	.w2(32'hbbb56a15),
	.w3(32'h3b87bf5b),
	.w4(32'hb91dd429),
	.w5(32'h3c776630),
	.w6(32'h3c2a65b0),
	.w7(32'h3b006f1f),
	.w8(32'h3bc2b33d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48410a),
	.w1(32'h3c0e0cef),
	.w2(32'hbc4fd77b),
	.w3(32'hbc46f24b),
	.w4(32'hbc40f174),
	.w5(32'h3c787250),
	.w6(32'hbb839dd5),
	.w7(32'hbb435357),
	.w8(32'h3c715e00),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23712a),
	.w1(32'hbc799278),
	.w2(32'h3c6f57fa),
	.w3(32'hba6c0c5c),
	.w4(32'h3c317892),
	.w5(32'hbbb602e7),
	.w6(32'hbc81cb61),
	.w7(32'h3c6ba03a),
	.w8(32'hbc56f415),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbce9d4),
	.w1(32'h3cb22521),
	.w2(32'h3a70d8ea),
	.w3(32'h3a82d7d2),
	.w4(32'hba2a2e3b),
	.w5(32'hba2a34a0),
	.w6(32'h3b2b439b),
	.w7(32'hbbd4b703),
	.w8(32'h3c7e8431),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e026),
	.w1(32'hbc0df9fe),
	.w2(32'hbc671303),
	.w3(32'hbc06d901),
	.w4(32'h3b27aadc),
	.w5(32'h3c35ca86),
	.w6(32'hbba7e13f),
	.w7(32'hbc1cf546),
	.w8(32'h3ad6c169),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e2b12),
	.w1(32'hbc429b40),
	.w2(32'h3c82122a),
	.w3(32'h3abd7f63),
	.w4(32'h3b06e811),
	.w5(32'hbc243e69),
	.w6(32'hbc87ac36),
	.w7(32'hbbca5935),
	.w8(32'hbd17ca79),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1ae76),
	.w1(32'hbc68d633),
	.w2(32'h3cb40f70),
	.w3(32'hbc683fc7),
	.w4(32'h3c767311),
	.w5(32'h3c4e7e5f),
	.w6(32'hbcb50c95),
	.w7(32'h3cb04979),
	.w8(32'h3c5157e0),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf7319),
	.w1(32'h3c792201),
	.w2(32'h3b532374),
	.w3(32'h3badad1c),
	.w4(32'h3b6fb626),
	.w5(32'h3ad2acdf),
	.w6(32'h3c04d081),
	.w7(32'hbaa66676),
	.w8(32'hba6c5bc5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3743),
	.w1(32'h3b8f33e4),
	.w2(32'hbb80e711),
	.w3(32'h3b114cd3),
	.w4(32'h3b866bd0),
	.w5(32'h38aba2ba),
	.w6(32'h3c1e7896),
	.w7(32'hbb8e798d),
	.w8(32'hbada0330),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b050),
	.w1(32'hb97812b8),
	.w2(32'h3816600b),
	.w3(32'hbae7da2e),
	.w4(32'h3a96b55e),
	.w5(32'hbae0c9f1),
	.w6(32'hbb10be4d),
	.w7(32'hbb57fdf3),
	.w8(32'hbb207880),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27ef13),
	.w1(32'h3a59ca6c),
	.w2(32'hbc3ee9cd),
	.w3(32'hbb3a92cc),
	.w4(32'hbbc13d9d),
	.w5(32'hbb16f35b),
	.w6(32'hbb1e7f40),
	.w7(32'hbbc17c04),
	.w8(32'hbc95664d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ae105),
	.w1(32'h3c51f3e8),
	.w2(32'h3c27fa02),
	.w3(32'h3b8c8545),
	.w4(32'h3c21e16d),
	.w5(32'hbbfe07f4),
	.w6(32'hbca60b41),
	.w7(32'h3b7aa135),
	.w8(32'h3b183e9b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8416bd),
	.w1(32'h3c3ba689),
	.w2(32'hbc239b4d),
	.w3(32'h3b735494),
	.w4(32'hbc3ad015),
	.w5(32'h39a559fe),
	.w6(32'hbb7d54d6),
	.w7(32'hbb5f6233),
	.w8(32'hbc1f8f88),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c496133),
	.w1(32'hb9a67510),
	.w2(32'h3c5941ab),
	.w3(32'hb943bd28),
	.w4(32'hbbd233dc),
	.w5(32'h3bcb3882),
	.w6(32'hbbbe1fa3),
	.w7(32'hbca1fb9e),
	.w8(32'hbc10b7bf),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f473f),
	.w1(32'h3a61c1ba),
	.w2(32'hbbb03e85),
	.w3(32'h3bb65b32),
	.w4(32'hbb8b0b17),
	.w5(32'hbd0cec9b),
	.w6(32'hbb9d5c6d),
	.w7(32'hbbe2064d),
	.w8(32'hbc47817b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c728b),
	.w1(32'hbc4ef9ae),
	.w2(32'h36facc2a),
	.w3(32'hbc48c7e0),
	.w4(32'hbb5f61b2),
	.w5(32'h3c1c491a),
	.w6(32'h3bdc48bf),
	.w7(32'hbc1a549c),
	.w8(32'hbd463de6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c061140),
	.w1(32'h3b86b4ab),
	.w2(32'hbc2908d5),
	.w3(32'hbbd932ca),
	.w4(32'hbc9e9907),
	.w5(32'hbb5ca764),
	.w6(32'hba5f22d9),
	.w7(32'h3cb71395),
	.w8(32'h3b03eb12),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce99b2c),
	.w1(32'h3c8dcd38),
	.w2(32'h3c31b454),
	.w3(32'h3bc35023),
	.w4(32'h3b8236b6),
	.w5(32'h3c2a9bcd),
	.w6(32'hbcb18985),
	.w7(32'hbb6c481c),
	.w8(32'hbcc4000e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca996a),
	.w1(32'h3aac0bdd),
	.w2(32'hbae83563),
	.w3(32'h3b1611eb),
	.w4(32'hbb95b7cb),
	.w5(32'hbadba379),
	.w6(32'h3b6d26f5),
	.w7(32'h3a0ed614),
	.w8(32'hb9420be2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d2fa1),
	.w1(32'hba1f788f),
	.w2(32'hbb4f292c),
	.w3(32'hba75aa74),
	.w4(32'hbba613f3),
	.w5(32'hbb76fa64),
	.w6(32'hbc032607),
	.w7(32'h3b0adf9d),
	.w8(32'hbbbf8194),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a497f9),
	.w1(32'hbaea1c8a),
	.w2(32'h3b838ac3),
	.w3(32'hb95048d0),
	.w4(32'hbbc02e82),
	.w5(32'h3c365d09),
	.w6(32'h399785bc),
	.w7(32'h3c4a888a),
	.w8(32'h3c9bed62),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f8d1a),
	.w1(32'h3c92d936),
	.w2(32'h3a88b97f),
	.w3(32'h3c1ad18b),
	.w4(32'hbc085d47),
	.w5(32'hbac90d7b),
	.w6(32'hbcd89e87),
	.w7(32'hbaea51a1),
	.w8(32'h3b9f47b6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfcc6c7),
	.w1(32'hbc124df1),
	.w2(32'hbcb7c002),
	.w3(32'h3cad3c4f),
	.w4(32'hbb5f466a),
	.w5(32'hbc98111d),
	.w6(32'h3c76a90e),
	.w7(32'hbd091e72),
	.w8(32'h3c65b269),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707d2f),
	.w1(32'h3c4c90b0),
	.w2(32'hbc62ca6b),
	.w3(32'hbc19ec56),
	.w4(32'hbc701a1b),
	.w5(32'hbd0e2664),
	.w6(32'hba26820a),
	.w7(32'hbc6aab5f),
	.w8(32'h3ccb7049),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbae754),
	.w1(32'h3a5b2b3f),
	.w2(32'hbc805618),
	.w3(32'h3c0b80c4),
	.w4(32'h3b93c1c2),
	.w5(32'h3d038186),
	.w6(32'hbbe225fc),
	.w7(32'h3cb364c9),
	.w8(32'hbd768b12),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48306c),
	.w1(32'h3beebb24),
	.w2(32'hba5ee89e),
	.w3(32'hbb3a22a6),
	.w4(32'hba840ab3),
	.w5(32'hbb740447),
	.w6(32'hbcac980c),
	.w7(32'hbb667b8c),
	.w8(32'hbba5abc9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb454ec1),
	.w1(32'hbb365dfa),
	.w2(32'hbccc18ab),
	.w3(32'hbb8009c3),
	.w4(32'hbb4a76b1),
	.w5(32'hbcaad42c),
	.w6(32'hbb48685b),
	.w7(32'hbc90995a),
	.w8(32'hbd0d8030),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc1b9b3),
	.w1(32'h3c3d81ab),
	.w2(32'h3cc18357),
	.w3(32'hbb1d38fa),
	.w4(32'h3addb378),
	.w5(32'h3c9ff74d),
	.w6(32'h3ba7b3be),
	.w7(32'hbb9400e4),
	.w8(32'hbc31312f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e07d5),
	.w1(32'hbc89aa3a),
	.w2(32'h399279d1),
	.w3(32'hbbd303d5),
	.w4(32'h3bfc7864),
	.w5(32'h3c4c1ad2),
	.w6(32'h3ae7b932),
	.w7(32'hbc186e9e),
	.w8(32'hbc098d5e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f42a3),
	.w1(32'h3b5d8c11),
	.w2(32'hbb9351bd),
	.w3(32'hbbfe6409),
	.w4(32'h3ad99267),
	.w5(32'hbb8b129f),
	.w6(32'h3c58ddee),
	.w7(32'h3a6f4d72),
	.w8(32'hbbc3dccf),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51e2fa),
	.w1(32'h3b0579e5),
	.w2(32'h3c1c631a),
	.w3(32'hb92431b0),
	.w4(32'hbc022a0b),
	.w5(32'hbbd9548e),
	.w6(32'h3c1e948e),
	.w7(32'h3c5108e0),
	.w8(32'h3c31dcfe),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5986),
	.w1(32'hbad06383),
	.w2(32'hbca44932),
	.w3(32'hbc2833d1),
	.w4(32'hbc801e91),
	.w5(32'hbc2ca757),
	.w6(32'h3c962a43),
	.w7(32'hbc234ae3),
	.w8(32'h3c29f494),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0dbc0),
	.w1(32'hbc05456d),
	.w2(32'hbacf7385),
	.w3(32'h3b20c73e),
	.w4(32'h3c6694a6),
	.w5(32'h3bb643a4),
	.w6(32'hbb93ed8c),
	.w7(32'hbb97fd2a),
	.w8(32'hbbdc9620),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d8efb),
	.w1(32'hbc102c97),
	.w2(32'hbcdd4d1b),
	.w3(32'h3c0e959c),
	.w4(32'hbc07f80e),
	.w5(32'hbcf79aa8),
	.w6(32'hbb697ab7),
	.w7(32'hbc782025),
	.w8(32'hbc7790a4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38751f),
	.w1(32'hbb6213f6),
	.w2(32'h3bc78429),
	.w3(32'hbc45593f),
	.w4(32'h3bf81934),
	.w5(32'h3aa4ed4c),
	.w6(32'hba97b6e0),
	.w7(32'h3c2dc206),
	.w8(32'h3bc80a08),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b93f3),
	.w1(32'h3c10552a),
	.w2(32'hba2298da),
	.w3(32'h3a1d09ac),
	.w4(32'hba7c4fa5),
	.w5(32'h3b5fba35),
	.w6(32'h3bfb1514),
	.w7(32'hbc0586bb),
	.w8(32'hbc81aa1e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf91691),
	.w1(32'h3b22aec6),
	.w2(32'hbc1e066c),
	.w3(32'h3b2c0a7e),
	.w4(32'hbccccbfa),
	.w5(32'h3bfc9211),
	.w6(32'hbc8ecf26),
	.w7(32'h3d12fc51),
	.w8(32'h3c1bd136),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba1aba),
	.w1(32'h3c2c8848),
	.w2(32'h3bcbe801),
	.w3(32'h3ab84614),
	.w4(32'h3b26f25d),
	.w5(32'hbc0c2a64),
	.w6(32'hbcf2c488),
	.w7(32'hbcee0f01),
	.w8(32'hbd2aa285),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfbc471),
	.w1(32'hbc783668),
	.w2(32'h3b7a6001),
	.w3(32'h3a004432),
	.w4(32'h3b09165d),
	.w5(32'h3b056e1f),
	.w6(32'h3d1623aa),
	.w7(32'hbba33498),
	.w8(32'hbb008cf8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696f21),
	.w1(32'h3b7711eb),
	.w2(32'h3b52c618),
	.w3(32'h3aafa59a),
	.w4(32'hbaf8332c),
	.w5(32'hbc8cceef),
	.w6(32'h3ac991af),
	.w7(32'hbc018a99),
	.w8(32'h3b89607f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc931345),
	.w1(32'h3baee809),
	.w2(32'h3b207575),
	.w3(32'h3b027da4),
	.w4(32'hbcb13e6f),
	.w5(32'hbb6f3778),
	.w6(32'hbc42e5ef),
	.w7(32'h3cb40fac),
	.w8(32'h3ca7373f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4ec4e),
	.w1(32'h3c0ce870),
	.w2(32'h3b8703b4),
	.w3(32'hbba2282d),
	.w4(32'hbb90d820),
	.w5(32'hbc608d4d),
	.w6(32'hbbab8d62),
	.w7(32'h3bb8d4be),
	.w8(32'h3cc1d565),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd02b02),
	.w1(32'hbc030857),
	.w2(32'h3b34433f),
	.w3(32'hbcf79ccd),
	.w4(32'hbc155174),
	.w5(32'hbc13105f),
	.w6(32'h3bcdb715),
	.w7(32'hba2c8c72),
	.w8(32'h3c44f039),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d426b),
	.w1(32'h3c3573d8),
	.w2(32'hba6b0dc2),
	.w3(32'h3cbb5ad8),
	.w4(32'hbbf03726),
	.w5(32'h3c0e3332),
	.w6(32'hbc64f204),
	.w7(32'hbc3cce63),
	.w8(32'h398163f1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9e782d),
	.w1(32'hbcdbe187),
	.w2(32'hbbeaaf0c),
	.w3(32'hbc07c9e8),
	.w4(32'hbc5384ed),
	.w5(32'hbbf62037),
	.w6(32'hbbe778bb),
	.w7(32'hbc1b00dd),
	.w8(32'hbbafdef8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e5764),
	.w1(32'hbc038a6b),
	.w2(32'hbaea3a2e),
	.w3(32'hbc2707a1),
	.w4(32'hbcac1e1a),
	.w5(32'h3aaf684c),
	.w6(32'hbc4d2817),
	.w7(32'h3bc9b967),
	.w8(32'h3c6015d9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07d5a6),
	.w1(32'h3ba74633),
	.w2(32'h3c48a7ae),
	.w3(32'h3c8557cb),
	.w4(32'h3caa5b09),
	.w5(32'h3cdf1326),
	.w6(32'hbd03c6a0),
	.w7(32'hbcaac53d),
	.w8(32'hbc28f09b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe64c02),
	.w1(32'hbb8083f9),
	.w2(32'hbb4647f1),
	.w3(32'h3c59fcdf),
	.w4(32'hbb310904),
	.w5(32'h3b5b9b50),
	.w6(32'hbbfc16c2),
	.w7(32'hbbc638a8),
	.w8(32'hbc0b3e3f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fe203),
	.w1(32'h3b8130a3),
	.w2(32'h3b108c13),
	.w3(32'hbc242d79),
	.w4(32'h3b033f62),
	.w5(32'h39f363bc),
	.w6(32'hbb2343d9),
	.w7(32'hbb010ba1),
	.w8(32'h3a0b57df),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3c19a),
	.w1(32'h3ad5ecb5),
	.w2(32'hbbb92fea),
	.w3(32'hb9651953),
	.w4(32'h3bd07ba8),
	.w5(32'hbb52766b),
	.w6(32'h3b5354f2),
	.w7(32'hbd02574c),
	.w8(32'h3d630a2e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d3878),
	.w1(32'hbc9a76a9),
	.w2(32'h3a9bcfc1),
	.w3(32'hbbcf5e41),
	.w4(32'hbc626daf),
	.w5(32'hbb4fce5e),
	.w6(32'h3c9787f5),
	.w7(32'hbc5496ff),
	.w8(32'h3b346eac),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f2c9d),
	.w1(32'hbbf55336),
	.w2(32'hbb197726),
	.w3(32'h3ba94757),
	.w4(32'hba452309),
	.w5(32'hbb9056d0),
	.w6(32'hbb81b883),
	.w7(32'hbc395f2c),
	.w8(32'hbbc722ae),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a0c16),
	.w1(32'hbafbb33b),
	.w2(32'hbc859d02),
	.w3(32'h39b566fc),
	.w4(32'hbbc7d3fe),
	.w5(32'h3bd3c4b0),
	.w6(32'hbc0ebd40),
	.w7(32'h3ce5db35),
	.w8(32'hbcf4e3cb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce86427),
	.w1(32'h3c02ebe7),
	.w2(32'h3b5c6f56),
	.w3(32'hbb214323),
	.w4(32'h3b3b9e1f),
	.w5(32'h3b26dc66),
	.w6(32'hbb32516e),
	.w7(32'hbb84bed6),
	.w8(32'h3a0a6c98),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ed3d3),
	.w1(32'h3ab33a2f),
	.w2(32'hbb0baa2e),
	.w3(32'hba99ec34),
	.w4(32'h3b163b41),
	.w5(32'hbc950019),
	.w6(32'h3b5f4579),
	.w7(32'hbcb0e657),
	.w8(32'h3cbb46de),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2940e1),
	.w1(32'hbcdd9a7a),
	.w2(32'hbb24f483),
	.w3(32'h3a4c2001),
	.w4(32'hbc7acd08),
	.w5(32'h3bbbdc41),
	.w6(32'h3ce911ce),
	.w7(32'h3be16eaa),
	.w8(32'hbc40e2d7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8f6c6),
	.w1(32'h3c599cd5),
	.w2(32'h39de7ab9),
	.w3(32'h3b4ac721),
	.w4(32'hbbfb7633),
	.w5(32'hbbe203f5),
	.w6(32'hbbcc6e9f),
	.w7(32'h3a2412e3),
	.w8(32'hbb259a42),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9650a5),
	.w1(32'hbadd0784),
	.w2(32'h3c0f170b),
	.w3(32'hbb93b905),
	.w4(32'h3adbff5a),
	.w5(32'h3acd0625),
	.w6(32'hbb8e3cab),
	.w7(32'hbceb85f1),
	.w8(32'h3bd8009f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc248175),
	.w1(32'hbc8642b6),
	.w2(32'hb94bd49b),
	.w3(32'hbc4770ec),
	.w4(32'h3b69f217),
	.w5(32'hbc1de831),
	.w6(32'hbba77ce9),
	.w7(32'hbbb497ba),
	.w8(32'hbb86ffac),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecf868),
	.w1(32'hbc004cf9),
	.w2(32'hba5aeeeb),
	.w3(32'hbb2e6424),
	.w4(32'hbc18324e),
	.w5(32'hba26c20a),
	.w6(32'h3c40e74b),
	.w7(32'hbbddafbb),
	.w8(32'h3c0aff54),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3b237),
	.w1(32'hbc8292d3),
	.w2(32'h3b4c98ae),
	.w3(32'hbb948f3e),
	.w4(32'h3bc4f350),
	.w5(32'h3ba33ec4),
	.w6(32'hba4c94e4),
	.w7(32'hb90090d2),
	.w8(32'hbc6b46a5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c84c7c6),
	.w1(32'h3c018745),
	.w2(32'hbb8e22fa),
	.w3(32'hbb6e0408),
	.w4(32'h3c2aa802),
	.w5(32'hbbda373b),
	.w6(32'h3b4d02f2),
	.w7(32'h3aa2ec8a),
	.w8(32'hba742cc2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf21ff3),
	.w1(32'hbb82cbfe),
	.w2(32'h3c24a9e6),
	.w3(32'hbc1e2827),
	.w4(32'hbb343c73),
	.w5(32'h3b69c985),
	.w6(32'h3c59cff1),
	.w7(32'hbc8a4785),
	.w8(32'hbd1be4a5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0f0e7),
	.w1(32'hba840fa1),
	.w2(32'hbba7f6f2),
	.w3(32'hbbb98c51),
	.w4(32'hbc9ccca4),
	.w5(32'hbb9894d4),
	.w6(32'h3b2354cc),
	.w7(32'h3be5cc5a),
	.w8(32'h3c8af2fa),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c190a31),
	.w1(32'hbba68a09),
	.w2(32'h3c135803),
	.w3(32'h3bab24f5),
	.w4(32'h3adfe8f2),
	.w5(32'h3cb473fe),
	.w6(32'hbc2f4882),
	.w7(32'hbbc5f277),
	.w8(32'hbcc7b5db),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4fc30),
	.w1(32'hbb28b240),
	.w2(32'h3c14429c),
	.w3(32'hbb608540),
	.w4(32'hbb02deb7),
	.w5(32'h3a30afc4),
	.w6(32'hbb2b227f),
	.w7(32'hbc44b60d),
	.w8(32'hbcdfc357),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b69d),
	.w1(32'hbb2d5857),
	.w2(32'hbc2576b6),
	.w3(32'hb9e9bd0b),
	.w4(32'hbb915519),
	.w5(32'hbbdd3cc9),
	.w6(32'hbaeb2e7e),
	.w7(32'hbc53ab66),
	.w8(32'hbc2cf977),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc095e08),
	.w1(32'hbc6dd913),
	.w2(32'h3b5b02bd),
	.w3(32'hbc431954),
	.w4(32'hba1ec1c0),
	.w5(32'hbb11bad4),
	.w6(32'hbbb2b3eb),
	.w7(32'hba7fa476),
	.w8(32'hbc2a32cf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df7fc),
	.w1(32'hbb71ac2a),
	.w2(32'h3c9a93c7),
	.w3(32'hbb9a3fa8),
	.w4(32'h3c4d43c8),
	.w5(32'hbcc14759),
	.w6(32'hbb02a984),
	.w7(32'hbd4aa47c),
	.w8(32'h3c51f898),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c348367),
	.w1(32'hbd1f8c9b),
	.w2(32'hbc215d9b),
	.w3(32'h3b7aea5e),
	.w4(32'hbccaccad),
	.w5(32'hbbfbed4a),
	.w6(32'h3d4c0c5c),
	.w7(32'h3bfac47e),
	.w8(32'h3c0c6616),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa76d6),
	.w1(32'hbb15c725),
	.w2(32'h3a93c2dd),
	.w3(32'hbc53e30b),
	.w4(32'hba5a7573),
	.w5(32'hbaa64dba),
	.w6(32'hbc85b380),
	.w7(32'hbc26aaaf),
	.w8(32'hbb342dbe),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4db64),
	.w1(32'hbac9a48a),
	.w2(32'hbba2ddb7),
	.w3(32'hbaa531c6),
	.w4(32'hbafa4691),
	.w5(32'hbbc1a94e),
	.w6(32'h3b9d1dc0),
	.w7(32'hbbd7d0c9),
	.w8(32'hbc5da9fe),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c496bbc),
	.w1(32'h3c9fae34),
	.w2(32'h3bbcef65),
	.w3(32'hbc1f5452),
	.w4(32'hbbc20335),
	.w5(32'h3ab37025),
	.w6(32'hbab9c7f9),
	.w7(32'hbc31d4c0),
	.w8(32'hbbce96b9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a3022),
	.w1(32'h3aa850cd),
	.w2(32'hbb243c93),
	.w3(32'hbb49230b),
	.w4(32'hbbd6a00c),
	.w5(32'hbb908219),
	.w6(32'h3c0b9280),
	.w7(32'hbbdaf915),
	.w8(32'hbbe59370),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac32d8),
	.w1(32'hbc0c330b),
	.w2(32'h39584a0c),
	.w3(32'hbacaae84),
	.w4(32'hbc507f52),
	.w5(32'h3b657327),
	.w6(32'hbac7cb6a),
	.w7(32'h3c440852),
	.w8(32'hbc15ec7f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cffc96d),
	.w1(32'h3cc9d942),
	.w2(32'h3b185bf0),
	.w3(32'h3be73182),
	.w4(32'h3b818682),
	.w5(32'h3bb05fa4),
	.w6(32'hbcc3081e),
	.w7(32'h3c074ff1),
	.w8(32'h3c871c84),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6740ff),
	.w1(32'hbc0500aa),
	.w2(32'hbc803baf),
	.w3(32'h3bcfae1d),
	.w4(32'h3b80c1a6),
	.w5(32'h3c34b499),
	.w6(32'h3a97fd52),
	.w7(32'h3b4df0ff),
	.w8(32'hbcd4587e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718173),
	.w1(32'h3c33f895),
	.w2(32'hbabeed5a),
	.w3(32'hbb957c1f),
	.w4(32'hbb558add),
	.w5(32'h3bed8915),
	.w6(32'hbb1e3cda),
	.w7(32'hba9dc2ba),
	.w8(32'hba9708e9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc305b2f),
	.w1(32'h3b5c892a),
	.w2(32'h3d19dfeb),
	.w3(32'hbbfbc046),
	.w4(32'h3c69c3c9),
	.w5(32'hbb6455dd),
	.w6(32'hbc22f926),
	.w7(32'hbc982598),
	.w8(32'hbcbfa141),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c0a17),
	.w1(32'hbcbedaf0),
	.w2(32'h3b96ecd3),
	.w3(32'hbbde4d3a),
	.w4(32'hbc892003),
	.w5(32'hbb859ac1),
	.w6(32'h3d1b7a05),
	.w7(32'hbc77d3bf),
	.w8(32'h3cb65c16),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52f8c8),
	.w1(32'h3be9e4ec),
	.w2(32'h3a6b35fc),
	.w3(32'h3c2b178b),
	.w4(32'hbaf11f56),
	.w5(32'h3c68a570),
	.w6(32'h3b99022d),
	.w7(32'hbae87ecb),
	.w8(32'h3bea084a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e62e8),
	.w1(32'h3c4aa386),
	.w2(32'h3a929d62),
	.w3(32'h3c251870),
	.w4(32'hbb3b2e7f),
	.w5(32'h3be62793),
	.w6(32'hbc1039b2),
	.w7(32'h3ad3bd99),
	.w8(32'h3c73b078),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb01c1),
	.w1(32'h3b8eb88f),
	.w2(32'hbc378b9a),
	.w3(32'h3bdbd767),
	.w4(32'hbc27681d),
	.w5(32'hbbce2e3e),
	.w6(32'hbbb4c31f),
	.w7(32'hbc17d649),
	.w8(32'hbb5cb0ff),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedbb0c),
	.w1(32'hbb493a09),
	.w2(32'hbc347061),
	.w3(32'h3a09b04c),
	.w4(32'h3b8fd0fe),
	.w5(32'h3bc59d19),
	.w6(32'h3ab912a0),
	.w7(32'h3b80a786),
	.w8(32'h3b17be92),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc993442),
	.w1(32'hbcb4eef2),
	.w2(32'h3c6451fd),
	.w3(32'h3b46f877),
	.w4(32'hba7eba86),
	.w5(32'h3c85cc20),
	.w6(32'hbc5763c3),
	.w7(32'h3c995dcc),
	.w8(32'h3da835c9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4931e6),
	.w1(32'hbd66ca2d),
	.w2(32'h3c639d06),
	.w3(32'h3ca85638),
	.w4(32'hbacd4350),
	.w5(32'hbc11325d),
	.w6(32'h3bfad532),
	.w7(32'hbcc1fb6a),
	.w8(32'hbcbd5505),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60081c),
	.w1(32'h3b4ec655),
	.w2(32'h3c6157f3),
	.w3(32'hbc818a68),
	.w4(32'h3a5e9db6),
	.w5(32'h3c11b2c6),
	.w6(32'h3c82f057),
	.w7(32'hbad6a7b9),
	.w8(32'h3b291cdc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f0a87),
	.w1(32'hbc61ad73),
	.w2(32'h3c9d2c34),
	.w3(32'h3b956ed7),
	.w4(32'h3c1b2b6a),
	.w5(32'h3b92893f),
	.w6(32'hbc4cbc83),
	.w7(32'h3cb9831e),
	.w8(32'h3a7573f0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba97ecc),
	.w1(32'h39c92e60),
	.w2(32'h3c1023a4),
	.w3(32'h3b9353ad),
	.w4(32'hbc08794a),
	.w5(32'hbc93d114),
	.w6(32'hbc441ef1),
	.w7(32'hbb4d9a48),
	.w8(32'hbc87597b),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c561f1e),
	.w1(32'h3b9b6e22),
	.w2(32'hbb5e942c),
	.w3(32'hbc2e5ca3),
	.w4(32'hbb20e9bc),
	.w5(32'hbb6c8fd5),
	.w6(32'h3a977348),
	.w7(32'hbb72a475),
	.w8(32'hbbaa2942),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4f6d0),
	.w1(32'hbc2e61b1),
	.w2(32'h3a96bb0c),
	.w3(32'hbb225fe5),
	.w4(32'hbc08c6f2),
	.w5(32'hbbe01520),
	.w6(32'hbbb698a4),
	.w7(32'hbc95d6df),
	.w8(32'hbd2f7d67),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d814bb4),
	.w1(32'h3d5d55a7),
	.w2(32'h3bfc8fd4),
	.w3(32'hb985d1a4),
	.w4(32'h3a9c1ad1),
	.w5(32'hbcd9f23d),
	.w6(32'hbc90422b),
	.w7(32'hbcfe9249),
	.w8(32'h3bc31735),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca609a9),
	.w1(32'hbbd6af2c),
	.w2(32'h37ff5aef),
	.w3(32'hbb3b5ba2),
	.w4(32'h3ba2deb2),
	.w5(32'h3c0f5932),
	.w6(32'h3c286234),
	.w7(32'h3c524d0b),
	.w8(32'h3b4c737d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9867f0),
	.w1(32'hbcbcbc2c),
	.w2(32'h3b89054b),
	.w3(32'h3b356977),
	.w4(32'h3bc78f8d),
	.w5(32'h3c06a0fa),
	.w6(32'h3c9fee9a),
	.w7(32'h3bf01123),
	.w8(32'h3c0dd6a2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23ee3b),
	.w1(32'hbc3128ea),
	.w2(32'h386ee8cb),
	.w3(32'h3bdb22f0),
	.w4(32'h3c071006),
	.w5(32'hbc2ed607),
	.w6(32'hbb735181),
	.w7(32'hbc8f8ccd),
	.w8(32'h3a7c4525),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befc972),
	.w1(32'h3c8496b3),
	.w2(32'hbbb72a13),
	.w3(32'hba7da1c4),
	.w4(32'hbba0d459),
	.w5(32'hba7d96dd),
	.w6(32'hbbf1ba1c),
	.w7(32'hbb25eb0b),
	.w8(32'hbc6526b3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bffb5),
	.w1(32'h3ca83a0f),
	.w2(32'hbb83ba3e),
	.w3(32'hbb87d541),
	.w4(32'hbbbc3657),
	.w5(32'h3c548766),
	.w6(32'hbc0d11e7),
	.w7(32'h3bf4d9dc),
	.w8(32'h3b84c95b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31704f),
	.w1(32'hbb039fcc),
	.w2(32'hbae997c9),
	.w3(32'h3cbed9e0),
	.w4(32'hbbc246b8),
	.w5(32'hbc0554c1),
	.w6(32'h3cc3266d),
	.w7(32'hbc2ed9a3),
	.w8(32'hbc8aada3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4efece),
	.w1(32'h3c11b6b3),
	.w2(32'h3b8ade9c),
	.w3(32'hbc132aa2),
	.w4(32'hbc6d17e7),
	.w5(32'hbc4ad474),
	.w6(32'hbc77b59b),
	.w7(32'hbafeeb4b),
	.w8(32'hba0291ba),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b267b),
	.w1(32'hb9c214f1),
	.w2(32'h3ca8e59e),
	.w3(32'hbc593f33),
	.w4(32'hbb3ac671),
	.w5(32'h392a966e),
	.w6(32'hbb661f7e),
	.w7(32'h3bb16f5d),
	.w8(32'hbd1b3b9f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6ff445),
	.w1(32'hbb8d1815),
	.w2(32'h3b303df3),
	.w3(32'hbb8d51cb),
	.w4(32'hb9d6d210),
	.w5(32'h3bf14bb7),
	.w6(32'h3d161326),
	.w7(32'hbcc5f09b),
	.w8(32'hbc6b2f6d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b2245),
	.w1(32'h3bbe412f),
	.w2(32'hbc671156),
	.w3(32'hbca7af29),
	.w4(32'h3bb63f37),
	.w5(32'h3b9ddb59),
	.w6(32'hbc4df400),
	.w7(32'h3b7ee337),
	.w8(32'hb9fa5d6b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced0a6e),
	.w1(32'h3b8703c3),
	.w2(32'hbbab2941),
	.w3(32'h3b1f6b86),
	.w4(32'hb72d8bfe),
	.w5(32'hbb962c0c),
	.w6(32'hbcfdf58c),
	.w7(32'hbba2fe5f),
	.w8(32'hbc689bc7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e8ccc),
	.w1(32'h3c8d39d4),
	.w2(32'h3bd0530f),
	.w3(32'hbc571030),
	.w4(32'hbbebab17),
	.w5(32'hbb809b8d),
	.w6(32'hbae68656),
	.w7(32'h3c70ac11),
	.w8(32'h3c6df268),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ba226),
	.w1(32'hbc0c3b1a),
	.w2(32'hbc128cd4),
	.w3(32'hbbb954ee),
	.w4(32'h3c0f0629),
	.w5(32'h3c01156d),
	.w6(32'hbbffa3e5),
	.w7(32'h3aabd0da),
	.w8(32'hbbff2142),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7b595),
	.w1(32'h3d0a0708),
	.w2(32'h3c507295),
	.w3(32'hbb965e73),
	.w4(32'h3ba48287),
	.w5(32'hbb18794f),
	.w6(32'hbcc71cbd),
	.w7(32'h3ccb4534),
	.w8(32'h3c8b9873),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca77ce4),
	.w1(32'hbbcc73e7),
	.w2(32'hba381ba6),
	.w3(32'h39a94dc0),
	.w4(32'h3c0af498),
	.w5(32'h3c156be1),
	.w6(32'hbc3dfe0a),
	.w7(32'h3bd9d753),
	.w8(32'h3c06e6bd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc669fd2),
	.w1(32'hbc5294d4),
	.w2(32'hbcb25a47),
	.w3(32'h3c96ba3b),
	.w4(32'h3ae59948),
	.w5(32'hbc42cc3a),
	.w6(32'h3c31edf8),
	.w7(32'hbc611f2d),
	.w8(32'hbd27a7c7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5205bd),
	.w1(32'h3cc1a719),
	.w2(32'hbcbeb997),
	.w3(32'hbcbd7fdf),
	.w4(32'hbd021ef1),
	.w5(32'hbcc9e265),
	.w6(32'h3a2abc28),
	.w7(32'hbd25a786),
	.w8(32'hbd18b356),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d122c95),
	.w1(32'h3d25c8ad),
	.w2(32'h3b785881),
	.w3(32'hbcb99785),
	.w4(32'hbbed3ac5),
	.w5(32'h3b2a35b9),
	.w6(32'h3c342910),
	.w7(32'h3c84be8b),
	.w8(32'h3d119b62),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9f8c1),
	.w1(32'h3b615ca7),
	.w2(32'h3b0f2bad),
	.w3(32'h3c41d7e1),
	.w4(32'h3aaa9ffa),
	.w5(32'h3c057ded),
	.w6(32'h3bdafa74),
	.w7(32'h3ca90991),
	.w8(32'h3d017c25),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbced6dc3),
	.w1(32'hbca55e29),
	.w2(32'hbbb97a78),
	.w3(32'h3a35dff8),
	.w4(32'hbbac0858),
	.w5(32'h3aaab78f),
	.w6(32'hbb3d2c69),
	.w7(32'hbbaa0f42),
	.w8(32'hbca4915b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc5a7a),
	.w1(32'h3c11c7c6),
	.w2(32'hb9d228df),
	.w3(32'hbc199ed6),
	.w4(32'hbb001166),
	.w5(32'hbb392972),
	.w6(32'h3cd8ec06),
	.w7(32'hbbf566f9),
	.w8(32'hbc397d68),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c184a24),
	.w1(32'h3c82e5a6),
	.w2(32'h38fab95a),
	.w3(32'hbc120f34),
	.w4(32'hbc1a8c63),
	.w5(32'hbba0e220),
	.w6(32'h3b0cf392),
	.w7(32'h3b83d9cf),
	.w8(32'h3cbf0555),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad7d07),
	.w1(32'hbbfcdb9f),
	.w2(32'hbb0ad1d6),
	.w3(32'hbb817905),
	.w4(32'hbb805053),
	.w5(32'hbc26d5b8),
	.w6(32'h3bb375f8),
	.w7(32'hbc614202),
	.w8(32'hbcd9d25f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2388ea),
	.w1(32'h3bc083fc),
	.w2(32'h3b9218e8),
	.w3(32'hbc2e6f5b),
	.w4(32'hbb7949cb),
	.w5(32'hbc3d306d),
	.w6(32'h3a52a30c),
	.w7(32'hbbe80758),
	.w8(32'hbb98cc68),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77f104),
	.w1(32'h3afa5594),
	.w2(32'h3c518ae0),
	.w3(32'hbb94cc6d),
	.w4(32'hbaf34f26),
	.w5(32'h3c90dc93),
	.w6(32'h3c542b5e),
	.w7(32'h3cb6c116),
	.w8(32'h3d4a0011),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1003fd),
	.w1(32'hbd29fdb7),
	.w2(32'hbb4fae5e),
	.w3(32'h3c58ac22),
	.w4(32'hba96730d),
	.w5(32'hbb966db4),
	.w6(32'hbc308c3c),
	.w7(32'hbbbfe1f4),
	.w8(32'hbc4cf53d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e2755),
	.w1(32'h3c7897d1),
	.w2(32'h3c2040da),
	.w3(32'hbc333ddc),
	.w4(32'h3a9b89f6),
	.w5(32'h3b31122e),
	.w6(32'hb97024ff),
	.w7(32'h3bb47be2),
	.w8(32'h3d2617a7),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1e32ac),
	.w1(32'h3b8b86c5),
	.w2(32'h3cf3449b),
	.w3(32'h3c0658f2),
	.w4(32'h3b0a04d6),
	.w5(32'hb9e1c8c7),
	.w6(32'hbcb83144),
	.w7(32'hbb3cc5d4),
	.w8(32'hbccc85a8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c7f64),
	.w1(32'hbcfd09c4),
	.w2(32'hb91d41d0),
	.w3(32'h3ba1065b),
	.w4(32'hba0a0fb1),
	.w5(32'h3a9535c0),
	.w6(32'h3c1ad43f),
	.w7(32'h3a3a64a1),
	.w8(32'h3b8961d0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e108),
	.w1(32'hbc2e13cb),
	.w2(32'h3bcbdbe5),
	.w3(32'h3af48816),
	.w4(32'hbc4a76cf),
	.w5(32'h39d126a2),
	.w6(32'hbb60b890),
	.w7(32'h3a02be01),
	.w8(32'h3a8b13ba),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e8806),
	.w1(32'hbbfe9f92),
	.w2(32'hbbb4ead6),
	.w3(32'h3af5b382),
	.w4(32'hb95d927c),
	.w5(32'hbc0e3472),
	.w6(32'h3c128e97),
	.w7(32'hbc843771),
	.w8(32'hbcd0acf5),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule