module layer_8_featuremap_125(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be72d),
	.w1(32'h3a94b122),
	.w2(32'hbb51fcf5),
	.w3(32'h387abaab),
	.w4(32'hbbc7f9f5),
	.w5(32'hbc0626ed),
	.w6(32'hbae7685e),
	.w7(32'hbbb9d59e),
	.w8(32'hbc19da6f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd36485),
	.w1(32'hbc045286),
	.w2(32'hb98dcd20),
	.w3(32'hbba516d8),
	.w4(32'hbb87064e),
	.w5(32'hbc2e5882),
	.w6(32'hbc0282d1),
	.w7(32'hbada85af),
	.w8(32'hbc3d0186),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c1534),
	.w1(32'hbb0f1575),
	.w2(32'h3b823801),
	.w3(32'h3bdbe84f),
	.w4(32'h3b97cf5c),
	.w5(32'h3b20faf0),
	.w6(32'h3b753e13),
	.w7(32'h3b97b23d),
	.w8(32'hbaa413fa),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8cf01),
	.w1(32'h3a6d02ed),
	.w2(32'hb8e59a36),
	.w3(32'hbb4c6c0e),
	.w4(32'hbbdf239f),
	.w5(32'hbc3c13fb),
	.w6(32'hba918371),
	.w7(32'h3b28cf3b),
	.w8(32'hba1efc44),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0966c),
	.w1(32'hbbb8d3dc),
	.w2(32'hbb9576e0),
	.w3(32'hbc08e0fd),
	.w4(32'h3994a776),
	.w5(32'hbb80a5f5),
	.w6(32'h3b4b6e2f),
	.w7(32'hbabc2081),
	.w8(32'hbb1ca7cb),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e080e),
	.w1(32'hbbcab73e),
	.w2(32'hbc01bbbc),
	.w3(32'h3afe0579),
	.w4(32'h3ae27965),
	.w5(32'h3ac9f885),
	.w6(32'hbb147270),
	.w7(32'hbba4545b),
	.w8(32'hbb89d072),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ecdf1),
	.w1(32'hbc203069),
	.w2(32'hbb291b64),
	.w3(32'hbb49bd74),
	.w4(32'hba8baeac),
	.w5(32'hbaf47a79),
	.w6(32'hbb4e93cf),
	.w7(32'hbb26a968),
	.w8(32'hbb47bed8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c1c42),
	.w1(32'hbbb45715),
	.w2(32'hbadb79e9),
	.w3(32'hbb1800fb),
	.w4(32'h3ba43fa1),
	.w5(32'h3acd5f4c),
	.w6(32'hbbaffe54),
	.w7(32'h3a2127b8),
	.w8(32'h3bd98ef0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8839e9a),
	.w1(32'hbba4e082),
	.w2(32'hbaefe79b),
	.w3(32'hbb599b61),
	.w4(32'hbb1c54b3),
	.w5(32'hbba59fb6),
	.w6(32'hbb600d8d),
	.w7(32'h3a1d100a),
	.w8(32'hbb8ea0de),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b6d0d),
	.w1(32'hbb462679),
	.w2(32'hbb8bfafb),
	.w3(32'hba773676),
	.w4(32'hbba214dc),
	.w5(32'hba941791),
	.w6(32'hbaa12866),
	.w7(32'hbb5e79c1),
	.w8(32'hba810903),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9270a3),
	.w1(32'h3bca5cc8),
	.w2(32'hba456be1),
	.w3(32'hbb190460),
	.w4(32'h3bda6226),
	.w5(32'h3c02d7cb),
	.w6(32'hbc00fe11),
	.w7(32'h3b0fbbd6),
	.w8(32'h3bd083ec),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf3f4d),
	.w1(32'hbc1e45c7),
	.w2(32'h3a9d0a42),
	.w3(32'hbb1f7424),
	.w4(32'hb98f3d1e),
	.w5(32'hbb1e6ed3),
	.w6(32'hbb7d16f0),
	.w7(32'hb7a1ed1c),
	.w8(32'hbb496644),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cbecc),
	.w1(32'hbbd7c876),
	.w2(32'hb9946ebe),
	.w3(32'h3a921047),
	.w4(32'h3aaf0431),
	.w5(32'h3a310e76),
	.w6(32'hbb9383fa),
	.w7(32'h3ab31467),
	.w8(32'h39060a03),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d983c),
	.w1(32'hbb238c76),
	.w2(32'hba341562),
	.w3(32'hbb163f12),
	.w4(32'h3a69ef4b),
	.w5(32'hba152b50),
	.w6(32'hbaef6edd),
	.w7(32'h3a88712e),
	.w8(32'hb9bc510a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9589837),
	.w1(32'hbb3b6a26),
	.w2(32'h3a345992),
	.w3(32'hbb732a53),
	.w4(32'h3ab4cf1c),
	.w5(32'h38858add),
	.w6(32'hbba3e0b7),
	.w7(32'h3afc7ab2),
	.w8(32'h3a20a085),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39375302),
	.w1(32'hbb0ffc47),
	.w2(32'h3b344350),
	.w3(32'hbb46e595),
	.w4(32'h3b7afead),
	.w5(32'hbacb0d9a),
	.w6(32'hbb2f8731),
	.w7(32'h3afafc8b),
	.w8(32'hbba494a7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d5028),
	.w1(32'h3aed2e12),
	.w2(32'h3b7e6402),
	.w3(32'hbbd4b906),
	.w4(32'h3bec3426),
	.w5(32'h3a9cbbcb),
	.w6(32'hbb7f4f1d),
	.w7(32'h3b3f704a),
	.w8(32'h3b1c8b96),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9892456),
	.w1(32'h3b344380),
	.w2(32'hbac29066),
	.w3(32'h3c0ad46c),
	.w4(32'h3c0d6b2d),
	.w5(32'hbaf20f2a),
	.w6(32'h3b1309b2),
	.w7(32'h3be3e74d),
	.w8(32'h3abc381b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13cda4),
	.w1(32'hbb8fb0f0),
	.w2(32'h3b98dbce),
	.w3(32'h3c142b8b),
	.w4(32'h3b8ac9ed),
	.w5(32'hba1aca48),
	.w6(32'hba8af9b9),
	.w7(32'hb6a59190),
	.w8(32'hb9365e23),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa78963),
	.w1(32'hbb5dd542),
	.w2(32'h3a135b04),
	.w3(32'h3a90ffd0),
	.w4(32'hbbad9f88),
	.w5(32'hbc051916),
	.w6(32'hbb80f4d0),
	.w7(32'hbb444499),
	.w8(32'hbba0802c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c2c39),
	.w1(32'h3b9f42c9),
	.w2(32'h3b912f69),
	.w3(32'hbb9a5d22),
	.w4(32'hb9c57d16),
	.w5(32'h3bfcf503),
	.w6(32'hbba353f6),
	.w7(32'h3a8647ce),
	.w8(32'h3b8cc119),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038467),
	.w1(32'h3bab641e),
	.w2(32'hbbcf7ac5),
	.w3(32'h3aa41722),
	.w4(32'h3b11ad89),
	.w5(32'h3bb097d2),
	.w6(32'h3b3ba24c),
	.w7(32'hba422202),
	.w8(32'h3a3faaef),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5aa6d),
	.w1(32'h3bc66e95),
	.w2(32'hbaa00e5f),
	.w3(32'h3c3d3eb2),
	.w4(32'hbb958114),
	.w5(32'hb9ffe8b6),
	.w6(32'h3c327e68),
	.w7(32'hbace2dd2),
	.w8(32'h3a53e5db),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e77d4),
	.w1(32'h3a850d85),
	.w2(32'h3ad59b43),
	.w3(32'hbb7b75d3),
	.w4(32'h3c078c22),
	.w5(32'hbadb2ff4),
	.w6(32'h3a4ed2d2),
	.w7(32'h3bc0e929),
	.w8(32'hbb2d70de),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a04a6),
	.w1(32'hbb75f326),
	.w2(32'hbab05d21),
	.w3(32'hbb53d09a),
	.w4(32'hbae743db),
	.w5(32'hbbc14962),
	.w6(32'hbb8a7217),
	.w7(32'hbb788825),
	.w8(32'hbb93cb41),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16842),
	.w1(32'hb9b1e737),
	.w2(32'h3bc4c71d),
	.w3(32'hbb3c70ce),
	.w4(32'hb8bf0cb0),
	.w5(32'h3ad9b961),
	.w6(32'hbb5e8a62),
	.w7(32'hba9fe2ba),
	.w8(32'h3ba5f2be),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d90ca),
	.w1(32'hbaa27ed9),
	.w2(32'h3a21c27d),
	.w3(32'h3c191cfa),
	.w4(32'h3a49f661),
	.w5(32'hbab6598a),
	.w6(32'hba02776a),
	.w7(32'h37426845),
	.w8(32'h3a16d85d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b909874),
	.w1(32'h3bf4f1db),
	.w2(32'h3ab5b7c6),
	.w3(32'hbb146c67),
	.w4(32'h3bf51d38),
	.w5(32'h3b8b3ed0),
	.w6(32'h39d33627),
	.w7(32'h39f87acb),
	.w8(32'h3b2169b3),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b343b3f),
	.w1(32'hbacc70ce),
	.w2(32'h3b8c1db6),
	.w3(32'h3bb93655),
	.w4(32'hbb65c5ff),
	.w5(32'h3a03f4e8),
	.w6(32'hba52de26),
	.w7(32'hbaa0fc32),
	.w8(32'hbb343ed7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97a8885),
	.w1(32'hbb96674b),
	.w2(32'h3b4dd8d6),
	.w3(32'h3abf39db),
	.w4(32'h3c154714),
	.w5(32'h3bb73516),
	.w6(32'hbbaa6ef5),
	.w7(32'h3bbd4298),
	.w8(32'h3b93a255),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6d6e0),
	.w1(32'hba8c69de),
	.w2(32'hba8d0fe8),
	.w3(32'h3ab58d9c),
	.w4(32'hb9f4903e),
	.w5(32'hba00c7bc),
	.w6(32'hb9752021),
	.w7(32'hb9629e08),
	.w8(32'hb80df139),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8de09e),
	.w1(32'hbadd6f17),
	.w2(32'h3b667162),
	.w3(32'hbaaabb5f),
	.w4(32'h3c2bdea0),
	.w5(32'h3c8a7bd5),
	.w6(32'hbabee3f7),
	.w7(32'h3c05c732),
	.w8(32'h3bccd5ee),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58ee81),
	.w1(32'hba734222),
	.w2(32'h3b5e5437),
	.w3(32'h3b93ed5d),
	.w4(32'h3a844fb8),
	.w5(32'hb92bbb10),
	.w6(32'h3b8bbd95),
	.w7(32'h3bb7a11c),
	.w8(32'h3c0b46ed),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af700f4),
	.w1(32'h3bf33df7),
	.w2(32'hbae953eb),
	.w3(32'h3b7fedf2),
	.w4(32'h3c3ea0a5),
	.w5(32'h3af4a675),
	.w6(32'h3ba9c404),
	.w7(32'h3b9be348),
	.w8(32'h3c132df7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b038886),
	.w1(32'h3b0e650d),
	.w2(32'h3ba33398),
	.w3(32'h3b6c72b3),
	.w4(32'h3b8de3e6),
	.w5(32'hbaa3b4a1),
	.w6(32'h39e44635),
	.w7(32'h3b99d189),
	.w8(32'hba7d9f2b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392418d7),
	.w1(32'h3ad41555),
	.w2(32'h3a42edd4),
	.w3(32'h3ad7698d),
	.w4(32'hbb433383),
	.w5(32'hbbc73121),
	.w6(32'h3ab2d2cd),
	.w7(32'hbb99bccb),
	.w8(32'hbb182714),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10f84d),
	.w1(32'hbb9293a2),
	.w2(32'h3b896a07),
	.w3(32'hbae00d48),
	.w4(32'hb99cdb32),
	.w5(32'h39866d94),
	.w6(32'hbc07f2c0),
	.w7(32'h3a86ce9d),
	.w8(32'h39a34181),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87127),
	.w1(32'h3b4d36a8),
	.w2(32'hbacd2724),
	.w3(32'h3b8bddbc),
	.w4(32'hbb816044),
	.w5(32'hbb8afbfb),
	.w6(32'h3b8d85c7),
	.w7(32'hbade2801),
	.w8(32'hbb4da075),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7224f),
	.w1(32'hbb205517),
	.w2(32'h3bcde6b2),
	.w3(32'hb800eea0),
	.w4(32'h3c2b0d14),
	.w5(32'h3c45a613),
	.w6(32'h39fa4f2a),
	.w7(32'h3c0f7359),
	.w8(32'h3b024d1a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b1290),
	.w1(32'h3bb16d7c),
	.w2(32'h38ad49ed),
	.w3(32'h3c0a1562),
	.w4(32'hbaa95e90),
	.w5(32'h3a4b3fc9),
	.w6(32'h3ba32149),
	.w7(32'hbafe311c),
	.w8(32'hbb1f942a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5af080),
	.w1(32'hba8ba499),
	.w2(32'h3b8355fb),
	.w3(32'hbaa07d8a),
	.w4(32'h3942bd9e),
	.w5(32'h3b8fd1a3),
	.w6(32'hba7849c3),
	.w7(32'h3b34ed3d),
	.w8(32'h3c2ed45c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c177f75),
	.w1(32'h3c48184c),
	.w2(32'hb80a691a),
	.w3(32'hbaa88153),
	.w4(32'h3aa35c46),
	.w5(32'hbb5d8ee0),
	.w6(32'h3c12087a),
	.w7(32'hba2f90dd),
	.w8(32'hbae835ac),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b4cc5),
	.w1(32'hb9f96688),
	.w2(32'h3c16b0b4),
	.w3(32'hb8fc13dc),
	.w4(32'hbacd5cc8),
	.w5(32'h3babca87),
	.w6(32'hbb30667f),
	.w7(32'h3bb07fdc),
	.w8(32'hbb8d60b6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b001c06),
	.w1(32'h3a2b7a11),
	.w2(32'hba35714f),
	.w3(32'h3a1d9a5b),
	.w4(32'h3a8aae73),
	.w5(32'h396df361),
	.w6(32'h3b874d47),
	.w7(32'h3ad2aac1),
	.w8(32'h3a6ab3fa),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba139f21),
	.w1(32'hbb61cad8),
	.w2(32'hbaf036ed),
	.w3(32'hbb60de31),
	.w4(32'hbba0878d),
	.w5(32'h3b71b906),
	.w6(32'hbb3d5e27),
	.w7(32'hbae9722f),
	.w8(32'h39ca4722),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae4d8a),
	.w1(32'h3a94f9d5),
	.w2(32'h3ba32a48),
	.w3(32'h3bde9ee4),
	.w4(32'h3bf4ffee),
	.w5(32'hbb7a8f3e),
	.w6(32'h3af5d3e3),
	.w7(32'h3c2a8b53),
	.w8(32'hba2327e8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39558a),
	.w1(32'h3b44063f),
	.w2(32'h3b15a407),
	.w3(32'h3c2422ce),
	.w4(32'hbabbaa07),
	.w5(32'hb8e3afd5),
	.w6(32'h3c3d03ee),
	.w7(32'h3b9d1f4b),
	.w8(32'hbb7470a0),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba5763),
	.w1(32'h3a8f50e4),
	.w2(32'hba4a158e),
	.w3(32'h3b916553),
	.w4(32'hbb7a8c32),
	.w5(32'hbbcd9a93),
	.w6(32'h3afe4c91),
	.w7(32'hbbd9e11f),
	.w8(32'hbb88259e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afed189),
	.w1(32'hbbb25b4e),
	.w2(32'h3b59849e),
	.w3(32'h3c14f7e5),
	.w4(32'h3c7a5a4e),
	.w5(32'h3b622884),
	.w6(32'h3a254270),
	.w7(32'h3bbc83ac),
	.w8(32'h3c115131),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf44952),
	.w1(32'h3c0e1f94),
	.w2(32'h3ba63336),
	.w3(32'h3c232ff2),
	.w4(32'h3bcdbc6f),
	.w5(32'h3ba22e11),
	.w6(32'h3ac963da),
	.w7(32'h3b01643e),
	.w8(32'hba16c8b8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b720f61),
	.w1(32'h3c209cc2),
	.w2(32'hb98ebc04),
	.w3(32'h3c018951),
	.w4(32'h3c0a560d),
	.w5(32'hbb937ea2),
	.w6(32'h3be4f0cf),
	.w7(32'h3b43bd45),
	.w8(32'h3b6dd786),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032a1a),
	.w1(32'h3acff58c),
	.w2(32'hbb356595),
	.w3(32'h3b757329),
	.w4(32'hbbb97429),
	.w5(32'hba88cc6c),
	.w6(32'h3c092f7f),
	.w7(32'hbc0989aa),
	.w8(32'hbb85bcfd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad35824),
	.w1(32'h3bab6f79),
	.w2(32'h3940479d),
	.w3(32'h3b3eeefd),
	.w4(32'h3a1933b1),
	.w5(32'h3c3aefa2),
	.w6(32'h3b4d5ed2),
	.w7(32'h3bc44dac),
	.w8(32'h3c340a99),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb377c9f),
	.w1(32'hbc1a2c69),
	.w2(32'hbad37959),
	.w3(32'h39de0d79),
	.w4(32'h3a78abbd),
	.w5(32'h3a2b661c),
	.w6(32'hbb41807f),
	.w7(32'h381cc07b),
	.w8(32'hb9f99f23),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3e70),
	.w1(32'hbb818d7d),
	.w2(32'h3c1a2d6f),
	.w3(32'hbb1780ca),
	.w4(32'h3a8333b0),
	.w5(32'hbb25b87d),
	.w6(32'hbb4f5252),
	.w7(32'h3a936834),
	.w8(32'hbbd53ec8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2cab7),
	.w1(32'hbb2bb510),
	.w2(32'h3b3f9a6a),
	.w3(32'h3bde17d7),
	.w4(32'h3b9cb38b),
	.w5(32'h3b696ed6),
	.w6(32'h3acfce2f),
	.w7(32'h399d2b04),
	.w8(32'h3ba68f0f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9a8f4),
	.w1(32'h3bc59f73),
	.w2(32'hbb84ad3b),
	.w3(32'h3ba13863),
	.w4(32'h3adf0d20),
	.w5(32'hbaee0a69),
	.w6(32'h3bc6e658),
	.w7(32'hbb1ca515),
	.w8(32'hbb83b6f6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9482c0),
	.w1(32'hbb923716),
	.w2(32'h3ba6d864),
	.w3(32'hbb36d0aa),
	.w4(32'h3b88001e),
	.w5(32'hbac7279a),
	.w6(32'hbb818fb8),
	.w7(32'hba98a823),
	.w8(32'hbb88c1db),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079f29),
	.w1(32'hbb2b2b70),
	.w2(32'hbac3e65e),
	.w3(32'hbb7bf39c),
	.w4(32'h3a97d07b),
	.w5(32'h3818d1f7),
	.w6(32'hbb2f70f6),
	.w7(32'h3a86e2bf),
	.w8(32'hb8a39af1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5cea),
	.w1(32'hbb773fac),
	.w2(32'h3c72a03d),
	.w3(32'hbb4dc198),
	.w4(32'h3a19e589),
	.w5(32'hbb5f5501),
	.w6(32'hbb702f1b),
	.w7(32'hb92b379a),
	.w8(32'h3ab7f886),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61ca6b),
	.w1(32'h378b7202),
	.w2(32'h39d00182),
	.w3(32'hba70ac80),
	.w4(32'hbb4870c2),
	.w5(32'hba79b045),
	.w6(32'h3b42648d),
	.w7(32'h3bbcb664),
	.w8(32'h3b5c0d5b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e29c),
	.w1(32'h3c0626b3),
	.w2(32'h38457d42),
	.w3(32'h3b13ee84),
	.w4(32'hbb1c7b90),
	.w5(32'hbba35842),
	.w6(32'h3c74ae97),
	.w7(32'hb8eb0913),
	.w8(32'hbba5cf87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbdc02),
	.w1(32'h3a446961),
	.w2(32'hbb635db4),
	.w3(32'hbb661697),
	.w4(32'hb92750cc),
	.w5(32'h3bfea7b9),
	.w6(32'hbb29e699),
	.w7(32'h3ade6ff1),
	.w8(32'h3bc88978),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7821b8),
	.w1(32'h3ac601d6),
	.w2(32'hbb6719b8),
	.w3(32'h3b8af123),
	.w4(32'hb9db0195),
	.w5(32'h3b954a7e),
	.w6(32'h3bd7a737),
	.w7(32'hbb795cdb),
	.w8(32'hb945386c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba48bc),
	.w1(32'hbaf78e65),
	.w2(32'hb9c7808d),
	.w3(32'h3b2bc0aa),
	.w4(32'hbb0a7028),
	.w5(32'hbaf85f6d),
	.w6(32'hba121e61),
	.w7(32'hbaf2f5d7),
	.w8(32'hbb23e18d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace1c09),
	.w1(32'h3912ffdc),
	.w2(32'hbbaf79a6),
	.w3(32'hb977fbaf),
	.w4(32'hba1fb530),
	.w5(32'hbb08699e),
	.w6(32'hbb33674f),
	.w7(32'hbb7bfd51),
	.w8(32'h3a89e27b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05d8c6),
	.w1(32'h3b30b028),
	.w2(32'h3b9d1df8),
	.w3(32'h3add56c2),
	.w4(32'h3bc92de1),
	.w5(32'h3bb02760),
	.w6(32'h3a7c3547),
	.w7(32'h3c607c0f),
	.w8(32'hb9bc5ed0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b921c47),
	.w1(32'hbbae3808),
	.w2(32'h3b9dff8c),
	.w3(32'hba6dd952),
	.w4(32'hba682acd),
	.w5(32'h3bb8c02b),
	.w6(32'hbbda5081),
	.w7(32'h3c04f8b4),
	.w8(32'h3b57f496),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33764c),
	.w1(32'hb9f4a28b),
	.w2(32'h3bc51569),
	.w3(32'h3a3b4ca9),
	.w4(32'h3b90fd0b),
	.w5(32'h3af61b1d),
	.w6(32'h3b8f54d4),
	.w7(32'hba0f6ee6),
	.w8(32'hb99964bf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a5353),
	.w1(32'hba429da3),
	.w2(32'hba794f43),
	.w3(32'h3bf0c6e6),
	.w4(32'h39be6a53),
	.w5(32'h3ac65449),
	.w6(32'h3b181228),
	.w7(32'hba1cb0d2),
	.w8(32'h3b1dedbf),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5bb340),
	.w1(32'h3ba130cb),
	.w2(32'hbb8dc974),
	.w3(32'hbb0d59c6),
	.w4(32'h3ad13be8),
	.w5(32'hbb41010c),
	.w6(32'h3adc207c),
	.w7(32'hbbcb2349),
	.w8(32'h3bfedba8),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b874878),
	.w1(32'h3c1e427c),
	.w2(32'hbbf54e06),
	.w3(32'hbb8f7547),
	.w4(32'h3b362bf2),
	.w5(32'h3b099b9e),
	.w6(32'hba21136b),
	.w7(32'hbaf9cb44),
	.w8(32'h3cac4cdf),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d593),
	.w1(32'h3c22e764),
	.w2(32'hbb5df691),
	.w3(32'h3b615e39),
	.w4(32'hbba4892b),
	.w5(32'hba48f81e),
	.w6(32'h3c203aa7),
	.w7(32'hbbf9ba32),
	.w8(32'hb987a6cb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0937b2),
	.w1(32'h3b82f834),
	.w2(32'h3b2a731c),
	.w3(32'h39cbca76),
	.w4(32'h3b603b6e),
	.w5(32'hbbfdd16f),
	.w6(32'h3b557d66),
	.w7(32'h3ae6e177),
	.w8(32'h3bc6ea3e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8a471),
	.w1(32'h39c8f39f),
	.w2(32'h3c4d89b4),
	.w3(32'hbbda40f9),
	.w4(32'h3c802634),
	.w5(32'h3bfe0650),
	.w6(32'hbae43ae7),
	.w7(32'h3c8abd10),
	.w8(32'h3b3e86c5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f0c5),
	.w1(32'h3a97af22),
	.w2(32'h3a99fd0a),
	.w3(32'h3b2c1ee1),
	.w4(32'h3b991147),
	.w5(32'h3b4c669b),
	.w6(32'hbab8f3d5),
	.w7(32'h3a543332),
	.w8(32'h3bbebbbd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae79a6c),
	.w1(32'h3c4e3427),
	.w2(32'hba035b13),
	.w3(32'h3c078d83),
	.w4(32'hb9e2badc),
	.w5(32'h3b5e7dee),
	.w6(32'h3c1a843e),
	.w7(32'h3ab070ce),
	.w8(32'h3c053c2d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0a99),
	.w1(32'h39d0d75d),
	.w2(32'hbaede786),
	.w3(32'h3ad97da1),
	.w4(32'hbb2b3723),
	.w5(32'h3b1ef983),
	.w6(32'h3b4d8128),
	.w7(32'h3b5fcc76),
	.w8(32'h3c5d2ddb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e964f),
	.w1(32'h3999989e),
	.w2(32'hba28ca48),
	.w3(32'hba53b2c1),
	.w4(32'hbaf99578),
	.w5(32'hb9f8b005),
	.w6(32'h3bbcf9b8),
	.w7(32'h3b240367),
	.w8(32'h3bc73d66),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebb9e8),
	.w1(32'h3a21b488),
	.w2(32'h3a172307),
	.w3(32'hbadf23c0),
	.w4(32'hbb81802d),
	.w5(32'h3a0dcd06),
	.w6(32'h3b622772),
	.w7(32'hba5863aa),
	.w8(32'h3b617e27),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80207c),
	.w1(32'hbb1520a9),
	.w2(32'hbae8d580),
	.w3(32'hbb2a7220),
	.w4(32'hbacd311b),
	.w5(32'hba9f68a7),
	.w6(32'h3b252224),
	.w7(32'hbb210db0),
	.w8(32'hbadde6f2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1849c2),
	.w1(32'h3a057c64),
	.w2(32'hbb44209b),
	.w3(32'h3a4a01ea),
	.w4(32'hbb8fca7f),
	.w5(32'hbb7a2dbf),
	.w6(32'h3b31bf04),
	.w7(32'hbb96b39e),
	.w8(32'hbb6e1d02),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aca1b),
	.w1(32'h3c2731d0),
	.w2(32'hbaa4098c),
	.w3(32'hbadec009),
	.w4(32'hbb4cba3b),
	.w5(32'h3aa898c8),
	.w6(32'h3c42a65c),
	.w7(32'hbada3b43),
	.w8(32'h3b4c3aa0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e739),
	.w1(32'hbaec1ef7),
	.w2(32'hba6826cf),
	.w3(32'h3b99ac42),
	.w4(32'hba87311e),
	.w5(32'hbb2a3042),
	.w6(32'h3bb16bad),
	.w7(32'h3c6a5d0d),
	.w8(32'h3cb885eb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca35f1),
	.w1(32'h3a037c36),
	.w2(32'h3b478b7d),
	.w3(32'h3a56194c),
	.w4(32'h3b9e19a3),
	.w5(32'h3c08997b),
	.w6(32'h3c90d691),
	.w7(32'hb8efbb22),
	.w8(32'h3b863549),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4266ac),
	.w1(32'h39861fb8),
	.w2(32'hbb187895),
	.w3(32'hbb1b089e),
	.w4(32'hba915b70),
	.w5(32'h3bfc3759),
	.w6(32'hbb8ce56d),
	.w7(32'hbaba1442),
	.w8(32'h3c207fef),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca604ba),
	.w1(32'h3b834f04),
	.w2(32'hbb91ea99),
	.w3(32'h3b06ff63),
	.w4(32'hbb3db3fd),
	.w5(32'hbad54a9c),
	.w6(32'h37676a86),
	.w7(32'h397e201d),
	.w8(32'h3a8e60d6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c76e2),
	.w1(32'hbb573bbf),
	.w2(32'h388f6116),
	.w3(32'hbb4868b4),
	.w4(32'h3a77299c),
	.w5(32'hbab1e9b2),
	.w6(32'hbb1ce535),
	.w7(32'h3a98dec8),
	.w8(32'h3a7dfe42),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a19cc),
	.w1(32'h3a2826e6),
	.w2(32'h3b415bf6),
	.w3(32'h38da9584),
	.w4(32'h3ba96da2),
	.w5(32'hba9a63bd),
	.w6(32'h3b40ecdd),
	.w7(32'h3b93d77c),
	.w8(32'hbb089133),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f5c31),
	.w1(32'hba01ee19),
	.w2(32'hba99fb57),
	.w3(32'h3a5e7644),
	.w4(32'hb9115000),
	.w5(32'hba0dcd5c),
	.w6(32'h388c3bd3),
	.w7(32'hba1ff182),
	.w8(32'hbb8f2875),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8323bc),
	.w1(32'hb9d73177),
	.w2(32'h3b92b808),
	.w3(32'h3ab82774),
	.w4(32'h3b7dba8a),
	.w5(32'h3aebd635),
	.w6(32'hb8847f81),
	.w7(32'h3c766989),
	.w8(32'h3c38605b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b216bfe),
	.w1(32'hb8e8a811),
	.w2(32'h3afcbcc1),
	.w3(32'h37232809),
	.w4(32'hb8955a0f),
	.w5(32'hbb6bc9fc),
	.w6(32'h3bd59900),
	.w7(32'hba9429e8),
	.w8(32'hbbb80a93),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2035),
	.w1(32'h3aa401e4),
	.w2(32'h39b7c03b),
	.w3(32'hbadd6260),
	.w4(32'hbb754619),
	.w5(32'hbb1bc0c2),
	.w6(32'hbc0c47d1),
	.w7(32'hbba31340),
	.w8(32'hbb7028bc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8b046),
	.w1(32'hbbcc2f84),
	.w2(32'hb7d6fd46),
	.w3(32'hbb656357),
	.w4(32'hbb0eb6af),
	.w5(32'hba21672e),
	.w6(32'hbc0629fe),
	.w7(32'hbab94284),
	.w8(32'h3abe32b8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88e5c5),
	.w1(32'h3b5be775),
	.w2(32'h3b1fe95b),
	.w3(32'h381eae3c),
	.w4(32'h3b525bca),
	.w5(32'h3c2849fd),
	.w6(32'h3a9296a8),
	.w7(32'h3c077d69),
	.w8(32'h3c8f44a4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dcf31),
	.w1(32'h3b3cd97d),
	.w2(32'h3ba31f37),
	.w3(32'h3b8d207b),
	.w4(32'hbb581910),
	.w5(32'hb9abd5f6),
	.w6(32'h3c1aabd4),
	.w7(32'hbc082c2e),
	.w8(32'hbba042cc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdb65a),
	.w1(32'h3b91714a),
	.w2(32'hbb0ef389),
	.w3(32'hbb6ee748),
	.w4(32'hbb246d94),
	.w5(32'hbb2ded30),
	.w6(32'hbbf9949d),
	.w7(32'h39c2de5d),
	.w8(32'h3b956a9c),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17610f),
	.w1(32'hbac96aad),
	.w2(32'h3b52160a),
	.w3(32'hb8d1081e),
	.w4(32'h3ab42177),
	.w5(32'h3abb39cf),
	.w6(32'h3b202ae2),
	.w7(32'h3a39ef2f),
	.w8(32'hb9ed6873),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa20199),
	.w1(32'hbb53e7c5),
	.w2(32'h3976be25),
	.w3(32'h3b73e394),
	.w4(32'hb9486ea1),
	.w5(32'h3a0dce18),
	.w6(32'h3bac66e3),
	.w7(32'hb94e6ca6),
	.w8(32'h3a4e2aa9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3ad7c),
	.w1(32'hb98a338f),
	.w2(32'hbbc6fe88),
	.w3(32'h396f104a),
	.w4(32'hba7aba7b),
	.w5(32'h3ac3910b),
	.w6(32'hba4e6d8c),
	.w7(32'hbb0f5789),
	.w8(32'h3b54c36a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf5a88),
	.w1(32'h3af0c0ab),
	.w2(32'h3b04b41e),
	.w3(32'h3b77c3ac),
	.w4(32'hbb3ff682),
	.w5(32'hb9084df5),
	.w6(32'hbb082dce),
	.w7(32'hb984cfb1),
	.w8(32'hba4b9b5d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb059284),
	.w1(32'h3ac5cbc8),
	.w2(32'h39178f84),
	.w3(32'hba1e107c),
	.w4(32'h3b0adfce),
	.w5(32'h3921ef4b),
	.w6(32'hbb2f3f21),
	.w7(32'h3a396861),
	.w8(32'hbb24e0de),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3da2af),
	.w1(32'hbb6c2f0f),
	.w2(32'h3b9230aa),
	.w3(32'h39b8b40d),
	.w4(32'hbabe2579),
	.w5(32'hbaee0443),
	.w6(32'hbb2c6f0a),
	.w7(32'h3ac3742a),
	.w8(32'h3a9daaa2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6648d),
	.w1(32'hbafa0265),
	.w2(32'h3b8064e9),
	.w3(32'hbaa923ac),
	.w4(32'h39bb8cae),
	.w5(32'hbabe71b2),
	.w6(32'h3c0b81ca),
	.w7(32'h3b82feb9),
	.w8(32'h3b04d555),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d3ee2),
	.w1(32'h3b0c488b),
	.w2(32'hbb79a306),
	.w3(32'hba34bff3),
	.w4(32'hbbbcc433),
	.w5(32'h3ae116ab),
	.w6(32'h3b114615),
	.w7(32'h3b87f197),
	.w8(32'h3c8831ee),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad6a2a),
	.w1(32'hbbddb4c8),
	.w2(32'hbb0358ab),
	.w3(32'hbaa62a95),
	.w4(32'h3a150273),
	.w5(32'hba9aec7c),
	.w6(32'h3b832324),
	.w7(32'hba6c43a0),
	.w8(32'hbbac9971),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd846fd),
	.w1(32'hbb61acbd),
	.w2(32'hb9d37f09),
	.w3(32'hba4e5a4a),
	.w4(32'h3a973124),
	.w5(32'h3b6b1df8),
	.w6(32'hbb85f30e),
	.w7(32'hbb34332e),
	.w8(32'hbbfea12e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba993574),
	.w1(32'h3b340aa3),
	.w2(32'hba2e213a),
	.w3(32'h3b4f2f2c),
	.w4(32'hb9a88e20),
	.w5(32'h3b94ff31),
	.w6(32'hbb9f8c90),
	.w7(32'h3b234164),
	.w8(32'h3c2f8d72),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c05af),
	.w1(32'h3a4d1eb1),
	.w2(32'h3b88a181),
	.w3(32'h3b4b3e84),
	.w4(32'h3b83858d),
	.w5(32'h3b281a4b),
	.w6(32'h3ba5b189),
	.w7(32'h3b4390b9),
	.w8(32'hbb023885),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c538),
	.w1(32'hb8bd949a),
	.w2(32'h3b7e69d9),
	.w3(32'h390bdf2c),
	.w4(32'h3b918e6c),
	.w5(32'hbba51ab2),
	.w6(32'hbb61fa2f),
	.w7(32'h3a0c92e6),
	.w8(32'hbbb020f8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf573dc),
	.w1(32'h39ad7067),
	.w2(32'h3aad66e4),
	.w3(32'hba80c62e),
	.w4(32'h3ac53243),
	.w5(32'hbb3ec995),
	.w6(32'hbb315962),
	.w7(32'h3a0d58c3),
	.w8(32'hbab5647c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb667aac),
	.w1(32'h3b5bb261),
	.w2(32'h3b2a4c71),
	.w3(32'h3a17f17c),
	.w4(32'h3b9c46b7),
	.w5(32'hba3dee42),
	.w6(32'hbaeb4382),
	.w7(32'h3b866eb6),
	.w8(32'hbb0cec68),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3492c6),
	.w1(32'h3a7289fa),
	.w2(32'h3b290a4d),
	.w3(32'h3b3cc6f0),
	.w4(32'h3b5a057f),
	.w5(32'hba4e6d62),
	.w6(32'hbb16702e),
	.w7(32'hbb65e80d),
	.w8(32'hbba4bef2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0325d6),
	.w1(32'h3b8479e5),
	.w2(32'h3b97a159),
	.w3(32'hbae33f4b),
	.w4(32'h3ae25940),
	.w5(32'hbb10f1be),
	.w6(32'hbae37dab),
	.w7(32'h3b2a847f),
	.w8(32'h3b6a79a2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a1e7b),
	.w1(32'h3b1e69c0),
	.w2(32'h3b57d318),
	.w3(32'hbb49625e),
	.w4(32'hbaf64084),
	.w5(32'hb9826fed),
	.w6(32'h3ac1005f),
	.w7(32'hba9e3e2f),
	.w8(32'hba97dd93),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7437f),
	.w1(32'hbabb9626),
	.w2(32'h3b630836),
	.w3(32'h3af26316),
	.w4(32'h3b5f46fd),
	.w5(32'h3a649fb9),
	.w6(32'hbb0915a2),
	.w7(32'h3b483653),
	.w8(32'hbb12318f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c34c8),
	.w1(32'h3ba0ef1d),
	.w2(32'h3b8e52ea),
	.w3(32'h3b8360cb),
	.w4(32'h3a921e2d),
	.w5(32'hba830d0d),
	.w6(32'h3b853930),
	.w7(32'hbae02b09),
	.w8(32'hbbb94fe8),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d5c00),
	.w1(32'hbade6f05),
	.w2(32'hba4892f0),
	.w3(32'h3b2b7af1),
	.w4(32'hba871de6),
	.w5(32'h3bbded50),
	.w6(32'hba629573),
	.w7(32'h3b32e0b4),
	.w8(32'h3c46ac57),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef4eb),
	.w1(32'h3a654668),
	.w2(32'h3a222278),
	.w3(32'h3b15e613),
	.w4(32'hbb7d13d2),
	.w5(32'hbbbdc62a),
	.w6(32'h3bb3ad56),
	.w7(32'h3a96ba01),
	.w8(32'hbba90522),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c5aac),
	.w1(32'hbb572bdb),
	.w2(32'h3b2070ba),
	.w3(32'hb94d5597),
	.w4(32'hba540f1f),
	.w5(32'hbb4c5a38),
	.w6(32'hbaabd50e),
	.w7(32'h3a072ed7),
	.w8(32'hba8b31c4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d78c5),
	.w1(32'hbafae18e),
	.w2(32'h3b5670fe),
	.w3(32'h39b39192),
	.w4(32'h3a2442b8),
	.w5(32'hb9e07633),
	.w6(32'hbb38559a),
	.w7(32'h3aea89f1),
	.w8(32'h397b4c3e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53b9b2),
	.w1(32'h3ba8ce36),
	.w2(32'hbaf9291a),
	.w3(32'h39ffdb84),
	.w4(32'h3a17cea0),
	.w5(32'h3ac85a8b),
	.w6(32'h3b0ec4ae),
	.w7(32'hba7ad978),
	.w8(32'hbb845e81),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97faa96),
	.w1(32'h3af01e0a),
	.w2(32'h398ddb71),
	.w3(32'h3b5b23f8),
	.w4(32'hb8bd3827),
	.w5(32'h3bda10d5),
	.w6(32'hbb512e10),
	.w7(32'h3b706921),
	.w8(32'h3c6600c1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1ee4e),
	.w1(32'h3ae49bd6),
	.w2(32'h3b85ea58),
	.w3(32'h3b71ca71),
	.w4(32'h3a3b26b5),
	.w5(32'hbac15901),
	.w6(32'h3be917b8),
	.w7(32'hba223a04),
	.w8(32'hbbcecc7b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c813),
	.w1(32'h3b549521),
	.w2(32'hbb0656c3),
	.w3(32'hb88a5d5c),
	.w4(32'hb9eab409),
	.w5(32'h3b614133),
	.w6(32'hbbc06b2d),
	.w7(32'h3acd7d1d),
	.w8(32'h3bd40c83),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4aeaa),
	.w1(32'hbb816852),
	.w2(32'h3acc8ea2),
	.w3(32'h3b09134a),
	.w4(32'h3b363d53),
	.w5(32'h3b52b48d),
	.w6(32'hbbb2643d),
	.w7(32'h3b04c0bc),
	.w8(32'hb936c855),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2255f0),
	.w1(32'hb9dfe608),
	.w2(32'hbb26bae2),
	.w3(32'h3acced8d),
	.w4(32'hba7d6ab9),
	.w5(32'hb8814e47),
	.w6(32'hb72d303c),
	.w7(32'hbb257f59),
	.w8(32'h3bc5e7f1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be25653),
	.w1(32'hbbd146ae),
	.w2(32'h3a34fd5b),
	.w3(32'hbb0b2b72),
	.w4(32'hba61fd3e),
	.w5(32'hbbcaf358),
	.w6(32'hbba80706),
	.w7(32'h3bcca776),
	.w8(32'h3b3a055a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule