module layer_8_featuremap_217(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c457f8e),
	.w1(32'h3b07b1f5),
	.w2(32'hbcb70954),
	.w3(32'h3c835735),
	.w4(32'h3c113f3d),
	.w5(32'hbccc42c8),
	.w6(32'h3c5df4b8),
	.w7(32'h3a43d84e),
	.w8(32'hbc1bbd15),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70edc5),
	.w1(32'h3b033e31),
	.w2(32'h3b69c17d),
	.w3(32'h38c8e235),
	.w4(32'h3b39e915),
	.w5(32'h3ba82946),
	.w6(32'h3a5529bc),
	.w7(32'h3a8d7990),
	.w8(32'h3bbb865c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e613),
	.w1(32'hbba5c619),
	.w2(32'hba78c9ac),
	.w3(32'hbb1f8382),
	.w4(32'hbb3065f7),
	.w5(32'h3aad4583),
	.w6(32'hbb875874),
	.w7(32'hbb73a1f7),
	.w8(32'h3abdc95e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c9aba),
	.w1(32'hbc862840),
	.w2(32'hbc1ff7a6),
	.w3(32'hbb98ed64),
	.w4(32'hbca246ee),
	.w5(32'hbc87883a),
	.w6(32'h393f9f6d),
	.w7(32'hbc3d7db8),
	.w8(32'hbc1ecc89),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c689dd),
	.w1(32'h3ace7242),
	.w2(32'h3af08133),
	.w3(32'hbb42d9d8),
	.w4(32'h3af8cc41),
	.w5(32'h3ad3ca00),
	.w6(32'h3b13bafa),
	.w7(32'h3bb579ee),
	.w8(32'h3b35ce29),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ba27e),
	.w1(32'hbc3a3e1e),
	.w2(32'h3bb20690),
	.w3(32'hbc2c6c8f),
	.w4(32'hbb715c89),
	.w5(32'h3b451ef2),
	.w6(32'hbad3a214),
	.w7(32'h3ca27a92),
	.w8(32'h3c89bdf1),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6019f3),
	.w1(32'hbaf0e9bf),
	.w2(32'hbb046edf),
	.w3(32'hb977165d),
	.w4(32'hbab61942),
	.w5(32'hbb0b37f8),
	.w6(32'hbacdec18),
	.w7(32'hbb01301d),
	.w8(32'hbabe1fb6),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4bbb6),
	.w1(32'h3a001cab),
	.w2(32'hbb80ea57),
	.w3(32'h3b61b245),
	.w4(32'hbab38669),
	.w5(32'hbbed94a1),
	.w6(32'hbb03ecb1),
	.w7(32'hbaf3ea4f),
	.w8(32'hbc03ac4c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24c2d3),
	.w1(32'h3b38488e),
	.w2(32'h3b6bd84e),
	.w3(32'hbb4ec3d7),
	.w4(32'h3b46c89f),
	.w5(32'h3b4cb8e2),
	.w6(32'h3bad589a),
	.w7(32'h3b9a3768),
	.w8(32'h3bd64a52),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8883af),
	.w1(32'h3a1679cb),
	.w2(32'hbc9a2d92),
	.w3(32'h3b9f264c),
	.w4(32'hbbceae2b),
	.w5(32'hbcacac60),
	.w6(32'hba188df9),
	.w7(32'hbca63b5e),
	.w8(32'hbc7653bb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a5f79),
	.w1(32'hbca31383),
	.w2(32'hbcd2f1ab),
	.w3(32'h3bd03433),
	.w4(32'hbb3aa72c),
	.w5(32'hbce03b6f),
	.w6(32'h3c28ad0f),
	.w7(32'h3bb3f994),
	.w8(32'hbc8327da),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9578ff),
	.w1(32'hb963f78c),
	.w2(32'hbc21aebc),
	.w3(32'h3b46d3fe),
	.w4(32'h3b19e6b5),
	.w5(32'hbc22b603),
	.w6(32'hbc1660da),
	.w7(32'hbc0fb503),
	.w8(32'h3a6d3716),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9349f2),
	.w1(32'h3af0073a),
	.w2(32'h3ba60db7),
	.w3(32'hb9ffd2af),
	.w4(32'hbae77d9f),
	.w5(32'h3b8da20f),
	.w6(32'hba426b17),
	.w7(32'hba68631f),
	.w8(32'h3b7aae63),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4a30),
	.w1(32'hbb751cdb),
	.w2(32'hbba741cb),
	.w3(32'hba08e9aa),
	.w4(32'hbac2004e),
	.w5(32'hbba59534),
	.w6(32'hbb175189),
	.w7(32'hbb8110e9),
	.w8(32'hba855f94),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29cbb3),
	.w1(32'h3b2b1820),
	.w2(32'h3ad89775),
	.w3(32'hbb57920d),
	.w4(32'h3b1ad528),
	.w5(32'h3ab57c6e),
	.w6(32'h3b2c283e),
	.w7(32'h3b03e329),
	.w8(32'h3b097246),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac95ddb),
	.w1(32'h3a06c10a),
	.w2(32'hbab94f6e),
	.w3(32'h3a91df69),
	.w4(32'h39baa353),
	.w5(32'hba0312fe),
	.w6(32'h3a95db42),
	.w7(32'hba09b58b),
	.w8(32'hba176fe2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd82fcb),
	.w1(32'h3bc04630),
	.w2(32'hbb22eeb2),
	.w3(32'h3c343a68),
	.w4(32'h3bc0ac7e),
	.w5(32'hbbaf6055),
	.w6(32'h3c350075),
	.w7(32'h3bf02715),
	.w8(32'hb825ad7c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2eb12e),
	.w1(32'h3ab51520),
	.w2(32'hbba88947),
	.w3(32'hbba88e85),
	.w4(32'hbaf8d44f),
	.w5(32'hbb897c0d),
	.w6(32'hbc58fdff),
	.w7(32'hbc51fc29),
	.w8(32'h3abe87fc),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d087b8f),
	.w1(32'hbc8420bd),
	.w2(32'hbd96979f),
	.w3(32'h3d894f39),
	.w4(32'h3cbfca88),
	.w5(32'hbd793d91),
	.w6(32'h3d506eea),
	.w7(32'h3b704738),
	.w8(32'hbd0abab6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85c6f0),
	.w1(32'h3c990c0f),
	.w2(32'h3c37a78b),
	.w3(32'hbbbc2a02),
	.w4(32'hba88a93a),
	.w5(32'h3b54d3b2),
	.w6(32'h3b9f4a55),
	.w7(32'h3a9a42a9),
	.w8(32'h3c4b7032),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbc15b),
	.w1(32'h3bbc8b70),
	.w2(32'hbc0a34ff),
	.w3(32'hbaa8b97b),
	.w4(32'h3cb20b62),
	.w5(32'hbb9430ba),
	.w6(32'h3bfba596),
	.w7(32'h3d037f4f),
	.w8(32'h3b96e65f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f83d5),
	.w1(32'h3badd325),
	.w2(32'h3c5cec15),
	.w3(32'h3aad75a9),
	.w4(32'h3bafa24e),
	.w5(32'h3c8b86fe),
	.w6(32'hbac2056d),
	.w7(32'hb879074f),
	.w8(32'h3c0f775f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c770efe),
	.w1(32'hbbc5d539),
	.w2(32'hbd91ed87),
	.w3(32'h3d11031a),
	.w4(32'h3b172d9d),
	.w5(32'hbda25c3a),
	.w6(32'h3cf61aec),
	.w7(32'h3c1e7b61),
	.w8(32'hbd1baf52),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90762c),
	.w1(32'h3ba2a8cf),
	.w2(32'h3c13b910),
	.w3(32'hbb0fb88b),
	.w4(32'h3ab1bf1b),
	.w5(32'h3b8bfdd2),
	.w6(32'h3b46f7e9),
	.w7(32'h3be08d93),
	.w8(32'h3b96a0e3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d93746),
	.w1(32'h3aff634e),
	.w2(32'h3ad53a23),
	.w3(32'hbb0cb759),
	.w4(32'h3a465dc6),
	.w5(32'h3aaf3b5a),
	.w6(32'h3b7c0679),
	.w7(32'h3b5c0213),
	.w8(32'h3b330a1a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba08051),
	.w1(32'h3b7d2e05),
	.w2(32'hbc79cddb),
	.w3(32'h3c35a6b4),
	.w4(32'h3b87866d),
	.w5(32'hbc9f4ac6),
	.w6(32'h3bbe0738),
	.w7(32'h3c0af110),
	.w8(32'hb7b62c76),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f9ec2),
	.w1(32'h3b7cb88e),
	.w2(32'h3b1de547),
	.w3(32'hbb753cb1),
	.w4(32'h3a4416ad),
	.w5(32'hb83bf645),
	.w6(32'h3bb1ad01),
	.w7(32'h3bc092cc),
	.w8(32'h3b825a4f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d398d30),
	.w1(32'hbc07e977),
	.w2(32'hbd234b3f),
	.w3(32'h3d9f5783),
	.w4(32'h3db2ebe7),
	.w5(32'hbd0579d5),
	.w6(32'h3dbb8b94),
	.w7(32'h3dc76047),
	.w8(32'h3b60d122),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c3418),
	.w1(32'h397efe86),
	.w2(32'hbc3a1e20),
	.w3(32'h3b6c8b0c),
	.w4(32'hbb9786c2),
	.w5(32'hbc84e371),
	.w6(32'hba6c3c7f),
	.w7(32'hbb8eff65),
	.w8(32'hbc1b8fff),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaec67),
	.w1(32'hba682f3e),
	.w2(32'hb8975aeb),
	.w3(32'hbb26bc02),
	.w4(32'hbb4823cb),
	.w5(32'hbb2b7769),
	.w6(32'h397b281d),
	.w7(32'h39c1a3a8),
	.w8(32'hbae7e7c4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc8975),
	.w1(32'hbb7d8600),
	.w2(32'hbbc47f2f),
	.w3(32'hbb503f97),
	.w4(32'hbb7d5305),
	.w5(32'hbbe454e0),
	.w6(32'hbb2c9109),
	.w7(32'hbb481fec),
	.w8(32'hbbcb8c09),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacbf1e2),
	.w1(32'h3a80ab68),
	.w2(32'hbb532ded),
	.w3(32'hbaf6fa68),
	.w4(32'h3b9cc6bc),
	.w5(32'h3b0edd4a),
	.w6(32'h3b3bdcf1),
	.w7(32'h3c118f3d),
	.w8(32'h3b08fab8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb904915),
	.w1(32'h3b1f74b7),
	.w2(32'h3b337d28),
	.w3(32'hbb5a9dd5),
	.w4(32'h3b307dfc),
	.w5(32'h3a9b8696),
	.w6(32'h3b8913e9),
	.w7(32'h3b356254),
	.w8(32'h3b829f85),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2acf58),
	.w1(32'h3a0a82e4),
	.w2(32'hba843f21),
	.w3(32'h3b84c64c),
	.w4(32'hb8f6fd17),
	.w5(32'hba9c6d04),
	.w6(32'hba5f945a),
	.w7(32'hba220d18),
	.w8(32'hba0bd4e2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd0cc0),
	.w1(32'h3bbe936f),
	.w2(32'h3c3ec327),
	.w3(32'hbbcebb85),
	.w4(32'hbb4f5d08),
	.w5(32'h3c5e6dc6),
	.w6(32'hbb516aba),
	.w7(32'hbb6a8277),
	.w8(32'h3c1d12d8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c599562),
	.w1(32'h3c5fce9b),
	.w2(32'hbc5b59df),
	.w3(32'h3cb0c472),
	.w4(32'h3cb839b8),
	.w5(32'hbbe8c564),
	.w6(32'h3c66a8d6),
	.w7(32'h3c4c7cfe),
	.w8(32'hbb884d19),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872012),
	.w1(32'h376dc9e7),
	.w2(32'h39b3fa93),
	.w3(32'h37f4fa2b),
	.w4(32'hba547a26),
	.w5(32'h3861eafc),
	.w6(32'h39081a93),
	.w7(32'h3a89179c),
	.w8(32'h3af0f1e6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07c4f),
	.w1(32'h3a359989),
	.w2(32'h3b010c88),
	.w3(32'hbae3705a),
	.w4(32'h3a1faa2b),
	.w5(32'h3ad9cf11),
	.w6(32'h3ab74166),
	.w7(32'h3aa0e283),
	.w8(32'h3b177870),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb83eb),
	.w1(32'hbb2a0eb9),
	.w2(32'hbb8f34b0),
	.w3(32'h3a18b937),
	.w4(32'hbb00be18),
	.w5(32'hbb66926a),
	.w6(32'hbb1a91d4),
	.w7(32'hbb8518aa),
	.w8(32'hbb0d565e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7cd19),
	.w1(32'hbb2c1537),
	.w2(32'hbb4ce755),
	.w3(32'hba0bd543),
	.w4(32'hbab41723),
	.w5(32'hbb0be5cf),
	.w6(32'h38fda6ac),
	.w7(32'hbac9facc),
	.w8(32'hbb15c3d5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a1ce8),
	.w1(32'hbcd9c373),
	.w2(32'hbc8029d5),
	.w3(32'hbc5ac72f),
	.w4(32'hbd26363e),
	.w5(32'hbd0d249f),
	.w6(32'hbcb023dc),
	.w7(32'hbd256e26),
	.w8(32'hbc367610),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f2aa6),
	.w1(32'h3c586f4c),
	.w2(32'h3bcf1266),
	.w3(32'h3caa56de),
	.w4(32'h3c5e8369),
	.w5(32'h3a7a792f),
	.w6(32'h3cc17234),
	.w7(32'h3c569f27),
	.w8(32'hb9a581e8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94799e),
	.w1(32'h3b163c62),
	.w2(32'h3b718964),
	.w3(32'h3ba3264d),
	.w4(32'h3b691bdd),
	.w5(32'h3baed2a9),
	.w6(32'h3a9c6bd0),
	.w7(32'h3b0941a9),
	.w8(32'h3ba25a20),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6cc58),
	.w1(32'hbbe8cfc5),
	.w2(32'hbc8c7351),
	.w3(32'h3b1b72c1),
	.w4(32'hb995c6d7),
	.w5(32'hbc9b332d),
	.w6(32'hbac5a2f1),
	.w7(32'hb9fdfec8),
	.w8(32'hbc049a27),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc70015),
	.w1(32'hbb6024ba),
	.w2(32'hbd040daf),
	.w3(32'h3c9356b0),
	.w4(32'h3ad54163),
	.w5(32'hbd1e1413),
	.w6(32'h3cb70ffd),
	.w7(32'h3c7f5441),
	.w8(32'hbca964da),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4e330),
	.w1(32'h3bcbdf6b),
	.w2(32'hbc886f45),
	.w3(32'h3cc06fea),
	.w4(32'h3b06600a),
	.w5(32'hbc8b4018),
	.w6(32'h3c53fd4b),
	.w7(32'hbbc4047e),
	.w8(32'hbc5cb927),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a258f),
	.w1(32'hbb251b59),
	.w2(32'hbb7ff53b),
	.w3(32'hbaea4076),
	.w4(32'hba9e02d8),
	.w5(32'hbb1976ff),
	.w6(32'hbb083c04),
	.w7(32'hbb60b321),
	.w8(32'hbb4561c4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c828fc1),
	.w1(32'h3bcd8cb1),
	.w2(32'hbcf53e00),
	.w3(32'h3d0ad9c8),
	.w4(32'h3cb57bb3),
	.w5(32'hbd0283ef),
	.w6(32'h3cf3f151),
	.w7(32'h3cb04844),
	.w8(32'hbc56ca99),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933e57),
	.w1(32'hba34774c),
	.w2(32'h3a737176),
	.w3(32'h3961f85e),
	.w4(32'hbad67b44),
	.w5(32'h3a6b1565),
	.w6(32'h3a9eab52),
	.w7(32'hb9d4003e),
	.w8(32'h3a800eb2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34b789),
	.w1(32'hbc859f4f),
	.w2(32'hbcc89eca),
	.w3(32'h3b49bcda),
	.w4(32'hbc5106af),
	.w5(32'hbcf79e90),
	.w6(32'hbb12d012),
	.w7(32'hbc694d55),
	.w8(32'hbc6a7b67),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e40eb),
	.w1(32'h3c8e40c1),
	.w2(32'h3b969c49),
	.w3(32'h3ad6d055),
	.w4(32'h3c62b7ff),
	.w5(32'h3c0992ef),
	.w6(32'hbb4c9060),
	.w7(32'h3bab7e74),
	.w8(32'h3c29506d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af34679),
	.w1(32'hbb5177da),
	.w2(32'hbcdacac3),
	.w3(32'h3cddcdae),
	.w4(32'hbbaefdf8),
	.w5(32'hbd247cc7),
	.w6(32'h3d30965b),
	.w7(32'h3c8b00a1),
	.w8(32'hbce8c414),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78f322),
	.w1(32'hbba23858),
	.w2(32'hbc3d122d),
	.w3(32'h3b08981e),
	.w4(32'hbb82c055),
	.w5(32'hbc2ca483),
	.w6(32'h3bae3b3e),
	.w7(32'h3ad137b8),
	.w8(32'hbb63e49d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c914f07),
	.w1(32'h3c988175),
	.w2(32'hbc5d8184),
	.w3(32'hb893ad2f),
	.w4(32'hbb41c0a4),
	.w5(32'hbcbee1ee),
	.w6(32'hbb49dcc0),
	.w7(32'hbca43800),
	.w8(32'hbc924fb7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61e2d2),
	.w1(32'h3aed50c1),
	.w2(32'hbb33116b),
	.w3(32'hbac6e0ed),
	.w4(32'h3af40390),
	.w5(32'hb9417299),
	.w6(32'h3a4e515c),
	.w7(32'hbac96515),
	.w8(32'hba9fd8f8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7d7142),
	.w1(32'h3d02b20f),
	.w2(32'hbd219846),
	.w3(32'h3d4420d7),
	.w4(32'h3d14206f),
	.w5(32'hbd02e4c2),
	.w6(32'h3ccc4baf),
	.w7(32'h3c0f924f),
	.w8(32'hbc5244c0),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd59d92),
	.w1(32'h3bc4b6f6),
	.w2(32'hbaf30b49),
	.w3(32'h3ad7363f),
	.w4(32'hbba6c4ea),
	.w5(32'hbc2accb6),
	.w6(32'h3bc9d7e5),
	.w7(32'h3ab46629),
	.w8(32'hbaa14032),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d4dc),
	.w1(32'h3b3c9b0c),
	.w2(32'hbb5e0815),
	.w3(32'h3c3d2d6f),
	.w4(32'h3a944a61),
	.w5(32'hbc177020),
	.w6(32'h3c623833),
	.w7(32'h3c34165d),
	.w8(32'hbc0d5cc8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b8a4),
	.w1(32'h3b54b833),
	.w2(32'hbc6cb9ff),
	.w3(32'h3c2dd33b),
	.w4(32'h3c14dd12),
	.w5(32'hbc824969),
	.w6(32'h3cadab9d),
	.w7(32'h3ca919f3),
	.w8(32'hbb85a237),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf108f7),
	.w1(32'hbb92273a),
	.w2(32'hbc0fd8c0),
	.w3(32'h3a81565d),
	.w4(32'hbc1be0f6),
	.w5(32'hbc0b034c),
	.w6(32'h3bdc535d),
	.w7(32'h3b5a878c),
	.w8(32'hbbcc034d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93f436),
	.w1(32'hb9ff8959),
	.w2(32'hbb39c658),
	.w3(32'hbb372334),
	.w4(32'hbab710f6),
	.w5(32'hbb7d46ca),
	.w6(32'h3b7d6bd0),
	.w7(32'hb92fc85e),
	.w8(32'hb9d98b6b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc563d),
	.w1(32'h3a42f85d),
	.w2(32'hbaabc223),
	.w3(32'hbac9e877),
	.w4(32'h3a8e12b4),
	.w5(32'hbab79697),
	.w6(32'h3ba09200),
	.w7(32'h3a3aefb9),
	.w8(32'hba3e0478),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c74b943),
	.w1(32'hb8d2488b),
	.w2(32'hbc56e9a3),
	.w3(32'h3c314aab),
	.w4(32'hbc4d5b0e),
	.w5(32'hbcff1661),
	.w6(32'hbc0204d9),
	.w7(32'hbcd3d866),
	.w8(32'hbc8dfb1f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2418e2),
	.w1(32'h3a5738f7),
	.w2(32'h3b15d2cb),
	.w3(32'hbb01c099),
	.w4(32'hb94e6c6f),
	.w5(32'h3b2c931d),
	.w6(32'h3ac7405d),
	.w7(32'h3ac69349),
	.w8(32'h3a84ed63),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b113a96),
	.w1(32'h3ac95f80),
	.w2(32'h3af7c718),
	.w3(32'h3b2b9524),
	.w4(32'h3ad27cc5),
	.w5(32'h3ad308b5),
	.w6(32'h3a7a10cc),
	.w7(32'h3af4aab4),
	.w8(32'h3aae7dcb),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc75ae0),
	.w1(32'h3b2b87a8),
	.w2(32'hba6cb3df),
	.w3(32'h3c36c564),
	.w4(32'h3c162232),
	.w5(32'h39d32fa1),
	.w6(32'h3bdd3029),
	.w7(32'h3bf0883f),
	.w8(32'h39a70c7f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572c3f),
	.w1(32'hbac662a6),
	.w2(32'h3b6624a3),
	.w3(32'hbaaa90fe),
	.w4(32'h3aa685ab),
	.w5(32'h3b7232f4),
	.w6(32'h3b5d62c5),
	.w7(32'h3bb5282b),
	.w8(32'h3bd98e5b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf168c1),
	.w1(32'h3c990aac),
	.w2(32'hbb04c579),
	.w3(32'h3c968ef8),
	.w4(32'h3c900c21),
	.w5(32'h3a26782a),
	.w6(32'h3bc33401),
	.w7(32'h3b095ed6),
	.w8(32'h3bb1d65c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb511e11),
	.w1(32'hb9f2cf1b),
	.w2(32'hbaa8e873),
	.w3(32'hbaacea67),
	.w4(32'h3a781c03),
	.w5(32'hbb47c832),
	.w6(32'hba96d049),
	.w7(32'hbb0e1c9c),
	.w8(32'h398f290f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04539d),
	.w1(32'hbc66c18d),
	.w2(32'hbd776d07),
	.w3(32'h3ca2b1ee),
	.w4(32'h3cf64ba6),
	.w5(32'hbd5249c4),
	.w6(32'h3d416205),
	.w7(32'h3d5be66e),
	.w8(32'hbc5e3ee8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86a7e2),
	.w1(32'h3b20b1b3),
	.w2(32'h3af9a89f),
	.w3(32'hbb2b0abb),
	.w4(32'h3acd0774),
	.w5(32'h3a6d8ad5),
	.w6(32'h3b896357),
	.w7(32'h3b545fe9),
	.w8(32'h3b41cda0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b133e78),
	.w1(32'hbbdaa0ab),
	.w2(32'hbba04efc),
	.w3(32'h3aedb7c1),
	.w4(32'hbb961746),
	.w5(32'hbbdcd31b),
	.w6(32'h3b97f82d),
	.w7(32'h3ac07558),
	.w8(32'h3b0e2f77),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a04b8),
	.w1(32'hba5cc0da),
	.w2(32'hba9510c4),
	.w3(32'hba4d3578),
	.w4(32'hbb33f629),
	.w5(32'hbb1a24af),
	.w6(32'hb970fb23),
	.w7(32'hba7bcd55),
	.w8(32'hba2be740),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39effd),
	.w1(32'h3bd17205),
	.w2(32'hbc774ced),
	.w3(32'hbc1f675b),
	.w4(32'h3a97c280),
	.w5(32'hbc3e752f),
	.w6(32'hbbffd5e8),
	.w7(32'hbc59d36e),
	.w8(32'hbbeea085),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d11a8),
	.w1(32'hbac08510),
	.w2(32'hbb4cd1ec),
	.w3(32'hba8e8356),
	.w4(32'hba8f3d7f),
	.w5(32'hbb34f62a),
	.w6(32'hb830e91c),
	.w7(32'hbb0a79f3),
	.w8(32'hbb02fc60),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b83b),
	.w1(32'hbb2f42ba),
	.w2(32'hbbbbf5bb),
	.w3(32'h3b0204bb),
	.w4(32'hbaceeec7),
	.w5(32'hbbc346b6),
	.w6(32'h3bc28ce4),
	.w7(32'h3bb207cf),
	.w8(32'hbb995b4f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9e79f),
	.w1(32'h3ab0f76f),
	.w2(32'hba785c76),
	.w3(32'hbb8f63d9),
	.w4(32'h3a912857),
	.w5(32'hba866054),
	.w6(32'h3b243575),
	.w7(32'h36fa3994),
	.w8(32'hba6a62fd),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8a0aa),
	.w1(32'hbbdf6713),
	.w2(32'hbcadfdde),
	.w3(32'h3c2f7c1e),
	.w4(32'h3c81fb34),
	.w5(32'hbc44c87b),
	.w6(32'h3ca37ea0),
	.w7(32'h3c724959),
	.w8(32'hba392593),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce8baea),
	.w1(32'h3c3008df),
	.w2(32'hbc8af205),
	.w3(32'h3c8ab2b0),
	.w4(32'hbb84911e),
	.w5(32'hbca6cd7b),
	.w6(32'h3c8c0cb7),
	.w7(32'hbc0474ba),
	.w8(32'hbc890ca6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a679041),
	.w1(32'hba42c73b),
	.w2(32'h3ad0b66f),
	.w3(32'h38f667dd),
	.w4(32'hb9eb9bc3),
	.w5(32'hb9c3c9df),
	.w6(32'h3980811a),
	.w7(32'hb98836c8),
	.w8(32'hba03fc39),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b97ee8),
	.w1(32'hbb3bb8b4),
	.w2(32'hbb785e3b),
	.w3(32'hbada17f5),
	.w4(32'hba065098),
	.w5(32'hbb05274b),
	.w6(32'hb9f2765c),
	.w7(32'hbaf10101),
	.w8(32'hbad852c5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7112d),
	.w1(32'hbc3a8aba),
	.w2(32'hbbd1cc28),
	.w3(32'hbc150523),
	.w4(32'hbb363cec),
	.w5(32'hbc2b5b14),
	.w6(32'h3ca4c661),
	.w7(32'h3cd3e4ac),
	.w8(32'hbb2805c3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c029da9),
	.w1(32'hbb105121),
	.w2(32'hbc872ee2),
	.w3(32'h3c522530),
	.w4(32'hb9d94846),
	.w5(32'hbcc43388),
	.w6(32'h3c04d40b),
	.w7(32'h3a9ccf9d),
	.w8(32'hbc333f44),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c5963),
	.w1(32'h3b81971b),
	.w2(32'hbc654264),
	.w3(32'hbc8d782c),
	.w4(32'hbd5b20c8),
	.w5(32'hbca81af8),
	.w6(32'hbc6cf9f6),
	.w7(32'hbd371ce8),
	.w8(32'hbc2b96e4),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b800ecf),
	.w1(32'hbbb1c20f),
	.w2(32'hbd3ec9db),
	.w3(32'h3cbb004c),
	.w4(32'hbb0a0989),
	.w5(32'hbd681651),
	.w6(32'h3b3063f0),
	.w7(32'hbac9a789),
	.w8(32'hbcc8faf2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc582b62),
	.w1(32'hbca8f8d1),
	.w2(32'hbc8936ef),
	.w3(32'h3ae755be),
	.w4(32'hbcc0ba94),
	.w5(32'hbd020cee),
	.w6(32'h3c50e43a),
	.w7(32'h3be5cd2b),
	.w8(32'hbc75fcfb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58e4f9),
	.w1(32'hbace5c4e),
	.w2(32'hbaaabb8b),
	.w3(32'hbb075715),
	.w4(32'hbaa55a4e),
	.w5(32'hbaa80d4d),
	.w6(32'hbb02c626),
	.w7(32'hbad61455),
	.w8(32'hbb1a5db2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8807f1),
	.w1(32'h37c8dbbc),
	.w2(32'h396081af),
	.w3(32'hba3a5ae3),
	.w4(32'h390dd972),
	.w5(32'h3aba1d3a),
	.w6(32'h3b48fd1e),
	.w7(32'h3b4cbec4),
	.w8(32'h3b864549),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888fb3),
	.w1(32'h3957835f),
	.w2(32'h377350b7),
	.w3(32'h3b032558),
	.w4(32'hb9b1ab88),
	.w5(32'hb9f28361),
	.w6(32'hb98cea4a),
	.w7(32'h388ace56),
	.w8(32'hb97e3d91),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8003f0),
	.w1(32'hb9d8a4ee),
	.w2(32'hbb7b4b8e),
	.w3(32'h3b9284f9),
	.w4(32'hbaebbdae),
	.w5(32'hbb872597),
	.w6(32'h3b5f22ed),
	.w7(32'h39426b71),
	.w8(32'hbba3c8a4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ad32f),
	.w1(32'hbb9f8cf3),
	.w2(32'hbb8b87fe),
	.w3(32'hbbb0e71c),
	.w4(32'hbbf40a48),
	.w5(32'hbc09b0d4),
	.w6(32'h3874ccd0),
	.w7(32'h3a92fc60),
	.w8(32'hbb60ec07),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048f27),
	.w1(32'hba4b95c0),
	.w2(32'hba3ef9d0),
	.w3(32'hba939fa3),
	.w4(32'hba81f2a7),
	.w5(32'hba3f3a61),
	.w6(32'hbaaf5929),
	.w7(32'hbaa8cb50),
	.w8(32'hba2602da),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79048d),
	.w1(32'hbb0132e3),
	.w2(32'h3c1b4b87),
	.w3(32'hbc918772),
	.w4(32'hbc129782),
	.w5(32'h3bc6fde3),
	.w6(32'hbb6e4e20),
	.w7(32'h3a480c67),
	.w8(32'h3bfa46b9),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d98d5),
	.w1(32'hbaa6dc93),
	.w2(32'hbbd33480),
	.w3(32'h3b2f8bc7),
	.w4(32'hbba313ba),
	.w5(32'hbc2b2517),
	.w6(32'hbae5b90c),
	.w7(32'hbbefaa0a),
	.w8(32'hbbfe4f7f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8308ec),
	.w1(32'h3c0a0831),
	.w2(32'h3b850215),
	.w3(32'h3bbdd701),
	.w4(32'h3ba11d58),
	.w5(32'h3bcf6044),
	.w6(32'h3ab0a0e8),
	.w7(32'h39928226),
	.w8(32'h3bddf8bd),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb9ede0),
	.w1(32'h3cb2fb7d),
	.w2(32'hbbba0670),
	.w3(32'h3cc78902),
	.w4(32'h3c85a10c),
	.w5(32'hbc05e8a3),
	.w6(32'h3cadc985),
	.w7(32'h3c1d86f1),
	.w8(32'hbc14df7e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170020),
	.w1(32'h3a5d7e74),
	.w2(32'hbbf05aab),
	.w3(32'h3c0ebdaa),
	.w4(32'hbb059b6e),
	.w5(32'hbc2ffef0),
	.w6(32'h3c5a6410),
	.w7(32'h3a713b67),
	.w8(32'hbbe4dc52),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea358e),
	.w1(32'hbba965b7),
	.w2(32'hbbf2e075),
	.w3(32'hbbb47adf),
	.w4(32'hbb94f0ab),
	.w5(32'hbbd98db0),
	.w6(32'hbb9fe8a0),
	.w7(32'hbbec91c5),
	.w8(32'hbb4b7431),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73ba2c),
	.w1(32'hba1c252d),
	.w2(32'hbb8869b0),
	.w3(32'hbb655f2a),
	.w4(32'hba0459c3),
	.w5(32'hbb749c6f),
	.w6(32'hba97e113),
	.w7(32'hbb346e1a),
	.w8(32'hba93c458),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb8da9),
	.w1(32'hbac12906),
	.w2(32'hba986e2f),
	.w3(32'hbaf90267),
	.w4(32'hbade291b),
	.w5(32'hbaf0f34d),
	.w6(32'hb9b8e825),
	.w7(32'h3ae9d40f),
	.w8(32'h3b0599ae),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a514782),
	.w1(32'h3a9fcd4e),
	.w2(32'h3a27ce2b),
	.w3(32'hbb037a00),
	.w4(32'h3b34ac6f),
	.w5(32'h3b8bea37),
	.w6(32'h3aaf0b1f),
	.w7(32'h3aa7bfbc),
	.w8(32'hbaaf5131),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba704ced),
	.w1(32'hbb1b53b6),
	.w2(32'h39a6dc72),
	.w3(32'h39e25148),
	.w4(32'hbaff125e),
	.w5(32'hba89eaeb),
	.w6(32'h3b0a848f),
	.w7(32'h3ae7099f),
	.w8(32'h3b2d7430),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ccf36),
	.w1(32'hba37c710),
	.w2(32'hbabeafac),
	.w3(32'h3a492186),
	.w4(32'hba3e5156),
	.w5(32'hbb01dca8),
	.w6(32'hba42621a),
	.w7(32'hba4317b2),
	.w8(32'hb96483cb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10447a),
	.w1(32'hba8b897e),
	.w2(32'h3c1b88db),
	.w3(32'hbc51723f),
	.w4(32'hbc29efe0),
	.w5(32'h3b18ffdd),
	.w6(32'h3baafa9e),
	.w7(32'h3c023151),
	.w8(32'h3bfc3b03),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab8371),
	.w1(32'hbabd41e4),
	.w2(32'h3bd030a1),
	.w3(32'hbbb77425),
	.w4(32'hbb9e45d6),
	.w5(32'h3b938f0b),
	.w6(32'hbafaecb9),
	.w7(32'h38a091bf),
	.w8(32'h3ad7954e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0867b8),
	.w1(32'hbbcef790),
	.w2(32'hbd059223),
	.w3(32'h3c349ec3),
	.w4(32'h3c594376),
	.w5(32'hbcfa830e),
	.w6(32'h3caf43b8),
	.w7(32'h3cd31188),
	.w8(32'hbc0b951c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d60ad6),
	.w1(32'h3b315053),
	.w2(32'hb981dc71),
	.w3(32'h3a3175d8),
	.w4(32'h3a20f51a),
	.w5(32'hba96b28d),
	.w6(32'h3b5647d8),
	.w7(32'h3b07f0e9),
	.w8(32'h3a13f79f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4939fa),
	.w1(32'h3c001f0c),
	.w2(32'h3c19ba6f),
	.w3(32'hbb401bac),
	.w4(32'h3b52051a),
	.w5(32'h3c0f1580),
	.w6(32'h3b32c58a),
	.w7(32'h3b1ac21f),
	.w8(32'h3bf190d6),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccdbd6),
	.w1(32'hbb016184),
	.w2(32'h39d4dee9),
	.w3(32'hbb5cbed5),
	.w4(32'hbb84cdba),
	.w5(32'hb8c5746d),
	.w6(32'hbb994989),
	.w7(32'hbb567a45),
	.w8(32'hba95a18d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0fec1),
	.w1(32'hbb8324b3),
	.w2(32'hbb59df40),
	.w3(32'h3a78dd87),
	.w4(32'hbb5e94c9),
	.w5(32'hbb3a3088),
	.w6(32'h39df1b79),
	.w7(32'hbb029120),
	.w8(32'hbabe386f),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7dc8cf),
	.w1(32'h3c91adc6),
	.w2(32'h3c582e50),
	.w3(32'h3b0c1dbc),
	.w4(32'h3c17fcc0),
	.w5(32'h3c0cfda0),
	.w6(32'hbb067f1a),
	.w7(32'h3ab9bdf2),
	.w8(32'h3c2c91c5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addec21),
	.w1(32'hbb0bbc5f),
	.w2(32'h3b34d0bc),
	.w3(32'h39d8e682),
	.w4(32'hb98e3e68),
	.w5(32'h3bc3bd29),
	.w6(32'hbbe3a74b),
	.w7(32'hbb66d7d1),
	.w8(32'h3b48cd59),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5c547),
	.w1(32'hbba1a256),
	.w2(32'hbac9086c),
	.w3(32'hbb616b56),
	.w4(32'hbb8724a8),
	.w5(32'h3acf357e),
	.w6(32'hbb25158d),
	.w7(32'hbbb36287),
	.w8(32'h3b0f088e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08cf1f),
	.w1(32'hba4dac83),
	.w2(32'hbacbc520),
	.w3(32'hbb5cbfae),
	.w4(32'hbace69f0),
	.w5(32'hbb006bdc),
	.w6(32'h3a10f779),
	.w7(32'hb90defba),
	.w8(32'hba69e50d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2dae1e),
	.w1(32'h3a7df021),
	.w2(32'hbafb6c45),
	.w3(32'h3adcd6ce),
	.w4(32'hbb533d8e),
	.w5(32'hbb43da28),
	.w6(32'h3b834a92),
	.w7(32'h397aa31c),
	.w8(32'hb7cd8c44),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac01df2),
	.w1(32'hba93303a),
	.w2(32'hbafd372c),
	.w3(32'hb93cfcb4),
	.w4(32'hbadb6f11),
	.w5(32'hbb327fd2),
	.w6(32'hbb0f151e),
	.w7(32'hbad8cb6a),
	.w8(32'hbb2cd59e),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4a723),
	.w1(32'h3bbffa47),
	.w2(32'h3bd76584),
	.w3(32'hbaf249b2),
	.w4(32'hba3bce6d),
	.w5(32'hb996e86b),
	.w6(32'h3bc0f796),
	.w7(32'h3baf1fc3),
	.w8(32'h3bb169f2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14baa5),
	.w1(32'h3b57f955),
	.w2(32'hbbef87e1),
	.w3(32'h3c1c6e45),
	.w4(32'h3b80c3bc),
	.w5(32'hbc4ac3e5),
	.w6(32'h3c03a241),
	.w7(32'hbb0d1689),
	.w8(32'hbb7d5121),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3050a6),
	.w1(32'hbb90c669),
	.w2(32'hbbbb9d46),
	.w3(32'hbb16b606),
	.w4(32'hbb993096),
	.w5(32'hbb8bbc94),
	.w6(32'hba9f40f1),
	.w7(32'hbb19d21e),
	.w8(32'hbb17df09),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947f50f),
	.w1(32'h3aa16516),
	.w2(32'hbb57993a),
	.w3(32'h3810c22d),
	.w4(32'h39d7b07b),
	.w5(32'hbb4ede30),
	.w6(32'h3af380c2),
	.w7(32'hbb15f989),
	.w8(32'hbb561e26),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15cf08),
	.w1(32'h3c38d0d7),
	.w2(32'hba4f83fb),
	.w3(32'hbc28fcf7),
	.w4(32'hbc89276f),
	.w5(32'hbc900068),
	.w6(32'h3bb727c5),
	.w7(32'hbb44a51e),
	.w8(32'hbbef5d83),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4641d2),
	.w1(32'hb9c466b3),
	.w2(32'h3a4bf565),
	.w3(32'h3bee6f26),
	.w4(32'h38d9b97d),
	.w5(32'h3b1980f8),
	.w6(32'h3bc25cdb),
	.w7(32'h3abedf8c),
	.w8(32'h3a84203a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe71f5),
	.w1(32'hba9b5813),
	.w2(32'hbacef3c0),
	.w3(32'h3915c304),
	.w4(32'hbaa58a55),
	.w5(32'hba673940),
	.w6(32'hbad8d6a5),
	.w7(32'hba8ef815),
	.w8(32'hba1f7b64),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51253e),
	.w1(32'hbb8d7d4a),
	.w2(32'hbb96bb00),
	.w3(32'hbb2eac87),
	.w4(32'hbb4437d4),
	.w5(32'hbb81b343),
	.w6(32'hbb97dd00),
	.w7(32'hbbb92797),
	.w8(32'hbb712b6e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77d80),
	.w1(32'hbaa498d5),
	.w2(32'hba150f40),
	.w3(32'hbb6dc67d),
	.w4(32'hb9a0d105),
	.w5(32'hb94173aa),
	.w6(32'hb9c9c60b),
	.w7(32'hbad089ec),
	.w8(32'hbafacbfd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2523e4),
	.w1(32'h3c811e53),
	.w2(32'h3a364ac3),
	.w3(32'h3b47ba6a),
	.w4(32'h3c773f22),
	.w5(32'h3b06ba7f),
	.w6(32'h3be2e814),
	.w7(32'h3bcaf147),
	.w8(32'hbaad8395),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5829cb),
	.w1(32'h3afed45c),
	.w2(32'hbb7e8d6d),
	.w3(32'h3be90930),
	.w4(32'h3b337a1f),
	.w5(32'h38d38242),
	.w6(32'h3b96f0ca),
	.w7(32'h3a4203c1),
	.w8(32'hba2b11dd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29a262),
	.w1(32'h3bf7e02b),
	.w2(32'hbca6bce4),
	.w3(32'h3c929f0d),
	.w4(32'h3bf888a6),
	.w5(32'hbc91ff5d),
	.w6(32'h3c72a842),
	.w7(32'h3bdb3663),
	.w8(32'hbbeed151),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule