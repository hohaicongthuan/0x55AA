module layer_10_featuremap_415(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3daf65),
	.w1(32'hbb5b1ec8),
	.w2(32'hba990240),
	.w3(32'hbbb6af51),
	.w4(32'hbc427450),
	.w5(32'hbc12aaf0),
	.w6(32'hbb83c3a9),
	.w7(32'h3b3cd6b6),
	.w8(32'h3c052a9f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1deed7),
	.w1(32'h3a227ce2),
	.w2(32'hbb249cd9),
	.w3(32'h3c446a88),
	.w4(32'hbb045cc5),
	.w5(32'h3be9bfd0),
	.w6(32'h3c1a926d),
	.w7(32'hb9680fec),
	.w8(32'hb8ce0506),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ffd6),
	.w1(32'hbb550136),
	.w2(32'hbaaee402),
	.w3(32'hbb9d51bb),
	.w4(32'h3b121a8f),
	.w5(32'hbb86d381),
	.w6(32'hbb6eec2d),
	.w7(32'h3bbf79cf),
	.w8(32'h3aa71939),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb03d25),
	.w1(32'h3bd32502),
	.w2(32'h3bd46b01),
	.w3(32'hb9af5020),
	.w4(32'hbb12d5b6),
	.w5(32'h3c9f0835),
	.w6(32'h3b83285c),
	.w7(32'h3b79ecab),
	.w8(32'hbb1b215c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb628b1),
	.w1(32'hb9363154),
	.w2(32'hbbe4c390),
	.w3(32'hbb202136),
	.w4(32'h3b04ac7a),
	.w5(32'hbc5c92e7),
	.w6(32'hbc1b4b19),
	.w7(32'h3b06c072),
	.w8(32'hbb7b7037),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb260013),
	.w1(32'hbb320bdb),
	.w2(32'hbb23162e),
	.w3(32'hbb5a1265),
	.w4(32'h3c004e20),
	.w5(32'h3bfde432),
	.w6(32'hbc20bd6c),
	.w7(32'hbbe16309),
	.w8(32'hbb2e0625),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04237f),
	.w1(32'h3b41f110),
	.w2(32'hb98b6e4b),
	.w3(32'hbc06dde5),
	.w4(32'hbbb3ad33),
	.w5(32'hbbf17e4a),
	.w6(32'hbc368295),
	.w7(32'hbb1fce86),
	.w8(32'h37a677e4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cb5f8),
	.w1(32'h3b48ef46),
	.w2(32'h3ab92f62),
	.w3(32'h3a4b61d0),
	.w4(32'h39569779),
	.w5(32'hba4ac092),
	.w6(32'h3b389b70),
	.w7(32'hbb0c387a),
	.w8(32'h3bb378b3),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f1a528),
	.w1(32'hbb04b3d5),
	.w2(32'h3ab05a7a),
	.w3(32'hb9558a10),
	.w4(32'h3a32e3dd),
	.w5(32'h3a25c913),
	.w6(32'h3be38d0c),
	.w7(32'h3b54b0f8),
	.w8(32'h3a27ff7d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30dace),
	.w1(32'hbb09460e),
	.w2(32'h3ac4b51c),
	.w3(32'hba414aa8),
	.w4(32'hb68c4586),
	.w5(32'h3bd82496),
	.w6(32'hbb0bf1b7),
	.w7(32'hbb9aabb0),
	.w8(32'hbaadbbd1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a67f9),
	.w1(32'hba4afdb2),
	.w2(32'hb9d4f07a),
	.w3(32'hbabdf46b),
	.w4(32'h3bc2a0d0),
	.w5(32'hba9ca959),
	.w6(32'hbb076626),
	.w7(32'hbb3b9888),
	.w8(32'hbb3ba0d2),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b301),
	.w1(32'hb9edfc36),
	.w2(32'hbbd4eab1),
	.w3(32'hbb5518fe),
	.w4(32'h3b6da8b8),
	.w5(32'hbcb8e63d),
	.w6(32'hbc0b9723),
	.w7(32'h3b9b3844),
	.w8(32'h3bb16226),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea682a),
	.w1(32'hba4724ba),
	.w2(32'hbbf5d90e),
	.w3(32'h3b4d9ff2),
	.w4(32'h3b38eb45),
	.w5(32'hb8be9cbf),
	.w6(32'h3c118a6f),
	.w7(32'hba828c89),
	.w8(32'hbb59c4b5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9486c4),
	.w1(32'h3ba97f1f),
	.w2(32'h3c108d4e),
	.w3(32'hbc082fd0),
	.w4(32'h3b1e5f18),
	.w5(32'h3a1bb256),
	.w6(32'hbbb3f870),
	.w7(32'hba818393),
	.w8(32'hbb8da71f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b072d25),
	.w1(32'hbbbc89e5),
	.w2(32'hbbc56545),
	.w3(32'hbb20a038),
	.w4(32'h3baeeb1c),
	.w5(32'h396e9862),
	.w6(32'hbba6248b),
	.w7(32'hbbc1fdaa),
	.w8(32'h3aa92e5d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b1961),
	.w1(32'hbbfc0d64),
	.w2(32'h3b6db302),
	.w3(32'hbbe5cbd0),
	.w4(32'hbbfd8630),
	.w5(32'hbc1d1163),
	.w6(32'h3b050427),
	.w7(32'hbb1845eb),
	.w8(32'h3c4372f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e7937),
	.w1(32'hba657982),
	.w2(32'hbb97e810),
	.w3(32'h3c86be0f),
	.w4(32'h3c61e459),
	.w5(32'h3c02bc68),
	.w6(32'h3c4805df),
	.w7(32'h3c064e86),
	.w8(32'h3c264190),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf710c7),
	.w1(32'hbbf7f123),
	.w2(32'h3b95f3dc),
	.w3(32'h3a6c10d4),
	.w4(32'hbc500cc4),
	.w5(32'h3c901279),
	.w6(32'h3b9f330f),
	.w7(32'hbbad6a10),
	.w8(32'hbb1b70b4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70c85c),
	.w1(32'hb9a388b5),
	.w2(32'hbc1e8d81),
	.w3(32'h3c73d61d),
	.w4(32'h3c298c9e),
	.w5(32'hbbc8732d),
	.w6(32'h3ba1bc38),
	.w7(32'h39d189fe),
	.w8(32'hbb123fcb),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffe27f),
	.w1(32'h398d0589),
	.w2(32'hba979eb4),
	.w3(32'hbc16ce60),
	.w4(32'hbba3223d),
	.w5(32'h3c6f8eb6),
	.w6(32'hbbb55253),
	.w7(32'h3c1dffde),
	.w8(32'h3b80ccf9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34eb69),
	.w1(32'hbc01fddf),
	.w2(32'hba6fa6c2),
	.w3(32'h394afc4d),
	.w4(32'hbbaf2f9b),
	.w5(32'h3a01fff8),
	.w6(32'h39e02e50),
	.w7(32'h3b3cbca9),
	.w8(32'h3b968392),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03267),
	.w1(32'hbc5e16b9),
	.w2(32'hbbb84428),
	.w3(32'hbc159541),
	.w4(32'hbbd6b86a),
	.w5(32'hbba1dae6),
	.w6(32'hbb69480e),
	.w7(32'hbb9e9731),
	.w8(32'hbbc37db6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4131be),
	.w1(32'hbafc66d4),
	.w2(32'hbafcfebe),
	.w3(32'hbc10b5ec),
	.w4(32'hb9efae2e),
	.w5(32'hbb2d846c),
	.w6(32'hbc1c4d8b),
	.w7(32'h3a7e07c9),
	.w8(32'hbc1a0b68),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada4d1e),
	.w1(32'h3664a06c),
	.w2(32'h3b66a356),
	.w3(32'hbc7e2a5f),
	.w4(32'hb9f69079),
	.w5(32'h3b9ec924),
	.w6(32'hbb82bb90),
	.w7(32'hbbf3ae0e),
	.w8(32'h399d5b95),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb580943),
	.w1(32'hbb36e3dc),
	.w2(32'hb91ad858),
	.w3(32'hbbdfa647),
	.w4(32'hbaed24d0),
	.w5(32'h3d1d873e),
	.w6(32'hbbb5d078),
	.w7(32'hbb8fd5b1),
	.w8(32'hbc499ae2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34a4d2),
	.w1(32'hbb648450),
	.w2(32'h3b673afe),
	.w3(32'hbb94fcdf),
	.w4(32'hbb3a0f18),
	.w5(32'hb925ae7c),
	.w6(32'hbb88cabc),
	.w7(32'hb81f20c7),
	.w8(32'hbb4f3a74),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99ff1e),
	.w1(32'h3abf173b),
	.w2(32'h3a0f97f9),
	.w3(32'hbbc53673),
	.w4(32'hbb57b5e5),
	.w5(32'h3b6c2e71),
	.w6(32'hbbd53f04),
	.w7(32'hbbb49027),
	.w8(32'h3a1d049b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba649365),
	.w1(32'hbaff6193),
	.w2(32'h3bcefc11),
	.w3(32'h3bd73de4),
	.w4(32'hbbd15fc0),
	.w5(32'h3c944f0c),
	.w6(32'hb86d9f32),
	.w7(32'hbbc8f60a),
	.w8(32'hbbd2b44c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc34d2d),
	.w1(32'h3a077a83),
	.w2(32'hbbe87fff),
	.w3(32'hbb9110c7),
	.w4(32'hbb2951bc),
	.w5(32'h3c5ab7c7),
	.w6(32'hbb6e8ae2),
	.w7(32'h3be4eead),
	.w8(32'h3ae258aa),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96c335),
	.w1(32'hbb82f4ab),
	.w2(32'hbc0c2eca),
	.w3(32'h3b1b14a3),
	.w4(32'h3b98d925),
	.w5(32'hbb9917c2),
	.w6(32'hbb39db90),
	.w7(32'h3b91301b),
	.w8(32'hba42f671),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb29a41),
	.w1(32'h3b73d08e),
	.w2(32'hbb1aff55),
	.w3(32'hbc1e6ebf),
	.w4(32'h3b0dbb50),
	.w5(32'h3c147144),
	.w6(32'hbb32fc97),
	.w7(32'hbb9fe32c),
	.w8(32'hba944341),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5cd49d),
	.w1(32'h3b2ac5b7),
	.w2(32'hba503a3f),
	.w3(32'h3c98eb05),
	.w4(32'h3bd74fe5),
	.w5(32'hbab0913a),
	.w6(32'h3afc3d9f),
	.w7(32'h3b90ff8e),
	.w8(32'hba843c5c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04f69a),
	.w1(32'hbb864ca6),
	.w2(32'hba73177a),
	.w3(32'h3b7f60d9),
	.w4(32'hbb2d174d),
	.w5(32'hbb635d98),
	.w6(32'h3b8c70e8),
	.w7(32'h3a5e3c70),
	.w8(32'hbacde2db),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b05a58),
	.w1(32'hbaa6f74f),
	.w2(32'h38b01099),
	.w3(32'h3b8b6226),
	.w4(32'h3a081859),
	.w5(32'h3b13111b),
	.w6(32'hbaeea8d2),
	.w7(32'hbaa78098),
	.w8(32'hbaa1ae83),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b41b033),
	.w1(32'h3b5fea9d),
	.w2(32'h3ba12a62),
	.w3(32'hbb155eb2),
	.w4(32'hbb11c523),
	.w5(32'h3b7d207c),
	.w6(32'hbb206735),
	.w7(32'hba58bd71),
	.w8(32'h3bcb80ac),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7541f),
	.w1(32'hbafe4cda),
	.w2(32'h3bf6b019),
	.w3(32'h3bac1db1),
	.w4(32'hbc4693af),
	.w5(32'h3c3d37f0),
	.w6(32'h3b612518),
	.w7(32'hbb29e433),
	.w8(32'h3b88b905),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2bfd5),
	.w1(32'h3a619361),
	.w2(32'hbac6812b),
	.w3(32'h3be24a4a),
	.w4(32'hb7e2c91f),
	.w5(32'hbbcd5ba3),
	.w6(32'hba2baa6b),
	.w7(32'hbb074a1e),
	.w8(32'hbbdee3c6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96d44a),
	.w1(32'hbaee58a6),
	.w2(32'hbbdb826c),
	.w3(32'hbaa59549),
	.w4(32'h3ae40a04),
	.w5(32'h3acbc978),
	.w6(32'hba9f1b2e),
	.w7(32'hbaaa796d),
	.w8(32'hbbd77c39),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad8d4c),
	.w1(32'hbad74786),
	.w2(32'hbad1795a),
	.w3(32'hba4b7081),
	.w4(32'hbc23b4b5),
	.w5(32'hba202465),
	.w6(32'hbb7834ac),
	.w7(32'h3ba0da0d),
	.w8(32'h39cf57f6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae06f58),
	.w1(32'hbb428880),
	.w2(32'h3bd13082),
	.w3(32'h3b38f76f),
	.w4(32'hbc0fc264),
	.w5(32'h3c738d62),
	.w6(32'h3a6f929e),
	.w7(32'hbba51b0a),
	.w8(32'hbb0c2b58),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab268),
	.w1(32'h3a0bdb06),
	.w2(32'hbc0751df),
	.w3(32'hbadc9945),
	.w4(32'hba135181),
	.w5(32'hbbdd92da),
	.w6(32'hb9261d8a),
	.w7(32'h3af8836b),
	.w8(32'hbb4840c2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafed683),
	.w1(32'hbb7dc706),
	.w2(32'hbb789f70),
	.w3(32'hbae5aa33),
	.w4(32'hba80f820),
	.w5(32'h3afb14be),
	.w6(32'hbc3bf24a),
	.w7(32'hbbe94a58),
	.w8(32'hbc09bff1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58008e),
	.w1(32'hb62df2c9),
	.w2(32'hbbd05f80),
	.w3(32'hbba3d8af),
	.w4(32'hbba66d56),
	.w5(32'hba5930d4),
	.w6(32'hbb87e847),
	.w7(32'hbbaa1a04),
	.w8(32'hbc26ee3f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4d92d),
	.w1(32'hbae7f4a9),
	.w2(32'h3b7c7d91),
	.w3(32'h3bfa8b71),
	.w4(32'hbc2136cf),
	.w5(32'h3bf825c9),
	.w6(32'h3aab2178),
	.w7(32'h3a4d4769),
	.w8(32'h3b21c79c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc050cee),
	.w1(32'hbb21f563),
	.w2(32'h3a9872d4),
	.w3(32'hbb05e4fd),
	.w4(32'hbb5d61b7),
	.w5(32'h3aeea262),
	.w6(32'hbb3560af),
	.w7(32'hbb348651),
	.w8(32'hbb1aa01a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3907fc),
	.w1(32'hba5ebcfd),
	.w2(32'h3c0b73f8),
	.w3(32'hba1434e3),
	.w4(32'hbbd0ce55),
	.w5(32'hbbaaddd1),
	.w6(32'h3aa14b88),
	.w7(32'hb9228b6e),
	.w8(32'h3c81da98),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14ab21),
	.w1(32'h3abbc2bb),
	.w2(32'hba9c7fd7),
	.w3(32'h3c6e1b68),
	.w4(32'hbc13e16c),
	.w5(32'hbc2b7a5d),
	.w6(32'h3c7c068e),
	.w7(32'hbc17ca9e),
	.w8(32'hbbfc8d3f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b048b67),
	.w1(32'hbb9bd16e),
	.w2(32'h3ad1f6cc),
	.w3(32'hbbaa3baa),
	.w4(32'hbc038877),
	.w5(32'h3c1e8327),
	.w6(32'hbb991c2a),
	.w7(32'hb90ffddd),
	.w8(32'h3b2e0884),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5475),
	.w1(32'h3b7594a3),
	.w2(32'h3be3722b),
	.w3(32'hbb105f6c),
	.w4(32'hbad3d4a6),
	.w5(32'h3c33aac4),
	.w6(32'hbab2f03c),
	.w7(32'h3a9d22f8),
	.w8(32'h3b730a34),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3a728),
	.w1(32'h3bb53b2b),
	.w2(32'h3b673eca),
	.w3(32'hbb49eb16),
	.w4(32'h3bec87d2),
	.w5(32'h3c3d5ba5),
	.w6(32'hba926d97),
	.w7(32'hbba0a582),
	.w8(32'hba1b7d0d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a5915),
	.w1(32'h3ba7b541),
	.w2(32'h3be88435),
	.w3(32'h3abc9caf),
	.w4(32'hbb915d71),
	.w5(32'h3c89f640),
	.w6(32'hbb7b7f41),
	.w7(32'hbc283b30),
	.w8(32'hba0636c2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8183a53),
	.w1(32'hbb5437f4),
	.w2(32'h3bde3e7a),
	.w3(32'hbb962499),
	.w4(32'hbb4f83b7),
	.w5(32'hbbc26cb4),
	.w6(32'hbb918354),
	.w7(32'h3bec4bed),
	.w8(32'hba96710c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7a96),
	.w1(32'h3a3cf74b),
	.w2(32'h3b3929f5),
	.w3(32'h3b638c0d),
	.w4(32'h3be8c7c4),
	.w5(32'h3bd3b0aa),
	.w6(32'hbb804f88),
	.w7(32'hbbd16848),
	.w8(32'h3b177026),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22619e),
	.w1(32'hbb6104f8),
	.w2(32'h3c21d2a1),
	.w3(32'h3ba15eb7),
	.w4(32'hbb19c145),
	.w5(32'h3ac03510),
	.w6(32'hba233522),
	.w7(32'hbaafd6b8),
	.w8(32'hbb08d26f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb274c39),
	.w1(32'hbbbab7d6),
	.w2(32'hbbb78ca4),
	.w3(32'hbb0f274d),
	.w4(32'h3ab82ea5),
	.w5(32'hbb91ae74),
	.w6(32'hbb99fa7c),
	.w7(32'hbaf6213a),
	.w8(32'hbb8f7780),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901efe4),
	.w1(32'h39b173b5),
	.w2(32'h3b6a226e),
	.w3(32'h3a0358d1),
	.w4(32'hb9817842),
	.w5(32'h3c47dbc3),
	.w6(32'h3b94dcdb),
	.w7(32'h3a3559ec),
	.w8(32'h3b3b345e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba906158),
	.w1(32'hbb028687),
	.w2(32'hbc22cf4d),
	.w3(32'h3c11946d),
	.w4(32'h3ba2db21),
	.w5(32'hbc589770),
	.w6(32'hb9901c36),
	.w7(32'hbad99371),
	.w8(32'h3abcf229),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb85c4),
	.w1(32'hbbf9e6ce),
	.w2(32'hbc07052d),
	.w3(32'hbba96950),
	.w4(32'hbb9e8c62),
	.w5(32'hbb96050c),
	.w6(32'hbbe9e12e),
	.w7(32'hbc373fe4),
	.w8(32'hbc3c485e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe294e),
	.w1(32'hb97a51cd),
	.w2(32'hbc26b110),
	.w3(32'hbb206e47),
	.w4(32'hbb08d40c),
	.w5(32'hbc683ddc),
	.w6(32'hbb154527),
	.w7(32'hbab8a024),
	.w8(32'hbc17d6af),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7183d),
	.w1(32'hbb58dea1),
	.w2(32'h3b446c32),
	.w3(32'hbb470e9b),
	.w4(32'hbbb33601),
	.w5(32'h3b92c637),
	.w6(32'h3a228db0),
	.w7(32'h3b9059b9),
	.w8(32'hbb128c3a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3de05e),
	.w1(32'hbb5f6c6d),
	.w2(32'h3ac499e2),
	.w3(32'hbc9d4557),
	.w4(32'hbbfbe5b1),
	.w5(32'hbb071ead),
	.w6(32'hbbf31deb),
	.w7(32'hbc13d442),
	.w8(32'hbb91c511),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3187b2),
	.w1(32'h3a5ad238),
	.w2(32'hbb3b8c98),
	.w3(32'h39985607),
	.w4(32'h3b30d8ce),
	.w5(32'h3a12c490),
	.w6(32'hbb065f9f),
	.w7(32'h3b5979ae),
	.w8(32'hb9ae62ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc7fff),
	.w1(32'hbb9ccd31),
	.w2(32'h3bb15045),
	.w3(32'hbb1e3975),
	.w4(32'hbc15ce3d),
	.w5(32'h3cd1d186),
	.w6(32'h3af771a9),
	.w7(32'hbb8d52cc),
	.w8(32'hbb9797e3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8381f2),
	.w1(32'h3b84f895),
	.w2(32'hbbebb063),
	.w3(32'h3bc37ebf),
	.w4(32'h3bc22ec4),
	.w5(32'hbcaec78d),
	.w6(32'hbb90a661),
	.w7(32'h3b22ff7b),
	.w8(32'h3bd58df9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc34957),
	.w1(32'h3a971eb3),
	.w2(32'hb85436eb),
	.w3(32'h3bc9a1a0),
	.w4(32'h3b050d82),
	.w5(32'h38943e15),
	.w6(32'h3c3fe30b),
	.w7(32'h3c212479),
	.w8(32'h3c18a9a3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11f401),
	.w1(32'h3b7f5910),
	.w2(32'hbabaf214),
	.w3(32'h3a8b271b),
	.w4(32'hbaf9f963),
	.w5(32'hbb124ef2),
	.w6(32'h3a880db2),
	.w7(32'hba1b3d4d),
	.w8(32'h3a167aa8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf060e),
	.w1(32'hb9aed908),
	.w2(32'h3a0bb62b),
	.w3(32'h3b546c4e),
	.w4(32'h39949a84),
	.w5(32'h3b60d6f6),
	.w6(32'h3a82d21e),
	.w7(32'hbbe4388f),
	.w8(32'hba922ff2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30b5d),
	.w1(32'h3c3ad3fc),
	.w2(32'h3c8f373f),
	.w3(32'hbc05afe9),
	.w4(32'h3b894878),
	.w5(32'h3ce7dcbc),
	.w6(32'hbb904d1f),
	.w7(32'h3b5b0893),
	.w8(32'h3bcf485e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63f8bc),
	.w1(32'h3a207a00),
	.w2(32'h3b97f2cb),
	.w3(32'h38810a4c),
	.w4(32'hbc146748),
	.w5(32'h3c1e8340),
	.w6(32'h3c543e5c),
	.w7(32'h3a832096),
	.w8(32'h38ed8f6e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81229f),
	.w1(32'hb954f3c4),
	.w2(32'hb8a9f49a),
	.w3(32'hba0f192f),
	.w4(32'hb91ceaf7),
	.w5(32'hb7811ae8),
	.w6(32'h3a3e192c),
	.w7(32'h377dd098),
	.w8(32'h398792b6),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36827414),
	.w1(32'hb61af22a),
	.w2(32'hb587f4af),
	.w3(32'h367dd78e),
	.w4(32'h360bd495),
	.w5(32'hb6f30c7a),
	.w6(32'hb62ea57f),
	.w7(32'h36dd8361),
	.w8(32'hb5c1aea6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79015be),
	.w1(32'h37134d73),
	.w2(32'h35dbb2b1),
	.w3(32'hb7839239),
	.w4(32'hb73ab5a4),
	.w5(32'hb6b58520),
	.w6(32'hb72058a3),
	.w7(32'hb7884e52),
	.w8(32'hb6f79fb5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3717328e),
	.w1(32'h3603ec56),
	.w2(32'h3680ca86),
	.w3(32'h3647b1e4),
	.w4(32'h36d9f545),
	.w5(32'h36b46594),
	.w6(32'hb764ec82),
	.w7(32'h360d3356),
	.w8(32'h3477fe0d),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881cd48),
	.w1(32'h3822753e),
	.w2(32'h3802a52e),
	.w3(32'h379837a5),
	.w4(32'hb78a4de6),
	.w5(32'hb5874e8e),
	.w6(32'h3706cf94),
	.w7(32'hb87f5568),
	.w8(32'hb84859dd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8690f02),
	.w1(32'hb81b408d),
	.w2(32'hb7067735),
	.w3(32'hb7984b36),
	.w4(32'hb771bcc4),
	.w5(32'hb52ab921),
	.w6(32'hb75cf413),
	.w7(32'h36f19c03),
	.w8(32'h36c52d8d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38015855),
	.w1(32'h37cc1cfe),
	.w2(32'hb71331e1),
	.w3(32'h389364ae),
	.w4(32'h38de8624),
	.w5(32'h38ae0cad),
	.w6(32'h38cba1bf),
	.w7(32'hb79ca4b4),
	.w8(32'hb8f5b7b7),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e0cc8),
	.w1(32'h396088dc),
	.w2(32'h387fdd55),
	.w3(32'h3945c212),
	.w4(32'h381b9460),
	.w5(32'h38f6a8cd),
	.w6(32'h3985320e),
	.w7(32'h38b0024d),
	.w8(32'hb89d77a0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848181c),
	.w1(32'hb7eceeb0),
	.w2(32'h39004248),
	.w3(32'h37f7ac81),
	.w4(32'h37f80651),
	.w5(32'h3939e050),
	.w6(32'h385e4aa2),
	.w7(32'h37f86970),
	.w8(32'h38f89dd7),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e92844),
	.w1(32'h3880b5f5),
	.w2(32'h38c05cad),
	.w3(32'h391f8914),
	.w4(32'h38aff511),
	.w5(32'h3822c6f0),
	.w6(32'h3912fafa),
	.w7(32'hb81ad7e0),
	.w8(32'h36ec2042),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c6ee25),
	.w1(32'h3874ed2a),
	.w2(32'h3819ea98),
	.w3(32'h38c69636),
	.w4(32'h395284af),
	.w5(32'h38fe4c6c),
	.w6(32'h39526a78),
	.w7(32'hb75b6482),
	.w8(32'hb8aefffa),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cce33f),
	.w1(32'hb825a151),
	.w2(32'h381ec694),
	.w3(32'h38e755aa),
	.w4(32'h37ccbfd6),
	.w5(32'h3889f618),
	.w6(32'h392593a9),
	.w7(32'h3879835b),
	.w8(32'h38f6d78c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a0f1ca),
	.w1(32'h37280676),
	.w2(32'h388efd49),
	.w3(32'h3830db76),
	.w4(32'h3846a0c2),
	.w5(32'h389a7e0a),
	.w6(32'h38520d7a),
	.w7(32'hb7dd3945),
	.w8(32'hb87852f1),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f78084),
	.w1(32'hb592ec47),
	.w2(32'hb6a4ed6d),
	.w3(32'hb6f800bb),
	.w4(32'h36578087),
	.w5(32'hb6919358),
	.w6(32'hb6832260),
	.w7(32'h36950277),
	.w8(32'h35e394ca),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ec9aa0),
	.w1(32'hb79e2656),
	.w2(32'h36982d6f),
	.w3(32'hb696def1),
	.w4(32'hb6888f29),
	.w5(32'h3712158d),
	.w6(32'h36d8f035),
	.w7(32'h368c90c8),
	.w8(32'h360c21bd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb706e48c),
	.w1(32'h37325cf3),
	.w2(32'h37761bf0),
	.w3(32'hb74dccf6),
	.w4(32'h37067585),
	.w5(32'h3760e78d),
	.w6(32'hb6f7aa6e),
	.w7(32'h360e79ec),
	.w8(32'h36a8b04d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364854bd),
	.w1(32'hb7632b81),
	.w2(32'hb47bbfe4),
	.w3(32'hb7a8116a),
	.w4(32'hb79bb365),
	.w5(32'hb645093b),
	.w6(32'hb75b696a),
	.w7(32'hb6cb4cdd),
	.w8(32'hb53ec253),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b048d),
	.w1(32'hb7eb377e),
	.w2(32'hb88c3ee7),
	.w3(32'h39038606),
	.w4(32'h371b6625),
	.w5(32'h38a79d8f),
	.w6(32'h37a433e5),
	.w7(32'h37fea1b4),
	.w8(32'h3822556e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3518c568),
	.w1(32'hb7e88594),
	.w2(32'hb6880e57),
	.w3(32'h374fdf6f),
	.w4(32'hb7b9c2c0),
	.w5(32'hb768ae31),
	.w6(32'h37084d01),
	.w7(32'h371b53f9),
	.w8(32'h37d9a97e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f26c7),
	.w1(32'h3920d2a9),
	.w2(32'h395773ba),
	.w3(32'h39600b38),
	.w4(32'h38bc306f),
	.w5(32'h38ff3125),
	.w6(32'h39549472),
	.w7(32'h39361ea9),
	.w8(32'h39803d7e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da621b),
	.w1(32'h3851aa1f),
	.w2(32'h37e62168),
	.w3(32'h38f559da),
	.w4(32'h37ec7977),
	.w5(32'hb78c3d2a),
	.w6(32'h391044e7),
	.w7(32'hb8417f00),
	.w8(32'hb913d147),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e116e9),
	.w1(32'hb9135ee4),
	.w2(32'hb891aa8b),
	.w3(32'hb8b0436f),
	.w4(32'hb93e91ae),
	.w5(32'hb7e3f91b),
	.w6(32'hb88485d0),
	.w7(32'hb8f9f14d),
	.w8(32'h381590dd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993572f),
	.w1(32'h3907439b),
	.w2(32'h389496c3),
	.w3(32'h39d8da39),
	.w4(32'h39ce62ff),
	.w5(32'h38ae4c01),
	.w6(32'h39ceb27c),
	.w7(32'h39237746),
	.w8(32'hb8769c5c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38355524),
	.w1(32'hb811314e),
	.w2(32'hb8575838),
	.w3(32'hb8a1375c),
	.w4(32'hb89d2e60),
	.w5(32'hb8acfa2c),
	.w6(32'hb85ea80e),
	.w7(32'hb8d9034f),
	.w8(32'hb8948a54),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dc020),
	.w1(32'h38a0b915),
	.w2(32'h38a43f16),
	.w3(32'h39fb8ec6),
	.w4(32'h393e1eea),
	.w5(32'h37fd7618),
	.w6(32'h39c82a22),
	.w7(32'hb876a826),
	.w8(32'hb86b50dc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2c6ec),
	.w1(32'h37b16e73),
	.w2(32'h3721c694),
	.w3(32'h3921257b),
	.w4(32'h391bc48d),
	.w5(32'h385e374d),
	.w6(32'h391d98f0),
	.w7(32'h38d8182f),
	.w8(32'h39078efe),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be8a63),
	.w1(32'h36a6cacf),
	.w2(32'h383095d4),
	.w3(32'h37f41207),
	.w4(32'h37f6b3c6),
	.w5(32'h381bfa4d),
	.w6(32'h38dcbe74),
	.w7(32'h3864646e),
	.w8(32'h3909ebfd),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ff21fa),
	.w1(32'hb8b5c345),
	.w2(32'hb90082d3),
	.w3(32'hb80198ef),
	.w4(32'hb8b365d9),
	.w5(32'hb8d5bf3f),
	.w6(32'hb81b4476),
	.w7(32'hb8e9cfac),
	.w8(32'hb8516850),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3738e407),
	.w1(32'hb8bc7c6d),
	.w2(32'h38450aaf),
	.w3(32'h3916e2bf),
	.w4(32'h37c416bc),
	.w5(32'hb8b66547),
	.w6(32'h394b0b24),
	.w7(32'hb7eed5cd),
	.w8(32'hb7aa6849),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8465c),
	.w1(32'hb8f53f7b),
	.w2(32'hb8ec1dda),
	.w3(32'hb7ca0abb),
	.w4(32'h39410833),
	.w5(32'h392a5971),
	.w6(32'h3980120d),
	.w7(32'h38af1b96),
	.w8(32'hb72a12ac),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37947be0),
	.w1(32'h39b045be),
	.w2(32'h3990c1a8),
	.w3(32'h399ec523),
	.w4(32'h389fd660),
	.w5(32'h3839f37a),
	.w6(32'h3982af36),
	.w7(32'h39a49f63),
	.w8(32'hb8d22379),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3701e650),
	.w1(32'hb9b75413),
	.w2(32'hb9834f5b),
	.w3(32'hb8aa4e4b),
	.w4(32'hb94a63da),
	.w5(32'hb72b8140),
	.w6(32'h391988bf),
	.w7(32'h38c3725b),
	.w8(32'h37e49887),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3753855f),
	.w1(32'h38b54698),
	.w2(32'h393b8438),
	.w3(32'h38e4cdf2),
	.w4(32'h393e3a04),
	.w5(32'h3922c421),
	.w6(32'h39183f68),
	.w7(32'h394a7c77),
	.w8(32'h39bad2f3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383b77c2),
	.w1(32'h39073338),
	.w2(32'h38641e39),
	.w3(32'h3943ae10),
	.w4(32'h39c105d5),
	.w5(32'h389c6adc),
	.w6(32'h39e01c1c),
	.w7(32'h39b92dc9),
	.w8(32'hb8d5f662),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb811fa63),
	.w1(32'hb92c38a8),
	.w2(32'hb97d5498),
	.w3(32'h37340ef9),
	.w4(32'hb854e164),
	.w5(32'hb9027345),
	.w6(32'h38ff95ef),
	.w7(32'h384b2047),
	.w8(32'hb877bfcb),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a69298),
	.w1(32'h396a6a82),
	.w2(32'h394b06f2),
	.w3(32'h39c5b053),
	.w4(32'h395530b3),
	.w5(32'h39ae742e),
	.w6(32'h3a241ff5),
	.w7(32'h3a0f179c),
	.w8(32'h37321e07),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914a1ae),
	.w1(32'hb8ab0d0a),
	.w2(32'h37933bd5),
	.w3(32'h37eb1132),
	.w4(32'hb89a846e),
	.w5(32'hb7054616),
	.w6(32'h38c26899),
	.w7(32'hb76d9dc0),
	.w8(32'hb7762474),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379e9105),
	.w1(32'h372c5906),
	.w2(32'h372b02c3),
	.w3(32'h371b1792),
	.w4(32'hb53cb460),
	.w5(32'hb5efb9a1),
	.w6(32'h374d3cb8),
	.w7(32'h36149081),
	.w8(32'hb5d9d21d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389880dd),
	.w1(32'h38ad7f55),
	.w2(32'h386bada1),
	.w3(32'h38084462),
	.w4(32'h38d6ea6f),
	.w5(32'h382a57d8),
	.w6(32'h37b5395c),
	.w7(32'h37cdb007),
	.w8(32'h3833d2ce),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aeb449),
	.w1(32'hb90ca184),
	.w2(32'h3720d8ab),
	.w3(32'h38745d4a),
	.w4(32'hb79c77bb),
	.w5(32'h37f45312),
	.w6(32'h392405ae),
	.w7(32'hb68614be),
	.w8(32'hb81f40dc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c764f),
	.w1(32'hb94a6247),
	.w2(32'hb75998be),
	.w3(32'hb89f2bd7),
	.w4(32'hb858a117),
	.w5(32'hb8937959),
	.w6(32'h36fa8dab),
	.w7(32'hb7b9bbf7),
	.w8(32'h385a2b61),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65fa396),
	.w1(32'hb913c735),
	.w2(32'hb8782b61),
	.w3(32'hb810c286),
	.w4(32'hb787ca09),
	.w5(32'h3874d1ff),
	.w6(32'h382a880c),
	.w7(32'hb880dbca),
	.w8(32'h372391a0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364c3b5e),
	.w1(32'hb7a31a79),
	.w2(32'h382ffb68),
	.w3(32'h3885ce66),
	.w4(32'h37b49328),
	.w5(32'h38a10c69),
	.w6(32'h386e3668),
	.w7(32'h38fa3e7b),
	.w8(32'h39026b56),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a76156),
	.w1(32'h393ddb7a),
	.w2(32'h38c56270),
	.w3(32'h3999a9e0),
	.w4(32'h37dd58dc),
	.w5(32'hb78439f0),
	.w6(32'h39486d03),
	.w7(32'h388a545a),
	.w8(32'h376aa2c5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393aaa3f),
	.w1(32'h38e342e6),
	.w2(32'h394a388d),
	.w3(32'h396b0dba),
	.w4(32'h3987c9fc),
	.w5(32'h393b46d9),
	.w6(32'h3928628e),
	.w7(32'hb89be1f1),
	.w8(32'hb80ec3cc),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36aeb2fa),
	.w1(32'hb82762ea),
	.w2(32'h389942e3),
	.w3(32'h3857b128),
	.w4(32'hb7df5215),
	.w5(32'h386146bb),
	.w6(32'h3883e698),
	.w7(32'h38231708),
	.w8(32'h38d0beca),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a9a374),
	.w1(32'hb6499c9b),
	.w2(32'hb4f5e0a8),
	.w3(32'h36d4b31b),
	.w4(32'h363e4bd8),
	.w5(32'hb671c76c),
	.w6(32'h36b71d3b),
	.w7(32'hb56e469e),
	.w8(32'hb54cebba),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3808af86),
	.w1(32'h3705ccc7),
	.w2(32'h37cfd977),
	.w3(32'h37b842fd),
	.w4(32'h352614fb),
	.w5(32'h37422868),
	.w6(32'hb7122edd),
	.w7(32'hb7ac9bbc),
	.w8(32'hb6977fdb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6eb6251),
	.w1(32'h368431f1),
	.w2(32'h3736fa52),
	.w3(32'hb70315cc),
	.w4(32'hb5c1daa5),
	.w5(32'h36830041),
	.w6(32'hb72258f9),
	.w7(32'hb5aebc47),
	.w8(32'h3566dabf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a19d85),
	.w1(32'h36b25bef),
	.w2(32'hb7ea0bca),
	.w3(32'h37ec51ce),
	.w4(32'h373c97a5),
	.w5(32'hb5f13b33),
	.w6(32'h36c0b690),
	.w7(32'h3699ca13),
	.w8(32'hb58825ba),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38089bc4),
	.w1(32'hb5bf86c9),
	.w2(32'h388bd721),
	.w3(32'h38cd6552),
	.w4(32'h37bd0cba),
	.w5(32'h381353e6),
	.w6(32'h3921c670),
	.w7(32'h38ff3c24),
	.w8(32'h390f3a1e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f0b9c5),
	.w1(32'h372c158e),
	.w2(32'hb66da75a),
	.w3(32'h377636b7),
	.w4(32'h362486fe),
	.w5(32'hb70fba74),
	.w6(32'h37144120),
	.w7(32'hb72f8e82),
	.w8(32'hb74bb927),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350717b1),
	.w1(32'h37ca9783),
	.w2(32'h360643f5),
	.w3(32'h37576bf2),
	.w4(32'h38934da0),
	.w5(32'h367018e6),
	.w6(32'h3873eb31),
	.w7(32'h3795ba84),
	.w8(32'hb8ed881d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3838fe13),
	.w1(32'hb8c96143),
	.w2(32'h36c71107),
	.w3(32'h381c126c),
	.w4(32'hb811b0b4),
	.w5(32'h3800973b),
	.w6(32'h382d3236),
	.w7(32'hb82fce77),
	.w8(32'h38db7563),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb781475e),
	.w1(32'h3722f286),
	.w2(32'hb5c170af),
	.w3(32'hb7a25b3e),
	.w4(32'h3702e2b2),
	.w5(32'hb6ae28d8),
	.w6(32'hb598bace),
	.w7(32'h371533c6),
	.w8(32'hb69c22c6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb712b67d),
	.w1(32'h36bae5f3),
	.w2(32'hb6db053e),
	.w3(32'hb79bde47),
	.w4(32'hb7ad3f84),
	.w5(32'hb783e509),
	.w6(32'hb6eaeee8),
	.w7(32'hb7b26d06),
	.w8(32'hb73e1720),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374967f2),
	.w1(32'h36f42ce5),
	.w2(32'h3731ab9f),
	.w3(32'h365d6ad8),
	.w4(32'h34886e5c),
	.w5(32'h36903fe8),
	.w6(32'hb73969d5),
	.w7(32'h34174479),
	.w8(32'h36d98f48),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ccb1cc),
	.w1(32'h36814e09),
	.w2(32'h37f8ffe2),
	.w3(32'h37a19ea7),
	.w4(32'h36c1ae57),
	.w5(32'h3707c87b),
	.w6(32'h37b9a613),
	.w7(32'h37814792),
	.w8(32'h37cd1861),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39890dbb),
	.w1(32'h39f09c3d),
	.w2(32'h391bf2c0),
	.w3(32'h395e368d),
	.w4(32'h36adbb80),
	.w5(32'hb92792d1),
	.w6(32'h397baa7f),
	.w7(32'h392b1a94),
	.w8(32'hb92be20c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38becd32),
	.w1(32'h3903a634),
	.w2(32'h39391fb6),
	.w3(32'h391e9637),
	.w4(32'h38be28de),
	.w5(32'h388924df),
	.w6(32'h3982393f),
	.w7(32'hb755c1ba),
	.w8(32'hb70b2ff3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ba6546),
	.w1(32'hb6c52d8e),
	.w2(32'h3785b24b),
	.w3(32'h3822ba57),
	.w4(32'h36fe421e),
	.w5(32'h37c0c9f5),
	.w6(32'h37db8887),
	.w7(32'hb7a15e40),
	.w8(32'hb777034c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4d939),
	.w1(32'h38346962),
	.w2(32'h37de5a2d),
	.w3(32'h388ba742),
	.w4(32'hb84da7dd),
	.w5(32'hb745d4e9),
	.w6(32'h388854ef),
	.w7(32'hb76a4ea5),
	.w8(32'hb7a0c389),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e4045e),
	.w1(32'hb80e6d72),
	.w2(32'hb65d3ce9),
	.w3(32'h366b0794),
	.w4(32'hb779545e),
	.w5(32'h378d1167),
	.w6(32'hb73513af),
	.w7(32'hb797f143),
	.w8(32'h37810fad),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb632ddee),
	.w1(32'h374bf90b),
	.w2(32'h383c6900),
	.w3(32'h38a6a167),
	.w4(32'h3772863d),
	.w5(32'hb624e886),
	.w6(32'h38d891a7),
	.w7(32'hb7d078d7),
	.w8(32'h37d58764),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fe5273),
	.w1(32'h38910afd),
	.w2(32'h391e1cf4),
	.w3(32'h38a39dff),
	.w4(32'h38e70169),
	.w5(32'h391bec77),
	.w6(32'h38ef8f50),
	.w7(32'h374d0e7d),
	.w8(32'h385e190c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c81b10),
	.w1(32'h3818e7ec),
	.w2(32'h3891a0df),
	.w3(32'h390c24a5),
	.w4(32'h38d916eb),
	.w5(32'h37a53f42),
	.w6(32'h398f5f7d),
	.w7(32'hb8871d8f),
	.w8(32'hb8f483c2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383132a9),
	.w1(32'h367d229c),
	.w2(32'h3834cf4d),
	.w3(32'h38ce540d),
	.w4(32'h38541c51),
	.w5(32'h38ca36f2),
	.w6(32'h3894ff18),
	.w7(32'h387659a2),
	.w8(32'h3904c814),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9569b),
	.w1(32'h37e4bf9e),
	.w2(32'h388fcc1d),
	.w3(32'h39225d00),
	.w4(32'h393b48e5),
	.w5(32'h3916debb),
	.w6(32'h391be9c8),
	.w7(32'h374fcae1),
	.w8(32'hb83725aa),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3922b4a2),
	.w1(32'h392a3b3b),
	.w2(32'h38afdfa2),
	.w3(32'h3978460a),
	.w4(32'h395dd87f),
	.w5(32'h38a737d6),
	.w6(32'h3989e1b8),
	.w7(32'h392694d9),
	.w8(32'hb868b56d),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe5efe),
	.w1(32'h384c804b),
	.w2(32'h3910cf30),
	.w3(32'h3916f8cf),
	.w4(32'h375aafb1),
	.w5(32'h387f0924),
	.w6(32'h38a9b35a),
	.w7(32'h37f19aca),
	.w8(32'h38a41159),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39566052),
	.w1(32'h38957448),
	.w2(32'h38c10e23),
	.w3(32'h39923ccc),
	.w4(32'h3944cb6e),
	.w5(32'h3896d8c4),
	.w6(32'h39a0b53e),
	.w7(32'h3909b968),
	.w8(32'h374721a9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fbc787),
	.w1(32'hb69c0df3),
	.w2(32'h383f843f),
	.w3(32'h377907a1),
	.w4(32'hb6d7b1f4),
	.w5(32'h37dc51b7),
	.w6(32'h381a9aa5),
	.w7(32'h368d9bcd),
	.w8(32'h37dcc2e6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377e8dde),
	.w1(32'hb79c71bf),
	.w2(32'h38c61274),
	.w3(32'h38ba27b6),
	.w4(32'h389726c4),
	.w5(32'h392e9c3d),
	.w6(32'h3942015c),
	.w7(32'h394d31ac),
	.w8(32'h398ef114),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bcf603),
	.w1(32'h382c0988),
	.w2(32'hb7dabc87),
	.w3(32'h38e3635a),
	.w4(32'h381811ad),
	.w5(32'hb79e08b1),
	.w6(32'h38b5a2f9),
	.w7(32'h37c090fb),
	.w8(32'h381318de),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ce9a50),
	.w1(32'h3716e1c3),
	.w2(32'h3638d8a9),
	.w3(32'h35e01c69),
	.w4(32'h3765e3a0),
	.w5(32'hb629f679),
	.w6(32'hb5fccd8a),
	.w7(32'h371b537e),
	.w8(32'h339feb79),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76da4db),
	.w1(32'h36ba36ed),
	.w2(32'h371084d3),
	.w3(32'hb6e316ed),
	.w4(32'h367bbd9d),
	.w5(32'h36b3ab18),
	.w6(32'hb6d66e40),
	.w7(32'hb70a97c8),
	.w8(32'h34dd173c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f1557),
	.w1(32'hb8189920),
	.w2(32'hb8060c13),
	.w3(32'h37caa7f6),
	.w4(32'hb6853395),
	.w5(32'hb40b1ea7),
	.w6(32'h37e93ce4),
	.w7(32'hb692c38b),
	.w8(32'hb79bef29),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e67bf3),
	.w1(32'hb6071f98),
	.w2(32'hb81da6bb),
	.w3(32'h38df0ad1),
	.w4(32'h385f3e7c),
	.w5(32'h389a6ab5),
	.w6(32'h379163bf),
	.w7(32'h38464048),
	.w8(32'h38bd08c0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f96564),
	.w1(32'h3839fb97),
	.w2(32'h38c403b4),
	.w3(32'h387c266d),
	.w4(32'h36b57bb6),
	.w5(32'h38a8c3fe),
	.w6(32'h362936d8),
	.w7(32'hb8ba0a98),
	.w8(32'hb8b6a3b9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6db5e1b),
	.w1(32'hb7384869),
	.w2(32'h36500d4f),
	.w3(32'hb705e999),
	.w4(32'hb670269c),
	.w5(32'h36c2f8e3),
	.w6(32'h36b08500),
	.w7(32'hb5918234),
	.w8(32'h369c56c5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379379d2),
	.w1(32'h366dab7d),
	.w2(32'h38caab1e),
	.w3(32'h391a4af4),
	.w4(32'h38f34c01),
	.w5(32'h38e54667),
	.w6(32'h395bd233),
	.w7(32'hb6ec0327),
	.w8(32'h3804a32f),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384c69a1),
	.w1(32'hb64b3cb9),
	.w2(32'hb691ea8c),
	.w3(32'h393053ab),
	.w4(32'h37b05f44),
	.w5(32'h38229a67),
	.w6(32'h392e7830),
	.w7(32'h39220135),
	.w8(32'h39260182),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886a8c0),
	.w1(32'h392b5713),
	.w2(32'h39271380),
	.w3(32'h3906ed20),
	.w4(32'h398d1b97),
	.w5(32'h394fcf5f),
	.w6(32'h3968f0c7),
	.w7(32'h388bbbc2),
	.w8(32'hb8874581),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8839b81),
	.w1(32'hb931f578),
	.w2(32'h38a3b486),
	.w3(32'h38f4dc52),
	.w4(32'hb70da42a),
	.w5(32'h39437b58),
	.w6(32'h392bfdb2),
	.w7(32'h37f3a4d9),
	.w8(32'h399456e3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38096800),
	.w1(32'hb70d8836),
	.w2(32'hb8b2dae9),
	.w3(32'h382b253c),
	.w4(32'h3717f9d3),
	.w5(32'hb93086f1),
	.w6(32'hb72ff432),
	.w7(32'hb88454e1),
	.w8(32'hb9001069),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88570b7),
	.w1(32'hb96b4282),
	.w2(32'hb91bfe7f),
	.w3(32'h375fe19f),
	.w4(32'h387b2ca3),
	.w5(32'hb8a3f339),
	.w6(32'h38d6c14b),
	.w7(32'h390fdc45),
	.w8(32'h36379c96),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882a245),
	.w1(32'hb9019c42),
	.w2(32'hb8998425),
	.w3(32'h37cfa586),
	.w4(32'hb6b5084f),
	.w5(32'h38a4744b),
	.w6(32'h38b968c3),
	.w7(32'h39049b6f),
	.w8(32'h3917da34),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f09e90),
	.w1(32'hb896d7cb),
	.w2(32'hb8d1fdde),
	.w3(32'hb7e125ed),
	.w4(32'hb8c53f7b),
	.w5(32'hb8699d9e),
	.w6(32'hb8c94d63),
	.w7(32'hb9071a33),
	.w8(32'hb794bb17),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3600f084),
	.w1(32'hb8b21fe0),
	.w2(32'hb80ee500),
	.w3(32'hb7e3a11a),
	.w4(32'hb8997d71),
	.w5(32'h3689f842),
	.w6(32'hb86c22ba),
	.w7(32'hb8af6ad3),
	.w8(32'h380e29a7),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3708d09a),
	.w1(32'h37713f2a),
	.w2(32'h34d161af),
	.w3(32'h379c445e),
	.w4(32'h37b5260f),
	.w5(32'h3707d474),
	.w6(32'h37db784f),
	.w7(32'h376aa93b),
	.w8(32'hb800c592),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h348467f9),
	.w1(32'h36fd3d2b),
	.w2(32'h3613c147),
	.w3(32'hb697070f),
	.w4(32'h36dfbaac),
	.w5(32'h358f6f9a),
	.w6(32'h36b9d57c),
	.w7(32'h3639281f),
	.w8(32'hb6804e05),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38da4500),
	.w1(32'h3884ced9),
	.w2(32'h38a74e4d),
	.w3(32'h39277f85),
	.w4(32'h38e65192),
	.w5(32'h38966818),
	.w6(32'h39599bb5),
	.w7(32'h389aecca),
	.w8(32'hb6135abd),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70b5572),
	.w1(32'h3665acd1),
	.w2(32'hb7d06dd7),
	.w3(32'hb7b78f17),
	.w4(32'h374c7864),
	.w5(32'hb6f3bd30),
	.w6(32'h37c693ec),
	.w7(32'h3745f62b),
	.w8(32'hb7d470ff),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b9ba87),
	.w1(32'hb709ebb5),
	.w2(32'h38a2c1fe),
	.w3(32'h391d33e8),
	.w4(32'h389be4ad),
	.w5(32'h38d7a280),
	.w6(32'h393d3b99),
	.w7(32'h390a3bdd),
	.w8(32'h3940e830),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ff598),
	.w1(32'hb7c1785a),
	.w2(32'h3646e6d3),
	.w3(32'hb7f86705),
	.w4(32'h36fe3a0a),
	.w5(32'h378f1f86),
	.w6(32'hb7ae9ea4),
	.w7(32'hb776bf6b),
	.w8(32'h361733c2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37564485),
	.w1(32'hb78f661a),
	.w2(32'hb844e0d8),
	.w3(32'hb7e840e2),
	.w4(32'hb91bfde4),
	.w5(32'hb8be918a),
	.w6(32'hb81bc583),
	.w7(32'hb94bc59d),
	.w8(32'hb961ea34),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377d16b4),
	.w1(32'hb7811977),
	.w2(32'h36c86618),
	.w3(32'h3751b4bf),
	.w4(32'hb7cc3170),
	.w5(32'hb67b2c3a),
	.w6(32'h377bba38),
	.w7(32'hb7bc6a16),
	.w8(32'hb78f024e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3520fb9b),
	.w1(32'hb73d9c10),
	.w2(32'hb6c789b1),
	.w3(32'h378bbfd9),
	.w4(32'h3688fe51),
	.w5(32'hb788a047),
	.w6(32'h37ec76d5),
	.w7(32'h382ab6a9),
	.w8(32'hb73c8185),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f68d5),
	.w1(32'hb7ac8d20),
	.w2(32'hb7395543),
	.w3(32'h390f8383),
	.w4(32'h38432050),
	.w5(32'h375104f6),
	.w6(32'h38aac759),
	.w7(32'h38f4c27d),
	.w8(32'h3887ae05),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7b0ff),
	.w1(32'h3956afe7),
	.w2(32'h38e37e68),
	.w3(32'h3957d395),
	.w4(32'h3938aba6),
	.w5(32'h382d5c24),
	.w6(32'h39b8ceb8),
	.w7(32'h39c4f2a7),
	.w8(32'h391347d7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389af439),
	.w1(32'hb75329b6),
	.w2(32'hb716f1bd),
	.w3(32'hb7485b56),
	.w4(32'hb88ba6bb),
	.w5(32'hb84a895a),
	.w6(32'h37803524),
	.w7(32'hb8050e99),
	.w8(32'hb8021258),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7bb77),
	.w1(32'h3864e269),
	.w2(32'h39160b7c),
	.w3(32'h38e94583),
	.w4(32'h371e8b83),
	.w5(32'h38f4b3ee),
	.w6(32'h396d6f9e),
	.w7(32'h392a57f8),
	.w8(32'h3954a5be),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d66e58),
	.w1(32'hb78ecf70),
	.w2(32'h37e213d0),
	.w3(32'hb79e2d39),
	.w4(32'hb8196b0e),
	.w5(32'h37ddfdd8),
	.w6(32'hb79987cd),
	.w7(32'hb82d6db1),
	.w8(32'h37c35e13),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9c17e),
	.w1(32'h36aaa7b9),
	.w2(32'h38d9a26e),
	.w3(32'h3945a007),
	.w4(32'h38146e91),
	.w5(32'h3907f841),
	.w6(32'h38f14cfd),
	.w7(32'hb9493045),
	.w8(32'hb857e715),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3824eaa4),
	.w1(32'hb82ceb09),
	.w2(32'hb87b2d39),
	.w3(32'h38f2e141),
	.w4(32'hb6bd1090),
	.w5(32'h37a421fc),
	.w6(32'h39276b7f),
	.w7(32'hb82c389a),
	.w8(32'h37cbd5b6),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38488205),
	.w1(32'h388d5b74),
	.w2(32'h38b88149),
	.w3(32'h3935c0b4),
	.w4(32'h390d0281),
	.w5(32'h388b5c00),
	.w6(32'h395fb814),
	.w7(32'h3915df71),
	.w8(32'h386a78a8),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3762c01b),
	.w1(32'h37314152),
	.w2(32'hb7e33856),
	.w3(32'hb7fbe7f0),
	.w4(32'h37434551),
	.w5(32'hb7d79c9e),
	.w6(32'hb7aa89e3),
	.w7(32'hb7187cd7),
	.w8(32'hb835ad6a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39171b47),
	.w1(32'h3902b14f),
	.w2(32'h38f318f6),
	.w3(32'h392939ba),
	.w4(32'h39358e4b),
	.w5(32'h384b66c1),
	.w6(32'h3932b96e),
	.w7(32'h3873c6c0),
	.w8(32'h38195bf0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ad584c),
	.w1(32'h379a11eb),
	.w2(32'h36935561),
	.w3(32'h3629a040),
	.w4(32'h378920aa),
	.w5(32'hb6841d98),
	.w6(32'h36324075),
	.w7(32'h37737704),
	.w8(32'h35f12834),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c2c0cd),
	.w1(32'hb774ddfc),
	.w2(32'h370baa0d),
	.w3(32'hb7dfed6d),
	.w4(32'hb77da221),
	.w5(32'h37dcacd9),
	.w6(32'h3643c65f),
	.w7(32'hb73657bb),
	.w8(32'h37bb2dd9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7854527),
	.w1(32'hb72cc9e8),
	.w2(32'h378b823f),
	.w3(32'h368ba0e5),
	.w4(32'h37c1d70e),
	.w5(32'h37d2e353),
	.w6(32'hb6f6a9d6),
	.w7(32'h37486ece),
	.w8(32'h34847993),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a76e00),
	.w1(32'h380b4ebd),
	.w2(32'h38cc1ade),
	.w3(32'h3954b89d),
	.w4(32'h3912168c),
	.w5(32'h391ce069),
	.w6(32'h389de154),
	.w7(32'hb8de9309),
	.w8(32'h381738b1),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75109c4),
	.w1(32'hb72448e5),
	.w2(32'hb7929825),
	.w3(32'hb707751f),
	.w4(32'h369c7121),
	.w5(32'h35d0d40d),
	.w6(32'hb61ca7c4),
	.w7(32'h367c938c),
	.w8(32'h3729441e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8116aa4),
	.w1(32'hb7e5a298),
	.w2(32'hb7844254),
	.w3(32'hb74cdfbb),
	.w4(32'hb7684a09),
	.w5(32'hb632a66a),
	.w6(32'hb63b0f46),
	.w7(32'hb7415144),
	.w8(32'hb606b10a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e5c2f7),
	.w1(32'hb80e39cf),
	.w2(32'h368cc49e),
	.w3(32'h37d7f3b8),
	.w4(32'hb7c2d54e),
	.w5(32'h376e9222),
	.w6(32'h37c30bb2),
	.w7(32'hb871cc77),
	.w8(32'h38028742),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3800f07d),
	.w1(32'hb79fde4b),
	.w2(32'h37eedd51),
	.w3(32'h38b454c0),
	.w4(32'h390fc6c6),
	.w5(32'h38f1fd4a),
	.w6(32'h392e53f1),
	.w7(32'h38ab2a4c),
	.w8(32'h38a21a5b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b88bda),
	.w1(32'hb8b8095e),
	.w2(32'hb7dbb8cd),
	.w3(32'h374c6f85),
	.w4(32'h38782bb5),
	.w5(32'h393f7185),
	.w6(32'h3946d77f),
	.w7(32'h3948cc38),
	.w8(32'hb75ad80b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37978cc3),
	.w1(32'h3823e894),
	.w2(32'h37a1153b),
	.w3(32'hb65ac6d1),
	.w4(32'h374e8f33),
	.w5(32'h38077562),
	.w6(32'h35125797),
	.w7(32'h372e126b),
	.w8(32'h381ff54f),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38974148),
	.w1(32'h37b91cac),
	.w2(32'h38015f19),
	.w3(32'h3923e764),
	.w4(32'hb84b1be7),
	.w5(32'hb7e2bc41),
	.w6(32'h395d4ebf),
	.w7(32'hb9633928),
	.w8(32'hb9b1b9bc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38096d5f),
	.w1(32'hb96f72ea),
	.w2(32'h37d9d1e4),
	.w3(32'h3988b0c2),
	.w4(32'h38aa3b26),
	.w5(32'h39636b1a),
	.w6(32'h38dfd181),
	.w7(32'hb7137722),
	.w8(32'h39678cce),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382c76d1),
	.w1(32'h3704c7dc),
	.w2(32'hb7f217b0),
	.w3(32'h37c5b584),
	.w4(32'h38545f68),
	.w5(32'h3841909c),
	.w6(32'h37a2d943),
	.w7(32'h37831260),
	.w8(32'hb7a4d2c2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e07d4b),
	.w1(32'hb671f6be),
	.w2(32'hb695baf5),
	.w3(32'h36978a60),
	.w4(32'h35041e8d),
	.w5(32'h3642c0ee),
	.w6(32'hb57bdc54),
	.w7(32'hb5569672),
	.w8(32'h36a164cb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76c523a),
	.w1(32'hb7a7723e),
	.w2(32'hb785726b),
	.w3(32'h37996b78),
	.w4(32'h382fa445),
	.w5(32'hb6f9ae13),
	.w6(32'hb78242d2),
	.w7(32'h388448dd),
	.w8(32'h38186fd8),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65a1679),
	.w1(32'h36fe0f60),
	.w2(32'h3623eb82),
	.w3(32'hb74812da),
	.w4(32'h363d888e),
	.w5(32'h3643d6cd),
	.w6(32'hb5751b3f),
	.w7(32'h363dec5d),
	.w8(32'h368b4a4d),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3865097a),
	.w1(32'h38d04092),
	.w2(32'hb801d63b),
	.w3(32'h3849fb69),
	.w4(32'h38d370bd),
	.w5(32'h380b52da),
	.w6(32'h3911b8aa),
	.w7(32'h38e6ca8b),
	.w8(32'hb840190c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39208e5e),
	.w1(32'h38218aef),
	.w2(32'h389dd09b),
	.w3(32'h3863697c),
	.w4(32'hb81f6b00),
	.w5(32'hb8887097),
	.w6(32'h38e2134f),
	.w7(32'h37b1a065),
	.w8(32'hb8191066),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37569b84),
	.w1(32'h383f4f02),
	.w2(32'h38c3cf6e),
	.w3(32'h38d46f18),
	.w4(32'h387d5c12),
	.w5(32'h38738a5b),
	.w6(32'h38af1d5b),
	.w7(32'h37fd2366),
	.w8(32'h3618769a),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38426cd9),
	.w1(32'h36a7d787),
	.w2(32'h3800f9f5),
	.w3(32'hb738f9ed),
	.w4(32'hb8389f22),
	.w5(32'h37a191f0),
	.w6(32'h38139329),
	.w7(32'h36f61d0f),
	.w8(32'h382a0edb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a46a64),
	.w1(32'h3b5c4f72),
	.w2(32'hbbc02104),
	.w3(32'h38df4a48),
	.w4(32'h3b24fc32),
	.w5(32'hbc297e7c),
	.w6(32'h390db64e),
	.w7(32'hbb68b85f),
	.w8(32'hbbaad399),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2fc43),
	.w1(32'hbb1b28eb),
	.w2(32'hbb4f9670),
	.w3(32'hbc341167),
	.w4(32'hba3a82ae),
	.w5(32'h3b2e0ffe),
	.w6(32'h3b48236b),
	.w7(32'h3ba9251b),
	.w8(32'hbb639875),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb35cd5),
	.w1(32'hbb42cfa8),
	.w2(32'hbc2eddf4),
	.w3(32'hbb295771),
	.w4(32'hbc2fb458),
	.w5(32'h3c4ebef4),
	.w6(32'hbb36f892),
	.w7(32'hbbdfa1d4),
	.w8(32'h3c08b9a3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c447c64),
	.w1(32'h3aab5c87),
	.w2(32'h3c3d0376),
	.w3(32'h3c2e05e7),
	.w4(32'h39738b5d),
	.w5(32'hbaee5312),
	.w6(32'h3ba1d2ae),
	.w7(32'h3b1687fd),
	.w8(32'h3ba992eb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd15bc),
	.w1(32'hb9441f76),
	.w2(32'hb9c0efda),
	.w3(32'h3bcdd127),
	.w4(32'h3b799fd8),
	.w5(32'hbc835c80),
	.w6(32'hbb12b4bd),
	.w7(32'h3aed1bfc),
	.w8(32'hbbda4e26),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb351752),
	.w1(32'hbbe8e159),
	.w2(32'hbb83e4c4),
	.w3(32'h3b9abdc6),
	.w4(32'hbbdbd38a),
	.w5(32'hbabab620),
	.w6(32'hbb115803),
	.w7(32'hbc37b239),
	.w8(32'hbb477f29),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1ed2db),
	.w1(32'h3b9277c0),
	.w2(32'h3b46bee7),
	.w3(32'h38e30689),
	.w4(32'hbb003cdb),
	.w5(32'h3a6cbd48),
	.w6(32'hbb09a093),
	.w7(32'hbc4cd866),
	.w8(32'hbb936565),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42b089),
	.w1(32'h3b701a98),
	.w2(32'hba9dc821),
	.w3(32'hbb13251e),
	.w4(32'hbbb380d5),
	.w5(32'h3b409683),
	.w6(32'h3b55bcce),
	.w7(32'h3ba020cc),
	.w8(32'hbb424d30),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c373c),
	.w1(32'hbc4978ef),
	.w2(32'hbb00f95d),
	.w3(32'hbacaa79b),
	.w4(32'hbc29470c),
	.w5(32'h3c33d939),
	.w6(32'h3b2b4dab),
	.w7(32'hbb9c855b),
	.w8(32'h3bb33eb9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5f44b),
	.w1(32'hbc3d7cf8),
	.w2(32'h3b2a708e),
	.w3(32'hbbc7c732),
	.w4(32'hbb811da5),
	.w5(32'h3d008c4f),
	.w6(32'h3b406471),
	.w7(32'hbc2e37f0),
	.w8(32'h3affbad0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc818dff),
	.w1(32'hbbdba698),
	.w2(32'hbbb07240),
	.w3(32'hbbf412aa),
	.w4(32'hbbed3ad4),
	.w5(32'hbba70e20),
	.w6(32'hbc0156de),
	.w7(32'hbae31c11),
	.w8(32'hbc83fadc),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94bb5e),
	.w1(32'h3ca5ae13),
	.w2(32'h3c453e69),
	.w3(32'hbb98871a),
	.w4(32'h3cc99da5),
	.w5(32'hbb5d12b0),
	.w6(32'hbb2e135f),
	.w7(32'h3cb26122),
	.w8(32'h3c4a8c30),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c224aff),
	.w1(32'h3991dd32),
	.w2(32'h3b8e8366),
	.w3(32'hbb165b6d),
	.w4(32'hbb0909bf),
	.w5(32'hbc1177d9),
	.w6(32'h3c29b57e),
	.w7(32'h3a2e0296),
	.w8(32'h3ab8b04b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bad00),
	.w1(32'h398caace),
	.w2(32'h389026af),
	.w3(32'h3bd99b77),
	.w4(32'h3b52a1c8),
	.w5(32'h3c56e153),
	.w6(32'h3c043703),
	.w7(32'h3b8354ce),
	.w8(32'h3b0bd87e),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0406),
	.w1(32'hbbbb0f2a),
	.w2(32'hbb8b5130),
	.w3(32'hbb12eb1e),
	.w4(32'h3b6a566c),
	.w5(32'hbc5d77af),
	.w6(32'hbb41ba7c),
	.w7(32'h3bcfbde9),
	.w8(32'hbae99ea9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82fa8d),
	.w1(32'hbb2fb78b),
	.w2(32'h3a673176),
	.w3(32'h3ba79db9),
	.w4(32'hbbccf1b2),
	.w5(32'hbb7ecb90),
	.w6(32'hb802e82a),
	.w7(32'hbbc7b2d5),
	.w8(32'h3c4471ef),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc4f7a),
	.w1(32'hbb83f132),
	.w2(32'hba2a81e7),
	.w3(32'h3c99fa0c),
	.w4(32'h3bde77b9),
	.w5(32'h3c06abe8),
	.w6(32'h3b45f6d2),
	.w7(32'h3bd9e579),
	.w8(32'h3a60e9a5),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0640a8),
	.w1(32'hbcc06996),
	.w2(32'hbb6ef554),
	.w3(32'hbbd31d82),
	.w4(32'hbb970e5a),
	.w5(32'h3c88647d),
	.w6(32'hbbf8db26),
	.w7(32'hba5607db),
	.w8(32'hbc44849d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b6202),
	.w1(32'hbc9ec581),
	.w2(32'h3c69d2d9),
	.w3(32'h3b780bf5),
	.w4(32'hbbfcff47),
	.w5(32'hbbc11379),
	.w6(32'h3bedd4b5),
	.w7(32'h3bb6b726),
	.w8(32'hbc1a7ebb),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3eb92),
	.w1(32'hbabeeeb5),
	.w2(32'hbb1d7f00),
	.w3(32'h3b805396),
	.w4(32'hbb11a7a7),
	.w5(32'h39b3bd84),
	.w6(32'h3af4822a),
	.w7(32'h3ba21121),
	.w8(32'h39154093),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d5c87),
	.w1(32'hbc37e0e8),
	.w2(32'hbb4d455d),
	.w3(32'hbb44cb4e),
	.w4(32'hbc3fe163),
	.w5(32'h3c94ac5a),
	.w6(32'hbb3c0c30),
	.w7(32'hbbd45be8),
	.w8(32'hba83afa6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f648),
	.w1(32'hbc1ca696),
	.w2(32'hbab5e861),
	.w3(32'h3b206158),
	.w4(32'hbc4d44e8),
	.w5(32'h3a59f775),
	.w6(32'hbab95923),
	.w7(32'hbbb52dfc),
	.w8(32'h3a26dee8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f95bb),
	.w1(32'hbb94e0c1),
	.w2(32'hbbc6815e),
	.w3(32'h3c1430df),
	.w4(32'h3be45754),
	.w5(32'h3b116931),
	.w6(32'hbaa0f35a),
	.w7(32'h396c4067),
	.w8(32'hbbb0cf3e),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd624e),
	.w1(32'h390cdc09),
	.w2(32'hbbb51b29),
	.w3(32'hbaeb815a),
	.w4(32'hbb74e301),
	.w5(32'hbc0263b0),
	.w6(32'hbbe4303e),
	.w7(32'h3b7a232e),
	.w8(32'h39b67cae),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a176060),
	.w1(32'h3a697e6d),
	.w2(32'hbb34c685),
	.w3(32'h3bb458c1),
	.w4(32'hb9d2af46),
	.w5(32'hbbd64352),
	.w6(32'hbb470158),
	.w7(32'h3b10c984),
	.w8(32'hbc241f6f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b728),
	.w1(32'h392721ca),
	.w2(32'hbb5f0223),
	.w3(32'h3ba9c9d7),
	.w4(32'hbb36d2f0),
	.w5(32'hbb12aea4),
	.w6(32'hbade15ad),
	.w7(32'h3b2003cf),
	.w8(32'hbc3e1e32),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf50af3),
	.w1(32'hbc04706a),
	.w2(32'hbb9b44e3),
	.w3(32'hbb55749d),
	.w4(32'hbbb85f6e),
	.w5(32'hbc9d94c7),
	.w6(32'hbb1e2260),
	.w7(32'hbb8bba9c),
	.w8(32'hbc1779e9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc871fdc),
	.w1(32'hbbf458c2),
	.w2(32'h3c015aad),
	.w3(32'h3c0444e6),
	.w4(32'hbaf996a1),
	.w5(32'hbc67f00e),
	.w6(32'hbc452520),
	.w7(32'h3c09032e),
	.w8(32'h3c0046de),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb380ab9),
	.w1(32'hbb0e98bc),
	.w2(32'hbb4608f1),
	.w3(32'h3bf34335),
	.w4(32'hbc13a9cb),
	.w5(32'h3c527cc4),
	.w6(32'h3a6ad2ce),
	.w7(32'hbb597b63),
	.w8(32'h3adb7e6d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8af74d),
	.w1(32'hbbebef7b),
	.w2(32'hbae16809),
	.w3(32'hbc1bd944),
	.w4(32'hbc317159),
	.w5(32'hbb7c5f66),
	.w6(32'hbb81c662),
	.w7(32'hbb74fcc3),
	.w8(32'h3c57d6c0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af95a71),
	.w1(32'h3c08914d),
	.w2(32'hbb006cae),
	.w3(32'hbb864e3f),
	.w4(32'h3bbd6871),
	.w5(32'h3c136465),
	.w6(32'h3b3febdd),
	.w7(32'h3a1debd6),
	.w8(32'h3be14b41),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b6bbf),
	.w1(32'hbc63272a),
	.w2(32'hbbd35bb1),
	.w3(32'h3abafa8b),
	.w4(32'hbc187dc3),
	.w5(32'hba820c2a),
	.w6(32'hba916d3b),
	.w7(32'hbbaea32b),
	.w8(32'h3b9a7d10),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6827a2),
	.w1(32'hbaf2ab4d),
	.w2(32'hbc4ffb7a),
	.w3(32'h3c02446b),
	.w4(32'hbc47510a),
	.w5(32'hba9bff46),
	.w6(32'h3c01a7b4),
	.w7(32'hbc3eca99),
	.w8(32'h3b82ee77),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085058),
	.w1(32'hbc0d20c5),
	.w2(32'hb9d932ac),
	.w3(32'h3b423db0),
	.w4(32'hbc1e0d64),
	.w5(32'hbb7fa051),
	.w6(32'hbbc3ba22),
	.w7(32'hbc545b8e),
	.w8(32'hbc0e1b0d),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed6d4e),
	.w1(32'hbbc7bea0),
	.w2(32'h3a952ba3),
	.w3(32'h3a5861f9),
	.w4(32'h39f58b14),
	.w5(32'h3c915648),
	.w6(32'hbae12835),
	.w7(32'hbc0dad24),
	.w8(32'h3c401845),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3e3cd),
	.w1(32'hbb3d7e1e),
	.w2(32'hbacb0963),
	.w3(32'h3c8754d0),
	.w4(32'h3b9b13c9),
	.w5(32'hba9566dc),
	.w6(32'h3abe1dc1),
	.w7(32'h3b842120),
	.w8(32'h3c149229),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ab516),
	.w1(32'hbbd72446),
	.w2(32'hbabed0ba),
	.w3(32'hbc69ea54),
	.w4(32'hbbb86731),
	.w5(32'h399ca323),
	.w6(32'hba63712e),
	.w7(32'h3aff99b6),
	.w8(32'h381cd2a0),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd86bf4),
	.w1(32'h3b5a0b0d),
	.w2(32'hbaf2e3da),
	.w3(32'h3b0e7e34),
	.w4(32'h3afeccb6),
	.w5(32'h3bd199b0),
	.w6(32'hbb7864f5),
	.w7(32'hbb170257),
	.w8(32'h3ae72159),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc9927),
	.w1(32'hbbb2ac02),
	.w2(32'h3b584058),
	.w3(32'hbc805ee7),
	.w4(32'h3bb1c1cc),
	.w5(32'hbbfe02e2),
	.w6(32'hba498f6a),
	.w7(32'h3c0381e0),
	.w8(32'hba9fb00d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac76662),
	.w1(32'h3b9477b6),
	.w2(32'h3af4fd9e),
	.w3(32'hbbe113c0),
	.w4(32'h3bca2de3),
	.w5(32'hbc1411b7),
	.w6(32'hbbb8b270),
	.w7(32'h3b9fc531),
	.w8(32'h3c2115e6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d5c88),
	.w1(32'h3b19a7ac),
	.w2(32'hbc0b55ff),
	.w3(32'hba9ed83d),
	.w4(32'hbb419f40),
	.w5(32'hbc408bba),
	.w6(32'hbadade38),
	.w7(32'hbb941dfa),
	.w8(32'h3b403d8c),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd57aa9),
	.w1(32'h3c09e6f9),
	.w2(32'h3bfc1ea3),
	.w3(32'h3bf530cb),
	.w4(32'h3bcebb2d),
	.w5(32'h3b2ecd08),
	.w6(32'hbb44cb01),
	.w7(32'h3b93036f),
	.w8(32'h3b978b30),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04df2d),
	.w1(32'h3b4e643a),
	.w2(32'h3c14a074),
	.w3(32'h399e887c),
	.w4(32'hba3597bb),
	.w5(32'hbbbb9478),
	.w6(32'h3c2649b4),
	.w7(32'h3bcf1f90),
	.w8(32'h3bf0968a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3beee5),
	.w1(32'h3c2d44fc),
	.w2(32'h3c22cf29),
	.w3(32'hb8ea55f5),
	.w4(32'hba025038),
	.w5(32'hbcc3b475),
	.w6(32'h3bfa2afa),
	.w7(32'h3c033beb),
	.w8(32'hbb053d55),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb197514),
	.w1(32'hbc084904),
	.w2(32'hbb114ba9),
	.w3(32'h3cc8c58f),
	.w4(32'hbbd863d3),
	.w5(32'h3c9cc541),
	.w6(32'h3c12cc88),
	.w7(32'hbc1bc78c),
	.w8(32'hbae84914),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b961ec8),
	.w1(32'hbc2c2bbf),
	.w2(32'hba6ff09b),
	.w3(32'h3c1e1a33),
	.w4(32'hbb6d519c),
	.w5(32'h3d066a66),
	.w6(32'h3aad0cb8),
	.w7(32'hba8cc40b),
	.w8(32'h3b834578),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b139),
	.w1(32'hbbc7f4d9),
	.w2(32'hbb6fef18),
	.w3(32'h3a259f9d),
	.w4(32'hbc006a85),
	.w5(32'h3b76a343),
	.w6(32'h3b227145),
	.w7(32'hbc02c072),
	.w8(32'h37dbb4f4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9b690),
	.w1(32'h3af16451),
	.w2(32'hbbee41c1),
	.w3(32'h3ae9049d),
	.w4(32'hbb181e66),
	.w5(32'hbc0fd11a),
	.w6(32'hbb782788),
	.w7(32'hb9bd974a),
	.w8(32'h39cc8669),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c5981),
	.w1(32'h3b50adbf),
	.w2(32'h3ba15e00),
	.w3(32'h3c7e1bee),
	.w4(32'hba0fca23),
	.w5(32'h3b2520b5),
	.w6(32'hbbb452da),
	.w7(32'h3be77f0c),
	.w8(32'hbbc3a5ad),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c76ea),
	.w1(32'hbc84e188),
	.w2(32'hbb5a0a31),
	.w3(32'hbbb68b77),
	.w4(32'hbca0e61b),
	.w5(32'hbcbe874c),
	.w6(32'hbb751872),
	.w7(32'hbacdecea),
	.w8(32'hbc6a9649),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cf7db),
	.w1(32'hbb29043d),
	.w2(32'hba5d094d),
	.w3(32'hbc2abe98),
	.w4(32'hbc3aac4b),
	.w5(32'h3c9fcd46),
	.w6(32'hbbf9d60e),
	.w7(32'hbc0c449a),
	.w8(32'h3b5b724e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdb39d),
	.w1(32'h3b64ec65),
	.w2(32'h36a29a4b),
	.w3(32'hbbe4bb7b),
	.w4(32'h3b66cf8f),
	.w5(32'hbb8a8efb),
	.w6(32'hbb68bc3c),
	.w7(32'h3b81dda3),
	.w8(32'h3a12828a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb33da),
	.w1(32'h3b8f123a),
	.w2(32'hb9a02ceb),
	.w3(32'hbbd53364),
	.w4(32'h3b86bf8c),
	.w5(32'hbc7546da),
	.w6(32'hbbc82e86),
	.w7(32'hb9d926cc),
	.w8(32'h3c0d4191),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb919eca),
	.w1(32'h3babbfa1),
	.w2(32'h3c0ce081),
	.w3(32'hbc258d21),
	.w4(32'h3b24d31f),
	.w5(32'hbc237afb),
	.w6(32'h3b495896),
	.w7(32'h3bd0f6d5),
	.w8(32'h3b5b6e46),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b465d10),
	.w1(32'h3c4226bb),
	.w2(32'h3b6582a8),
	.w3(32'h3c72c92d),
	.w4(32'h3c0e2f94),
	.w5(32'hbd2176d2),
	.w6(32'h3aa3ecc2),
	.w7(32'h3c5047d5),
	.w8(32'h37bfa019),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3adf62),
	.w1(32'h3c3a65bc),
	.w2(32'hba074f23),
	.w3(32'h3c92b8e6),
	.w4(32'h3b44c860),
	.w5(32'hbbd027db),
	.w6(32'h3b7f4602),
	.w7(32'hbc044ad6),
	.w8(32'h3c2d6161),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e1d09),
	.w1(32'hbc0abee6),
	.w2(32'hbc53d7d5),
	.w3(32'h3bbe277c),
	.w4(32'hbc334856),
	.w5(32'h3c5fe56c),
	.w6(32'h3bec5b82),
	.w7(32'hbc82644d),
	.w8(32'h3b2657a3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a6830),
	.w1(32'h3a2aacdb),
	.w2(32'hbb2d745c),
	.w3(32'hba665341),
	.w4(32'hbc0c39d3),
	.w5(32'h3bb5d6e8),
	.w6(32'h3be1ed5b),
	.w7(32'h3a16e6a5),
	.w8(32'hbbce373c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86b32b),
	.w1(32'hbc20ae25),
	.w2(32'hbbd7c229),
	.w3(32'hbb699815),
	.w4(32'h3bb3b829),
	.w5(32'h3abddb30),
	.w6(32'hbc12b871),
	.w7(32'h3b9b6b8f),
	.w8(32'h3ba6c0e8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule