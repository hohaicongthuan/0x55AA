module layer_8_featuremap_64(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a444ca2),
	.w1(32'hba75c7d1),
	.w2(32'hba9354d0),
	.w3(32'h3a6e36d1),
	.w4(32'hbaa33d3b),
	.w5(32'hba5337fd),
	.w6(32'hb9b83381),
	.w7(32'hb829392f),
	.w8(32'hb9b689b6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d63e2),
	.w1(32'hba0d4d17),
	.w2(32'hba021e31),
	.w3(32'hb95a2903),
	.w4(32'hba4849c2),
	.w5(32'hba16501c),
	.w6(32'hba0eb690),
	.w7(32'hba22734b),
	.w8(32'h39e05362),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39662a62),
	.w1(32'hb9423850),
	.w2(32'hb8cc2ed5),
	.w3(32'h39f214f8),
	.w4(32'hb924e8ca),
	.w5(32'hb8b58f2d),
	.w6(32'hb9018b10),
	.w7(32'hb88faf2b),
	.w8(32'h391c8b87),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41788c),
	.w1(32'hbabda37f),
	.w2(32'h3adb956d),
	.w3(32'hb9cf40cf),
	.w4(32'hba723503),
	.w5(32'hb99129e1),
	.w6(32'hba24bc2b),
	.w7(32'hb9979171),
	.w8(32'h3a88d607),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a866cc4),
	.w1(32'h3a1e21cc),
	.w2(32'hb90c52e6),
	.w3(32'h3a3d2d4e),
	.w4(32'h39c666dd),
	.w5(32'hb999509d),
	.w6(32'h3a983def),
	.w7(32'h3a2c880d),
	.w8(32'h3b669738),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b264bd2),
	.w1(32'hba5e4595),
	.w2(32'hb94f4731),
	.w3(32'h3b50e31d),
	.w4(32'hba668bfa),
	.w5(32'hba6df28b),
	.w6(32'hb57ac835),
	.w7(32'h39be83c7),
	.w8(32'h3a5ac6f2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89526c),
	.w1(32'hb9594b19),
	.w2(32'hba5b381f),
	.w3(32'h3a6f36c9),
	.w4(32'h37f76d34),
	.w5(32'hba12fb07),
	.w6(32'h39bf3343),
	.w7(32'h3805c24b),
	.w8(32'h3a78203f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bccb4),
	.w1(32'h3a3ce498),
	.w2(32'hb6a13925),
	.w3(32'h3a0ea345),
	.w4(32'h3934ac8c),
	.w5(32'hba1c48aa),
	.w6(32'h3aaacc46),
	.w7(32'h3a0b7424),
	.w8(32'h3a790b9d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a970d5e),
	.w1(32'h39640850),
	.w2(32'hba793645),
	.w3(32'h3a3995ae),
	.w4(32'hb9b6dd5c),
	.w5(32'hba8c0197),
	.w6(32'h3a02a4eb),
	.w7(32'hb99b1529),
	.w8(32'h3a65a095),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4b39a),
	.w1(32'hba019387),
	.w2(32'h3a6d5f1a),
	.w3(32'hbbaa445f),
	.w4(32'hba89c393),
	.w5(32'hb9a96ce5),
	.w6(32'h3ad139bf),
	.w7(32'hbb3dec03),
	.w8(32'h3a63519c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58e429),
	.w1(32'h3a6b0784),
	.w2(32'hb9ffc5e2),
	.w3(32'hb935f01b),
	.w4(32'h39ab02cb),
	.w5(32'hba49c39e),
	.w6(32'h3ab10dae),
	.w7(32'h3a0f65f2),
	.w8(32'h394fa718),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a343e42),
	.w1(32'hb929b926),
	.w2(32'hba1fcb7b),
	.w3(32'h3a35918e),
	.w4(32'hb9385d18),
	.w5(32'hba091bc1),
	.w6(32'h38b75ba5),
	.w7(32'hb928f468),
	.w8(32'h3a74fff8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49b591),
	.w1(32'hb9a6acd1),
	.w2(32'hba0995b4),
	.w3(32'hb8bc42c9),
	.w4(32'hba33716d),
	.w5(32'hba0fcfdf),
	.w6(32'h39811b9b),
	.w7(32'hb9da7a28),
	.w8(32'h3b8f7ca5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b541fe0),
	.w1(32'hba8ae26b),
	.w2(32'hb96312da),
	.w3(32'h3b87c78f),
	.w4(32'hba4834f8),
	.w5(32'hba4cfcd8),
	.w6(32'hb8afdec0),
	.w7(32'h39c79f1e),
	.w8(32'h3afffd5f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0c57b),
	.w1(32'hba5cb3c5),
	.w2(32'h389e7b9f),
	.w3(32'h3b1179d1),
	.w4(32'hb99b5dfe),
	.w5(32'hba07f308),
	.w6(32'h395dd8fe),
	.w7(32'h3a06afbc),
	.w8(32'hb98887a5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24e2e6),
	.w1(32'hbad2d293),
	.w2(32'hba12be22),
	.w3(32'hba589a83),
	.w4(32'hbb0d2576),
	.w5(32'hba04f52e),
	.w6(32'hbab45c8a),
	.w7(32'hba4563ed),
	.w8(32'h362ccf3e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1af97),
	.w1(32'hbb51bac6),
	.w2(32'h3adee640),
	.w3(32'hbba2c121),
	.w4(32'h396a2bb2),
	.w5(32'h3b37cd4f),
	.w6(32'hbb819d2c),
	.w7(32'hbb805c76),
	.w8(32'h39fab25d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10d5db),
	.w1(32'hb9880e9a),
	.w2(32'hba54be10),
	.w3(32'hb884c46b),
	.w4(32'hba3136e9),
	.w5(32'hba660a9f),
	.w6(32'hb81ceeb5),
	.w7(32'hba642b26),
	.w8(32'h39bcf3fb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a552964),
	.w1(32'hb9879bdb),
	.w2(32'hbab42199),
	.w3(32'hba352a5d),
	.w4(32'hbac45139),
	.w5(32'hbb1cbcc0),
	.w6(32'h3ab59db0),
	.w7(32'h39d18435),
	.w8(32'hbb930d65),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d2ca0),
	.w1(32'h3be576dc),
	.w2(32'h3b3e71b6),
	.w3(32'hba38e2fc),
	.w4(32'hba479a85),
	.w5(32'hbaa82f59),
	.w6(32'h3b0d1d7d),
	.w7(32'hb97b4db4),
	.w8(32'hb9896fa3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a531d2),
	.w1(32'h3a96911b),
	.w2(32'h3a8c3b35),
	.w3(32'h3ad687a1),
	.w4(32'h3b1e8a1b),
	.w5(32'h3aeabc17),
	.w6(32'h3a712417),
	.w7(32'h3a8e6273),
	.w8(32'h3aa506b5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94651d2),
	.w1(32'hb91d8733),
	.w2(32'h381703b2),
	.w3(32'hb6932c0b),
	.w4(32'hb98033c5),
	.w5(32'hb904e423),
	.w6(32'hb8a9ed31),
	.w7(32'hb9d60b60),
	.w8(32'h3a78a5b7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b388697),
	.w1(32'h3ab5e408),
	.w2(32'h3aaa781e),
	.w3(32'h3b83fbf6),
	.w4(32'h3b88555e),
	.w5(32'h3b7c855d),
	.w6(32'h399c257b),
	.w7(32'h3a69cd7b),
	.w8(32'h3b1a8ebb),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af552ec),
	.w1(32'h3a60c6e7),
	.w2(32'h39a18dde),
	.w3(32'h3ab4e060),
	.w4(32'hb9a40199),
	.w5(32'hb9517f3b),
	.w6(32'h3a51d8d8),
	.w7(32'h3a5262e1),
	.w8(32'hbbcc829e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe208c1),
	.w1(32'hbb22972e),
	.w2(32'hbb218989),
	.w3(32'hbbed7d42),
	.w4(32'hbb9f9a52),
	.w5(32'hbb83f136),
	.w6(32'hbba80eae),
	.w7(32'hbb679f2a),
	.w8(32'h3ad908b5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa7403),
	.w1(32'h3a3a17be),
	.w2(32'h3a459603),
	.w3(32'h3b5b610a),
	.w4(32'h3b6d1c59),
	.w5(32'h3b601a7b),
	.w6(32'hb9b6debf),
	.w7(32'h398b9ac6),
	.w8(32'h3a8fedd6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5d5f8),
	.w1(32'h3a35a4ee),
	.w2(32'h3a5be640),
	.w3(32'h3b2fab92),
	.w4(32'h3b3a3e1a),
	.w5(32'h3b46b6ab),
	.w6(32'hb98e73f9),
	.w7(32'hb846896b),
	.w8(32'hba2a8734),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4c5c4),
	.w1(32'h3b56a143),
	.w2(32'hba337a40),
	.w3(32'h3afadb76),
	.w4(32'h3b45f612),
	.w5(32'h3ac3ebb8),
	.w6(32'h3af98fa4),
	.w7(32'h3ad0a1b4),
	.w8(32'h3b023760),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba416388),
	.w1(32'h3a83686d),
	.w2(32'h3ac7aacf),
	.w3(32'h3a966dcd),
	.w4(32'hbb2c2302),
	.w5(32'h3a11135c),
	.w6(32'h39147b9e),
	.w7(32'h3aa5e4de),
	.w8(32'h39828a0e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399dc76e),
	.w1(32'hb892539c),
	.w2(32'h38d81a85),
	.w3(32'h3987d17f),
	.w4(32'hb8c894ad),
	.w5(32'hb884c62e),
	.w6(32'h35a0fd31),
	.w7(32'h38c5af99),
	.w8(32'h3a48895e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58ed28),
	.w1(32'h3a8f45e9),
	.w2(32'h3badb8fc),
	.w3(32'hbac142e3),
	.w4(32'hba6a30e2),
	.w5(32'hbb3e6206),
	.w6(32'h39ae26b1),
	.w7(32'h3b403466),
	.w8(32'hbae9315d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba518fcd),
	.w1(32'h39b66eef),
	.w2(32'h3a30aa13),
	.w3(32'h39f47943),
	.w4(32'h3ac16efc),
	.w5(32'h3b0cf2f1),
	.w6(32'h39d01e85),
	.w7(32'h3a8ef73f),
	.w8(32'h3b6a0a6c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae23634),
	.w1(32'hbb42ad5b),
	.w2(32'h3b50a681),
	.w3(32'h3b1eeb02),
	.w4(32'h3a1f8e89),
	.w5(32'h3a933c3f),
	.w6(32'h3a3543b8),
	.w7(32'h3b209bf7),
	.w8(32'h38a16eb8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dbdca),
	.w1(32'h3c34885f),
	.w2(32'h3b6b94bc),
	.w3(32'hbb0ad3e4),
	.w4(32'hbb837856),
	.w5(32'hb9424a0b),
	.w6(32'h3bb2569b),
	.w7(32'h3b6d97a3),
	.w8(32'h3b78e337),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3622ba),
	.w1(32'hba6bc8a1),
	.w2(32'hb94bc078),
	.w3(32'h3b63df42),
	.w4(32'hba364f80),
	.w5(32'hba3e8223),
	.w6(32'hb96f9429),
	.w7(32'h3995c030),
	.w8(32'h3a8f26fc),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac26dd),
	.w1(32'h38833322),
	.w2(32'hba81725b),
	.w3(32'h3a82f0df),
	.w4(32'hbaa7b2a6),
	.w5(32'hba8c0a00),
	.w6(32'h3a5232a3),
	.w7(32'h39071f19),
	.w8(32'hbb953ec3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252712),
	.w1(32'h3a9676b2),
	.w2(32'hbb120018),
	.w3(32'hbb6ef4dc),
	.w4(32'hbb0bb0cb),
	.w5(32'hbb2cc7b6),
	.w6(32'hb9c9ae95),
	.w7(32'hbabb02e6),
	.w8(32'h39da57cc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7bbb3),
	.w1(32'hb87f49cc),
	.w2(32'h39890571),
	.w3(32'h3a3b338a),
	.w4(32'h368c4857),
	.w5(32'h397817dc),
	.w6(32'hb5f6696c),
	.w7(32'h3948b765),
	.w8(32'h3b486306),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cb59e),
	.w1(32'hbae51134),
	.w2(32'h3a24c281),
	.w3(32'h3b8c984a),
	.w4(32'h38fb6ee5),
	.w5(32'hba038ecc),
	.w6(32'h3894409d),
	.w7(32'h3a8f660e),
	.w8(32'hbb082a1a),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe1f2),
	.w1(32'h3a5ce5ff),
	.w2(32'h36aaf9f8),
	.w3(32'hba9feeed),
	.w4(32'h39dd3c00),
	.w5(32'h39d716a6),
	.w6(32'h396ea1f8),
	.w7(32'h39a7f207),
	.w8(32'h39a0fc3b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39edea6d),
	.w1(32'h391fc3e1),
	.w2(32'h394db5ba),
	.w3(32'h3a8b65b2),
	.w4(32'h3ab358f7),
	.w5(32'h3ab5cbfd),
	.w6(32'hb949d7b4),
	.w7(32'hb86bc97d),
	.w8(32'hbb0a1f44),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd4ba7),
	.w1(32'hbaad0204),
	.w2(32'hba69c2df),
	.w3(32'hba2d32eb),
	.w4(32'hbb2122dc),
	.w5(32'hba324f4c),
	.w6(32'hbb6ce3f5),
	.w7(32'hbb8a96ff),
	.w8(32'hbc0d0648),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84de63),
	.w1(32'h3b9852d4),
	.w2(32'hb9d1b1b0),
	.w3(32'hbc6353ce),
	.w4(32'h3cd58298),
	.w5(32'hbc114573),
	.w6(32'hbc9347d2),
	.w7(32'h3a6bfce9),
	.w8(32'h3aa372ac),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39764f62),
	.w1(32'hba96c25c),
	.w2(32'h3b4bd70b),
	.w3(32'h3a2507cc),
	.w4(32'hbae24c65),
	.w5(32'h3b2159ca),
	.w6(32'h3b8726a5),
	.w7(32'hbb201d85),
	.w8(32'hbb0d34f8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a533c7),
	.w1(32'hbb655906),
	.w2(32'h39c7e19b),
	.w3(32'h3a0c65c5),
	.w4(32'hbaa02096),
	.w5(32'h3b09684d),
	.w6(32'hbb9e4378),
	.w7(32'hbbb9008e),
	.w8(32'h3b2080ee),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bdd53),
	.w1(32'hbb7021d4),
	.w2(32'h3bca162b),
	.w3(32'hbb746357),
	.w4(32'hbb0519ac),
	.w5(32'h3b3cfec8),
	.w6(32'h3a682fb0),
	.w7(32'hbbf1bd57),
	.w8(32'h3b58dc52),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c612bfb),
	.w1(32'hbbbdd8e3),
	.w2(32'h3c34b14a),
	.w3(32'h3a05a25f),
	.w4(32'hbc88a8e0),
	.w5(32'h3bdff478),
	.w6(32'hbccb9e18),
	.w7(32'hbbe6492f),
	.w8(32'hbb9ce3b8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926bad6),
	.w1(32'hbb5a5d1e),
	.w2(32'h3b85694d),
	.w3(32'hbb2ac90a),
	.w4(32'hbbcf2541),
	.w5(32'hbc45ed9b),
	.w6(32'h3c287b04),
	.w7(32'h3b9169ea),
	.w8(32'h3b3c698e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b077b0d),
	.w1(32'h3a592411),
	.w2(32'hbbea698c),
	.w3(32'hbb782248),
	.w4(32'h3b812530),
	.w5(32'hbaef547e),
	.w6(32'hbbd59dd9),
	.w7(32'h3b1f5eb0),
	.w8(32'hbb04d13a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a373f2),
	.w1(32'hbac618c8),
	.w2(32'h3af320df),
	.w3(32'h39f2546c),
	.w4(32'hba0bb411),
	.w5(32'h3b06ae3e),
	.w6(32'hbae05745),
	.w7(32'hbbb3bb3c),
	.w8(32'hb77b1c7a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ffa16),
	.w1(32'h3a109f7c),
	.w2(32'h3b3cf70e),
	.w3(32'hb913398e),
	.w4(32'hbab6638e),
	.w5(32'h3b112ccb),
	.w6(32'h398d7233),
	.w7(32'hbaf62937),
	.w8(32'h391c8bc9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab08e0),
	.w1(32'hb98a9cfd),
	.w2(32'h3b77ee8d),
	.w3(32'h3a439df9),
	.w4(32'hbb5e69b4),
	.w5(32'h3ae5d4a1),
	.w6(32'h3b6bbb2c),
	.w7(32'hbb5e3a4d),
	.w8(32'hb91acb86),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e955d),
	.w1(32'h3cc636c6),
	.w2(32'hbc1946f3),
	.w3(32'hbb5022b1),
	.w4(32'hbc5d29fd),
	.w5(32'h3c3cc8c5),
	.w6(32'hbc9369e2),
	.w7(32'hbb6d664f),
	.w8(32'hbab75d6f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61d652),
	.w1(32'hbbaadf69),
	.w2(32'hbb494e42),
	.w3(32'hbb3addd8),
	.w4(32'h39d2a18e),
	.w5(32'h3a1b78b2),
	.w6(32'hbc1082fc),
	.w7(32'hbb20191c),
	.w8(32'hbc3cf898),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdcbaff),
	.w1(32'hbcb7552f),
	.w2(32'hbb6402db),
	.w3(32'h3c01ff44),
	.w4(32'h3bd2e0ac),
	.w5(32'hbb128777),
	.w6(32'hbbdcdc4f),
	.w7(32'h3ab1ba73),
	.w8(32'hbc3cb072),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5ae33),
	.w1(32'hbc75dc04),
	.w2(32'hbac7f8ed),
	.w3(32'hba9a5078),
	.w4(32'hbc1a2a68),
	.w5(32'hbbe0972a),
	.w6(32'hbb98cef2),
	.w7(32'hbae3e999),
	.w8(32'h3a9857d6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bec3a),
	.w1(32'h3b2feb15),
	.w2(32'hb9e899fa),
	.w3(32'h3bd94dd0),
	.w4(32'h3c5b1c02),
	.w5(32'h3c1030eb),
	.w6(32'h3c9eda1f),
	.w7(32'h3b2650ce),
	.w8(32'hbc99e848),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5390a3),
	.w1(32'hbb936fc7),
	.w2(32'hbc707135),
	.w3(32'hbc872e68),
	.w4(32'hbc275906),
	.w5(32'hbc54c1b5),
	.w6(32'hbc4e2f6c),
	.w7(32'hbc1dac22),
	.w8(32'h3a4d01dd),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745cfd),
	.w1(32'hbba4e413),
	.w2(32'hbb4b7294),
	.w3(32'h3ae01281),
	.w4(32'h3a7f0b33),
	.w5(32'hbb014182),
	.w6(32'h3b9331ea),
	.w7(32'h3adfcc35),
	.w8(32'h3b19fdc1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be44b47),
	.w1(32'h3bf4f78a),
	.w2(32'hba8ff5a4),
	.w3(32'hbaa234a6),
	.w4(32'hb525fe6b),
	.w5(32'hbb68704e),
	.w6(32'hbbf5dfb6),
	.w7(32'h3b5a1186),
	.w8(32'h3b8cb013),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fddc0),
	.w1(32'hbbeb4220),
	.w2(32'h3c979e0a),
	.w3(32'h3c971cbf),
	.w4(32'h3b4f7459),
	.w5(32'h3bab387c),
	.w6(32'hbc68b501),
	.w7(32'hbb145b50),
	.w8(32'h3a8da8f5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa1e2),
	.w1(32'h3ab0369e),
	.w2(32'hb5875306),
	.w3(32'hbb0abfbc),
	.w4(32'h3b4945df),
	.w5(32'hbbcc8137),
	.w6(32'h3c837a57),
	.w7(32'h39828187),
	.w8(32'hbb9dc46d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30e433),
	.w1(32'hbc0e5e46),
	.w2(32'hbb498b5c),
	.w3(32'hba0d29ef),
	.w4(32'hbb3ab98b),
	.w5(32'hb9f2233b),
	.w6(32'hbc245260),
	.w7(32'hbc39e823),
	.w8(32'hbc996146),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4809bf),
	.w1(32'h3c41ff88),
	.w2(32'hbc8639b0),
	.w3(32'hbaf2c1a7),
	.w4(32'hbac2fe06),
	.w5(32'hbc7310c7),
	.w6(32'hbcb6717e),
	.w7(32'hbc060266),
	.w8(32'h3a80c401),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a14e72),
	.w1(32'hbb02fc0a),
	.w2(32'h37c60acd),
	.w3(32'h392c9f3a),
	.w4(32'hbad9686e),
	.w5(32'h3b32a72d),
	.w6(32'h39a2a694),
	.w7(32'hbb556d0c),
	.w8(32'h39298066),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff9492),
	.w1(32'hb9ceced6),
	.w2(32'h3ae94eb8),
	.w3(32'h39cd2114),
	.w4(32'hb9fe4343),
	.w5(32'h3aa15dcf),
	.w6(32'h3accc447),
	.w7(32'hba498007),
	.w8(32'hb93ca99f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5d853),
	.w1(32'h391c108b),
	.w2(32'h3a860bb5),
	.w3(32'hb8e689d7),
	.w4(32'hba038b40),
	.w5(32'h3abbc07d),
	.w6(32'hba3dad28),
	.w7(32'hbafc6f03),
	.w8(32'hbb82ada9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c87c3),
	.w1(32'h3c5fc37e),
	.w2(32'h3a219031),
	.w3(32'hbaa7affc),
	.w4(32'hbb28a178),
	.w5(32'hbbe1914f),
	.w6(32'h3cac72e1),
	.w7(32'h3a018a31),
	.w8(32'hbb1468e1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9990bd4),
	.w1(32'hbad9edf7),
	.w2(32'h39c8c303),
	.w3(32'h3aab781f),
	.w4(32'hba260adb),
	.w5(32'h3b0f0773),
	.w6(32'hbb09fcf2),
	.w7(32'hbb8f7f6e),
	.w8(32'hbb1e9dc8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe29ad),
	.w1(32'hbc000977),
	.w2(32'h3b26ebe7),
	.w3(32'h3bd4ffdb),
	.w4(32'hbb39159b),
	.w5(32'hbaa2d543),
	.w6(32'h3c76e314),
	.w7(32'hba2be288),
	.w8(32'hba826e46),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66454c),
	.w1(32'hbae59282),
	.w2(32'hb9b1f3d9),
	.w3(32'hba677399),
	.w4(32'hbb168a68),
	.w5(32'h39031e3d),
	.w6(32'hbb594487),
	.w7(32'hbbca1d3e),
	.w8(32'hbad8a5a3),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39912ebb),
	.w1(32'hb9c7fd81),
	.w2(32'h3a36e2a0),
	.w3(32'h39f7aafc),
	.w4(32'hb9df4735),
	.w5(32'h3acb0e40),
	.w6(32'hbae00d00),
	.w7(32'hbb97244d),
	.w8(32'h38629fcb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a924381),
	.w1(32'hba4f09ef),
	.w2(32'h38a5094d),
	.w3(32'hb8ffde00),
	.w4(32'hbb1257a2),
	.w5(32'h3b33dddb),
	.w6(32'hbb6b57de),
	.w7(32'hbbd834eb),
	.w8(32'hbc9a31df),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3338d5),
	.w1(32'h3d283169),
	.w2(32'hbc6d2101),
	.w3(32'hbb65857b),
	.w4(32'hbc55560c),
	.w5(32'hbcdbbf27),
	.w6(32'hbb333efe),
	.w7(32'hbbfbd80c),
	.w8(32'hbb92f8ee),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a0173),
	.w1(32'hba110d01),
	.w2(32'hbbae41ea),
	.w3(32'hbafe9b54),
	.w4(32'hbb359080),
	.w5(32'hb8f808d2),
	.w6(32'hbbec4abd),
	.w7(32'hbbe737c4),
	.w8(32'h38a3307b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a380),
	.w1(32'hba54d1b5),
	.w2(32'h3aea601f),
	.w3(32'h3a1277d7),
	.w4(32'hba92804b),
	.w5(32'h3a899729),
	.w6(32'h3ab9c12b),
	.w7(32'hbb3e3ecf),
	.w8(32'hbb24f191),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94669f),
	.w1(32'hba3c0b45),
	.w2(32'hba59eea5),
	.w3(32'hba328db9),
	.w4(32'hba1320eb),
	.w5(32'h397c854d),
	.w6(32'hbb0f1428),
	.w7(32'hbb2b770f),
	.w8(32'hbb2cf1e1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24171a),
	.w1(32'hbc2452b7),
	.w2(32'h3b13bbf9),
	.w3(32'h3be022fa),
	.w4(32'hbb540eac),
	.w5(32'hbabc27de),
	.w6(32'h3c89954e),
	.w7(32'hba6b8362),
	.w8(32'hbaf278fe),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85814),
	.w1(32'hbbcea1cc),
	.w2(32'h3bb31ab7),
	.w3(32'h3b6c99de),
	.w4(32'hbb95c27e),
	.w5(32'hbab39cc1),
	.w6(32'h3c3c746f),
	.w7(32'hbaec4947),
	.w8(32'hba832b5c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8de44be),
	.w1(32'hbb212ef8),
	.w2(32'h38a43467),
	.w3(32'hba0b9552),
	.w4(32'hbb48dcd9),
	.w5(32'h3a19210b),
	.w6(32'h3bad3641),
	.w7(32'hb9d25829),
	.w8(32'hbc804a15),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60767a),
	.w1(32'h3d226444),
	.w2(32'hbcee93ed),
	.w3(32'hba9b1902),
	.w4(32'h3cc09379),
	.w5(32'hbbdacc72),
	.w6(32'hbad1cd49),
	.w7(32'h3b9bc874),
	.w8(32'hbabf8a28),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc3bfd),
	.w1(32'hba887723),
	.w2(32'hba7ca213),
	.w3(32'hbab639a4),
	.w4(32'hba751b76),
	.w5(32'h3a87a438),
	.w6(32'hbb1600ae),
	.w7(32'hbb03f737),
	.w8(32'hba98e0bf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8a665),
	.w1(32'hbb00c3d4),
	.w2(32'h3bf1f867),
	.w3(32'hbb83e9fb),
	.w4(32'hbabe85e6),
	.w5(32'h3b995b30),
	.w6(32'h3b46c348),
	.w7(32'hbb9c9b2d),
	.w8(32'hbb198e71),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3039c2),
	.w1(32'h3b1c554c),
	.w2(32'hbcaa7fd5),
	.w3(32'h3ba58ba7),
	.w4(32'h3cb402f6),
	.w5(32'h3abec9fa),
	.w6(32'h3c043bf8),
	.w7(32'hbc57e4ad),
	.w8(32'h3ad0770b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285e25),
	.w1(32'hb9f96a0e),
	.w2(32'h3ac02741),
	.w3(32'hbac74879),
	.w4(32'h38d09392),
	.w5(32'hb805121b),
	.w6(32'hbaac87dd),
	.w7(32'h3b1cca9f),
	.w8(32'hbb83cb5c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39d7bb),
	.w1(32'hbb467dba),
	.w2(32'hbaae17d9),
	.w3(32'h3a98bdee),
	.w4(32'hba110bce),
	.w5(32'h396f1698),
	.w6(32'hbb968607),
	.w7(32'hbbdd7f97),
	.w8(32'h3b6f0c16),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30e98c),
	.w1(32'h3a8f236b),
	.w2(32'hbc1b9007),
	.w3(32'hbba317ef),
	.w4(32'h3bad89fa),
	.w5(32'hbb19ffa1),
	.w6(32'hbc0cc850),
	.w7(32'h3b545997),
	.w8(32'h3abde83a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0987fd),
	.w1(32'hbb8c2c6c),
	.w2(32'h3aa710ca),
	.w3(32'h3b321b49),
	.w4(32'hbb40112d),
	.w5(32'h3b960bca),
	.w6(32'h38b83051),
	.w7(32'hbba18b9b),
	.w8(32'hbb1c0fa7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab94bed),
	.w1(32'h3bef7411),
	.w2(32'hbc0215fb),
	.w3(32'hbb5fc77f),
	.w4(32'h3bfa8b72),
	.w5(32'hbbe3b3f1),
	.w6(32'hbb3a0fe1),
	.w7(32'hb9c02bcf),
	.w8(32'h3b5f21c1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef0f0),
	.w1(32'h3a87d008),
	.w2(32'hbc138e4b),
	.w3(32'hbb96c908),
	.w4(32'h3ba1e73a),
	.w5(32'hbb19cb16),
	.w6(32'hbc03add2),
	.w7(32'h3b4a45bf),
	.w8(32'h3b3f7be6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0eb3f7),
	.w1(32'h3a7257af),
	.w2(32'hbbf80942),
	.w3(32'hbb83b9f0),
	.w4(32'h3b8a88d0),
	.w5(32'hbaf6d72c),
	.w6(32'hbbe2ba94),
	.w7(32'h3b2abcc0),
	.w8(32'h39b051ac),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fe48d),
	.w1(32'hbae6c7fa),
	.w2(32'hba2c3c5c),
	.w3(32'hbbc6fb5a),
	.w4(32'h383b1edb),
	.w5(32'hbae38ecd),
	.w6(32'hbbb7b79a),
	.w7(32'hb98030a8),
	.w8(32'hbb601030),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacf19b),
	.w1(32'hbc6dd9e3),
	.w2(32'h388c3ccc),
	.w3(32'hbb18651a),
	.w4(32'hbc82910a),
	.w5(32'h3b45971d),
	.w6(32'h3c86eb62),
	.w7(32'hbb8ff231),
	.w8(32'hb966f1ec),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ac5e2),
	.w1(32'h391f229e),
	.w2(32'h3a466234),
	.w3(32'hb9ef2629),
	.w4(32'hbabeb0d5),
	.w5(32'hb88cfad8),
	.w6(32'h3a4b4df7),
	.w7(32'hbac399e1),
	.w8(32'hbc2527e4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12dc99),
	.w1(32'hbb6e172f),
	.w2(32'hbc6fd1f1),
	.w3(32'hbc4b8ce8),
	.w4(32'h3c0bf711),
	.w5(32'hbcb5f7c4),
	.w6(32'hbb045912),
	.w7(32'hbba4372e),
	.w8(32'h3b4e58e8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e48f5),
	.w1(32'h3b434fcb),
	.w2(32'h3b628deb),
	.w3(32'hbc1307b3),
	.w4(32'hbb1e5a1b),
	.w5(32'hbbc79d02),
	.w6(32'hbacc2a86),
	.w7(32'h3b94e3b3),
	.w8(32'hbc946c65),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31d4d7),
	.w1(32'hbbcc9ebc),
	.w2(32'hbbe7ede1),
	.w3(32'hbb86d4fa),
	.w4(32'hbb0e1866),
	.w5(32'hbc437301),
	.w6(32'h3ad2fbe7),
	.w7(32'hbbbd8e49),
	.w8(32'hbb6259d8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb68a2),
	.w1(32'h3a2d5a75),
	.w2(32'hba5e9e75),
	.w3(32'hbb83547b),
	.w4(32'hba8ea329),
	.w5(32'hbc034cec),
	.w6(32'h3bc0a642),
	.w7(32'h3b20a4f0),
	.w8(32'hbb18578e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119dbf),
	.w1(32'hbc0e6195),
	.w2(32'h3b14add0),
	.w3(32'h3bc29502),
	.w4(32'hbb399fad),
	.w5(32'hba8708c0),
	.w6(32'h3c6f1e32),
	.w7(32'hba80a0be),
	.w8(32'h3a8a58f4),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77287c),
	.w1(32'hbb838610),
	.w2(32'h3b9a4099),
	.w3(32'h3a56ea2f),
	.w4(32'hb86fa6d5),
	.w5(32'h3c0ac8e7),
	.w6(32'h3ae7af08),
	.w7(32'hbb138871),
	.w8(32'hbb1138d5),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a797019),
	.w1(32'h3a7b4f7b),
	.w2(32'hbba47259),
	.w3(32'hb8e548af),
	.w4(32'h3aecd641),
	.w5(32'hbc068118),
	.w6(32'hbbf8c2ef),
	.w7(32'h3b44f027),
	.w8(32'h383cca10),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec4a0),
	.w1(32'h39635630),
	.w2(32'h3af41664),
	.w3(32'hb9888ce4),
	.w4(32'hbac3dd55),
	.w5(32'h3affbb70),
	.w6(32'hba1c9504),
	.w7(32'hbb12ee91),
	.w8(32'hbb9f7d94),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56964b),
	.w1(32'hbc939df5),
	.w2(32'h3c39b33c),
	.w3(32'h3c125a63),
	.w4(32'hbc0a6823),
	.w5(32'hbba91eda),
	.w6(32'h3cb8e650),
	.w7(32'hbb28a331),
	.w8(32'h3aedf36f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee0349),
	.w1(32'h3b4f7193),
	.w2(32'h3aa13a35),
	.w3(32'hbb8bcff4),
	.w4(32'h3b21d5a2),
	.w5(32'hbb3c7be2),
	.w6(32'hbac060fd),
	.w7(32'h3ab760c8),
	.w8(32'h3ac19e17),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa740f6),
	.w1(32'h3a36b349),
	.w2(32'hbb61351d),
	.w3(32'hbb05cd4d),
	.w4(32'h3b008f99),
	.w5(32'hba570a53),
	.w6(32'hbb6b309e),
	.w7(32'h3a9f842b),
	.w8(32'h3930f2b0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89437b),
	.w1(32'h394525bf),
	.w2(32'hb928583f),
	.w3(32'h3a9100a6),
	.w4(32'h3a09d642),
	.w5(32'hb7acdf40),
	.w6(32'h3aa72bc1),
	.w7(32'h3a823517),
	.w8(32'hbb6fa004),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e1d19),
	.w1(32'hbb13962c),
	.w2(32'h3afce43a),
	.w3(32'h3a62639c),
	.w4(32'hb87e81b5),
	.w5(32'h393e6087),
	.w6(32'hbb60c76d),
	.w7(32'hb78ddb6b),
	.w8(32'hba5bce95),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f82055),
	.w1(32'hb9cf9e7b),
	.w2(32'hb9975103),
	.w3(32'hba3277b4),
	.w4(32'hb9e9fe45),
	.w5(32'hb986d56c),
	.w6(32'hb9c943d3),
	.w7(32'hba1d2a1b),
	.w8(32'hb838fbc9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902758f),
	.w1(32'hba145f0e),
	.w2(32'h388859c3),
	.w3(32'hb9803d75),
	.w4(32'hb9f1a728),
	.w5(32'hb9978c00),
	.w6(32'hb9a83b49),
	.w7(32'hb9079dff),
	.w8(32'hb95e9c96),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0df59),
	.w1(32'hb9b5eb93),
	.w2(32'h39aba413),
	.w3(32'h38e50f51),
	.w4(32'h3a498e04),
	.w5(32'h3a8a255a),
	.w6(32'hbada61f7),
	.w7(32'h39254f42),
	.w8(32'hbad6f872),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0379bf),
	.w1(32'h3bf30157),
	.w2(32'h3adfc7f5),
	.w3(32'h3b3f32e2),
	.w4(32'h3b7f3255),
	.w5(32'h3b02e6fe),
	.w6(32'hbaaf0b59),
	.w7(32'h3a3e3008),
	.w8(32'hbae48bf1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaaddd2),
	.w1(32'hba88592c),
	.w2(32'h3963db9d),
	.w3(32'hbaf1af5b),
	.w4(32'hb99ba976),
	.w5(32'hb7b7c181),
	.w6(32'hbb094fd1),
	.w7(32'hb9d90abb),
	.w8(32'h3a97e8b6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fcb7dc),
	.w1(32'h388ddc7b),
	.w2(32'h3a0bdca1),
	.w3(32'hb9edf20a),
	.w4(32'hb90ba4cd),
	.w5(32'hb8f22b21),
	.w6(32'h3a135912),
	.w7(32'h3b0d127c),
	.w8(32'hb9b4e01d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa430a),
	.w1(32'hba2b1031),
	.w2(32'h3939993f),
	.w3(32'hb88fe016),
	.w4(32'hb8e2b148),
	.w5(32'h38bca024),
	.w6(32'hba1d5788),
	.w7(32'h381c31a6),
	.w8(32'hb9d5c7cf),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9938b48),
	.w1(32'hb9836f51),
	.w2(32'hb98497c5),
	.w3(32'hb8f56cbe),
	.w4(32'hb8fa0bf1),
	.w5(32'hb8a96881),
	.w6(32'hb9253e33),
	.w7(32'hb9f7f185),
	.w8(32'hba465692),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389003fb),
	.w1(32'h38d2b64e),
	.w2(32'hb8f58bf0),
	.w3(32'h3929f4a0),
	.w4(32'h395962d5),
	.w5(32'hb8e20dfa),
	.w6(32'h3942baf8),
	.w7(32'hba15d5aa),
	.w8(32'h3b4953f8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dec804),
	.w1(32'hbb129128),
	.w2(32'h3a88b9d9),
	.w3(32'hbaa61b8f),
	.w4(32'h3969cda7),
	.w5(32'h3b55318a),
	.w6(32'hb9df2469),
	.w7(32'hbb8a65f2),
	.w8(32'hb7a4a822),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba356cf9),
	.w1(32'hb8d5da1f),
	.w2(32'h3aafea27),
	.w3(32'hb9b00d35),
	.w4(32'h3a3a92e6),
	.w5(32'h3ac61c80),
	.w6(32'hb94da984),
	.w7(32'h3abc37e9),
	.w8(32'hba0d3aff),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb170dea),
	.w1(32'h3ab99564),
	.w2(32'h3b194195),
	.w3(32'h39e8df3d),
	.w4(32'h3b460517),
	.w5(32'h3b58cf60),
	.w6(32'hbb04d3da),
	.w7(32'h39e7c1f7),
	.w8(32'hbb9f0fd2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce90d),
	.w1(32'h3ad08098),
	.w2(32'h399bd863),
	.w3(32'hbab26196),
	.w4(32'h3b495181),
	.w5(32'hb9b5defa),
	.w6(32'hbb627bb2),
	.w7(32'hbb45fa33),
	.w8(32'hb9ae8cbe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a67cf),
	.w1(32'hbb193a9a),
	.w2(32'hba194fb4),
	.w3(32'hba3a62a8),
	.w4(32'hbac8d1bc),
	.w5(32'h3aaa04fc),
	.w6(32'hba31b207),
	.w7(32'hb9eb990b),
	.w8(32'h3afbe23b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88365e),
	.w1(32'hb908ed17),
	.w2(32'hbb1d6824),
	.w3(32'h3ae1f81d),
	.w4(32'h3b6b4809),
	.w5(32'h3a12cfd1),
	.w6(32'h3a1a70e5),
	.w7(32'hb974ad9f),
	.w8(32'hb96858a5),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ea08b),
	.w1(32'hb9c4fc52),
	.w2(32'h39478e8a),
	.w3(32'hb935258d),
	.w4(32'h395b85b4),
	.w5(32'h3a23088e),
	.w6(32'h3972a6ee),
	.w7(32'h39b3f13a),
	.w8(32'h3b42c645),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f57e30),
	.w1(32'hbb17ac16),
	.w2(32'hb92cd06c),
	.w3(32'hba9adb93),
	.w4(32'hbb148878),
	.w5(32'hba9a3a73),
	.w6(32'h3a885c89),
	.w7(32'h3a71e3e4),
	.w8(32'h399bcebb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb646249),
	.w1(32'hbb194954),
	.w2(32'hba1301a9),
	.w3(32'h3b472404),
	.w4(32'h3b366ffc),
	.w5(32'h3b63756d),
	.w6(32'hbb5323d6),
	.w7(32'hb922731c),
	.w8(32'hbac6265a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3a440),
	.w1(32'h3aca6c46),
	.w2(32'h39aaf2d1),
	.w3(32'h39aa673a),
	.w4(32'hb8a74ca8),
	.w5(32'hb6c8fe38),
	.w6(32'hbb15eab1),
	.w7(32'hba13243d),
	.w8(32'hbb0acef9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc2468),
	.w1(32'hbaeb4cfc),
	.w2(32'hba878ac8),
	.w3(32'hba962131),
	.w4(32'hba7922e9),
	.w5(32'hb8eb0ef9),
	.w6(32'hbacee65f),
	.w7(32'hba949484),
	.w8(32'h39b93018),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f1454),
	.w1(32'hbb1888a1),
	.w2(32'hbb461c10),
	.w3(32'hbb4a9e1d),
	.w4(32'hbaf185c3),
	.w5(32'hbb83da7a),
	.w6(32'hbadad44d),
	.w7(32'hbb3a9abc),
	.w8(32'hb9c8c65c),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule