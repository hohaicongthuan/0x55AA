module layer_8_featuremap_8(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fa935),
	.w1(32'h3ba13b0d),
	.w2(32'h3b34cc28),
	.w3(32'hba0b2a86),
	.w4(32'h3b8f8d95),
	.w5(32'hbaa7423a),
	.w6(32'h3be0d3a5),
	.w7(32'h3ba305da),
	.w8(32'hbb956896),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92664d),
	.w1(32'hba180456),
	.w2(32'hbb9b85ec),
	.w3(32'h3acac15c),
	.w4(32'hbb227f19),
	.w5(32'hbb9d08d2),
	.w6(32'h3aa7385a),
	.w7(32'hb9872600),
	.w8(32'hbb6fa83e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb814cd3),
	.w1(32'hbb9a9f8b),
	.w2(32'h392fe2fb),
	.w3(32'hbb5d9bc9),
	.w4(32'hbc0c8d95),
	.w5(32'hbba40f02),
	.w6(32'hbb968cff),
	.w7(32'hbc1944ef),
	.w8(32'hbba5197d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc11b0f),
	.w1(32'hbb3556ad),
	.w2(32'h3b9e9cdf),
	.w3(32'h39f00c65),
	.w4(32'hbc3801c1),
	.w5(32'hbb8b17ad),
	.w6(32'hbb5a5112),
	.w7(32'hbc62ace7),
	.w8(32'hbc1a3e66),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c66bd5b),
	.w1(32'h3ad757d6),
	.w2(32'h3b2aabae),
	.w3(32'h3b92e9d7),
	.w4(32'h3a653656),
	.w5(32'h37131055),
	.w6(32'hba759735),
	.w7(32'h3b0e82fd),
	.w8(32'hbb14cdea),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92269ed),
	.w1(32'h39a2eba0),
	.w2(32'h39a2c01b),
	.w3(32'h3b0a8cc6),
	.w4(32'hbb52fc55),
	.w5(32'hbbb9f09e),
	.w6(32'hbaabb53d),
	.w7(32'h3b393cdd),
	.w8(32'h3aaf751f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49ecbf),
	.w1(32'h3b0d9695),
	.w2(32'hbae13bb5),
	.w3(32'hbad530ba),
	.w4(32'hbb88bddc),
	.w5(32'hbbd62e3f),
	.w6(32'h3a7e6150),
	.w7(32'hbc08cda4),
	.w8(32'hbc3f2b59),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01bd22),
	.w1(32'hbad22c63),
	.w2(32'hbba97cac),
	.w3(32'hbbdd3a4a),
	.w4(32'hbc059df3),
	.w5(32'hbc39b530),
	.w6(32'hbc1230bf),
	.w7(32'hba30550d),
	.w8(32'hbbd321d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf209c7),
	.w1(32'hbba97039),
	.w2(32'hbc836fe6),
	.w3(32'hbc81ce8a),
	.w4(32'hbc3be7f1),
	.w5(32'hbcc2fe05),
	.w6(32'hb8c85b5a),
	.w7(32'hbb37e324),
	.w8(32'hbc60b16c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b140009),
	.w1(32'h39e5abd9),
	.w2(32'hbbf7dc10),
	.w3(32'hbbbd1010),
	.w4(32'hbac19191),
	.w5(32'hbbc5fe28),
	.w6(32'hbb45a314),
	.w7(32'hbac9079c),
	.w8(32'h3a6b8b16),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992ee24),
	.w1(32'hba8ac02e),
	.w2(32'hbb833a9e),
	.w3(32'h3b2f4161),
	.w4(32'hbb61c652),
	.w5(32'hbb9241ec),
	.w6(32'h3bb882e8),
	.w7(32'hbb43bb48),
	.w8(32'hbb5f027d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a6ee3),
	.w1(32'h3b4ba8b5),
	.w2(32'hbaef6bef),
	.w3(32'hbb83610d),
	.w4(32'h3bb50128),
	.w5(32'hba6b6d17),
	.w6(32'hbaa51322),
	.w7(32'h3b8078b3),
	.w8(32'hbace6b5d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9271e0),
	.w1(32'h3ad55c7d),
	.w2(32'h3aaaebc4),
	.w3(32'h39654494),
	.w4(32'hbaadd2e1),
	.w5(32'h3a77a5ca),
	.w6(32'h3bc36c5f),
	.w7(32'hbc0961b7),
	.w8(32'hbb63984d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a9c9),
	.w1(32'h3b52a3bf),
	.w2(32'hbc477e95),
	.w3(32'h395b6458),
	.w4(32'hbbbe31ff),
	.w5(32'hbcb46cb0),
	.w6(32'hbbeaecbe),
	.w7(32'hbc05e7d7),
	.w8(32'hbcae780a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fa910),
	.w1(32'hbc088d34),
	.w2(32'hbc08b37d),
	.w3(32'hbcc50470),
	.w4(32'hbc3dab00),
	.w5(32'hbc56c62a),
	.w6(32'hbcad0c1f),
	.w7(32'hbc2f8e47),
	.w8(32'hbc1cd2b0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb6140),
	.w1(32'hba81438e),
	.w2(32'hba8bfa34),
	.w3(32'hbc0de8dc),
	.w4(32'hbbf553af),
	.w5(32'hbc113782),
	.w6(32'hbbfda90b),
	.w7(32'hb99ef3d9),
	.w8(32'hb8dba858),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f94093),
	.w1(32'h3bd57fea),
	.w2(32'h3b940a3d),
	.w3(32'hbbf885d2),
	.w4(32'h3a441cd4),
	.w5(32'hbaee9e74),
	.w6(32'h3aeb9ecd),
	.w7(32'hbaad6cd7),
	.w8(32'hbc06d455),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3b4fb),
	.w1(32'hbb4879d5),
	.w2(32'hbaa714cd),
	.w3(32'hbbc7c1d7),
	.w4(32'hbb548c5c),
	.w5(32'hbad5e570),
	.w6(32'hbc0d148c),
	.w7(32'hbb7268b1),
	.w8(32'hbb602f92),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e3d8e),
	.w1(32'h3c566de7),
	.w2(32'h3c534884),
	.w3(32'h3ba1b5dd),
	.w4(32'h3bc5fac7),
	.w5(32'h3bcf6f38),
	.w6(32'h3bbe8822),
	.w7(32'h3ca7b5d9),
	.w8(32'h3c63a9f4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d90a4),
	.w1(32'hbbb80066),
	.w2(32'hbc8d3c68),
	.w3(32'h3c7729ca),
	.w4(32'hbc8eedc3),
	.w5(32'hbd028bd3),
	.w6(32'h3cba50ef),
	.w7(32'hbb19726b),
	.w8(32'hbc66e8ae),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17d3b7),
	.w1(32'hbafa4d8d),
	.w2(32'h3c1fa7f5),
	.w3(32'hbcbd620f),
	.w4(32'h3c830add),
	.w5(32'h3d0c0ce6),
	.w6(32'hbc8f577a),
	.w7(32'h3c58eb13),
	.w8(32'h3cf4830e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb53ded),
	.w1(32'hbc00796b),
	.w2(32'hbb9cfe23),
	.w3(32'h3cb75883),
	.w4(32'hbc32ad0d),
	.w5(32'hbc007dab),
	.w6(32'h3ca8220f),
	.w7(32'h3add9f3f),
	.w8(32'hbb708faa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c532fcd),
	.w1(32'h3c036a61),
	.w2(32'h3c50c44c),
	.w3(32'h3bd1ca21),
	.w4(32'h3b965cfd),
	.w5(32'h39277ba1),
	.w6(32'h3bffb44c),
	.w7(32'h3c36458d),
	.w8(32'h3c162e42),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00cfbc),
	.w1(32'hbb48cbf5),
	.w2(32'h3b833b9a),
	.w3(32'h3bb4b7b1),
	.w4(32'h3b498c65),
	.w5(32'h3c691f70),
	.w6(32'h3b35f40f),
	.w7(32'h39b7c9be),
	.w8(32'h3c38681b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5660a),
	.w1(32'hb7b2ddaf),
	.w2(32'hba4d6876),
	.w3(32'h3c1af831),
	.w4(32'h3a6c5f41),
	.w5(32'hbbabc789),
	.w6(32'h3bfab82b),
	.w7(32'hbb92301f),
	.w8(32'hbbd706e2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7db3d),
	.w1(32'h3bb70c86),
	.w2(32'h3bd8b082),
	.w3(32'h3be84383),
	.w4(32'h3bb1525a),
	.w5(32'h3b6484d9),
	.w6(32'h3ba48cbb),
	.w7(32'h3c4eb4d1),
	.w8(32'h3c3944d8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca3a7f),
	.w1(32'hbcaa616e),
	.w2(32'hbc4a2075),
	.w3(32'h3bd2a8ed),
	.w4(32'hbc62c55e),
	.w5(32'h3bc2ced3),
	.w6(32'h3bfad09e),
	.w7(32'hbc566c8e),
	.w8(32'h3b36ead9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74749b),
	.w1(32'hbb9acdc4),
	.w2(32'hbc47a845),
	.w3(32'hba2d497a),
	.w4(32'h3a2be67f),
	.w5(32'hbb9b3dcf),
	.w6(32'hbaa3fdea),
	.w7(32'h3c432875),
	.w8(32'h3bc8fa74),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbef21),
	.w1(32'hbab88e70),
	.w2(32'hbb9852e5),
	.w3(32'hbbd21f34),
	.w4(32'hbb1d0b4b),
	.w5(32'hbbe42a7d),
	.w6(32'hbb368d5d),
	.w7(32'h3925197c),
	.w8(32'hbb27d76a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd37b2d),
	.w1(32'hbc2d1c70),
	.w2(32'hbc707119),
	.w3(32'hbc146692),
	.w4(32'hbc6ceabc),
	.w5(32'hbc9f502f),
	.w6(32'hbb9854be),
	.w7(32'hbc3941ca),
	.w8(32'hbc574f7a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed835),
	.w1(32'h3a137e1c),
	.w2(32'h3a00bd23),
	.w3(32'hbc537b07),
	.w4(32'h3b2e12b4),
	.w5(32'hbaf5912c),
	.w6(32'hbc1fb58b),
	.w7(32'h3a5f9f46),
	.w8(32'hba28e014),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e2171),
	.w1(32'h3c81ac16),
	.w2(32'h3cda5dc6),
	.w3(32'h3a807a65),
	.w4(32'h3cb0e3f9),
	.w5(32'h3d08d510),
	.w6(32'h3b89f05b),
	.w7(32'h3ca2ec32),
	.w8(32'h3d05da05),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc22605),
	.w1(32'h3bc29249),
	.w2(32'hbbac93e0),
	.w3(32'h3cff5a7e),
	.w4(32'hbb886548),
	.w5(32'hbc911591),
	.w6(32'h3ce4cc87),
	.w7(32'hbbed1a68),
	.w8(32'hbc9d76bc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b4090),
	.w1(32'h3b0d058c),
	.w2(32'h3992682d),
	.w3(32'hbc6adf1d),
	.w4(32'h3b34c396),
	.w5(32'h3ae30a10),
	.w6(32'hbc77145a),
	.w7(32'h3b953ae5),
	.w8(32'hb7e1dafd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e514c),
	.w1(32'hbbd25bb1),
	.w2(32'hbbb3e52a),
	.w3(32'hba1e325d),
	.w4(32'hbbb09c12),
	.w5(32'hbbafa12a),
	.w6(32'hba98954a),
	.w7(32'hbb16202b),
	.w8(32'h3a6b57a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28692e),
	.w1(32'hbba3d74d),
	.w2(32'hbb993e31),
	.w3(32'hb9cf3de4),
	.w4(32'hbbdbfcb6),
	.w5(32'hbb89b805),
	.w6(32'h3b216460),
	.w7(32'hbbf782d8),
	.w8(32'hbbaa28a8),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf51794),
	.w1(32'h3c1aa09a),
	.w2(32'h3b62fd1f),
	.w3(32'hbba8f246),
	.w4(32'h3be7f735),
	.w5(32'hb9f3cfae),
	.w6(32'hbba8f487),
	.w7(32'h3c0b9539),
	.w8(32'h3bb9ae73),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a6d9c),
	.w1(32'hb9cc0571),
	.w2(32'hbbc6ba8a),
	.w3(32'h3adf0019),
	.w4(32'hbb6f2bfb),
	.w5(32'hbb361f0a),
	.w6(32'h3c0459c2),
	.w7(32'hbb4af6c9),
	.w8(32'hba9520cd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1253f9),
	.w1(32'h3b2aa5ce),
	.w2(32'h3b374d05),
	.w3(32'hbb9140d5),
	.w4(32'h39e6071f),
	.w5(32'hbbb54c14),
	.w6(32'hbb9ba708),
	.w7(32'hbab41a47),
	.w8(32'hbbac4b32),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269197),
	.w1(32'h3b9dd174),
	.w2(32'h3ba3a175),
	.w3(32'hba0513d7),
	.w4(32'h3ba3dbea),
	.w5(32'h3b21b629),
	.w6(32'hbb48976b),
	.w7(32'h3b98af7c),
	.w8(32'h3ae37101),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c9fe),
	.w1(32'hba348f5e),
	.w2(32'h3b65c86b),
	.w3(32'h3b7dec7c),
	.w4(32'hbb1c021e),
	.w5(32'h3ba78d53),
	.w6(32'h3bbfeb23),
	.w7(32'hbb7265c5),
	.w8(32'hbb47ad93),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdf93e),
	.w1(32'hbb896f0c),
	.w2(32'hbc2a479c),
	.w3(32'h3b8af3d8),
	.w4(32'hbbe008e4),
	.w5(32'hbc4a3a7d),
	.w6(32'hb9dcaa0b),
	.w7(32'hbb6f8e2a),
	.w8(32'hbbaf686e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc270f),
	.w1(32'hbc572b34),
	.w2(32'hbc9e6b39),
	.w3(32'hbbfb3990),
	.w4(32'hbc9611b2),
	.w5(32'hbcdf36a8),
	.w6(32'hbb2ce6db),
	.w7(32'hbc8781aa),
	.w8(32'hbcc6f7fe),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73c719),
	.w1(32'h3aedf9c6),
	.w2(32'h3b3aef76),
	.w3(32'hbcb19a12),
	.w4(32'h3b167abd),
	.w5(32'h3921b8c6),
	.w6(32'hbc928c5d),
	.w7(32'h3ab1ca45),
	.w8(32'h3b6bc6c3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7fc55),
	.w1(32'hbaf65b1d),
	.w2(32'hbb6165ec),
	.w3(32'h3b2356e5),
	.w4(32'hbad8a1cd),
	.w5(32'hbbb68be6),
	.w6(32'h3c05ca15),
	.w7(32'h3b9f8adc),
	.w8(32'h3ba9bf3a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc4799),
	.w1(32'h3bceef33),
	.w2(32'h3b6a6c97),
	.w3(32'hbbfcda22),
	.w4(32'h3b74a7ca),
	.w5(32'h3bb0bd1f),
	.w6(32'h3a7266ee),
	.w7(32'h3bb422e0),
	.w8(32'h3c000b75),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed000),
	.w1(32'h3aaa677f),
	.w2(32'h3ab086ef),
	.w3(32'h3bb8adc2),
	.w4(32'hbaff9a22),
	.w5(32'hbb3f9408),
	.w6(32'h3c4e7dee),
	.w7(32'hba12b959),
	.w8(32'hbae3cf89),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eeba4),
	.w1(32'h3a693974),
	.w2(32'h3af8318e),
	.w3(32'h3bff8ca6),
	.w4(32'h3c004c8b),
	.w5(32'h3b566991),
	.w6(32'h3c8f9fb0),
	.w7(32'h3bfea21c),
	.w8(32'h3bb9f3d0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39002edb),
	.w1(32'h3b5eee56),
	.w2(32'hba7191b9),
	.w3(32'h3c033d87),
	.w4(32'hba910ff3),
	.w5(32'hbba99444),
	.w6(32'h3b80fc89),
	.w7(32'hba8bb732),
	.w8(32'hbbe5777f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ef1df),
	.w1(32'h3c1a4b4a),
	.w2(32'h3c016c68),
	.w3(32'hbabe849e),
	.w4(32'h3be5c707),
	.w5(32'h3ab0a53c),
	.w6(32'hbb2d9d9e),
	.w7(32'h3bedc107),
	.w8(32'hbc2b56a3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9e9e),
	.w1(32'h3b45424e),
	.w2(32'h3c2cf725),
	.w3(32'h3b3c4261),
	.w4(32'h3c5d9b4c),
	.w5(32'h3cd65c8e),
	.w6(32'h3b7efea9),
	.w7(32'h3c8c325e),
	.w8(32'h3cf611b2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9907a4),
	.w1(32'h3ae548c8),
	.w2(32'h3a184095),
	.w3(32'h3d1fb39f),
	.w4(32'h3b658551),
	.w5(32'h3af64c31),
	.w6(32'h3d165506),
	.w7(32'h3bfe4ce1),
	.w8(32'h3bf142be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e7dfb),
	.w1(32'h3af03e11),
	.w2(32'h3afc642e),
	.w3(32'h3b876d71),
	.w4(32'hba2d8a23),
	.w5(32'hbad26a23),
	.w6(32'h3c04cefc),
	.w7(32'hbb1fb369),
	.w8(32'hbb30a7b3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b18c),
	.w1(32'hba6a3b45),
	.w2(32'hbb9862c0),
	.w3(32'hbb8b66bf),
	.w4(32'h39a737f5),
	.w5(32'hbc56715f),
	.w6(32'hba48935a),
	.w7(32'h3ab52e53),
	.w8(32'hbbb1059e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944a71),
	.w1(32'h3b08af1c),
	.w2(32'h3be73fa2),
	.w3(32'hbbc14c79),
	.w4(32'h3aca9e57),
	.w5(32'hba398ea1),
	.w6(32'hbbc1c9d4),
	.w7(32'hbaedce72),
	.w8(32'hba2046fe),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b6619),
	.w1(32'hbad10fe1),
	.w2(32'hbb37f0e8),
	.w3(32'h3c4b22ff),
	.w4(32'hbb09020c),
	.w5(32'hbb005498),
	.w6(32'h3c6a5a90),
	.w7(32'h3b5ee177),
	.w8(32'h3b84f8c6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe7e57),
	.w1(32'h3b0d8c94),
	.w2(32'h3bd44897),
	.w3(32'hbab33a1e),
	.w4(32'h3b961fa5),
	.w5(32'h3c3569b9),
	.w6(32'h3b2ec6e1),
	.w7(32'h3bc013d1),
	.w8(32'h3c7793ad),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe16aa),
	.w1(32'h3b4e5c9b),
	.w2(32'hbac27aab),
	.w3(32'h3c6606be),
	.w4(32'hbb2475d0),
	.w5(32'hbb1d86f2),
	.w6(32'h3c8f3d88),
	.w7(32'hba94fadd),
	.w8(32'hba78ed9d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75ce34),
	.w1(32'h3adce4b4),
	.w2(32'hbb085eaf),
	.w3(32'h3ab09490),
	.w4(32'hbba6b593),
	.w5(32'hbc200e7f),
	.w6(32'h3ae998ce),
	.w7(32'hbb51db6b),
	.w8(32'hbc06dad7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290ec0),
	.w1(32'h3c05740e),
	.w2(32'h3b99cce8),
	.w3(32'hbc106929),
	.w4(32'h3b7a75bf),
	.w5(32'hbb3a8c7a),
	.w6(32'hbbe87158),
	.w7(32'h38273446),
	.w8(32'hb9a3a07e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45358d),
	.w1(32'hbaccddc0),
	.w2(32'hbb92b033),
	.w3(32'hbabcf8f6),
	.w4(32'hbbcd30ee),
	.w5(32'hbbe36045),
	.w6(32'h3b681251),
	.w7(32'hb7e74ba2),
	.w8(32'hba3d4c25),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24b71f),
	.w1(32'hbb834ec0),
	.w2(32'hbbf37be2),
	.w3(32'hbae1d08b),
	.w4(32'hbc000b73),
	.w5(32'hbc4d90b8),
	.w6(32'h3b9793a8),
	.w7(32'hbaf626d3),
	.w8(32'hbc1c331a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4d99),
	.w1(32'hbb6f82da),
	.w2(32'hbcaa3734),
	.w3(32'h3b85f098),
	.w4(32'hbcbee585),
	.w5(32'hbd41208e),
	.w6(32'h3c2530f9),
	.w7(32'hbc9c6d40),
	.w8(32'hbd2ef852),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5be5a2),
	.w1(32'h3baae390),
	.w2(32'h3ad33e97),
	.w3(32'hbd185218),
	.w4(32'hbc0c6633),
	.w5(32'hbb9bde79),
	.w6(32'hbd1159e4),
	.w7(32'hb75162c7),
	.w8(32'hba3803ee),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f94c9),
	.w1(32'hbb531728),
	.w2(32'hbb39280c),
	.w3(32'hbb6fcdb0),
	.w4(32'h39a34af3),
	.w5(32'h38d0fb54),
	.w6(32'h3b597b2f),
	.w7(32'h3aeb0c6a),
	.w8(32'h39a8ff7a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1312e3),
	.w1(32'hba88e420),
	.w2(32'hbb8b9a2f),
	.w3(32'h3b67e7a1),
	.w4(32'hba0121d8),
	.w5(32'hbb88368d),
	.w6(32'h3b81a4b5),
	.w7(32'h3b5202fa),
	.w8(32'h3b424784),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f2526),
	.w1(32'hbc0d76e1),
	.w2(32'hbd11093d),
	.w3(32'h396c5b9f),
	.w4(32'hbd0dc724),
	.w5(32'hbd89fb58),
	.w6(32'h3bb0f163),
	.w7(32'hbcdba861),
	.w8(32'hbd6b0c81),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca74174),
	.w1(32'hbb550aa5),
	.w2(32'hbd15fe4b),
	.w3(32'hbd4afe42),
	.w4(32'hbd335f2a),
	.w5(32'hbdace0af),
	.w6(32'hbd298086),
	.w7(32'hbce9eebe),
	.w8(32'hbd859a7b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e933e),
	.w1(32'h3bb08469),
	.w2(32'h3b6972a2),
	.w3(32'hbd7c3aff),
	.w4(32'h3aa8210b),
	.w5(32'h3a0d73a7),
	.w6(32'hbd3f05f9),
	.w7(32'h3b44a8d3),
	.w8(32'hbaa8248b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c590f39),
	.w1(32'h3a365b7f),
	.w2(32'hbab50b6c),
	.w3(32'h3bdbd355),
	.w4(32'h3bd66dd4),
	.w5(32'h3bc37420),
	.w6(32'h3bc1385d),
	.w7(32'h3bc91c3c),
	.w8(32'hbbc0a91a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ba89c),
	.w1(32'hbb928235),
	.w2(32'h3b5e5d91),
	.w3(32'h3aa1c67c),
	.w4(32'hbb4cff66),
	.w5(32'h3b449c37),
	.w6(32'hbc677e34),
	.w7(32'hbb0ebb27),
	.w8(32'h3b51c992),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a52c0),
	.w1(32'hbb8e3b61),
	.w2(32'hbbe9e831),
	.w3(32'h3c1787bc),
	.w4(32'h3b06d58f),
	.w5(32'hbc0de8d5),
	.w6(32'h3c1e527e),
	.w7(32'h3c13099e),
	.w8(32'h3c07b0d2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea2da4),
	.w1(32'hbb17ff70),
	.w2(32'hbb204efd),
	.w3(32'hba5388de),
	.w4(32'hbb275987),
	.w5(32'hbaf0e915),
	.w6(32'hbb9a0525),
	.w7(32'hba1cfe9d),
	.w8(32'h3a5d3495),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be9deda),
	.w1(32'h3b6d1d82),
	.w2(32'hba99fe5c),
	.w3(32'h3bc66e8c),
	.w4(32'h3bb7e6bc),
	.w5(32'h3b0c68b2),
	.w6(32'h3c3a062a),
	.w7(32'hbc0c9b28),
	.w8(32'hbb3fde91),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa41249),
	.w1(32'h3b1b2172),
	.w2(32'h3a3f7c53),
	.w3(32'h3c0b4adc),
	.w4(32'h3ac9ab65),
	.w5(32'hb9368119),
	.w6(32'h3c6e4d02),
	.w7(32'h3b6f749e),
	.w8(32'h3b0141b9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ba360),
	.w1(32'hba9fab11),
	.w2(32'hbc1cbab2),
	.w3(32'h3bea106f),
	.w4(32'hbbe67d0e),
	.w5(32'hbc899097),
	.w6(32'h3c472472),
	.w7(32'hbb48f776),
	.w8(32'hbc467bea),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f085),
	.w1(32'hbba758d8),
	.w2(32'h388d5907),
	.w3(32'hbacc7b06),
	.w4(32'hbc42571f),
	.w5(32'h3bcd229d),
	.w6(32'hba077afc),
	.w7(32'hbb98b7ea),
	.w8(32'h3bfe9e2d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1af10e),
	.w1(32'hbb93fc9c),
	.w2(32'h3b360188),
	.w3(32'h3c8bf24e),
	.w4(32'h392bd99e),
	.w5(32'h3bf1b882),
	.w6(32'h3cd20764),
	.w7(32'h3b11620f),
	.w8(32'h3bed5f79),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f2fa5),
	.w1(32'hbbc7404d),
	.w2(32'h3b24d0fb),
	.w3(32'h3b1621c2),
	.w4(32'hbbad1e20),
	.w5(32'h3a44705d),
	.w6(32'h3b3007a7),
	.w7(32'hbb3af1ea),
	.w8(32'h3b68452e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fe75f),
	.w1(32'h3a34071d),
	.w2(32'hbb0e7aba),
	.w3(32'h39cb0235),
	.w4(32'hbc275237),
	.w5(32'hbc245783),
	.w6(32'h3b212caa),
	.w7(32'h3c2b5044),
	.w8(32'h3c8629d0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0fded),
	.w1(32'h3a607cc1),
	.w2(32'h3b7ca945),
	.w3(32'hbc06c8a9),
	.w4(32'h3a4957ee),
	.w5(32'h3ace8f06),
	.w6(32'h3c9b7baa),
	.w7(32'hbb66f0f2),
	.w8(32'h3ad3c4f0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e6902),
	.w1(32'h3b13732f),
	.w2(32'h3b015695),
	.w3(32'h3b22b33d),
	.w4(32'h3adeb74d),
	.w5(32'h3b1c9862),
	.w6(32'hbb42b3c7),
	.w7(32'h3b793ffe),
	.w8(32'h3baed043),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06e9b),
	.w1(32'hbbfa86fa),
	.w2(32'hbb09fa8e),
	.w3(32'h3bfa544f),
	.w4(32'hbc396eb5),
	.w5(32'h3bdc931f),
	.w6(32'h3c2b8264),
	.w7(32'hbb1a2fe5),
	.w8(32'h3c07373b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fac846),
	.w1(32'hbb8ef8e2),
	.w2(32'h3a0a46da),
	.w3(32'h3c4c9cfb),
	.w4(32'hbb9c44b7),
	.w5(32'hba40347f),
	.w6(32'h3c421a72),
	.w7(32'h3ad96493),
	.w8(32'h3be37ea6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8aae9a),
	.w1(32'h3c106c33),
	.w2(32'h3c4e95db),
	.w3(32'h3c84ced7),
	.w4(32'h3c2c1187),
	.w5(32'h3c68f9cc),
	.w6(32'h3cb34819),
	.w7(32'h3c5bd715),
	.w8(32'h3c8752f0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc5da4),
	.w1(32'hbc1b7118),
	.w2(32'h3c21bc7b),
	.w3(32'h3b3f6b73),
	.w4(32'hbb31147d),
	.w5(32'hbaaf4791),
	.w6(32'h3b5bbd53),
	.w7(32'h3bb24402),
	.w8(32'h3b3dd601),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd24951),
	.w1(32'hbc094bed),
	.w2(32'h398bedf1),
	.w3(32'h3b37b85d),
	.w4(32'hbc19c962),
	.w5(32'hbb2ef75f),
	.w6(32'h3c1767a9),
	.w7(32'h386efe17),
	.w8(32'h3c229603),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb77172),
	.w1(32'hbbb7538c),
	.w2(32'hbaa50ec2),
	.w3(32'hbc0cad16),
	.w4(32'hbbb4fa8c),
	.w5(32'hbb13ce6f),
	.w6(32'h3a84b17a),
	.w7(32'hbb85f8a4),
	.w8(32'hbaefa397),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061709),
	.w1(32'h39880367),
	.w2(32'h3c519ea1),
	.w3(32'hbb3b445b),
	.w4(32'h3b43aa2b),
	.w5(32'h3ca97eb8),
	.w6(32'hbb182f2a),
	.w7(32'h3bdb8dcf),
	.w8(32'h3c3f61af),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc76bff),
	.w1(32'h3c003eb5),
	.w2(32'h3b66f988),
	.w3(32'h3bbd7468),
	.w4(32'h3c258dc4),
	.w5(32'h3b373fd3),
	.w6(32'h3bbbe325),
	.w7(32'h3c8872c3),
	.w8(32'hbc555372),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c441d85),
	.w1(32'h3bb8d13a),
	.w2(32'h3c5d3897),
	.w3(32'hbba4b46b),
	.w4(32'h3a7e0dd8),
	.w5(32'h3bed109f),
	.w6(32'hbcc8d07f),
	.w7(32'h3b887112),
	.w8(32'h3c4acb9c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad657af),
	.w1(32'hbb951cf6),
	.w2(32'hbbf16054),
	.w3(32'hb9bd0b7b),
	.w4(32'hbabc5b1d),
	.w5(32'hbc00bef4),
	.w6(32'h3af85ffa),
	.w7(32'hb9cc6ddb),
	.w8(32'hba944d08),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd183),
	.w1(32'hba6af540),
	.w2(32'h3b979042),
	.w3(32'h3b7f6436),
	.w4(32'hbafcbbf5),
	.w5(32'h3b997a85),
	.w6(32'h3c3ed337),
	.w7(32'h3ab30828),
	.w8(32'h3badc366),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f5ec3),
	.w1(32'hb7d7b7f5),
	.w2(32'h3b4eb419),
	.w3(32'h3b34b8ea),
	.w4(32'hb90eb1ab),
	.w5(32'h3ae631a4),
	.w6(32'h3c387113),
	.w7(32'h3aab1111),
	.w8(32'h3b45c8dc),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61242d),
	.w1(32'h3ad07522),
	.w2(32'hbc257a16),
	.w3(32'h3b7548e7),
	.w4(32'h3a8066dc),
	.w5(32'hbc234bca),
	.w6(32'h3b9491ed),
	.w7(32'h3bdbdf27),
	.w8(32'hbae70b19),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4be16),
	.w1(32'h39c045ef),
	.w2(32'h3ba6176c),
	.w3(32'h3bdae7f8),
	.w4(32'h39f5935b),
	.w5(32'h3b0aa13c),
	.w6(32'h3c02c009),
	.w7(32'h3b0c1fee),
	.w8(32'h3aeb9861),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dc7a6),
	.w1(32'h3bd4a940),
	.w2(32'h3c03d1e2),
	.w3(32'h3c4405c0),
	.w4(32'h3c075a6d),
	.w5(32'h3c3ac2e8),
	.w6(32'h3c948042),
	.w7(32'h3c94b136),
	.w8(32'h3c9bf2d5),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a604c),
	.w1(32'h3ba2a582),
	.w2(32'h3c151c2e),
	.w3(32'h3b8071fb),
	.w4(32'h3ab1f3e4),
	.w5(32'h3bd691a9),
	.w6(32'h3be12831),
	.w7(32'hb9a56022),
	.w8(32'h3b470c1b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90f25f),
	.w1(32'h3ac38257),
	.w2(32'h3723e3b2),
	.w3(32'h3bd29391),
	.w4(32'h3b06627a),
	.w5(32'h3a911cde),
	.w6(32'h3c5044f4),
	.w7(32'h3b809515),
	.w8(32'h3b87f926),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ff8464),
	.w1(32'h3ae00ccd),
	.w2(32'hb9b63a43),
	.w3(32'h3b831e86),
	.w4(32'h3a011d12),
	.w5(32'hba0e449f),
	.w6(32'h3bd9eb89),
	.w7(32'hbb940c5a),
	.w8(32'hbbb92998),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94fb4c),
	.w1(32'hbbd35698),
	.w2(32'hbb886816),
	.w3(32'h3bbdf5d0),
	.w4(32'hbbdc282a),
	.w5(32'hbc66a938),
	.w6(32'hbb66920e),
	.w7(32'hbb3f3274),
	.w8(32'hbbceac85),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d989b),
	.w1(32'h3a3f18c9),
	.w2(32'h3be66ffa),
	.w3(32'hbc157bd6),
	.w4(32'hbac1afd9),
	.w5(32'hbacc0d1d),
	.w6(32'hbaec97bf),
	.w7(32'h3bfa92e5),
	.w8(32'h3bedc335),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f445),
	.w1(32'h3b25fbd1),
	.w2(32'h3b631971),
	.w3(32'h3b286a4f),
	.w4(32'hbc33f0ad),
	.w5(32'hbbbcc2e2),
	.w6(32'hbaacc07a),
	.w7(32'h3b1cddd3),
	.w8(32'h3b171905),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e6dd),
	.w1(32'hbac5a7c0),
	.w2(32'hbc04b0f1),
	.w3(32'hbcbc6a2d),
	.w4(32'hbb8cd01a),
	.w5(32'hbc0875f5),
	.w6(32'hbbd4654f),
	.w7(32'hbb9ae21d),
	.w8(32'hbc1570e4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dc3a0),
	.w1(32'hba8aaf61),
	.w2(32'hba74370b),
	.w3(32'hbb019100),
	.w4(32'hba97a80d),
	.w5(32'h3a0170af),
	.w6(32'hbb9cc131),
	.w7(32'h3b0efbe4),
	.w8(32'h3b997350),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1fb07),
	.w1(32'h3b95700c),
	.w2(32'h3c1ecb02),
	.w3(32'h3b8b9848),
	.w4(32'h3bc47938),
	.w5(32'h3c25264d),
	.w6(32'h3c23b0f9),
	.w7(32'h3bbc21af),
	.w8(32'h3c1e6549),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39927de8),
	.w1(32'h3b078d32),
	.w2(32'h3a58fd0a),
	.w3(32'h3b34c0f4),
	.w4(32'h3b31bb7e),
	.w5(32'h396cd1c9),
	.w6(32'h3b968df2),
	.w7(32'h3b75e30d),
	.w8(32'h3a8de286),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f105d),
	.w1(32'h3a391a4f),
	.w2(32'h3adba979),
	.w3(32'h3b8c8576),
	.w4(32'hbb1d5477),
	.w5(32'hbc05f0fc),
	.w6(32'h3c01efb0),
	.w7(32'hbb72bbcf),
	.w8(32'hbc200358),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe01cd9),
	.w1(32'hbbdac823),
	.w2(32'h3bbd434f),
	.w3(32'hbc567595),
	.w4(32'hbc084c5b),
	.w5(32'h3bdba371),
	.w6(32'hbc33db96),
	.w7(32'hbc7bca35),
	.w8(32'h3c1e8d88),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cacbbda),
	.w1(32'hbb861cb2),
	.w2(32'h3a51d014),
	.w3(32'h3ca35ca3),
	.w4(32'hbb17455e),
	.w5(32'h3c188c28),
	.w6(32'h3c8f2436),
	.w7(32'h3bc24975),
	.w8(32'h3c8ffd42),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f1e83),
	.w1(32'h3abe3ea8),
	.w2(32'h3be54df6),
	.w3(32'h3bf7e0b6),
	.w4(32'hbb1fe8d5),
	.w5(32'h3b42a056),
	.w6(32'h3caf3dd8),
	.w7(32'hbc010b71),
	.w8(32'h3acaa4d8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba295153),
	.w1(32'h3ba47bcf),
	.w2(32'hbaf71da6),
	.w3(32'hbb4fe5ea),
	.w4(32'h3b0af5da),
	.w5(32'hbb87db7a),
	.w6(32'hbc81351d),
	.w7(32'hbaef7b4d),
	.w8(32'hbbe2790a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a8b61),
	.w1(32'hbb9b900c),
	.w2(32'hbbd1d00b),
	.w3(32'hbb93d718),
	.w4(32'hbb9e87c1),
	.w5(32'hbbb53821),
	.w6(32'hbbdfc092),
	.w7(32'hbb22e80f),
	.w8(32'hbb6dc292),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e374),
	.w1(32'hbb4e85fa),
	.w2(32'hbb9583c0),
	.w3(32'h3b54258a),
	.w4(32'hbb9a4007),
	.w5(32'hbc1c9eb9),
	.w6(32'h3b771235),
	.w7(32'hb9940748),
	.w8(32'hbb491815),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb108bf9),
	.w1(32'h39f930d1),
	.w2(32'h3be74b92),
	.w3(32'hbc0181a7),
	.w4(32'h3a95d55b),
	.w5(32'h3c01c1c6),
	.w6(32'hbaed4c17),
	.w7(32'h3a0ef492),
	.w8(32'h3c0f864f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90fefd),
	.w1(32'h3aaa8187),
	.w2(32'h3abdab12),
	.w3(32'h3bb51fe9),
	.w4(32'h3b33f5b2),
	.w5(32'h3b4f0940),
	.w6(32'h3c028263),
	.w7(32'h3b2f75c4),
	.w8(32'h3b2db8e5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10f63f),
	.w1(32'hbbebac98),
	.w2(32'hbbcb5229),
	.w3(32'h3a71b38f),
	.w4(32'hbc2a8980),
	.w5(32'hbb9470b3),
	.w6(32'h3b0733a4),
	.w7(32'hbb1abf55),
	.w8(32'hbb98f9c5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba420c1),
	.w1(32'hbb911a44),
	.w2(32'hbbf8e6d1),
	.w3(32'hb7e251cf),
	.w4(32'hbb25dcad),
	.w5(32'hbbbcb7c5),
	.w6(32'hbbfa5a4b),
	.w7(32'hbbfd8089),
	.w8(32'hbbf051de),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e7556),
	.w1(32'hbbacd081),
	.w2(32'hbca0c4f8),
	.w3(32'h3bdf1038),
	.w4(32'hbb417e20),
	.w5(32'hbc98f276),
	.w6(32'h3c31fc78),
	.w7(32'h3bdf41ea),
	.w8(32'h3b3e2359),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5a9f8e),
	.w1(32'h3b0caf14),
	.w2(32'h3b2ea314),
	.w3(32'hbca2cc21),
	.w4(32'h3aed42bb),
	.w5(32'h3b5b5522),
	.w6(32'hbc02d7b9),
	.w7(32'h3af65d3a),
	.w8(32'h3b869542),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca7b0),
	.w1(32'hbab3e594),
	.w2(32'hba35f720),
	.w3(32'h3b9d1089),
	.w4(32'hbb7f1924),
	.w5(32'hbb744d3e),
	.w6(32'h3ba63aca),
	.w7(32'hbaf3cb4e),
	.w8(32'hbafac9ad),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba998c36),
	.w1(32'h3b2e5a95),
	.w2(32'h3bfc8843),
	.w3(32'hbc2e833f),
	.w4(32'hbb24488f),
	.w5(32'h3b0360f5),
	.w6(32'hbc346c92),
	.w7(32'hbbfe6c86),
	.w8(32'hbac9a358),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b268f),
	.w1(32'hb9f423eb),
	.w2(32'hba949b45),
	.w3(32'hbc26af12),
	.w4(32'hb90b9884),
	.w5(32'h3a008b04),
	.w6(32'hbbfae72f),
	.w7(32'hb9e4e51f),
	.w8(32'hba2e1b33),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1038c),
	.w1(32'hbb704960),
	.w2(32'hbbd8479d),
	.w3(32'hbaaa7a67),
	.w4(32'hbaf8f927),
	.w5(32'hbbf16a6e),
	.w6(32'hbb2848ad),
	.w7(32'hbb7e408c),
	.w8(32'hbc10c234),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd6e11),
	.w1(32'hbb3b6d5f),
	.w2(32'hbc8f2bdd),
	.w3(32'h3b28152c),
	.w4(32'hbc21d459),
	.w5(32'hbca8310c),
	.w6(32'h3bcc8082),
	.w7(32'h3d268967),
	.w8(32'h3d87385e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45ea08),
	.w1(32'hbbb6d0a3),
	.w2(32'h3c128117),
	.w3(32'h3cd38670),
	.w4(32'hbb92e33c),
	.w5(32'h3bde85bc),
	.w6(32'h3e051e45),
	.w7(32'hbc280e87),
	.w8(32'h3ad780cc),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6cb85),
	.w1(32'hbaf67aa5),
	.w2(32'hbb3d4c4d),
	.w3(32'hbc17bc18),
	.w4(32'hba80b1a3),
	.w5(32'hbac96ae2),
	.w6(32'hbc485fe8),
	.w7(32'h3b360522),
	.w8(32'h3ae01e83),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b582e),
	.w1(32'hbc2120e9),
	.w2(32'hbb8bab13),
	.w3(32'h3b53814f),
	.w4(32'hbbe23276),
	.w5(32'hbb090424),
	.w6(32'h3bc717f2),
	.w7(32'h3bb68281),
	.w8(32'h3cab90fa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule