module layer_8_featuremap_84(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c14255),
	.w1(32'hb97ee2d7),
	.w2(32'hb8f9efdd),
	.w3(32'hb92759b2),
	.w4(32'hb8082f5b),
	.w5(32'h385d4cc4),
	.w6(32'h380a5b99),
	.w7(32'h3903a753),
	.w8(32'h39071ca0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa3abb),
	.w1(32'h3820ddf8),
	.w2(32'h37745400),
	.w3(32'h39b0ea16),
	.w4(32'h39273c9e),
	.w5(32'hb8d10bee),
	.w6(32'h39f24c64),
	.w7(32'h377e4223),
	.w8(32'h3950a032),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38846e65),
	.w1(32'hb9013d43),
	.w2(32'h37c1c3f5),
	.w3(32'h3a149616),
	.w4(32'h39569549),
	.w5(32'h38dda735),
	.w6(32'h3a69f499),
	.w7(32'h39c2e054),
	.w8(32'h39d24992),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35909e34),
	.w1(32'h36a1c157),
	.w2(32'h374d6ed5),
	.w3(32'hb6fd5963),
	.w4(32'h36cb1996),
	.w5(32'h37009549),
	.w6(32'hb669df32),
	.w7(32'hb4be263f),
	.w8(32'hb76cdc3b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94598d1),
	.w1(32'hb9b7ea3f),
	.w2(32'hb9b15654),
	.w3(32'hb6f35ed8),
	.w4(32'hb64b87e5),
	.w5(32'hb91b0575),
	.w6(32'h39045e19),
	.w7(32'h385d3056),
	.w8(32'hb7c02192),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ec546),
	.w1(32'hb9944816),
	.w2(32'hb9d8cf39),
	.w3(32'h398ed605),
	.w4(32'h390a51d7),
	.w5(32'h36ec9a1c),
	.w6(32'h39caedcc),
	.w7(32'h39651d7e),
	.w8(32'h38f82c84),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b4914c),
	.w1(32'h36cbf441),
	.w2(32'h37039b3d),
	.w3(32'hb72b9a80),
	.w4(32'hb664627f),
	.w5(32'hb565dc96),
	.w6(32'hb782503d),
	.w7(32'hb7121f61),
	.w8(32'hb70858a3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98a863f),
	.w1(32'hb9bc98af),
	.w2(32'hba1a7f2c),
	.w3(32'hb7eed0a7),
	.w4(32'hb9a4a9a6),
	.w5(32'hb9bf0eb4),
	.w6(32'hb7ea48b7),
	.w7(32'hb98671d2),
	.w8(32'hb9fef3bd),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8904639),
	.w1(32'hb7546c42),
	.w2(32'h389f3594),
	.w3(32'h395de463),
	.w4(32'h38b650f0),
	.w5(32'hb8ce7511),
	.w6(32'h39813419),
	.w7(32'hb80fb06c),
	.w8(32'h38cb669a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883da85),
	.w1(32'hb7bd4021),
	.w2(32'h39143627),
	.w3(32'h3a07f6b3),
	.w4(32'h38da9fc9),
	.w5(32'hb8db0075),
	.w6(32'h39edd5d5),
	.w7(32'h3882249f),
	.w8(32'h39b4c551),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915ce35),
	.w1(32'hb9e666d0),
	.w2(32'hb9bf76df),
	.w3(32'hb8e0acc9),
	.w4(32'h391d308d),
	.w5(32'h3954224b),
	.w6(32'h39bd019d),
	.w7(32'h39e972a1),
	.w8(32'h39b1bf6f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d128bc),
	.w1(32'hb9393560),
	.w2(32'hb949f2c5),
	.w3(32'h38360e99),
	.w4(32'hb8145f94),
	.w5(32'hb7930f12),
	.w6(32'h38cbd979),
	.w7(32'h388373d4),
	.w8(32'h3889db2f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bbee1),
	.w1(32'hb96dd982),
	.w2(32'hb980c2d6),
	.w3(32'h399f1f18),
	.w4(32'h37a50a0f),
	.w5(32'hb8d6e866),
	.w6(32'h39dd5a50),
	.w7(32'h3840be56),
	.w8(32'h38b75b61),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6336ac8),
	.w1(32'h36ad5733),
	.w2(32'h370c3cfb),
	.w3(32'hb787ddd0),
	.w4(32'hb6cfffc1),
	.w5(32'hb70a85b5),
	.w6(32'hb7d35ef6),
	.w7(32'hb793bfe0),
	.w8(32'hb771be51),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362f86f2),
	.w1(32'h36ed9fbd),
	.w2(32'h370977da),
	.w3(32'hb6bd6ec8),
	.w4(32'h3563f505),
	.w5(32'h35ea9398),
	.w6(32'hb72ad7dc),
	.w7(32'hb6ae7a15),
	.w8(32'hb6abfcac),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370f3a95),
	.w1(32'h375a2659),
	.w2(32'h3742081c),
	.w3(32'hb755dd8b),
	.w4(32'hb68f4161),
	.w5(32'hb56deac9),
	.w6(32'hb7724899),
	.w7(32'hb6bd5990),
	.w8(32'hb63d4fa8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394eea59),
	.w1(32'hb96c21de),
	.w2(32'hb91819ed),
	.w3(32'h38ae907f),
	.w4(32'hb8bc8fda),
	.w5(32'hb91184c6),
	.w6(32'h38ec0c47),
	.w7(32'h3885eda0),
	.w8(32'h39c0ec2e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a14dec),
	.w1(32'hb991019a),
	.w2(32'hb992fe63),
	.w3(32'h3a13e050),
	.w4(32'h390295b2),
	.w5(32'hb88c0e28),
	.w6(32'h3a1a6c50),
	.w7(32'h39632031),
	.w8(32'h390b3976),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac06715),
	.w1(32'hbb13370e),
	.w2(32'hbaa9ad7e),
	.w3(32'hba4c4d27),
	.w4(32'h39dcf9ac),
	.w5(32'h3945191c),
	.w6(32'h3a73560e),
	.w7(32'h3ab8518c),
	.w8(32'h39737bb1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdd93f),
	.w1(32'hba49f42a),
	.w2(32'hba2c7547),
	.w3(32'h39faf5e1),
	.w4(32'h38989168),
	.w5(32'h39149143),
	.w6(32'h3a8db075),
	.w7(32'h3a46e01d),
	.w8(32'h3a575a33),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98decf4),
	.w1(32'hb947ec6f),
	.w2(32'hb9bd84ad),
	.w3(32'hb84c4b2a),
	.w4(32'h39648f0e),
	.w5(32'hb7d90d0e),
	.w6(32'hb97fe3d6),
	.w7(32'hb8f7feda),
	.w8(32'hb99a0e9e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac4599),
	.w1(32'hb83bd6b1),
	.w2(32'h38de5b0d),
	.w3(32'h3a1cd1b3),
	.w4(32'h39173a02),
	.w5(32'hb79d56e9),
	.w6(32'h3a6beade),
	.w7(32'h395e0508),
	.w8(32'h39aa5501),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab91ca1),
	.w1(32'hbb165448),
	.w2(32'hbaec2b24),
	.w3(32'hbaafc024),
	.w4(32'hba8574b8),
	.w5(32'hb96eb40c),
	.w6(32'hb9970894),
	.w7(32'h397998d0),
	.w8(32'hb99304b8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3888bcfd),
	.w1(32'hb8d752f9),
	.w2(32'hb8598cb1),
	.w3(32'h39774b85),
	.w4(32'h38993f57),
	.w5(32'hb983209e),
	.w6(32'h3998f826),
	.w7(32'hb7e3a7b1),
	.w8(32'h398588a3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64d05e4),
	.w1(32'h36ad58a0),
	.w2(32'h3700c5f8),
	.w3(32'hb753b833),
	.w4(32'hb7a75e1c),
	.w5(32'hb7a5939e),
	.w6(32'hb7b4f569),
	.w7(32'hb7cecb04),
	.w8(32'hb7833200),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2896ca),
	.w1(32'hba831dad),
	.w2(32'hba3e0e46),
	.w3(32'hba01c181),
	.w4(32'hb98fbd5e),
	.w5(32'h38cba399),
	.w6(32'hb73c6d12),
	.w7(32'h394c6cc1),
	.w8(32'h38b427d2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374dc55c),
	.w1(32'h374df4de),
	.w2(32'h375f6d9d),
	.w3(32'h36e483d9),
	.w4(32'h36b0d359),
	.w5(32'h36f8aa3f),
	.w6(32'hb5daf3a6),
	.w7(32'h36419635),
	.w8(32'h362f298e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65f5be),
	.w1(32'hbc00b91a),
	.w2(32'hbc3251f7),
	.w3(32'hbb3338a1),
	.w4(32'hbbc8d617),
	.w5(32'h3bb96b5d),
	.w6(32'hbb41e672),
	.w7(32'h3b7c35af),
	.w8(32'h3b082a2e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca83f0),
	.w1(32'hba269cb0),
	.w2(32'hba0ab3c2),
	.w3(32'hb9713961),
	.w4(32'hb8596c53),
	.w5(32'h382f9432),
	.w6(32'h39424a67),
	.w7(32'h398ae5bf),
	.w8(32'h391fe1fe),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f7ad52),
	.w1(32'hb92bd98a),
	.w2(32'hb91866fc),
	.w3(32'h383dd451),
	.w4(32'hb8640116),
	.w5(32'hb88d0992),
	.w6(32'h39006c9b),
	.w7(32'h36ed67eb),
	.w8(32'h36445503),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8556086),
	.w1(32'hb88c3048),
	.w2(32'hb7a77c3c),
	.w3(32'h369de67f),
	.w4(32'hb69f2da2),
	.w5(32'h380cb636),
	.w6(32'h381ac59d),
	.w7(32'h38ae1625),
	.w8(32'h388502af),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1bc38),
	.w1(32'hb9012257),
	.w2(32'hb9830ab7),
	.w3(32'h37ee5417),
	.w4(32'hb8f7ee4b),
	.w5(32'hb8b485ac),
	.w6(32'h388a403d),
	.w7(32'h38ce96be),
	.w8(32'h3947d713),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371146ee),
	.w1(32'h3791d584),
	.w2(32'h378abc2b),
	.w3(32'hb744a43a),
	.w4(32'hb47717a1),
	.w5(32'h356642da),
	.w6(32'hb7c94fb5),
	.w7(32'hb7743e3e),
	.w8(32'hb724b39c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36da0994),
	.w1(32'h377bc677),
	.w2(32'h378921c0),
	.w3(32'hb72608c8),
	.w4(32'hb54ecd69),
	.w5(32'h349479b9),
	.w6(32'hb77542fa),
	.w7(32'hb6c17593),
	.w8(32'hb72e8082),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903958f),
	.w1(32'h393fc594),
	.w2(32'h39ad9ea1),
	.w3(32'h3a019d3b),
	.w4(32'h38ef1dfc),
	.w5(32'h37ec577d),
	.w6(32'h3a0111af),
	.w7(32'h38d62be8),
	.w8(32'h39c1845c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b84752),
	.w1(32'hba29c35b),
	.w2(32'hb9a60023),
	.w3(32'hb91083c2),
	.w4(32'hb8c49035),
	.w5(32'h39011908),
	.w6(32'h392ea821),
	.w7(32'h38d8dd99),
	.w8(32'hb95c3546),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355639cf),
	.w1(32'h369d1e92),
	.w2(32'h36ab033f),
	.w3(32'hb729f390),
	.w4(32'hb5ee2817),
	.w5(32'hb525e330),
	.w6(32'hb732af1c),
	.w7(32'hb6dd8417),
	.w8(32'hb6fcb393),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9305301),
	.w1(32'hb909cf36),
	.w2(32'h37c37c18),
	.w3(32'h36e9dd9f),
	.w4(32'hb82563f2),
	.w5(32'hb949691b),
	.w6(32'h3918f271),
	.w7(32'hb8f3c525),
	.w8(32'hb981b89f),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37562b3d),
	.w1(32'h37cdf6b1),
	.w2(32'h37c855f0),
	.w3(32'hb722c88d),
	.w4(32'h3603aac2),
	.w5(32'h3674700f),
	.w6(32'hb7db1d48),
	.w7(32'hb7846034),
	.w8(32'hb723673d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c030b),
	.w1(32'h37af09cd),
	.w2(32'h37784d2a),
	.w3(32'hb755bb1e),
	.w4(32'hb64e447d),
	.w5(32'h361647e3),
	.w6(32'hb7cd132e),
	.w7(32'hb711e6f8),
	.w8(32'hb71ce5f3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c5247),
	.w1(32'hba3c6439),
	.w2(32'hb9e2587e),
	.w3(32'h398bb101),
	.w4(32'h388120b5),
	.w5(32'hb8d2f6e5),
	.w6(32'h3a097701),
	.w7(32'hb9156c51),
	.w8(32'h38ee45c4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc6057),
	.w1(32'h383de5d8),
	.w2(32'h384cd8d6),
	.w3(32'hb91d06b1),
	.w4(32'hb7801306),
	.w5(32'h3925c4b4),
	.w6(32'hba1cb96f),
	.w7(32'hba8d69bd),
	.w8(32'hb8cd143c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d552f),
	.w1(32'hbb00d5cd),
	.w2(32'h3aca2c9e),
	.w3(32'hba2e79ec),
	.w4(32'hbaa3772c),
	.w5(32'hbb0dda1f),
	.w6(32'h3b0bce10),
	.w7(32'h3af60b77),
	.w8(32'hb9b61533),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20de8b),
	.w1(32'hb9ef518b),
	.w2(32'hb9af72ff),
	.w3(32'hba566756),
	.w4(32'hb9bafbc6),
	.w5(32'h37b51c46),
	.w6(32'hba1417e9),
	.w7(32'hba45f8b4),
	.w8(32'h3934ae91),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d55ee),
	.w1(32'hbaeaa264),
	.w2(32'hbab26d43),
	.w3(32'hba748092),
	.w4(32'hb9af3459),
	.w5(32'hb8aceb22),
	.w6(32'hba41b99a),
	.w7(32'h38c67ebf),
	.w8(32'h3ab4219c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f6459),
	.w1(32'hba0e7d2e),
	.w2(32'h3a6cf0b3),
	.w3(32'h39d32e49),
	.w4(32'h38c78306),
	.w5(32'h3a5a3bbd),
	.w6(32'h3901431b),
	.w7(32'hb8d24587),
	.w8(32'hbb95b9e6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec8c4f),
	.w1(32'hbbcb40b9),
	.w2(32'hbb09a494),
	.w3(32'hbbb547e2),
	.w4(32'hbb332fa7),
	.w5(32'hbbc4a14d),
	.w6(32'hbaabb08e),
	.w7(32'hb9c1de85),
	.w8(32'hb297e195),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec56b6),
	.w1(32'hb7e61dd4),
	.w2(32'h3a72a6ec),
	.w3(32'h38129431),
	.w4(32'h3a660c2c),
	.w5(32'h3a920773),
	.w6(32'h396c750d),
	.w7(32'h3a2b3309),
	.w8(32'h37c9130b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857ed37),
	.w1(32'hbaa4b2d5),
	.w2(32'hb9b16e72),
	.w3(32'hb9162fe7),
	.w4(32'hbac35e8d),
	.w5(32'hb98e6250),
	.w6(32'h3802fc32),
	.w7(32'h39b51a3e),
	.w8(32'h39d03ac5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96f8d1),
	.w1(32'hbaa8dff6),
	.w2(32'hb9d7676e),
	.w3(32'hba643f77),
	.w4(32'hba09096a),
	.w5(32'hb7f1d1ab),
	.w6(32'hba45664d),
	.w7(32'hb9f2527a),
	.w8(32'h39c8c523),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a34d53),
	.w1(32'hb8a043af),
	.w2(32'hb8bf9a4d),
	.w3(32'hb92f5f9a),
	.w4(32'hb90b263f),
	.w5(32'h391a9ffb),
	.w6(32'hb9bec295),
	.w7(32'hb993ce65),
	.w8(32'h3a69020e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb194e),
	.w1(32'hbb87bd1a),
	.w2(32'hbb4afa00),
	.w3(32'hbaf214d4),
	.w4(32'hba9d9fde),
	.w5(32'hb9906319),
	.w6(32'hb9a4403e),
	.w7(32'h39825602),
	.w8(32'h3b4254b3),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92713d),
	.w1(32'hbb87c4c8),
	.w2(32'hbb7a5b2c),
	.w3(32'h3b488b36),
	.w4(32'hbb7922b6),
	.w5(32'hbb9b9799),
	.w6(32'hba897f0c),
	.w7(32'h3a395103),
	.w8(32'h3abb480d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddb065),
	.w1(32'hba98346a),
	.w2(32'hbabc2263),
	.w3(32'hb818cce0),
	.w4(32'hba0dec55),
	.w5(32'hb8fec5df),
	.w6(32'h3969c864),
	.w7(32'hb9dcbe2e),
	.w8(32'h3a886437),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2da66),
	.w1(32'hbb0760d1),
	.w2(32'hbb3bb29b),
	.w3(32'hba5e8267),
	.w4(32'hbb356575),
	.w5(32'hbbc16176),
	.w6(32'h3b2442b8),
	.w7(32'hb9fe0889),
	.w8(32'h3ad699f7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a112e35),
	.w1(32'hbb996ca8),
	.w2(32'hba9f4aea),
	.w3(32'hb9ff08a7),
	.w4(32'hbbaa9cb8),
	.w5(32'hbad076b1),
	.w6(32'h3b01b0fb),
	.w7(32'h3b48ac18),
	.w8(32'hbafaeb11),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00cfa4),
	.w1(32'hbadbd392),
	.w2(32'hbaa68b84),
	.w3(32'hbaa9727d),
	.w4(32'hbb0f2fb2),
	.w5(32'hbb081c48),
	.w6(32'h3acdc76e),
	.w7(32'hba197edb),
	.w8(32'hba7ed816),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7aeda),
	.w1(32'hb9918aa0),
	.w2(32'hbb47b9ca),
	.w3(32'h3a732eae),
	.w4(32'h39558264),
	.w5(32'hbb403f43),
	.w6(32'h39dbc12d),
	.w7(32'hbb29e261),
	.w8(32'hb8d78b37),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e1447d),
	.w1(32'h39afd004),
	.w2(32'h3ab193ad),
	.w3(32'hba8129f5),
	.w4(32'hba95401a),
	.w5(32'h3a3743be),
	.w6(32'h3a583070),
	.w7(32'h3b20506f),
	.w8(32'hb9b826b9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0e3ce),
	.w1(32'hbaa21405),
	.w2(32'hba1e2aa6),
	.w3(32'h39e8b1e6),
	.w4(32'hb9a48dc7),
	.w5(32'hba50baa6),
	.w6(32'hba048292),
	.w7(32'hba53f5de),
	.w8(32'h3b11e3d1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacec31f),
	.w1(32'hbb81ec2c),
	.w2(32'h3ba174c5),
	.w3(32'hbb3fc6fb),
	.w4(32'h3a096d8d),
	.w5(32'h3a32a222),
	.w6(32'h3b977f49),
	.w7(32'h3b2703b8),
	.w8(32'h3a1bae95),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b935c8),
	.w1(32'hb9cbc2ff),
	.w2(32'h3a301ead),
	.w3(32'h3b01a72d),
	.w4(32'h3a33b1e7),
	.w5(32'h3a21fb60),
	.w6(32'h3a3b5136),
	.w7(32'h36204d83),
	.w8(32'h3aac91a7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f37c9),
	.w1(32'hba3b4832),
	.w2(32'hba087713),
	.w3(32'h3a4c8b45),
	.w4(32'h39d72457),
	.w5(32'h3a8c9605),
	.w6(32'h3a0b71af),
	.w7(32'h3a1ac118),
	.w8(32'hbb06d1d1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba494cda),
	.w1(32'h3a67b262),
	.w2(32'hbb194370),
	.w3(32'h3b433ef7),
	.w4(32'h3ba1af53),
	.w5(32'h397148c4),
	.w6(32'hba8a5d68),
	.w7(32'h3aa3bcee),
	.w8(32'hba2b863f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e0f20),
	.w1(32'hba8c5ff0),
	.w2(32'hb9e8dbf6),
	.w3(32'hba895904),
	.w4(32'hba058e14),
	.w5(32'hb910cf47),
	.w6(32'hba8c363c),
	.w7(32'hba4d309e),
	.w8(32'hb97528b1),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03c6d7),
	.w1(32'hba0f570c),
	.w2(32'hb9d0be5c),
	.w3(32'hb9a2b52c),
	.w4(32'hb94865c1),
	.w5(32'hb836af62),
	.w6(32'h38f58290),
	.w7(32'hb9ddb2da),
	.w8(32'h3a08917a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364f5316),
	.w1(32'hba2f742b),
	.w2(32'hba13e722),
	.w3(32'hb839e597),
	.w4(32'hb97c06ec),
	.w5(32'hb7067418),
	.w6(32'h38baf1cd),
	.w7(32'hb95ca831),
	.w8(32'hbab9ec35),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb009a1c),
	.w1(32'h3aad5b48),
	.w2(32'h3a775a31),
	.w3(32'h3acdd84a),
	.w4(32'h3af701e1),
	.w5(32'h3a9a4a87),
	.w6(32'hb962504b),
	.w7(32'h37c52945),
	.w8(32'h39ce10b1),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0a657),
	.w1(32'hba2c9c3b),
	.w2(32'hb941252b),
	.w3(32'hb9606635),
	.w4(32'hb986efd8),
	.w5(32'h38a1cf87),
	.w6(32'hba0fd3f6),
	.w7(32'hb9ba0af9),
	.w8(32'h3a72b684),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a4abab),
	.w1(32'h3a72e1d7),
	.w2(32'h3b079ade),
	.w3(32'hbab2dfc0),
	.w4(32'hb9995b74),
	.w5(32'h3aeeedf8),
	.w6(32'h3ade9441),
	.w7(32'h3b8ace6e),
	.w8(32'h3a413973),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a7e09),
	.w1(32'hb96ded83),
	.w2(32'hba081e51),
	.w3(32'hba0c847a),
	.w4(32'hb87c5e9f),
	.w5(32'h39689987),
	.w6(32'hba800572),
	.w7(32'hba88ee01),
	.w8(32'h39bdf6e7),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edbbbb),
	.w1(32'hba497c01),
	.w2(32'hb9e43fe3),
	.w3(32'h38c9cee4),
	.w4(32'hb9c19364),
	.w5(32'h381303d0),
	.w6(32'hb93dcdbb),
	.w7(32'hb76b9975),
	.w8(32'h3a0f17d1),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9016e13),
	.w1(32'hba4a52bd),
	.w2(32'hba855d7d),
	.w3(32'hba040a29),
	.w4(32'hb9f836e8),
	.w5(32'hb929bc0b),
	.w6(32'hbaa63b87),
	.w7(32'hbab60f21),
	.w8(32'hbb9a22cf),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef6139),
	.w1(32'h3b8095dc),
	.w2(32'hbb79f22b),
	.w3(32'hba96b927),
	.w4(32'h3a208d9d),
	.w5(32'h39aa7f98),
	.w6(32'hbbdeceb1),
	.w7(32'hbb1142bb),
	.w8(32'h3ab497f8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a0ecf),
	.w1(32'h37df3b99),
	.w2(32'h390529ed),
	.w3(32'h3a9e0fde),
	.w4(32'h3a34a060),
	.w5(32'h39ea3f19),
	.w6(32'h38997e13),
	.w7(32'h3980dfa3),
	.w8(32'hb6ae7391),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba511abb),
	.w1(32'hbab46495),
	.w2(32'hba98f629),
	.w3(32'hba3c6e44),
	.w4(32'hb656e904),
	.w5(32'h3829f37f),
	.w6(32'h396def80),
	.w7(32'hb9a5b103),
	.w8(32'h391853a1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a79b8),
	.w1(32'h38528eb1),
	.w2(32'h38b61eae),
	.w3(32'h39b9df3c),
	.w4(32'h39821580),
	.w5(32'h39b1648a),
	.w6(32'hb96e68e7),
	.w7(32'hb9c7190a),
	.w8(32'h3a8c0bfa),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f39c45),
	.w1(32'h3af5e527),
	.w2(32'h3b59aedc),
	.w3(32'hbad1ad43),
	.w4(32'hb9d523c5),
	.w5(32'h3aa0d404),
	.w6(32'h3affb72c),
	.w7(32'h3b7af49c),
	.w8(32'h39ff72c0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907eccb),
	.w1(32'h3aa8aff1),
	.w2(32'h3aaa6aa5),
	.w3(32'hba865e4a),
	.w4(32'hb839f4b5),
	.w5(32'h399c3d1d),
	.w6(32'h38f34cd4),
	.w7(32'h3a2a3df7),
	.w8(32'hba8d9899),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84ac20),
	.w1(32'hb9d6b1f4),
	.w2(32'hb9c5464e),
	.w3(32'hba16e486),
	.w4(32'hb96b00ba),
	.w5(32'h388edee7),
	.w6(32'hba2967cc),
	.w7(32'hb90b7ec4),
	.w8(32'hba28910a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa228ba),
	.w1(32'h3b4eb384),
	.w2(32'h3b014da9),
	.w3(32'hb9f66d52),
	.w4(32'h3b4e1c4a),
	.w5(32'h3afe4b26),
	.w6(32'h3b6ce6d3),
	.w7(32'h3b55fbec),
	.w8(32'h3a603a2b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a31575a),
	.w1(32'hb9c7055a),
	.w2(32'h38c2bfb5),
	.w3(32'h3a9d7f39),
	.w4(32'h3a76b994),
	.w5(32'h3a3d20e8),
	.w6(32'h3a1f4321),
	.w7(32'h39cec0d8),
	.w8(32'h3a6aa7cd),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a2e88),
	.w1(32'hba6e8304),
	.w2(32'hb7b70041),
	.w3(32'hb9933d17),
	.w4(32'hb995b0ac),
	.w5(32'h396ff22f),
	.w6(32'h3a478442),
	.w7(32'h3a4f246d),
	.w8(32'hbb19315b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a20df),
	.w1(32'hbc31fe6a),
	.w2(32'hbc07d21f),
	.w3(32'hbb512938),
	.w4(32'hbbecb0ce),
	.w5(32'hbbd43b3d),
	.w6(32'h3abb7c80),
	.w7(32'hbb1a8ab4),
	.w8(32'h3a855934),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bfc284),
	.w1(32'hba486833),
	.w2(32'hba10b79a),
	.w3(32'h3a43abcc),
	.w4(32'h3a530a39),
	.w5(32'h3aca1ee9),
	.w6(32'h3930df9a),
	.w7(32'h3a06cb8f),
	.w8(32'h3a333318),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3788cb22),
	.w1(32'hba837a94),
	.w2(32'hba4350da),
	.w3(32'hb9b2fea9),
	.w4(32'hb9667be9),
	.w5(32'hb8aa58c1),
	.w6(32'hba1ee203),
	.w7(32'hba114372),
	.w8(32'hb97dde5a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7112c),
	.w1(32'hba8a7d49),
	.w2(32'h392cbc1b),
	.w3(32'hb97dacc7),
	.w4(32'hbaf22e74),
	.w5(32'hb97d997f),
	.w6(32'hb9b456a4),
	.w7(32'h39564546),
	.w8(32'hb9d3c962),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac49765),
	.w1(32'hba8f2f16),
	.w2(32'hb83d73f1),
	.w3(32'hba64a92a),
	.w4(32'hba62bbf2),
	.w5(32'hba0207f1),
	.w6(32'hba8ba2cb),
	.w7(32'hba177363),
	.w8(32'hbac827a8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397fe277),
	.w1(32'hb848f529),
	.w2(32'hba6dfe64),
	.w3(32'h3afdf0c5),
	.w4(32'h3b24a00e),
	.w5(32'h3a85cbfe),
	.w6(32'hb98fec31),
	.w7(32'hb9bcc45d),
	.w8(32'hb9be43e4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a408724),
	.w1(32'hba77d645),
	.w2(32'h39bd3416),
	.w3(32'hb9a474f9),
	.w4(32'hbad16f54),
	.w5(32'h38e32a4f),
	.w6(32'hb98ab3f2),
	.w7(32'h3a04e010),
	.w8(32'hb8cea471),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39097d32),
	.w1(32'hbaafc3b4),
	.w2(32'hb9bd1771),
	.w3(32'hb97a6f99),
	.w4(32'hbacbdfd2),
	.w5(32'hb9438859),
	.w6(32'hb98584f0),
	.w7(32'h39c0e3ed),
	.w8(32'h39c9478c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd94ef),
	.w1(32'hba3b7a1f),
	.w2(32'hba4ddde8),
	.w3(32'h38121982),
	.w4(32'h391be693),
	.w5(32'h38bf1947),
	.w6(32'hba300eb0),
	.w7(32'hba8ae2e8),
	.w8(32'hbb26b24d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010050),
	.w1(32'hbb6b104d),
	.w2(32'hbb9fc98a),
	.w3(32'hbbc51cd6),
	.w4(32'hbb956fdb),
	.w5(32'hbbd4dd9c),
	.w6(32'hbaf7fbce),
	.w7(32'hba815bd0),
	.w8(32'h38ae6014),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372bc70e),
	.w1(32'hb988c094),
	.w2(32'hb98ef74f),
	.w3(32'h3902abfc),
	.w4(32'h3785d5e3),
	.w5(32'h391fdf39),
	.w6(32'h394555fe),
	.w7(32'h37b04075),
	.w8(32'hbb07c22a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb777983),
	.w1(32'hbafd6dc4),
	.w2(32'hbaed82bc),
	.w3(32'hba4f6a39),
	.w4(32'hba9370ad),
	.w5(32'hbb3f7c47),
	.w6(32'hb971f9f3),
	.w7(32'hba73050a),
	.w8(32'h38e89920),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2642a),
	.w1(32'hb97bc960),
	.w2(32'hb9d17ccd),
	.w3(32'h3acbdf46),
	.w4(32'h3b4065d6),
	.w5(32'h3b5dde94),
	.w6(32'hba54be4d),
	.w7(32'hba383b26),
	.w8(32'hbb44557d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205178),
	.w1(32'h3aaa1e1e),
	.w2(32'h39d8ee5e),
	.w3(32'hbac255ab),
	.w4(32'h3a520921),
	.w5(32'hba953043),
	.w6(32'hbb261d85),
	.w7(32'hbb7964e8),
	.w8(32'h39cc43ad),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a48a3),
	.w1(32'hbbcc8dd9),
	.w2(32'hbb1bf59d),
	.w3(32'h3a933ef4),
	.w4(32'hbb21122c),
	.w5(32'hbafd54fc),
	.w6(32'h3b853999),
	.w7(32'h3b6a142f),
	.w8(32'h3a742ece),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398436db),
	.w1(32'h3b086304),
	.w2(32'h3b4edf2f),
	.w3(32'hbaaa9301),
	.w4(32'hb9eb4610),
	.w5(32'h3a6c1630),
	.w6(32'h3abc8f1c),
	.w7(32'h3b42edbc),
	.w8(32'hb99c1769),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba708ee3),
	.w1(32'hba1b15b2),
	.w2(32'hb799a857),
	.w3(32'hb9d38baa),
	.w4(32'hb90bd5ad),
	.w5(32'hb92774cf),
	.w6(32'hb9cc5529),
	.w7(32'hba39b853),
	.w8(32'hb8a690e4),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a440f81),
	.w1(32'hbabc2c67),
	.w2(32'hbabc2bc6),
	.w3(32'h39fea1a4),
	.w4(32'h39dbfbca),
	.w5(32'hba409b42),
	.w6(32'hb93ba02b),
	.w7(32'hbacd4e5f),
	.w8(32'h3a4d09b0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0952d6),
	.w1(32'h388d9733),
	.w2(32'h396fe865),
	.w3(32'h399315f8),
	.w4(32'h39b3f3b0),
	.w5(32'h39ca41e8),
	.w6(32'h3927a509),
	.w7(32'hb8880908),
	.w8(32'h3a4325a4),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cc136f),
	.w1(32'h3b4c0732),
	.w2(32'h3b39f378),
	.w3(32'hbaa7541f),
	.w4(32'h3a52be0a),
	.w5(32'h3a96af2c),
	.w6(32'h39d0f33a),
	.w7(32'h3ab4437a),
	.w8(32'h389eee46),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d0bb6),
	.w1(32'hb8829644),
	.w2(32'hb9a23238),
	.w3(32'h3a95d7c6),
	.w4(32'h3a9f57ce),
	.w5(32'h3a9b6985),
	.w6(32'h39cea4fc),
	.w7(32'hba2cac13),
	.w8(32'h38245294),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3840e8ce),
	.w1(32'hba10fd92),
	.w2(32'hb979f441),
	.w3(32'hb83a246e),
	.w4(32'hba5c0e94),
	.w5(32'hb99b22e1),
	.w6(32'hb95c016f),
	.w7(32'hb8958e62),
	.w8(32'hb91df13b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80442cd),
	.w1(32'hba09e609),
	.w2(32'hba015e04),
	.w3(32'hb9338c1f),
	.w4(32'hb91e2bc1),
	.w5(32'h391f8ea7),
	.w6(32'h399ce6ff),
	.w7(32'h3ab61407),
	.w8(32'hba1b2242),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1584d3),
	.w1(32'hbb0e4a28),
	.w2(32'h3ac80a86),
	.w3(32'hbacf89cf),
	.w4(32'hba948ff8),
	.w5(32'h39fc00b9),
	.w6(32'h3a9aff79),
	.w7(32'h3a71816a),
	.w8(32'hb8949ea9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0171aa),
	.w1(32'h39a7b3f7),
	.w2(32'h38f29ea4),
	.w3(32'h3a310463),
	.w4(32'h38a14a7e),
	.w5(32'hb9a96272),
	.w6(32'h39c9447f),
	.w7(32'h3a45679d),
	.w8(32'h3a17ea01),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74db63),
	.w1(32'h3a23b649),
	.w2(32'h3a654e06),
	.w3(32'h3a516bdc),
	.w4(32'h3985af79),
	.w5(32'h39a14ef1),
	.w6(32'h39b6e8d4),
	.w7(32'h3a81b1d7),
	.w8(32'hb919f9a9),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38724b1c),
	.w1(32'hbaf200c8),
	.w2(32'hbacadb79),
	.w3(32'hba75cf1c),
	.w4(32'hba8e0e1a),
	.w5(32'hba9b5fe1),
	.w6(32'hba341aac),
	.w7(32'hba2d8ce4),
	.w8(32'hbb60cfae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae61795),
	.w1(32'h398b781c),
	.w2(32'hbb0c7aad),
	.w3(32'hbb1dc7b0),
	.w4(32'h3b19f661),
	.w5(32'h3a9ae876),
	.w6(32'hba5c772a),
	.w7(32'hbb419353),
	.w8(32'hba13f650),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd8560),
	.w1(32'hbb64fbbd),
	.w2(32'hbabc66e4),
	.w3(32'hba0f6383),
	.w4(32'hbb0d4242),
	.w5(32'hba958cb8),
	.w6(32'hba93cfe4),
	.w7(32'hba279eff),
	.w8(32'h3971d0c6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61fb87),
	.w1(32'hba970c49),
	.w2(32'hb96452be),
	.w3(32'hba3617ec),
	.w4(32'hba6ae013),
	.w5(32'h39637b28),
	.w6(32'hba015f0b),
	.w7(32'h379d5f07),
	.w8(32'h3a0952e2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8efe2d),
	.w1(32'h3a01efc3),
	.w2(32'h3a64fcd9),
	.w3(32'h3a5917cd),
	.w4(32'h399935c4),
	.w5(32'h3a1d1aa5),
	.w6(32'h396f8199),
	.w7(32'h3a8ec773),
	.w8(32'hb9c813eb),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc6fe7),
	.w1(32'hb8ddb6f6),
	.w2(32'h37ca7923),
	.w3(32'h387fa0d7),
	.w4(32'hb93e841c),
	.w5(32'hb9a58cc2),
	.w6(32'hb9a1cf80),
	.w7(32'h38100cae),
	.w8(32'hba133114),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c799ab),
	.w1(32'h397da281),
	.w2(32'h3994c9bb),
	.w3(32'h39c2d6b4),
	.w4(32'h386fd091),
	.w5(32'hb9525084),
	.w6(32'hb9aea0f9),
	.w7(32'h3a0ea6e1),
	.w8(32'h3a4ca386),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad396c5),
	.w1(32'hba9e3156),
	.w2(32'hba86094c),
	.w3(32'h3a6df74c),
	.w4(32'hba276a14),
	.w5(32'hb9609a68),
	.w6(32'h3b19c9b4),
	.w7(32'h397c52f4),
	.w8(32'h397445fc),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de1d52),
	.w1(32'hba2f4313),
	.w2(32'h35b9d788),
	.w3(32'h3a03ce49),
	.w4(32'hb9bb6048),
	.w5(32'h39d3ca16),
	.w6(32'h3838127b),
	.w7(32'h3a94d5e5),
	.w8(32'h3b3b6979),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180e53),
	.w1(32'hba6593a8),
	.w2(32'hbab94dc0),
	.w3(32'h3a941ade),
	.w4(32'h3b267bcf),
	.w5(32'h39899c4a),
	.w6(32'h3a744d46),
	.w7(32'hbaeb8c67),
	.w8(32'hbb25907d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29ad2f),
	.w1(32'hbb3e4207),
	.w2(32'hbb3feeaa),
	.w3(32'hbb48b9ae),
	.w4(32'hbb065555),
	.w5(32'hbb0176b0),
	.w6(32'hbb4b7414),
	.w7(32'hbb337f8b),
	.w8(32'h389b4737),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807e604),
	.w1(32'hb9537d5d),
	.w2(32'hbab8f610),
	.w3(32'h38508b59),
	.w4(32'hbaddeb03),
	.w5(32'h3886d9a1),
	.w6(32'h3952cc8a),
	.w7(32'hba206913),
	.w8(32'h3ad2686b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae94d90),
	.w1(32'hbb24ee8e),
	.w2(32'h38dbcc02),
	.w3(32'h3931c141),
	.w4(32'h391d7c8f),
	.w5(32'hb980d6cc),
	.w6(32'h3ab3ab29),
	.w7(32'hba6301d9),
	.w8(32'h38b08899),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39881ef3),
	.w1(32'h3991e489),
	.w2(32'h3a1a8ec8),
	.w3(32'h39964a1e),
	.w4(32'h39295d95),
	.w5(32'h39f47fd5),
	.w6(32'h3a29e609),
	.w7(32'h3a974d03),
	.w8(32'hb9af0c48),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9543eb4),
	.w1(32'h396db0df),
	.w2(32'hba90e8e0),
	.w3(32'hba55c72d),
	.w4(32'hba6a8342),
	.w5(32'hb99c3a73),
	.w6(32'hba916eda),
	.w7(32'hbac0579a),
	.w8(32'hba5b3da5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84bba8),
	.w1(32'hba25480a),
	.w2(32'hbbaf82dc),
	.w3(32'hbb7c1400),
	.w4(32'hbad11ba8),
	.w5(32'hbaab83a6),
	.w6(32'hbb1079fd),
	.w7(32'hbb46fb96),
	.w8(32'hb9cde44a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83a22b),
	.w1(32'hba8ee6da),
	.w2(32'hba2d13da),
	.w3(32'hb935b45d),
	.w4(32'hba21ef48),
	.w5(32'h38717ddd),
	.w6(32'hbab7923b),
	.w7(32'hba3e0225),
	.w8(32'h3a35c031),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9361eb),
	.w1(32'h3a59394a),
	.w2(32'h3a306cb0),
	.w3(32'h3ace274a),
	.w4(32'h3a0da854),
	.w5(32'hb7b1c66a),
	.w6(32'h3a9c0870),
	.w7(32'h3abc464f),
	.w8(32'hb93a5872),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5baba),
	.w1(32'hbb891063),
	.w2(32'h3ae425de),
	.w3(32'hbb268233),
	.w4(32'hbb74aa7e),
	.w5(32'hbb1287b8),
	.w6(32'h3a9a5f48),
	.w7(32'h3a5d6da9),
	.w8(32'h38abe70e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule