module layer_10_featuremap_93(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39219b75),
	.w1(32'h38e42bf5),
	.w2(32'h399f37f0),
	.w3(32'h3948ab0d),
	.w4(32'hb9d944c8),
	.w5(32'hb9b7eab0),
	.w6(32'h391b6f2d),
	.w7(32'h3a0c2ac4),
	.w8(32'h3aa1ec2b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c485b3a),
	.w1(32'h3b83eaf1),
	.w2(32'h3bafd592),
	.w3(32'h3c1195b3),
	.w4(32'hba7a26b1),
	.w5(32'hbab8f4d7),
	.w6(32'h3bfb37d2),
	.w7(32'h3b6cf271),
	.w8(32'h3bae0c20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37766378),
	.w1(32'hb7f9b3b8),
	.w2(32'h39135419),
	.w3(32'h384261f1),
	.w4(32'h393e7f3a),
	.w5(32'h3988d095),
	.w6(32'hb95cbac3),
	.w7(32'hb92143d4),
	.w8(32'hb8d5eb5e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0729b1),
	.w1(32'hbb184d32),
	.w2(32'hbb6776e9),
	.w3(32'h39b0bf6f),
	.w4(32'h3a869f8e),
	.w5(32'h39e47cc7),
	.w6(32'h39b1c85e),
	.w7(32'h3a237bbf),
	.w8(32'h3a4bbc00),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6428b),
	.w1(32'h3a20f2ee),
	.w2(32'h39be8588),
	.w3(32'h38334c49),
	.w4(32'h3a332eb5),
	.w5(32'h3a24e4c1),
	.w6(32'hb896043e),
	.w7(32'hb94c040f),
	.w8(32'hb8870bb8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392b51d3),
	.w1(32'h37cd8b90),
	.w2(32'hb8e66415),
	.w3(32'h391da91b),
	.w4(32'h38c4f87a),
	.w5(32'hb949aa20),
	.w6(32'hb8bcde6a),
	.w7(32'hb85121c6),
	.w8(32'hb913cb63),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0de522),
	.w1(32'hbb078a43),
	.w2(32'h3bfb0f71),
	.w3(32'hbbddf0c2),
	.w4(32'h3b27d715),
	.w5(32'h3c48da15),
	.w6(32'hbb673fc6),
	.w7(32'hbafc6edf),
	.w8(32'h3c4abf2a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd355df),
	.w1(32'h3cda18ac),
	.w2(32'h3c9b8e7c),
	.w3(32'h3cc7d20a),
	.w4(32'h3ca398b6),
	.w5(32'h3c699989),
	.w6(32'h3ca23c0a),
	.w7(32'h3cd908e4),
	.w8(32'h3bd9876f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b518c),
	.w1(32'hba7d0b8e),
	.w2(32'h3919bbce),
	.w3(32'h39b09119),
	.w4(32'hba593a58),
	.w5(32'hba7e9b76),
	.w6(32'hba0da8d2),
	.w7(32'hba4c765e),
	.w8(32'hb9ba5962),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6abcd),
	.w1(32'hb9446254),
	.w2(32'h3c485e0e),
	.w3(32'hbbdbf7c5),
	.w4(32'hbb2b5000),
	.w5(32'h3b9e4031),
	.w6(32'h3c3ebe91),
	.w7(32'h3c12cd9c),
	.w8(32'h3ca663a4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cd7fd),
	.w1(32'h3a958383),
	.w2(32'h3ad187af),
	.w3(32'h3a1c724a),
	.w4(32'h39bc1997),
	.w5(32'h3a683add),
	.w6(32'h39b0ee2a),
	.w7(32'h3936bf40),
	.w8(32'h39ef3db1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e7fe),
	.w1(32'hbc446f5a),
	.w2(32'h3b89ce1b),
	.w3(32'hbc849ff7),
	.w4(32'hbc14630d),
	.w5(32'h3c178d0b),
	.w6(32'hbb8fb5d5),
	.w7(32'hbbafa906),
	.w8(32'h3c251a3d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38f724),
	.w1(32'h39657442),
	.w2(32'h3bed44a0),
	.w3(32'hbc3132a0),
	.w4(32'hbb820998),
	.w5(32'h3b3860ed),
	.w6(32'h3bb62581),
	.w7(32'h3bdc1d3e),
	.w8(32'h3c8b4af7),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91ff4c),
	.w1(32'h3b5b9111),
	.w2(32'h3c2d2b7e),
	.w3(32'hbbbd5c0e),
	.w4(32'hbaf6660a),
	.w5(32'h3bf584fd),
	.w6(32'hba58fe3b),
	.w7(32'h3ac4e485),
	.w8(32'h3c06384a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5279f),
	.w1(32'hb9f5d96f),
	.w2(32'hba8a57bc),
	.w3(32'h3b25e35d),
	.w4(32'hbba8acdb),
	.w5(32'hbbccdec3),
	.w6(32'h3bb97806),
	.w7(32'h3b5c3d77),
	.w8(32'h3b9b7007),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89c6f0),
	.w1(32'h3c3dea1a),
	.w2(32'h3bd12402),
	.w3(32'h3bb9f6c9),
	.w4(32'h3ba2e392),
	.w5(32'hba3ddc3d),
	.w6(32'h3c9a2335),
	.w7(32'h3c43481d),
	.w8(32'h3c8e4cb9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1a4db),
	.w1(32'hba05356b),
	.w2(32'hba327903),
	.w3(32'hb84f0d1f),
	.w4(32'hba4f3ed5),
	.w5(32'hba4e6c81),
	.w6(32'hb9453eef),
	.w7(32'hba87094b),
	.w8(32'hba724c91),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98baf3),
	.w1(32'h3b428bd1),
	.w2(32'h3c67221e),
	.w3(32'h3b973381),
	.w4(32'h3b8374ec),
	.w5(32'h3ca01768),
	.w6(32'h3c873da6),
	.w7(32'h3ba78356),
	.w8(32'h3cb33ba4),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb596d00),
	.w1(32'hbb18ca73),
	.w2(32'h3b481eef),
	.w3(32'hbb9f61c4),
	.w4(32'hbad99894),
	.w5(32'h3b91b9ed),
	.w6(32'h3bd41b30),
	.w7(32'h3b54e1b6),
	.w8(32'h3c3f5d4b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39786d9d),
	.w1(32'hba0fe683),
	.w2(32'hba088c71),
	.w3(32'hb8aafb26),
	.w4(32'hba61b737),
	.w5(32'hba4c040b),
	.w6(32'hb73bddc8),
	.w7(32'hb9847090),
	.w8(32'hb98d7ba0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990b903),
	.w1(32'hb941e700),
	.w2(32'hb9ac6699),
	.w3(32'hb8a2f077),
	.w4(32'h3957b219),
	.w5(32'h395bcdf0),
	.w6(32'h3927ee31),
	.w7(32'h389254fe),
	.w8(32'hb9969237),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5544),
	.w1(32'hbb5cd34b),
	.w2(32'h39fccb11),
	.w3(32'hbbad7912),
	.w4(32'hbb59cc71),
	.w5(32'h39d2caf6),
	.w6(32'hbba69274),
	.w7(32'hba73eb8b),
	.w8(32'h3a98b8f2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c892de1),
	.w1(32'h3c6ad2d0),
	.w2(32'h3c75199e),
	.w3(32'hbb810eb1),
	.w4(32'h3ac7cbbc),
	.w5(32'h3c16116b),
	.w6(32'h3d469015),
	.w7(32'h3c97dce1),
	.w8(32'h3d35666e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb818d2f8),
	.w1(32'h39940995),
	.w2(32'h3c35882d),
	.w3(32'hbb451891),
	.w4(32'hbbaee3b8),
	.w5(32'h3b3d8234),
	.w6(32'h3c4c9e84),
	.w7(32'h3c142d4b),
	.w8(32'h3c8f0b69),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef3982),
	.w1(32'hbb9e58d0),
	.w2(32'h3a20d85d),
	.w3(32'h3c0ef1d5),
	.w4(32'hbb878acb),
	.w5(32'hbbc55b38),
	.w6(32'h3c50a5cc),
	.w7(32'h3c2ffc5d),
	.w8(32'h3c8076f2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf7311),
	.w1(32'h391de25a),
	.w2(32'h3a2fe03a),
	.w3(32'h391aedc8),
	.w4(32'hb91c0b25),
	.w5(32'h391e6067),
	.w6(32'hb959acc3),
	.w7(32'h3889f3a7),
	.w8(32'h38da82c1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b67493),
	.w1(32'hb998efe8),
	.w2(32'hb9f8918e),
	.w3(32'hba20b24c),
	.w4(32'hb93806ef),
	.w5(32'hba07e63a),
	.w6(32'hb9ee94d4),
	.w7(32'hb9ad3e76),
	.w8(32'hba308198),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd852864),
	.w1(32'h3ca0cadc),
	.w2(32'h3c5a688f),
	.w3(32'hbd5756be),
	.w4(32'h3cfeaa1e),
	.w5(32'h3ca3f9f0),
	.w6(32'hbd82e9f1),
	.w7(32'h3c8f08af),
	.w8(32'h3c86529a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb215c68),
	.w1(32'hbb7f7602),
	.w2(32'h3a9592e6),
	.w3(32'hbb3ba46f),
	.w4(32'hbb90c3e2),
	.w5(32'h369fad0c),
	.w6(32'hbb2c4931),
	.w7(32'hbb73a993),
	.w8(32'hba755d99),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd398ef4),
	.w1(32'hba034e0b),
	.w2(32'h3b156442),
	.w3(32'hbccd0fb5),
	.w4(32'h3c721366),
	.w5(32'h3c8136ac),
	.w6(32'hbd00395e),
	.w7(32'h3c21dd89),
	.w8(32'h3c97c1cf),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aec849),
	.w1(32'hb8e512b6),
	.w2(32'hb9703dae),
	.w3(32'hb84bbd4b),
	.w4(32'hb7d42da2),
	.w5(32'hb8f6f526),
	.w6(32'hb87f2afb),
	.w7(32'hb8cea592),
	.w8(32'hb8eed837),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c379c8),
	.w1(32'hb8843cb6),
	.w2(32'hb936da11),
	.w3(32'hb896c9ae),
	.w4(32'hb62da8a8),
	.w5(32'hb9466365),
	.w6(32'h37bcb20f),
	.w7(32'hb885f680),
	.w8(32'hb9124c7b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d41bb),
	.w1(32'hbaa806d7),
	.w2(32'h3b705d1d),
	.w3(32'hbb1f4833),
	.w4(32'hbb228f8c),
	.w5(32'h3b269f03),
	.w6(32'h3bd5a0d3),
	.w7(32'h3b982562),
	.w8(32'h3c37c3d1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933004),
	.w1(32'h3a417593),
	.w2(32'h3b50ecf9),
	.w3(32'h3ba731e3),
	.w4(32'hb8aa7126),
	.w5(32'hb9d4e870),
	.w6(32'h3b872498),
	.w7(32'h3b85cb16),
	.w8(32'h3b7c4221),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb228df8),
	.w1(32'hba935088),
	.w2(32'hbade2d99),
	.w3(32'hbb897a14),
	.w4(32'hbb0709a0),
	.w5(32'hba2e120c),
	.w6(32'hba96b130),
	.w7(32'hb920cf72),
	.w8(32'h3ab252a6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d6271),
	.w1(32'h3ac9b803),
	.w2(32'h3b849b12),
	.w3(32'hbb5f600d),
	.w4(32'h3b2b4ab3),
	.w5(32'h3bbc1cad),
	.w6(32'h3b7ffcff),
	.w7(32'hb8c64c1a),
	.w8(32'h3b298c4f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d17f679),
	.w1(32'h3aa542cb),
	.w2(32'h3cdd5e89),
	.w3(32'hbc01c143),
	.w4(32'hbcc882a6),
	.w5(32'hbc5c4692),
	.w6(32'h3c493ced),
	.w7(32'hbc72d4d9),
	.w8(32'h3b13f6e8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb106ac),
	.w1(32'hbbccfa72),
	.w2(32'h3c3fc562),
	.w3(32'hbc88c9b8),
	.w4(32'hbc1ea07f),
	.w5(32'h3bd28f1c),
	.w6(32'hbc44d133),
	.w7(32'h3c2e982c),
	.w8(32'h3ccb5660),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd7e4f3c),
	.w1(32'h3b0444bb),
	.w2(32'h3cdb175d),
	.w3(32'hbd4454de),
	.w4(32'h3c52a25f),
	.w5(32'h3d08f9ee),
	.w6(32'hbd411b4a),
	.w7(32'h3c8746b1),
	.w8(32'h3d23d8f1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804938),
	.w1(32'hbb32951b),
	.w2(32'hbb201015),
	.w3(32'h3b03df0d),
	.w4(32'hbb2e7ee5),
	.w5(32'hbb54cae2),
	.w6(32'h3adba7b1),
	.w7(32'h3a38d5a7),
	.w8(32'h3a54d19d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3914ec40),
	.w1(32'hb78fba67),
	.w2(32'hb8aba9ae),
	.w3(32'h398fc42c),
	.w4(32'hb9298cbf),
	.w5(32'hb901e18b),
	.w6(32'hb9eac13c),
	.w7(32'hb84077e4),
	.w8(32'hba031474),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02abb1),
	.w1(32'hb9f62f87),
	.w2(32'hba1c2401),
	.w3(32'hb9a3ea89),
	.w4(32'hb9aa275e),
	.w5(32'hba184e51),
	.w6(32'hba59605f),
	.w7(32'hba4de59a),
	.w8(32'hba70795c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4489fd),
	.w1(32'hbb951ece),
	.w2(32'h3a050e9f),
	.w3(32'hbb232289),
	.w4(32'hbb8e0baf),
	.w5(32'h3aedc9e1),
	.w6(32'hbab01a01),
	.w7(32'hbb60a44a),
	.w8(32'hb97db29c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6c950),
	.w1(32'h3b9e54d4),
	.w2(32'h3c6d9886),
	.w3(32'hbc041459),
	.w4(32'h3986a41e),
	.w5(32'h3c089748),
	.w6(32'h3c29d068),
	.w7(32'h3c4fa5a1),
	.w8(32'h3cfe7a58),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaede35e),
	.w1(32'h3a9fccb5),
	.w2(32'h3c09367b),
	.w3(32'h3a0d5764),
	.w4(32'hbb40de70),
	.w5(32'h3b29d83b),
	.w6(32'h3bd0181d),
	.w7(32'h3c0a446d),
	.w8(32'h3c8efd2f),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad10ba3),
	.w1(32'hb864bc66),
	.w2(32'h3bbc56d9),
	.w3(32'h3ad0b4ee),
	.w4(32'hbbc85d4f),
	.w5(32'hbb2af25d),
	.w6(32'h3cbb03d7),
	.w7(32'h3c4ae0b2),
	.w8(32'h3c9c17e5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb98657),
	.w1(32'h3aad6547),
	.w2(32'h3bec7a90),
	.w3(32'h38aa9f1d),
	.w4(32'hbb2bda6b),
	.w5(32'h3b8f3d5c),
	.w6(32'h3c4333af),
	.w7(32'h3c2893f7),
	.w8(32'h3c9238ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3223b8),
	.w1(32'hbb41de42),
	.w2(32'h3c6d0e7a),
	.w3(32'hbc3df1a0),
	.w4(32'hbafa0c66),
	.w5(32'h3ca29bff),
	.w6(32'h3c61a2bc),
	.w7(32'h3c008c8f),
	.w8(32'h3d01536e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dff86d),
	.w1(32'hb995ab0b),
	.w2(32'h392f4e9f),
	.w3(32'hba22abf6),
	.w4(32'hb9d11eaf),
	.w5(32'hb876a5d2),
	.w6(32'hba132e1c),
	.w7(32'hb8ba9be4),
	.w8(32'hb979ff69),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db3a67),
	.w1(32'hb971b2d5),
	.w2(32'hb9d77930),
	.w3(32'hb9adace1),
	.w4(32'h39cca6bf),
	.w5(32'hb9045933),
	.w6(32'h3a3f00bc),
	.w7(32'h3a5328ba),
	.w8(32'h3a4b9010),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3807da12),
	.w1(32'h39cf1ea7),
	.w2(32'h39f23f6c),
	.w3(32'h399e5bb1),
	.w4(32'h3a121eb7),
	.w5(32'h39c4781a),
	.w6(32'h39536f32),
	.w7(32'h396b1014),
	.w8(32'h3a0d6397),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a559676),
	.w1(32'h3c2bc8c9),
	.w2(32'h3c1570bd),
	.w3(32'hba566433),
	.w4(32'h3bd8f48e),
	.w5(32'h3bcd9130),
	.w6(32'h3beac426),
	.w7(32'h3bf7476f),
	.w8(32'h3c8abd9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b090cf1),
	.w1(32'h3aa9b364),
	.w2(32'h3b557599),
	.w3(32'h3abffaa2),
	.w4(32'h3aaaa92f),
	.w5(32'h3b02149f),
	.w6(32'h3b8fd8b0),
	.w7(32'h3b413403),
	.w8(32'h3b959e95),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b485d63),
	.w1(32'h3b1ed368),
	.w2(32'h3c54e18f),
	.w3(32'hbbcaa23a),
	.w4(32'h3ac1e100),
	.w5(32'h3c626194),
	.w6(32'h3c340495),
	.w7(32'h3c12133b),
	.w8(32'h3ccd05e0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b66a6),
	.w1(32'h3ba30f24),
	.w2(32'h3b80760d),
	.w3(32'hbabc1c77),
	.w4(32'h3b13b87b),
	.w5(32'h3baf54b6),
	.w6(32'hbab24db1),
	.w7(32'h3a11b96d),
	.w8(32'h3bcc8fc3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d4101),
	.w1(32'hba082a25),
	.w2(32'hb935ea5a),
	.w3(32'h39d4797e),
	.w4(32'hba8d57ff),
	.w5(32'hba9dcec6),
	.w6(32'hb9542900),
	.w7(32'hb9ec0060),
	.w8(32'hba688440),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd1f6d),
	.w1(32'hb9b2774d),
	.w2(32'hb9f90899),
	.w3(32'h399b326e),
	.w4(32'hb98bbd79),
	.w5(32'hb9c910cf),
	.w6(32'hb9b6be07),
	.w7(32'hb9c76b4d),
	.w8(32'hb9f2cb0e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48335a),
	.w1(32'hba3c6c51),
	.w2(32'h3a267b59),
	.w3(32'hbadf7523),
	.w4(32'h3a97c39e),
	.w5(32'h3b1693e4),
	.w6(32'hbaee77df),
	.w7(32'h39df2d4b),
	.w8(32'h3b4c8a2b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02e30c),
	.w1(32'hbb1a12a6),
	.w2(32'hba345225),
	.w3(32'hbaa6ea57),
	.w4(32'hbaafaf73),
	.w5(32'h388dacf9),
	.w6(32'hbabfae63),
	.w7(32'hbaa969bd),
	.w8(32'hb81cce35),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23e5e5),
	.w1(32'hba66b779),
	.w2(32'hba7cc338),
	.w3(32'hbb14f92c),
	.w4(32'hb894aeb3),
	.w5(32'h3a9b2dbd),
	.w6(32'hba922325),
	.w7(32'h38930a1a),
	.w8(32'h3a71c175),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390e0d15),
	.w1(32'h3ac4d097),
	.w2(32'h3b85312a),
	.w3(32'hbb6df929),
	.w4(32'hb9bf9587),
	.w5(32'h3baf2d11),
	.w6(32'h3ba40171),
	.w7(32'h3b44fda6),
	.w8(32'h3c3b2735),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62f252),
	.w1(32'h3c3f24f1),
	.w2(32'h3bd028a5),
	.w3(32'hbbeca612),
	.w4(32'h3c0d52c5),
	.w5(32'h3c1f3034),
	.w6(32'hbbcc8340),
	.w7(32'h3a68a4ea),
	.w8(32'h3c6adfc4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f28cee),
	.w1(32'hb9c5de6f),
	.w2(32'hba3b7b9f),
	.w3(32'h396bf939),
	.w4(32'hba1b2efe),
	.w5(32'hba5e658a),
	.w6(32'hb9d04768),
	.w7(32'hba5286c0),
	.w8(32'hba23ed1d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e57c4c),
	.w1(32'h39014b3d),
	.w2(32'hb9ad2ace),
	.w3(32'hba08c6c9),
	.w4(32'h3968d0f8),
	.w5(32'hb920ec07),
	.w6(32'hb82f5d33),
	.w7(32'hb9265c54),
	.w8(32'hb82589bc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894e8b4),
	.w1(32'hb98b4925),
	.w2(32'hb8c641c1),
	.w3(32'h389c946b),
	.w4(32'hb9927ca8),
	.w5(32'hb95a131e),
	.w6(32'hb96ced48),
	.w7(32'hb99ef63e),
	.w8(32'hb9b62d90),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a542be),
	.w1(32'hb9f6ee0c),
	.w2(32'hba0a2fe4),
	.w3(32'h38f0b2f5),
	.w4(32'hb963721d),
	.w5(32'hb9f99094),
	.w6(32'hba1bedf1),
	.w7(32'hba0636fa),
	.w8(32'hb85fa3d5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79148b),
	.w1(32'h3c065dfb),
	.w2(32'h3c28e270),
	.w3(32'hbc8706be),
	.w4(32'hbc6de08d),
	.w5(32'hbbdbfd38),
	.w6(32'h3bd1129e),
	.w7(32'h3c2a90ab),
	.w8(32'h3ca1be78),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eabee),
	.w1(32'hbaa819ba),
	.w2(32'h3ba52a0d),
	.w3(32'h3be1fa1f),
	.w4(32'h3ae5df5d),
	.w5(32'h3bcb8224),
	.w6(32'h3d1d714b),
	.w7(32'h3cbae56a),
	.w8(32'h3cf9471c),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0a927),
	.w1(32'h3bc99c72),
	.w2(32'h3ca2a208),
	.w3(32'h3b053eb7),
	.w4(32'h3adf823a),
	.w5(32'h3c76e2d7),
	.w6(32'h3ca9b99a),
	.w7(32'h3c36c976),
	.w8(32'h3d055682),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc761502),
	.w1(32'hbbae7078),
	.w2(32'h3b42dadd),
	.w3(32'hbaa1ba97),
	.w4(32'hbb5aebab),
	.w5(32'h3a18ecf6),
	.w6(32'h3c6e1829),
	.w7(32'h3cd181bb),
	.w8(32'h3d0e894b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1e1f0),
	.w1(32'hb7e54659),
	.w2(32'hb97fe129),
	.w3(32'h3a19f381),
	.w4(32'hb889ac05),
	.w5(32'hb9e5cc3e),
	.w6(32'hb9460946),
	.w7(32'hb943b9b7),
	.w8(32'hba039fdc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f42e3a),
	.w1(32'h392a9782),
	.w2(32'hb986b329),
	.w3(32'hb8a7d494),
	.w4(32'h39bcfd9d),
	.w5(32'hb94b84e5),
	.w6(32'hb930bca7),
	.w7(32'hb8ec0695),
	.w8(32'hb9c683e2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b948aa),
	.w1(32'h3962fc91),
	.w2(32'hb9688adb),
	.w3(32'hb8a3913f),
	.w4(32'h398da59b),
	.w5(32'hb92ba7d7),
	.w6(32'hb9647ede),
	.w7(32'hb9112ae2),
	.w8(32'hb9ecb39c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8830f2),
	.w1(32'hba53597c),
	.w2(32'hba1e2101),
	.w3(32'hbafb4ded),
	.w4(32'hbb08d9aa),
	.w5(32'h375aa7e4),
	.w6(32'h3a86f4f0),
	.w7(32'h39b3c150),
	.w8(32'h3b3e7e61),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98828d6),
	.w1(32'hb899dfcd),
	.w2(32'hb9b6741f),
	.w3(32'hb92078fa),
	.w4(32'h3935f608),
	.w5(32'hb91763df),
	.w6(32'hb928694b),
	.w7(32'hb94fe98a),
	.w8(32'hb99beec7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1105c2),
	.w1(32'h3b68e4fd),
	.w2(32'h3b6de03f),
	.w3(32'hba97f26f),
	.w4(32'h3ae2af70),
	.w5(32'h3bcf65f4),
	.w6(32'h3b8569bb),
	.w7(32'h3bd46720),
	.w8(32'h3c48e040),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04e8c9),
	.w1(32'h3b16d8c2),
	.w2(32'h3bf1df1c),
	.w3(32'hbab42f27),
	.w4(32'h3accf96e),
	.w5(32'h3c2d6dfd),
	.w6(32'h3c64704e),
	.w7(32'h3bd3ce5f),
	.w8(32'h3c7405c7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bcea6),
	.w1(32'h3b3eed1f),
	.w2(32'h3ac487a2),
	.w3(32'h3aa1e6b6),
	.w4(32'hbb048e0e),
	.w5(32'hbb847a7f),
	.w6(32'h3b98669e),
	.w7(32'h3bf68d59),
	.w8(32'h3c113024),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2731bf),
	.w1(32'h3b0c5d42),
	.w2(32'h3c046856),
	.w3(32'h3b0fb299),
	.w4(32'h3a1e814c),
	.w5(32'h3b9a9f1c),
	.w6(32'h3bf7e002),
	.w7(32'h3b9cb5ce),
	.w8(32'h3c2678be),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda6a6e),
	.w1(32'h3ba3aa08),
	.w2(32'h3b82a734),
	.w3(32'hbbc3859c),
	.w4(32'hbb871e4a),
	.w5(32'hbad6ef7c),
	.w6(32'h3b9850c1),
	.w7(32'h3b9605e4),
	.w8(32'h3bb542eb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8823d8),
	.w1(32'h3b53a0e7),
	.w2(32'h3bb34d5d),
	.w3(32'hba1cfb44),
	.w4(32'h3adbf9a0),
	.w5(32'h3b19f920),
	.w6(32'hba75443a),
	.w7(32'h3b2e60a6),
	.w8(32'h3bdcbb89),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c6d2c),
	.w1(32'hb7463771),
	.w2(32'h3bd0d322),
	.w3(32'hbb43701e),
	.w4(32'h3a727582),
	.w5(32'h3c033e9b),
	.w6(32'h3ba42477),
	.w7(32'h3b8b9ee2),
	.w8(32'h3c49e86b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d11a0b),
	.w1(32'hb96ee1f0),
	.w2(32'hb94dda2b),
	.w3(32'h39789e3c),
	.w4(32'hb94ff8e2),
	.w5(32'hb93732a6),
	.w6(32'hb9510d93),
	.w7(32'hb97bab8d),
	.w8(32'hb94a464b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39241b69),
	.w1(32'h397a154d),
	.w2(32'h39385624),
	.w3(32'h38b0e334),
	.w4(32'h392cf9d0),
	.w5(32'h3919829c),
	.w6(32'h390350fd),
	.w7(32'h37bb86c5),
	.w8(32'h39018392),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88061f2),
	.w1(32'hb7c219c4),
	.w2(32'hb8c12b49),
	.w3(32'h38ddded0),
	.w4(32'hb9e3f4ca),
	.w5(32'hb9cd201e),
	.w6(32'hba2a6e50),
	.w7(32'hba2d9a2d),
	.w8(32'hba52022d),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54dcfb),
	.w1(32'hbaae6906),
	.w2(32'hb9795376),
	.w3(32'hbab2af96),
	.w4(32'h3a3d6375),
	.w5(32'h3b0de7a6),
	.w6(32'hbb38c57e),
	.w7(32'h39e9e660),
	.w8(32'h3ac440c2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeb749),
	.w1(32'hbb568cae),
	.w2(32'h3b3cf962),
	.w3(32'h3c1375cc),
	.w4(32'hbbde0c75),
	.w5(32'hbb519ff0),
	.w6(32'h3c3eb556),
	.w7(32'h3bb54aad),
	.w8(32'h3bceb6f8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e0445),
	.w1(32'hbb50d48a),
	.w2(32'hbad22456),
	.w3(32'hbaae90bd),
	.w4(32'hbb2e2344),
	.w5(32'hba87efa6),
	.w6(32'h3a05446b),
	.w7(32'hbab4ea64),
	.w8(32'hb9cc7048),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90d13d),
	.w1(32'hbb0cb807),
	.w2(32'hbbec0b78),
	.w3(32'h3c217c80),
	.w4(32'h382d0b29),
	.w5(32'hbb8d8e48),
	.w6(32'h3c5d8e04),
	.w7(32'h3c142261),
	.w8(32'h3b9829ff),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fb525),
	.w1(32'h3b625e9a),
	.w2(32'h3c3fa35f),
	.w3(32'h3b4d7313),
	.w4(32'h3bc9a7d6),
	.w5(32'h3c9314ec),
	.w6(32'h3cb7d913),
	.w7(32'h3c725b5a),
	.w8(32'h3cec5af8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccc07e1),
	.w1(32'hbb87fd33),
	.w2(32'h3bbdbd40),
	.w3(32'hbc962763),
	.w4(32'h3bb9a2cb),
	.w5(32'h3c456ade),
	.w6(32'hbcb1abaa),
	.w7(32'h3bb15311),
	.w8(32'h3c5e938f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92bb64),
	.w1(32'h3bfebc4e),
	.w2(32'h3b7bb7c6),
	.w3(32'hbc3667c9),
	.w4(32'hbb3b8f26),
	.w5(32'hbc17cef6),
	.w6(32'h3ca730eb),
	.w7(32'h3c060c06),
	.w8(32'h3c956b51),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc081054),
	.w1(32'hb9ac30d3),
	.w2(32'h3bf21301),
	.w3(32'hbb8a1198),
	.w4(32'h3b5a5eb4),
	.w5(32'h3c36370c),
	.w6(32'h3b7a6e95),
	.w7(32'h3c05d10a),
	.w8(32'h3c65b091),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd0f0),
	.w1(32'h3b24bd6c),
	.w2(32'h3c17f674),
	.w3(32'h3b424d30),
	.w4(32'hbb11d617),
	.w5(32'hbb3811cd),
	.w6(32'h3cbcde14),
	.w7(32'h3c57621c),
	.w8(32'h3c8824d9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c465c32),
	.w1(32'h3c22c948),
	.w2(32'h3b2ccdf9),
	.w3(32'hba9b7bbd),
	.w4(32'h39eb13c2),
	.w5(32'hbb084006),
	.w6(32'h3bf3d3ca),
	.w7(32'h3bfc99df),
	.w8(32'h3c188a10),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d017a),
	.w1(32'hb9e809ca),
	.w2(32'h3a58e967),
	.w3(32'hbbd53ac3),
	.w4(32'h390838a1),
	.w5(32'hb8eddfca),
	.w6(32'hbc29521b),
	.w7(32'h3be20def),
	.w8(32'h3c4d8fd7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99151a0),
	.w1(32'hba1cce28),
	.w2(32'hba118071),
	.w3(32'hba7fe5f0),
	.w4(32'hba4ffd32),
	.w5(32'hba80ceca),
	.w6(32'hba825b08),
	.w7(32'hba841862),
	.w8(32'hbaba911a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c131),
	.w1(32'hbac777f0),
	.w2(32'h3c126ac1),
	.w3(32'hbbaa6c1d),
	.w4(32'hbb85b442),
	.w5(32'h3bad3046),
	.w6(32'h3c61daa1),
	.w7(32'h3c118449),
	.w8(32'h3cae05fb),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94225f),
	.w1(32'h3bc956c6),
	.w2(32'h3c17fdd4),
	.w3(32'hbc9456e7),
	.w4(32'hbb1287af),
	.w5(32'h3bc397e8),
	.w6(32'h3b274786),
	.w7(32'h3c619e02),
	.w8(32'h3cb50e03),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cee5f19),
	.w1(32'hbaef2368),
	.w2(32'h3ca06906),
	.w3(32'h3b95e540),
	.w4(32'h3a159ff2),
	.w5(32'hbb0edcf6),
	.w6(32'h3d186140),
	.w7(32'hbbad0c34),
	.w8(32'h3bf784b8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1b3a1),
	.w1(32'hbc1cebdf),
	.w2(32'h3c048f77),
	.w3(32'hbb44ef69),
	.w4(32'hbc4b74c6),
	.w5(32'hbbc4cba7),
	.w6(32'hbb62a378),
	.w7(32'hbb04e447),
	.w8(32'h3b46f4bd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4d7bd),
	.w1(32'hbaf4acf8),
	.w2(32'h3b84356f),
	.w3(32'h3a8de827),
	.w4(32'hbb6b003f),
	.w5(32'hbb23215b),
	.w6(32'h3c34ea06),
	.w7(32'h3c2624dc),
	.w8(32'h3c4a021f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c76ce9b),
	.w1(32'hbb0222b3),
	.w2(32'h3c838a30),
	.w3(32'hbc408cf2),
	.w4(32'hbbf31db2),
	.w5(32'hbbb428c0),
	.w6(32'h3c555718),
	.w7(32'hbc43ff94),
	.w8(32'h3c488357),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9992c1a),
	.w1(32'hba9a5065),
	.w2(32'hba1b9cae),
	.w3(32'hba183043),
	.w4(32'hb9a3f36d),
	.w5(32'hba22bd28),
	.w6(32'hba068ceb),
	.w7(32'hbaa55f31),
	.w8(32'hb9d13a73),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20a157),
	.w1(32'h3bafecf4),
	.w2(32'h3ca412ec),
	.w3(32'h3bf7c031),
	.w4(32'hbbd59b49),
	.w5(32'h3bcac6b5),
	.w6(32'h3c7774e9),
	.w7(32'h3b817298),
	.w8(32'h3c41801c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7163c3),
	.w1(32'hbc08b836),
	.w2(32'h3c840807),
	.w3(32'hbbcc976d),
	.w4(32'hbbba8c55),
	.w5(32'h3c3c9787),
	.w6(32'hbac3984d),
	.w7(32'h3b4189e3),
	.w8(32'h3be8d264),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45985),
	.w1(32'h39d575e9),
	.w2(32'h3a465d3f),
	.w3(32'hbad37e1f),
	.w4(32'h39a75a87),
	.w5(32'h3a30389f),
	.w6(32'hbb1060a9),
	.w7(32'hba545800),
	.w8(32'hb9a10052),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0baf2),
	.w1(32'h3b01b65a),
	.w2(32'hbab3eb09),
	.w3(32'h3be7966b),
	.w4(32'h3b14a505),
	.w5(32'hba92dc44),
	.w6(32'h3c0c75dd),
	.w7(32'h3bcb5440),
	.w8(32'h3b86c859),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc153a6e),
	.w1(32'hbb90d4f9),
	.w2(32'h3be5bd17),
	.w3(32'hbc3387a6),
	.w4(32'hbbcba006),
	.w5(32'h3b6c8f02),
	.w6(32'h3bc1f714),
	.w7(32'h3ba25277),
	.w8(32'h3c8276ce),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe48c90),
	.w1(32'hb9743749),
	.w2(32'h3b88a25f),
	.w3(32'hba9d1408),
	.w4(32'h3a0bd767),
	.w5(32'h3aa37bb1),
	.w6(32'h3a07d5b7),
	.w7(32'h3bac116c),
	.w8(32'h3c0dbef7),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e98c3),
	.w1(32'h3b12f5c3),
	.w2(32'h3bc90943),
	.w3(32'hbc5467d3),
	.w4(32'h3aff27ba),
	.w5(32'h3c011944),
	.w6(32'hbc941a41),
	.w7(32'h3bc2099d),
	.w8(32'h3c5a2f15),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39502800),
	.w1(32'h3a09c5c6),
	.w2(32'h3a067f14),
	.w3(32'hbaef9d0a),
	.w4(32'hbb9efd85),
	.w5(32'hbb0943b2),
	.w6(32'h3a234ed6),
	.w7(32'h3b8a4b6b),
	.w8(32'h3c048b73),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa6ce),
	.w1(32'hbc53036b),
	.w2(32'hbc50dbdf),
	.w3(32'h3b7a6214),
	.w4(32'h394b2edc),
	.w5(32'hbb503d95),
	.w6(32'h3c9f6d41),
	.w7(32'h3c143ebf),
	.w8(32'h3be5dae2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad4652),
	.w1(32'h3c58cc17),
	.w2(32'h3c07809f),
	.w3(32'h3ba069bc),
	.w4(32'h3b1d0bb5),
	.w5(32'hbae05cec),
	.w6(32'h3c77fb16),
	.w7(32'h3bafd247),
	.w8(32'h3bbf567d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57b22a),
	.w1(32'hb9fc4cb7),
	.w2(32'h3b582d0d),
	.w3(32'h3a10b724),
	.w4(32'hbab189e3),
	.w5(32'h3ab6aa34),
	.w6(32'h3bb0a34f),
	.w7(32'h3baa1bc5),
	.w8(32'h3c105ab0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a100fdd),
	.w1(32'h39cba15d),
	.w2(32'h39768748),
	.w3(32'h39d496be),
	.w4(32'h3a00a699),
	.w5(32'h3929b6ac),
	.w6(32'h3a3494e5),
	.w7(32'h39992855),
	.w8(32'h39a318d3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8404e2),
	.w1(32'h3b0e5999),
	.w2(32'h3a12a8a3),
	.w3(32'h3b1fd1f8),
	.w4(32'h3a00113c),
	.w5(32'hba8e2d0e),
	.w6(32'h3b1fa80f),
	.w7(32'h3b01491d),
	.w8(32'hb8de2232),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d65f44),
	.w1(32'hb42bd49a),
	.w2(32'hb744bfe6),
	.w3(32'h3984eb37),
	.w4(32'h396bfa5a),
	.w5(32'h38795174),
	.w6(32'h38c872ad),
	.w7(32'h384f58cf),
	.w8(32'h38105f1b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38118635),
	.w1(32'h39397ba0),
	.w2(32'h3a361900),
	.w3(32'h391ae0ef),
	.w4(32'h38d5f5a5),
	.w5(32'h39c4a5fd),
	.w6(32'hb972e504),
	.w7(32'hb96fc13c),
	.w8(32'hb92748e3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06540c),
	.w1(32'hbacb2b99),
	.w2(32'h3b29cb29),
	.w3(32'hba2364da),
	.w4(32'hbb723542),
	.w5(32'hba8f2063),
	.w6(32'h3baa5609),
	.w7(32'h3b932f67),
	.w8(32'h3bf66c63),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c01b3),
	.w1(32'h3a611807),
	.w2(32'h3a5b257b),
	.w3(32'h393f5dee),
	.w4(32'h398dd4b0),
	.w5(32'h3a8020f4),
	.w6(32'h3823b1ce),
	.w7(32'hb7ebc85e),
	.w8(32'h3a71d5ee),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aedd2b4),
	.w1(32'h3986c277),
	.w2(32'h3b1cb501),
	.w3(32'hbb8a5468),
	.w4(32'h392b3b67),
	.w5(32'h3ad5bb82),
	.w6(32'h3b4483aa),
	.w7(32'h3b2ada8b),
	.w8(32'h3bdff4f9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8df2e),
	.w1(32'hba549911),
	.w2(32'h3badf7f6),
	.w3(32'hbc04a22e),
	.w4(32'hba9669e8),
	.w5(32'h3b78ce66),
	.w6(32'hbc0a36b6),
	.w7(32'h3bdc462b),
	.w8(32'h3c8cc7dc),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398995dd),
	.w1(32'h398f3db3),
	.w2(32'h3a0ccbff),
	.w3(32'h38c9b332),
	.w4(32'hb9065e56),
	.w5(32'hb93b4f7a),
	.w6(32'h385c26cf),
	.w7(32'h3a14f302),
	.w8(32'h39dc4fcb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945513d),
	.w1(32'h39bb48b9),
	.w2(32'h3a580cbf),
	.w3(32'h3956b497),
	.w4(32'hb7e82316),
	.w5(32'hb8d426d1),
	.w6(32'h399269de),
	.w7(32'h3888b8ac),
	.w8(32'h39fdf53c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3926804a),
	.w1(32'hb98780b6),
	.w2(32'hb9b366e1),
	.w3(32'hb912b559),
	.w4(32'hb92ecab6),
	.w5(32'hb9711219),
	.w6(32'hb926bf47),
	.w7(32'hb95ace75),
	.w8(32'hb902016c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e270c),
	.w1(32'hbadbaa67),
	.w2(32'hbb121e2e),
	.w3(32'hba7cfe0d),
	.w4(32'hbaad4029),
	.w5(32'hbb02441e),
	.w6(32'h3980a020),
	.w7(32'hb9bd8b9b),
	.w8(32'hb8e7403b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb63df0),
	.w1(32'hbaa0402b),
	.w2(32'hbbab2a38),
	.w3(32'h3ad57365),
	.w4(32'h3c19e145),
	.w5(32'h3bae7d12),
	.w6(32'h3cbbf028),
	.w7(32'h3c0fb83b),
	.w8(32'h3c6ee866),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb923db1),
	.w1(32'hbaa5fd4b),
	.w2(32'h3bfb408c),
	.w3(32'hbbb4eda5),
	.w4(32'hbb6a889e),
	.w5(32'h3ba70b94),
	.w6(32'h3b95b029),
	.w7(32'h3be065f4),
	.w8(32'h3ca05787),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6591d2),
	.w1(32'hba17c63f),
	.w2(32'h3a234823),
	.w3(32'h38341229),
	.w4(32'hbab972f2),
	.w5(32'hba3b6ecc),
	.w6(32'h390fade8),
	.w7(32'h39851a42),
	.w8(32'h3aee4f56),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b577aa2),
	.w1(32'h3b9db3e7),
	.w2(32'h3b9a19d8),
	.w3(32'h3b0d85a8),
	.w4(32'hba40ac0a),
	.w5(32'h3ab66efb),
	.w6(32'h3bd03ba9),
	.w7(32'h3b9ea63c),
	.w8(32'h3bbc3e56),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adde7d6),
	.w1(32'h3b6ac450),
	.w2(32'h3b092957),
	.w3(32'hbb02ebae),
	.w4(32'h3a798e1b),
	.w5(32'h3aa04cf1),
	.w6(32'h3b2fb070),
	.w7(32'h3b20a644),
	.w8(32'h3b64585b),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ca190),
	.w1(32'h3b695a2c),
	.w2(32'h3b4cf8ff),
	.w3(32'hba06bd60),
	.w4(32'hbaac8372),
	.w5(32'hb9f61916),
	.w6(32'h3bb0d243),
	.w7(32'h3b51eb9a),
	.w8(32'h3afee700),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c625535),
	.w1(32'h3c7b0d6f),
	.w2(32'h3c1d7452),
	.w3(32'h3bb27ab7),
	.w4(32'h3ba35d58),
	.w5(32'h3a847c44),
	.w6(32'h3be4b25f),
	.w7(32'h3c03cb43),
	.w8(32'h3c3ca8f4),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bcb9b),
	.w1(32'h3b91de9d),
	.w2(32'h3c602c1c),
	.w3(32'hbc027ebe),
	.w4(32'h3b5d69c6),
	.w5(32'h3c423a06),
	.w6(32'h3bda86e0),
	.w7(32'h3c0dd928),
	.w8(32'h3cd456d1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a1024),
	.w1(32'hbb82a5f4),
	.w2(32'hba7f02b5),
	.w3(32'h3a18b3a0),
	.w4(32'hbb4369a9),
	.w5(32'hbabd9bd7),
	.w6(32'hb61e10dc),
	.w7(32'h3b1353dd),
	.w8(32'h3bbe2c64),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8f6bc),
	.w1(32'h3b49bd49),
	.w2(32'hba7f5962),
	.w3(32'hbb831324),
	.w4(32'hbb4f7f11),
	.w5(32'hbba029bd),
	.w6(32'h3c6bf921),
	.w7(32'h3ba8f465),
	.w8(32'h3bddd59e),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3152ca),
	.w1(32'h3bbbd791),
	.w2(32'h3bca59f3),
	.w3(32'h3a414c2f),
	.w4(32'h3ba2d6da),
	.w5(32'h3c0e9fc2),
	.w6(32'h3c23e762),
	.w7(32'h3b4522ce),
	.w8(32'h3c4b0269),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d21be),
	.w1(32'h3ac944fc),
	.w2(32'h3b06444c),
	.w3(32'h3bf958ad),
	.w4(32'h3a1f6de7),
	.w5(32'hbb621489),
	.w6(32'h3c9c21e1),
	.w7(32'h3c1d2f7b),
	.w8(32'h3bd3a727),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37d6a),
	.w1(32'hb9e0c74f),
	.w2(32'h3ae9d747),
	.w3(32'hbb2accb9),
	.w4(32'hbabf371b),
	.w5(32'h3b41e6d3),
	.w6(32'h3c07e600),
	.w7(32'h3b9615ab),
	.w8(32'h3c1f21b0),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03160c),
	.w1(32'h39aad707),
	.w2(32'h3afa1538),
	.w3(32'h3a7edec6),
	.w4(32'hb946de31),
	.w5(32'h3a68c3ed),
	.w6(32'h3b067b82),
	.w7(32'h3b368102),
	.w8(32'h3b8a026d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3f6f62),
	.w1(32'h3b9f4af4),
	.w2(32'hbbcdb3c8),
	.w3(32'hbce247c6),
	.w4(32'h3c8a69d6),
	.w5(32'h3c79e6d4),
	.w6(32'hbd06ab15),
	.w7(32'h3c9901d0),
	.w8(32'h3cc89b65),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd944f),
	.w1(32'h3a109cc6),
	.w2(32'h3a8c83de),
	.w3(32'h3b97be90),
	.w4(32'hbaae3a43),
	.w5(32'h3b008b43),
	.w6(32'h3c310064),
	.w7(32'h3b93f289),
	.w8(32'h3b9bf842),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1875c),
	.w1(32'h3a976354),
	.w2(32'hb98d8458),
	.w3(32'h399cf406),
	.w4(32'h3a2c9f32),
	.w5(32'hba2bb4fa),
	.w6(32'h3abc7218),
	.w7(32'hb8e22787),
	.w8(32'hb9746b50),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3092af),
	.w1(32'h3b70f93a),
	.w2(32'h3b798a3d),
	.w3(32'hb99e3bb2),
	.w4(32'h3ab9df83),
	.w5(32'h39e25bf5),
	.w6(32'h3b888859),
	.w7(32'h3b9bb231),
	.w8(32'hbadbcd62),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019aaf),
	.w1(32'hbb0bbaff),
	.w2(32'h3b451246),
	.w3(32'hbbeebb3a),
	.w4(32'hbb592615),
	.w5(32'h3acf885f),
	.w6(32'h3b57f5e7),
	.w7(32'h3a916c01),
	.w8(32'h3b815957),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be757c7),
	.w1(32'hb93dd286),
	.w2(32'h39530ac9),
	.w3(32'h3c232358),
	.w4(32'hbb8809db),
	.w5(32'hbba04eec),
	.w6(32'h3c2e463d),
	.w7(32'h3c0fdcdc),
	.w8(32'h3befa671),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba55d9d),
	.w1(32'hbb80b073),
	.w2(32'h3b045c01),
	.w3(32'hbbc01538),
	.w4(32'hbb83473f),
	.w5(32'hba86e0f4),
	.w6(32'h3bfece0d),
	.w7(32'h3bbbf5d6),
	.w8(32'h3c3d1db1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e97018),
	.w1(32'h3a363304),
	.w2(32'hba951ddd),
	.w3(32'h38bedfb5),
	.w4(32'h390834a6),
	.w5(32'hbacc05c4),
	.w6(32'h3ab4a4ea),
	.w7(32'hba362640),
	.w8(32'h3a814b0d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae69f49),
	.w1(32'h3bc0a90d),
	.w2(32'h3c4ef8d4),
	.w3(32'hbb85413e),
	.w4(32'h388e8788),
	.w5(32'h3b06633c),
	.w6(32'h3c19194b),
	.w7(32'h3c865f51),
	.w8(32'h3cca47c8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5849dd),
	.w1(32'hbaa5238e),
	.w2(32'h3b1e380d),
	.w3(32'hbbb1496f),
	.w4(32'hb774b641),
	.w5(32'h3a98e577),
	.w6(32'h3bf6e51b),
	.w7(32'h3bcb6987),
	.w8(32'h3be9f6f5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46a710),
	.w1(32'h3b181755),
	.w2(32'h3b05babd),
	.w3(32'hbb4c59bf),
	.w4(32'hb90419ae),
	.w5(32'hbc0db712),
	.w6(32'h3c21ab87),
	.w7(32'h3b331104),
	.w8(32'h3c4280e3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd067c36),
	.w1(32'h3c75b477),
	.w2(32'h3bd581c8),
	.w3(32'hbcfbfc9d),
	.w4(32'h3c30af3f),
	.w5(32'h3bc9012d),
	.w6(32'hbcf53ea2),
	.w7(32'h3ca101f0),
	.w8(32'h3ceb4e3e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d152),
	.w1(32'h3ac992f6),
	.w2(32'h3bd932a5),
	.w3(32'h3b856a57),
	.w4(32'hb94c8569),
	.w5(32'h3a1d2ef6),
	.w6(32'h3bae3e09),
	.w7(32'h3b73299d),
	.w8(32'h3b44f561),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abe539),
	.w1(32'hbb0acadc),
	.w2(32'hbb20c5d0),
	.w3(32'hbb8ebda3),
	.w4(32'hbad02d1f),
	.w5(32'hbb208c72),
	.w6(32'hbb17b71a),
	.w7(32'hbb44b2c6),
	.w8(32'hbb24b516),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b57ab),
	.w1(32'hbbc9a8fa),
	.w2(32'hbb5e5d9b),
	.w3(32'hbbf7a5de),
	.w4(32'hbb82c7e9),
	.w5(32'hbad2be8e),
	.w6(32'hbb2c85fa),
	.w7(32'h3aee4a5e),
	.w8(32'h3bd91161),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f25ad),
	.w1(32'h3bd085f6),
	.w2(32'h3c1d72a5),
	.w3(32'h3ada729a),
	.w4(32'hb996cb5e),
	.w5(32'h3b56317c),
	.w6(32'h3c1cfb79),
	.w7(32'h3bb3b0f1),
	.w8(32'h3be2bb58),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf138ab),
	.w1(32'hba8d799a),
	.w2(32'h3b82e653),
	.w3(32'hbb89398f),
	.w4(32'hbb74fe00),
	.w5(32'h3aaaf1a6),
	.w6(32'h3a76806e),
	.w7(32'h3bb2e7f4),
	.w8(32'h3b883810),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b4547),
	.w1(32'h3a52850a),
	.w2(32'h3a89101c),
	.w3(32'hbb6d0c01),
	.w4(32'hb9b88ead),
	.w5(32'h3a57d8ab),
	.w6(32'h3b4ca048),
	.w7(32'h39843ad4),
	.w8(32'h3ba416c6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b536b),
	.w1(32'h39a486ac),
	.w2(32'hba5dcf2d),
	.w3(32'h39c85c3d),
	.w4(32'h3988bfb9),
	.w5(32'hba81d9c5),
	.w6(32'h3a8259b4),
	.w7(32'hb7783f4e),
	.w8(32'h39bce38e),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39429fe6),
	.w1(32'hbaebb85a),
	.w2(32'h3b6de94c),
	.w3(32'hbbc2ff7c),
	.w4(32'hbaafaa22),
	.w5(32'h3971b9b2),
	.w6(32'h3c1538f3),
	.w7(32'h3b84e9c6),
	.w8(32'h3c1a428d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0c1e5),
	.w1(32'hbb7747e1),
	.w2(32'h3b828284),
	.w3(32'hba114010),
	.w4(32'hbb376849),
	.w5(32'h3b1b9ef7),
	.w6(32'hbba0025e),
	.w7(32'h3addea48),
	.w8(32'h3a9605f0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b9d7c),
	.w1(32'hbaa9ed2c),
	.w2(32'hbb3935f3),
	.w3(32'hbb80930a),
	.w4(32'h3bce08b5),
	.w5(32'h3bbb1c64),
	.w6(32'hbae8f6b8),
	.w7(32'h3bbedd4e),
	.w8(32'h3c22ba22),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aafc4d),
	.w1(32'h3889483d),
	.w2(32'hb9dba63f),
	.w3(32'h399567a5),
	.w4(32'hba05cd92),
	.w5(32'hba8ad827),
	.w6(32'h3993c217),
	.w7(32'hbaa098a1),
	.w8(32'hb9a55979),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45d82d),
	.w1(32'hbbf38571),
	.w2(32'hba4c5b05),
	.w3(32'hbc174af9),
	.w4(32'h3a8f5e4a),
	.w5(32'h3c28f825),
	.w6(32'hbb24732b),
	.w7(32'h3b0a1353),
	.w8(32'h3c43480d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34586e),
	.w1(32'h3af5953f),
	.w2(32'h3b27a967),
	.w3(32'hbab22613),
	.w4(32'h3a3b43bd),
	.w5(32'h3abdfc6c),
	.w6(32'h3a984969),
	.w7(32'h3af42a82),
	.w8(32'h39ec4c6f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa2e77a),
	.w1(32'h3a9386ae),
	.w2(32'h3936e8af),
	.w3(32'h392f32f4),
	.w4(32'h3a4d32d9),
	.w5(32'h38a67700),
	.w6(32'h3aaff1ea),
	.w7(32'h390033d1),
	.w8(32'h3a296b2a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8abb1d),
	.w1(32'hbb5cbb3a),
	.w2(32'h3a552be7),
	.w3(32'hbadae3df),
	.w4(32'hbb8eb605),
	.w5(32'hbae8a6b9),
	.w6(32'hba083038),
	.w7(32'h38accb95),
	.w8(32'h3b6223a4),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01d056),
	.w1(32'hbb9b6251),
	.w2(32'h3c08b009),
	.w3(32'hbba38385),
	.w4(32'hbb7927b4),
	.w5(32'h3c483111),
	.w6(32'h3cdfc2e7),
	.w7(32'h3c61e9ed),
	.w8(32'h3cc5ad89),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb987fa8a),
	.w1(32'hbb6d0b35),
	.w2(32'hb9ebb86a),
	.w3(32'hbb2eb9a0),
	.w4(32'hbb35abc2),
	.w5(32'h3ac03c3b),
	.w6(32'hbb024864),
	.w7(32'hbb2b1e81),
	.w8(32'h3a308f88),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd709cb),
	.w1(32'hbb13a655),
	.w2(32'h3af8ca43),
	.w3(32'hb992a273),
	.w4(32'hba943b02),
	.w5(32'h3aa4a339),
	.w6(32'hba499164),
	.w7(32'h3bcc0ad3),
	.w8(32'h3c108308),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e854f),
	.w1(32'h3b406a7f),
	.w2(32'h3b5368e5),
	.w3(32'hbc2cde4e),
	.w4(32'h3b81a775),
	.w5(32'h3bf3dad7),
	.w6(32'hbc2ec99e),
	.w7(32'h3aeabde3),
	.w8(32'h39b52e2f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8f587),
	.w1(32'h3bf503be),
	.w2(32'h3c18de2f),
	.w3(32'hbbad98e1),
	.w4(32'h3b1be977),
	.w5(32'h3b7e2856),
	.w6(32'h3c09257e),
	.w7(32'h3c10a1a7),
	.w8(32'h3ca8c629),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c129794),
	.w1(32'h3b97cb9c),
	.w2(32'h3c84e82e),
	.w3(32'h3abb4c8a),
	.w4(32'hba19539b),
	.w5(32'h3b3927eb),
	.w6(32'h3c17fcc1),
	.w7(32'h3bf9ecdd),
	.w8(32'h3c72ac11),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60e845),
	.w1(32'h3ab20365),
	.w2(32'h3bd0160f),
	.w3(32'hbb061784),
	.w4(32'h3aa6fca6),
	.w5(32'h3bee384b),
	.w6(32'h3c3b4e87),
	.w7(32'h3bdcff00),
	.w8(32'h3c9961d7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18a2ef),
	.w1(32'h3ba22c22),
	.w2(32'h3b9feff0),
	.w3(32'h3b0721a1),
	.w4(32'h3b5a530d),
	.w5(32'h3b8d58dc),
	.w6(32'h3af1809d),
	.w7(32'h3b1260e1),
	.w8(32'hbb5315a4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5f754),
	.w1(32'h3bf76b8f),
	.w2(32'h3b19fc13),
	.w3(32'hbb20ff4a),
	.w4(32'h39b4bade),
	.w5(32'hbb3f2f84),
	.w6(32'h3b292b6f),
	.w7(32'h3b464e5f),
	.w8(32'h3b8d3fd8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72cce6b),
	.w1(32'hba36e833),
	.w2(32'hbaad1d9b),
	.w3(32'hb8652c0e),
	.w4(32'hb9a9ea0b),
	.w5(32'hba99cf3b),
	.w6(32'hba6f6339),
	.w7(32'hbab22412),
	.w8(32'hba18d68a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5429f),
	.w1(32'h3b0837d0),
	.w2(32'h3b167d8a),
	.w3(32'hbb165547),
	.w4(32'h3aa22501),
	.w5(32'h3ae59e08),
	.w6(32'h3b3030ee),
	.w7(32'h3b95a2cb),
	.w8(32'h3b9a104a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad33602),
	.w1(32'hba9021f6),
	.w2(32'hbb0d727a),
	.w3(32'h3aefcb06),
	.w4(32'h3ab4f227),
	.w5(32'h3a77b7f6),
	.w6(32'hbade5bbe),
	.w7(32'hba1f98d5),
	.w8(32'h3b2c5155),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86de49),
	.w1(32'h3b941974),
	.w2(32'h3b7a2e2c),
	.w3(32'h3c0c2887),
	.w4(32'h3b5087cb),
	.w5(32'hbb222dff),
	.w6(32'h3c6ca757),
	.w7(32'h3b942200),
	.w8(32'h3c19e9f8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfe3de),
	.w1(32'h3b1ac4d7),
	.w2(32'hb70cf762),
	.w3(32'hbac9743d),
	.w4(32'h3af1bdae),
	.w5(32'hb9d92838),
	.w6(32'h3b01cf29),
	.w7(32'h3a3b4c9e),
	.w8(32'hba5a9064),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd90b8),
	.w1(32'h3b9609fe),
	.w2(32'h3bac618f),
	.w3(32'hba6a3702),
	.w4(32'h3b373b85),
	.w5(32'h3b72dd2a),
	.w6(32'h3ba07a80),
	.w7(32'h3bbdd15e),
	.w8(32'hb8537deb),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03bef),
	.w1(32'h3b91076a),
	.w2(32'h39b67e6c),
	.w3(32'hbb763678),
	.w4(32'hb9819a84),
	.w5(32'hbb76cece),
	.w6(32'h3b84bfb5),
	.w7(32'h3be173de),
	.w8(32'h3c30983d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c98e46a),
	.w1(32'h3b9f1bad),
	.w2(32'h3c80c069),
	.w3(32'h3bd95b6a),
	.w4(32'hbb09e08c),
	.w5(32'h3b626049),
	.w6(32'h3c41ded7),
	.w7(32'h3b1ba616),
	.w8(32'h3c41ec69),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87f320),
	.w1(32'h3b9c09d7),
	.w2(32'h3bff4929),
	.w3(32'h3b551d5a),
	.w4(32'h3ba66ef6),
	.w5(32'hbae9fcb0),
	.w6(32'h3ba03e71),
	.w7(32'h3b873aeb),
	.w8(32'h3b68de9b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f4f52),
	.w1(32'hb9bb8141),
	.w2(32'h38e8eb79),
	.w3(32'hbab826fd),
	.w4(32'h398d896f),
	.w5(32'h3a94d646),
	.w6(32'h3aea096c),
	.w7(32'h3abd4069),
	.w8(32'h3b276896),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc788f48),
	.w1(32'h3a858a22),
	.w2(32'h3bb8a5d8),
	.w3(32'hbc8a8167),
	.w4(32'hbc25c143),
	.w5(32'h3b5d6029),
	.w6(32'h3c7b1156),
	.w7(32'h3bb6f63d),
	.w8(32'h3cc4bcf6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85aedb),
	.w1(32'h3bc98511),
	.w2(32'h3aa479af),
	.w3(32'hbcb25a80),
	.w4(32'hbb81c357),
	.w5(32'hbc035987),
	.w6(32'hbc9da9ef),
	.w7(32'h3c13049f),
	.w8(32'h3c58116d),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d233),
	.w1(32'h3a163af3),
	.w2(32'h3b1f8045),
	.w3(32'hbb9dd81a),
	.w4(32'hbb3933de),
	.w5(32'h3adaafc7),
	.w6(32'hbb4344c6),
	.w7(32'h3b5b9747),
	.w8(32'h3b911fc6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83c8b2c),
	.w1(32'hbb2180a2),
	.w2(32'hbb57b367),
	.w3(32'hb8924a55),
	.w4(32'hbacee281),
	.w5(32'hbade77a8),
	.w6(32'h3978a088),
	.w7(32'hbaca5beb),
	.w8(32'hbb1230c2),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391af722),
	.w1(32'h3a1dde1c),
	.w2(32'h3a856fd1),
	.w3(32'h3a9f4762),
	.w4(32'h3a9ff157),
	.w5(32'h3b07f4f0),
	.w6(32'hba8893fb),
	.w7(32'hba02cfb8),
	.w8(32'hbb00d345),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba611783),
	.w1(32'hb9b668e1),
	.w2(32'hba533137),
	.w3(32'h39bbe502),
	.w4(32'hba06b5bb),
	.w5(32'hb9c57ad1),
	.w6(32'hb632586e),
	.w7(32'hb9f8f7a7),
	.w8(32'hbaac356c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf59660),
	.w1(32'hbbbc413c),
	.w2(32'h3a7e93ed),
	.w3(32'hbbb7d968),
	.w4(32'h394d9708),
	.w5(32'h3b4a2d54),
	.w6(32'hbae09810),
	.w7(32'h39ac32c0),
	.w8(32'h3b6156f5),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e92afa),
	.w1(32'h3b5a51fc),
	.w2(32'h3b8f8721),
	.w3(32'hbbbebd75),
	.w4(32'hbb51f549),
	.w5(32'h3b0c7504),
	.w6(32'h3c3b1f35),
	.w7(32'h3c0425a1),
	.w8(32'h3c474a3c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfcda9),
	.w1(32'h3ab3e669),
	.w2(32'h3bcf04f2),
	.w3(32'h3bc5aa0d),
	.w4(32'hbbb3ae89),
	.w5(32'hbb98b8f8),
	.w6(32'h3c0db5e9),
	.w7(32'h3c260578),
	.w8(32'h3bba9a12),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03c91f),
	.w1(32'hba003f5d),
	.w2(32'hba94bbfd),
	.w3(32'hbb58ec1b),
	.w4(32'hba77d164),
	.w5(32'hbac0e7c6),
	.w6(32'h3b0fec94),
	.w7(32'hb97313fb),
	.w8(32'h3ad92b35),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba642ab),
	.w1(32'hbb9aafff),
	.w2(32'h3bc42894),
	.w3(32'hbc360ffc),
	.w4(32'hbc07ce1c),
	.w5(32'h3ab3fb3b),
	.w6(32'h3c053278),
	.w7(32'h3b8f3a83),
	.w8(32'h3c796ea6),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0285),
	.w1(32'h3997be9d),
	.w2(32'h3bfe946f),
	.w3(32'hbb16279b),
	.w4(32'hb94fccab),
	.w5(32'h3bb95f34),
	.w6(32'h3b087d02),
	.w7(32'hba150eb2),
	.w8(32'h3aa1cd1c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b5bbd8),
	.w1(32'h3a8db8dd),
	.w2(32'hb9a6699c),
	.w3(32'h39e4a312),
	.w4(32'h3a5ba319),
	.w5(32'hba1dd193),
	.w6(32'h3a74f88d),
	.w7(32'hb604b9ea),
	.w8(32'h3923ec52),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28c18e),
	.w1(32'h3b9d5c26),
	.w2(32'h3b863da5),
	.w3(32'h3a964453),
	.w4(32'h3ae1ce16),
	.w5(32'h39d49f12),
	.w6(32'h3afff7de),
	.w7(32'h3a98ea82),
	.w8(32'hbaeb6562),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3161e),
	.w1(32'h3a0a5e96),
	.w2(32'hba97f238),
	.w3(32'h39129051),
	.w4(32'hb8d2e287),
	.w5(32'hbabd80fd),
	.w6(32'h394207f7),
	.w7(32'hba6e6bf2),
	.w8(32'hba144ef0),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01db76),
	.w1(32'hbb42e775),
	.w2(32'h3c1fb84d),
	.w3(32'hbc2626c9),
	.w4(32'hbb0926ae),
	.w5(32'h3c1e0d87),
	.w6(32'h3b59ed76),
	.w7(32'h3b9f3b34),
	.w8(32'h3c998219),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b333d04),
	.w1(32'hbb77f630),
	.w2(32'h3bade1f1),
	.w3(32'h3b95eb30),
	.w4(32'hbb658168),
	.w5(32'h3b9f9140),
	.w6(32'h3bf6152f),
	.w7(32'h3b89dda9),
	.w8(32'h3c698c38),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc249e),
	.w1(32'hb9df8d7f),
	.w2(32'h3ba7d398),
	.w3(32'h3ba99220),
	.w4(32'hbb2bd7be),
	.w5(32'h3b323e9d),
	.w6(32'h3bf1342f),
	.w7(32'h3bb63661),
	.w8(32'h3c424f13),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb298821),
	.w1(32'hbb89f97a),
	.w2(32'h399263c2),
	.w3(32'hbb2ba9bc),
	.w4(32'hbb520dc0),
	.w5(32'h3a9eb8c2),
	.w6(32'hbb3043cd),
	.w7(32'hbae580e6),
	.w8(32'h3b0587f0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13c1be),
	.w1(32'h3c15c272),
	.w2(32'h3c4d4405),
	.w3(32'hbb0fe2da),
	.w4(32'h3ad786c6),
	.w5(32'h3b9d4a6a),
	.w6(32'h3bcec610),
	.w7(32'h3c5ecae1),
	.w8(32'h3c828f47),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abbf061),
	.w1(32'h3adf4863),
	.w2(32'h3b8c150b),
	.w3(32'hbb947354),
	.w4(32'hba383abe),
	.w5(32'hba87a3e2),
	.w6(32'h3bf8a744),
	.w7(32'h3b6a0c24),
	.w8(32'h3b967492),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd4d9),
	.w1(32'hba646058),
	.w2(32'h3bbea0c1),
	.w3(32'hbb9d9ea6),
	.w4(32'hbb8b05e8),
	.w5(32'h3aa90bd2),
	.w6(32'h3c395165),
	.w7(32'h3c2c40b4),
	.w8(32'h3c509b3f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cfdaf),
	.w1(32'hba59168d),
	.w2(32'h394a2987),
	.w3(32'hb99a78c1),
	.w4(32'hba8095f6),
	.w5(32'hba37d550),
	.w6(32'hbac5ad36),
	.w7(32'hba3a9e15),
	.w8(32'h381ac654),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f8ada2),
	.w1(32'h3b121d01),
	.w2(32'h3ab1bda0),
	.w3(32'h3786a22a),
	.w4(32'h3b099e4f),
	.w5(32'h3b1bf3f3),
	.w6(32'h3ab2fb6a),
	.w7(32'h3a6dd60f),
	.w8(32'h3a960797),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c9404),
	.w1(32'hbbc368e2),
	.w2(32'h3b8e331f),
	.w3(32'hbb59c110),
	.w4(32'hbc2c2691),
	.w5(32'hbaf837ac),
	.w6(32'h3c99454b),
	.w7(32'h3bc266aa),
	.w8(32'h3c4c74e8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5361),
	.w1(32'h3bb3a818),
	.w2(32'h3c86bbc2),
	.w3(32'hbbbf2561),
	.w4(32'h3b93d088),
	.w5(32'h3c9b81e0),
	.w6(32'h3cb74e52),
	.w7(32'h3c6c8d4e),
	.w8(32'h3c9ee97d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2d151),
	.w1(32'h3b8ebad7),
	.w2(32'h3bfc9b5d),
	.w3(32'h3bf5fd74),
	.w4(32'hbb94d2ed),
	.w5(32'hba6a30ea),
	.w6(32'h3c83fa24),
	.w7(32'h3c36e4d0),
	.w8(32'h3c45f079),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19e4c1),
	.w1(32'h3a7b1a30),
	.w2(32'hbbb577bf),
	.w3(32'hbc70cbb7),
	.w4(32'hba058ca6),
	.w5(32'hbb15914d),
	.w6(32'hbb76e1cf),
	.w7(32'h3ab57217),
	.w8(32'h3c2a8635),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03d2e9),
	.w1(32'h39960a57),
	.w2(32'hba1cb6e1),
	.w3(32'h3b5f82e1),
	.w4(32'hb9dbea11),
	.w5(32'hba6dea90),
	.w6(32'h3b83e3bb),
	.w7(32'h3ac7ad5d),
	.w8(32'h3aef333c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b058f71),
	.w1(32'h3bd6123b),
	.w2(32'h3bc1e7b8),
	.w3(32'hb9be5f49),
	.w4(32'h3b0f3ccf),
	.w5(32'h3af43d6a),
	.w6(32'h3bd4f09b),
	.w7(32'h3bb46e83),
	.w8(32'h3a24a665),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2e688),
	.w1(32'hbb7eb7cf),
	.w2(32'h3c5b2237),
	.w3(32'hbb8f829b),
	.w4(32'h3b5d14b9),
	.w5(32'h3c7b4ec9),
	.w6(32'h3c67d603),
	.w7(32'hbba756a0),
	.w8(32'h3c3f00f1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf24a5),
	.w1(32'hb9ad2cdf),
	.w2(32'h3bd015cf),
	.w3(32'hbbd57e53),
	.w4(32'hb98b3698),
	.w5(32'h3bd26b5f),
	.w6(32'h3c7bb7b3),
	.w7(32'h3c0ae30b),
	.w8(32'h3c8fdaee),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1df2ff),
	.w1(32'hbacceb29),
	.w2(32'h3bf4a1d2),
	.w3(32'hbb991db1),
	.w4(32'hbba69a91),
	.w5(32'h3aa0098d),
	.w6(32'h3c8a2487),
	.w7(32'h3a2310e5),
	.w8(32'h3c45f005),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9a4c),
	.w1(32'hbbc0d5e4),
	.w2(32'hba481ef9),
	.w3(32'hbbbbfd34),
	.w4(32'hbaaa10a8),
	.w5(32'h3b7a4a44),
	.w6(32'hbb9e31fb),
	.w7(32'h3bde42ea),
	.w8(32'h3c0b4a5e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3885a9db),
	.w1(32'h3c065db3),
	.w2(32'h3c315814),
	.w3(32'hbb13bcf8),
	.w4(32'h39c52c52),
	.w5(32'h3b7583b7),
	.w6(32'h3b343e53),
	.w7(32'h3c4a9e6d),
	.w8(32'h3c86d47d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35dab0),
	.w1(32'hb99b9cda),
	.w2(32'hb9d628c6),
	.w3(32'h39c44f9e),
	.w4(32'hba9f90e7),
	.w5(32'hbababec1),
	.w6(32'hb9aeb21d),
	.w7(32'hb98a77e0),
	.w8(32'h37a8d576),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d64ce4),
	.w1(32'h3ae30f30),
	.w2(32'hba5e8c0d),
	.w3(32'hbae88964),
	.w4(32'h3b46cff7),
	.w5(32'hb907096f),
	.w6(32'h3a647438),
	.w7(32'hb9bb6e40),
	.w8(32'hbaad2f45),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc244d07),
	.w1(32'hbbfe0c89),
	.w2(32'hbbe7cab2),
	.w3(32'hbb396f79),
	.w4(32'h3a02a41b),
	.w5(32'h3b283875),
	.w6(32'h3a770d38),
	.w7(32'h3b6c227c),
	.w8(32'h3a2b24f4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a64b),
	.w1(32'hb99268f0),
	.w2(32'hba216d49),
	.w3(32'hbb21abe5),
	.w4(32'h3a2bd5f3),
	.w5(32'h3a371ee0),
	.w6(32'h38b951b3),
	.w7(32'h3a0038f1),
	.w8(32'h3ac02f99),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19f7c8),
	.w1(32'hbb9473e5),
	.w2(32'h3b619a1b),
	.w3(32'hba79a267),
	.w4(32'hbb042b39),
	.w5(32'h3b4306bf),
	.w6(32'hbb60e6af),
	.w7(32'hb9ec4b42),
	.w8(32'h3b2d828f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3883a5),
	.w1(32'h3baf2bfd),
	.w2(32'h3ac3c26b),
	.w3(32'hba5a327f),
	.w4(32'hb99c9674),
	.w5(32'h3b0c5127),
	.w6(32'h3ca21299),
	.w7(32'h3c236e24),
	.w8(32'h3c4af859),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb584448),
	.w1(32'hbb51aa03),
	.w2(32'h3ab0b68d),
	.w3(32'hba70041c),
	.w4(32'hbaca3c3e),
	.w5(32'h3984f8dd),
	.w6(32'h3bedf1b4),
	.w7(32'h3bb936c7),
	.w8(32'h3bb1dd5f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65c1de),
	.w1(32'h3ba0aba6),
	.w2(32'h3b87d588),
	.w3(32'hbb61bcfb),
	.w4(32'h3bd18286),
	.w5(32'h3b2a2f17),
	.w6(32'h3ab06fc1),
	.w7(32'h3b4a539e),
	.w8(32'h3a8882b8),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd63c9f),
	.w1(32'hbb4ca489),
	.w2(32'h3c4703a2),
	.w3(32'hba35fe23),
	.w4(32'hbbb236be),
	.w5(32'h3b88c182),
	.w6(32'h3ca51995),
	.w7(32'hbb3dcaae),
	.w8(32'h3c223ee5),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40175c),
	.w1(32'h3aa381a8),
	.w2(32'h3a907c74),
	.w3(32'hbbd6104f),
	.w4(32'hba27301a),
	.w5(32'h3a7f9fb6),
	.w6(32'h3baa45c9),
	.w7(32'h3b0f000f),
	.w8(32'h3c02611d),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e396f),
	.w1(32'h3a080064),
	.w2(32'hba279e28),
	.w3(32'h39a4729e),
	.w4(32'h3a6aff58),
	.w5(32'hb9d8b590),
	.w6(32'hb945c23b),
	.w7(32'hba7a24d9),
	.w8(32'hbab21246),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5ef30),
	.w1(32'hbb405811),
	.w2(32'h3b312a74),
	.w3(32'hbbdbd85a),
	.w4(32'hbafbb544),
	.w5(32'h3b04cdfe),
	.w6(32'h3ba5f12d),
	.w7(32'h3b4f4054),
	.w8(32'h3bf7f558),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba200b30),
	.w1(32'hb98b9162),
	.w2(32'h3998c89d),
	.w3(32'hb96fcc5e),
	.w4(32'hba8d8013),
	.w5(32'hba712d19),
	.w6(32'hba2aba6d),
	.w7(32'hb778ff65),
	.w8(32'hb8ff3404),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b270b),
	.w1(32'h3acf48f4),
	.w2(32'hb9cd0040),
	.w3(32'hbaba5fe9),
	.w4(32'hb98e51cb),
	.w5(32'hbabe39dd),
	.w6(32'h3b279bdc),
	.w7(32'h39b85a51),
	.w8(32'h3ad543cc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc7894),
	.w1(32'h39ada2b2),
	.w2(32'hba3d591a),
	.w3(32'h394832d2),
	.w4(32'h39fb230f),
	.w5(32'hba1f162f),
	.w6(32'hb9f8e251),
	.w7(32'hba8b877a),
	.w8(32'hbac7bfe5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab541d),
	.w1(32'hb9dc0e71),
	.w2(32'h3a042e33),
	.w3(32'hbaacd76a),
	.w4(32'h39066d10),
	.w5(32'h3a77c723),
	.w6(32'hba22ba81),
	.w7(32'h3a098db2),
	.w8(32'h3b0c4ae9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba938afb),
	.w1(32'hbaad7613),
	.w2(32'h391fd24c),
	.w3(32'h3b90e2a3),
	.w4(32'h3b7a841d),
	.w5(32'h3b3d3f4d),
	.w6(32'h3ba379f5),
	.w7(32'h3b8d9bbf),
	.w8(32'h3bac4667),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd82a6e),
	.w1(32'h3b44d179),
	.w2(32'h3bb489fd),
	.w3(32'hbb628ed4),
	.w4(32'h3ae95c29),
	.w5(32'h3b3d1bb4),
	.w6(32'h3c203659),
	.w7(32'h3bf6f296),
	.w8(32'h3c99adb3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab89753),
	.w1(32'h3b287bce),
	.w2(32'h3c16577c),
	.w3(32'h3af389c1),
	.w4(32'h3ad512bd),
	.w5(32'h3b988068),
	.w6(32'h3bd6ccf0),
	.w7(32'h3b52ff8d),
	.w8(32'h3c208bf7),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb670bdf),
	.w1(32'h39baa917),
	.w2(32'h3b74e71b),
	.w3(32'hbc1b2dc6),
	.w4(32'hb94c956e),
	.w5(32'hb9a8b5a2),
	.w6(32'h3b1fcdc9),
	.w7(32'h3b895ff4),
	.w8(32'h3c536bce),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87a889),
	.w1(32'hb8a0e89c),
	.w2(32'h3ae53d5c),
	.w3(32'h3a0bf185),
	.w4(32'hb9a30ecd),
	.w5(32'h3ac723bc),
	.w6(32'h39ec21d6),
	.w7(32'h3ae6a97c),
	.w8(32'h3b04d6b4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9369),
	.w1(32'h39af8940),
	.w2(32'hba2c5946),
	.w3(32'h3ad2b2d0),
	.w4(32'h3ab8bedc),
	.w5(32'hba27b9bb),
	.w6(32'hb846ded8),
	.w7(32'hbad94a6e),
	.w8(32'hbae476e6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaa473),
	.w1(32'h39d84ae6),
	.w2(32'hba87ed28),
	.w3(32'hbac33d9b),
	.w4(32'h39db6795),
	.w5(32'hba6e5426),
	.w6(32'hb6bc54ea),
	.w7(32'hba963e85),
	.w8(32'hba9af9aa),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cb80f),
	.w1(32'h3a36c47d),
	.w2(32'hba80f10b),
	.w3(32'hba80fa46),
	.w4(32'h3a3b82d7),
	.w5(32'hba2a0310),
	.w6(32'h39200029),
	.w7(32'hba91602f),
	.w8(32'hbab47196),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c115cb8),
	.w1(32'h3c14be42),
	.w2(32'h3c11149e),
	.w3(32'h3a647199),
	.w4(32'hba31a5bb),
	.w5(32'h3b8cd36c),
	.w6(32'h3c4127f4),
	.w7(32'h3c0e65ee),
	.w8(32'h3c8d5678),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e3ea6),
	.w1(32'hbae9abd1),
	.w2(32'h39e8431d),
	.w3(32'hba5878de),
	.w4(32'hbabe6042),
	.w5(32'h3a2ce173),
	.w6(32'hbafaa709),
	.w7(32'h3a4fd544),
	.w8(32'hba4da7f2),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c2616),
	.w1(32'hba4a2aae),
	.w2(32'h39814407),
	.w3(32'hbb426fb3),
	.w4(32'hba2d431d),
	.w5(32'h3a29e7be),
	.w6(32'h3a439037),
	.w7(32'hbb323dee),
	.w8(32'hb9d25de0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf98de),
	.w1(32'h3ba545d3),
	.w2(32'h3b89d102),
	.w3(32'h3b4df1f4),
	.w4(32'h3b6826b7),
	.w5(32'h3b2de5a9),
	.w6(32'h3aead469),
	.w7(32'h3a039714),
	.w8(32'h3aa41c90),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f23c4),
	.w1(32'h39e3d9c4),
	.w2(32'hb9dbcabb),
	.w3(32'hb9893b09),
	.w4(32'h39ba3b53),
	.w5(32'hb9f4a55a),
	.w6(32'h397bac36),
	.w7(32'hb9e093d1),
	.w8(32'hb6bab7fc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb272109),
	.w1(32'h3a4823be),
	.w2(32'h3b32bfa7),
	.w3(32'hbb7deae1),
	.w4(32'hb9b046e2),
	.w5(32'hba58f023),
	.w6(32'h3a64fc93),
	.w7(32'h3a7caa93),
	.w8(32'h3b932e9e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fab35f),
	.w1(32'h3b47360f),
	.w2(32'hb80a7535),
	.w3(32'hba2f14f1),
	.w4(32'h3aeef1d6),
	.w5(32'hba0da86f),
	.w6(32'h3b39b353),
	.w7(32'h39727064),
	.w8(32'hbabc8736),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84507),
	.w1(32'h3c3a8229),
	.w2(32'h3bdbc2fb),
	.w3(32'hbbad8d28),
	.w4(32'hb99343a6),
	.w5(32'hbbf4fcc7),
	.w6(32'h3be1cd9e),
	.w7(32'h3bbb05fb),
	.w8(32'h3c37b177),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f92479),
	.w1(32'hb9a917d4),
	.w2(32'hb8996855),
	.w3(32'hba004018),
	.w4(32'h38b04158),
	.w5(32'h397eabae),
	.w6(32'hb8f6a824),
	.w7(32'h380de071),
	.w8(32'h39bd8e5b),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7158d8),
	.w1(32'hbc28e8f0),
	.w2(32'hbc0500b1),
	.w3(32'h3b988bdb),
	.w4(32'hbb586183),
	.w5(32'hbbd1e12e),
	.w6(32'h3c759a36),
	.w7(32'h3bbab8e4),
	.w8(32'h3b3dd487),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule