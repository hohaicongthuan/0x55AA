module layer_10_featuremap_235(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eb698),
	.w1(32'h3b417d02),
	.w2(32'h3c618be3),
	.w3(32'h3b84b582),
	.w4(32'h3bf95fe5),
	.w5(32'h3b80488f),
	.w6(32'hb9cbc7d1),
	.w7(32'hbb3b23b7),
	.w8(32'hbadd7c4f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0dc8),
	.w1(32'h3c537cac),
	.w2(32'h3b0b9ad7),
	.w3(32'hbab6347b),
	.w4(32'h3d3909d5),
	.w5(32'hbbdbb424),
	.w6(32'h3baf497a),
	.w7(32'hbbb7f9f1),
	.w8(32'hbc488a97),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093e12),
	.w1(32'h3a044532),
	.w2(32'h3ae858b3),
	.w3(32'h3c1acb07),
	.w4(32'hbca4ee80),
	.w5(32'h3bba06a7),
	.w6(32'hbb8a8bd6),
	.w7(32'hbae65c88),
	.w8(32'h3b684827),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1bea1),
	.w1(32'hba460f03),
	.w2(32'h3b8928aa),
	.w3(32'hbc302fbf),
	.w4(32'hbb7ca675),
	.w5(32'h3c883206),
	.w6(32'h3b6141eb),
	.w7(32'h3b934e5d),
	.w8(32'hbc12a27c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc17f38),
	.w1(32'h3c462ff8),
	.w2(32'hbae1f52d),
	.w3(32'h3c0b34ad),
	.w4(32'hbbcc969d),
	.w5(32'hb8806971),
	.w6(32'h3c47405a),
	.w7(32'hbb972476),
	.w8(32'hbb81c854),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04eaed),
	.w1(32'h3cd47fb2),
	.w2(32'h3b6976be),
	.w3(32'hbb509bb4),
	.w4(32'h3aa2bd86),
	.w5(32'h3b1e3a76),
	.w6(32'hba9a0a94),
	.w7(32'hbb4ae96d),
	.w8(32'h3c53d822),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0387aa),
	.w1(32'hbc5fe4f2),
	.w2(32'h3caca725),
	.w3(32'hbb4112fd),
	.w4(32'hbbc5bb8c),
	.w5(32'h3b0a26e0),
	.w6(32'hbbe33077),
	.w7(32'h3c027d30),
	.w8(32'hbc4eece9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d334b67),
	.w1(32'h3baf5180),
	.w2(32'hbab84b25),
	.w3(32'hbbffef82),
	.w4(32'hba9633ed),
	.w5(32'h3b05e42f),
	.w6(32'hbbfbbdd0),
	.w7(32'h3c0ef448),
	.w8(32'hbba9b06c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f1825),
	.w1(32'hbbfe4aa0),
	.w2(32'h3abb585d),
	.w3(32'h3c1e2158),
	.w4(32'hbb21a3a1),
	.w5(32'hbb8c4e42),
	.w6(32'h3be75b96),
	.w7(32'hbacec9c2),
	.w8(32'hbac34e38),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943d4b),
	.w1(32'hb80f2df4),
	.w2(32'h3b570d37),
	.w3(32'hbb5bccdb),
	.w4(32'h3aa2d7dc),
	.w5(32'h3bc67533),
	.w6(32'h3bbcd3c6),
	.w7(32'hbb3306b2),
	.w8(32'hbc549dd1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacaaed),
	.w1(32'hbb0f902f),
	.w2(32'h3ba32969),
	.w3(32'h3ca26402),
	.w4(32'h37f19af8),
	.w5(32'h3c05e194),
	.w6(32'hbc089408),
	.w7(32'hbba79f96),
	.w8(32'h38ed1d32),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17160a),
	.w1(32'h3c36aa9f),
	.w2(32'h3bf631ea),
	.w3(32'h38c7b085),
	.w4(32'hbb988721),
	.w5(32'hba859ce4),
	.w6(32'hba9956b9),
	.w7(32'h3658ee65),
	.w8(32'hbb8e48bd),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6e5d6),
	.w1(32'hbba77880),
	.w2(32'hbc4ec2f9),
	.w3(32'hbb556bbb),
	.w4(32'h3ad73cb1),
	.w5(32'hbab65cc4),
	.w6(32'h3c451b8b),
	.w7(32'hbaed5468),
	.w8(32'hbc22dbf5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ead5e),
	.w1(32'h3be807fe),
	.w2(32'h3b75ff10),
	.w3(32'h3b7c242a),
	.w4(32'h3951f177),
	.w5(32'h3c224368),
	.w6(32'h3bcb5e1b),
	.w7(32'h3bf65134),
	.w8(32'h3a3229cb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed7fb),
	.w1(32'hbb17919b),
	.w2(32'hbc0742ca),
	.w3(32'h3b69e655),
	.w4(32'hbb677e76),
	.w5(32'hbbba8bff),
	.w6(32'h3a805fd2),
	.w7(32'h3c423c15),
	.w8(32'h39b6e1ec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f36f8),
	.w1(32'hbb399185),
	.w2(32'hbb6255bd),
	.w3(32'hbbcb663e),
	.w4(32'h390940c6),
	.w5(32'h3bfe9673),
	.w6(32'h3bfbe015),
	.w7(32'h39d11096),
	.w8(32'hbbd22bdc),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80ac27),
	.w1(32'hbbf8ed04),
	.w2(32'h3baefce1),
	.w3(32'h38c83274),
	.w4(32'hb443b8e2),
	.w5(32'h3b442c36),
	.w6(32'hbb342e71),
	.w7(32'h3a03f1c6),
	.w8(32'h3be54e9c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934655),
	.w1(32'h3aeb2689),
	.w2(32'hbc46c60e),
	.w3(32'hbaf0c8d2),
	.w4(32'hba374357),
	.w5(32'hb9eb93e8),
	.w6(32'hbb2d2f71),
	.w7(32'hbb3d0135),
	.w8(32'h3b910310),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e5ac0),
	.w1(32'hb951487c),
	.w2(32'hbab98185),
	.w3(32'hbbed0920),
	.w4(32'h3ba539f6),
	.w5(32'hbb879843),
	.w6(32'h3c66dff6),
	.w7(32'h3b5e30bd),
	.w8(32'h3a97301f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d2a7b),
	.w1(32'hbba2ca52),
	.w2(32'h3c07056f),
	.w3(32'hbb725656),
	.w4(32'h3aca3044),
	.w5(32'hbc0e0e44),
	.w6(32'hba0fbbff),
	.w7(32'hba6ccfd4),
	.w8(32'h3bc7c591),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb88689),
	.w1(32'hbada601b),
	.w2(32'h3c76ac8e),
	.w3(32'h3bdbebdf),
	.w4(32'h39ef48fb),
	.w5(32'h3c2b3650),
	.w6(32'hbbbea2cb),
	.w7(32'h3a9ef2bb),
	.w8(32'h3ca47d61),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a691d),
	.w1(32'hbac645ef),
	.w2(32'h3ba4430c),
	.w3(32'hbb427997),
	.w4(32'hbab9eb00),
	.w5(32'hba085669),
	.w6(32'h3bb0238e),
	.w7(32'h3945fabc),
	.w8(32'hbbc67f72),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3fa6f),
	.w1(32'hba1874bf),
	.w2(32'h3c0215e6),
	.w3(32'h3b7bb2f8),
	.w4(32'h3b58aafb),
	.w5(32'h3c4b9836),
	.w6(32'hbae171b3),
	.w7(32'hbb7ad948),
	.w8(32'h3c591b12),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a8bfd),
	.w1(32'h3c4cc9f3),
	.w2(32'h3c1603bf),
	.w3(32'h3ba9bced),
	.w4(32'h3c7b14a4),
	.w5(32'hbb58fd39),
	.w6(32'h3c8bab03),
	.w7(32'h3bc09b63),
	.w8(32'h3b4d7600),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb832f93),
	.w1(32'h3b9a2ed9),
	.w2(32'h3bf6ef6f),
	.w3(32'hbc0be817),
	.w4(32'hbc0e98fd),
	.w5(32'h3b971c25),
	.w6(32'h3c4743de),
	.w7(32'h3badde33),
	.w8(32'h3c03f36d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcfa5f),
	.w1(32'hbbb0f0a1),
	.w2(32'h3c1f52fa),
	.w3(32'h3b2fec12),
	.w4(32'h3c5cdc10),
	.w5(32'h3c7fb7a2),
	.w6(32'h3c0a8978),
	.w7(32'h3c83cf35),
	.w8(32'h3b66f604),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b9e61),
	.w1(32'h3822934a),
	.w2(32'hba1991c0),
	.w3(32'hbafaaa18),
	.w4(32'h3c26e3bc),
	.w5(32'hba61af99),
	.w6(32'h3b42069c),
	.w7(32'hb904ac14),
	.w8(32'h3c36fcae),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a0c0a),
	.w1(32'hb9ba6872),
	.w2(32'hbba169bc),
	.w3(32'hbc0683e2),
	.w4(32'h3b8cce32),
	.w5(32'h3c27a40b),
	.w6(32'h3ad3371d),
	.w7(32'hbc529b3e),
	.w8(32'hbb66ad67),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9adf8),
	.w1(32'h3bf0d304),
	.w2(32'hbb1b497e),
	.w3(32'h3b98258f),
	.w4(32'h3a14a2f9),
	.w5(32'hbb152c9f),
	.w6(32'hbc4efe5d),
	.w7(32'h3aa22cc5),
	.w8(32'hbbea1994),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c464a96),
	.w1(32'hbb11e64a),
	.w2(32'hbc09631e),
	.w3(32'h3c1a5072),
	.w4(32'h3a68e0c4),
	.w5(32'h3b67ab2a),
	.w6(32'h3c2eb3d2),
	.w7(32'hbc2edd9a),
	.w8(32'h3b48df04),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d6b0d),
	.w1(32'h3b83fe8e),
	.w2(32'h3c4afff3),
	.w3(32'h3c3945de),
	.w4(32'hbb968d6b),
	.w5(32'hbbca19c6),
	.w6(32'h3c08731a),
	.w7(32'h3bad1329),
	.w8(32'hbc15123d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084360),
	.w1(32'hbb949edb),
	.w2(32'h3c481177),
	.w3(32'hbd38dd6d),
	.w4(32'hbb8ca8ee),
	.w5(32'hbc305cc6),
	.w6(32'hbcacdae1),
	.w7(32'h3a7fe2d0),
	.w8(32'h3c096505),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba151c12),
	.w1(32'hbc9698f2),
	.w2(32'hbbf95ab1),
	.w3(32'hbb740968),
	.w4(32'hba881a65),
	.w5(32'hbc0b8fb4),
	.w6(32'hbb6d67f5),
	.w7(32'hbbe51f23),
	.w8(32'hbc3ee257),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a1e56),
	.w1(32'h3c05857e),
	.w2(32'hbb2e0085),
	.w3(32'h3bec4243),
	.w4(32'h3c1734ce),
	.w5(32'hbc105766),
	.w6(32'hba5364b9),
	.w7(32'hbc22b18e),
	.w8(32'hbad543dd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86eafd),
	.w1(32'h3c2a4905),
	.w2(32'h3a958cc5),
	.w3(32'hbb1e770b),
	.w4(32'hbb60ec5c),
	.w5(32'h3c55d1a4),
	.w6(32'hbbd54d82),
	.w7(32'hbc0834f7),
	.w8(32'h3b895f1e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a500),
	.w1(32'h3a852fc4),
	.w2(32'hbc3c0b73),
	.w3(32'h3b8f5157),
	.w4(32'h3c2c539a),
	.w5(32'h3b8f7a7a),
	.w6(32'h3c02385a),
	.w7(32'h3c281c92),
	.w8(32'hbbf0d672),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14220a),
	.w1(32'h3cd29744),
	.w2(32'hbc3107b5),
	.w3(32'hb70e818e),
	.w4(32'hba1cb4a7),
	.w5(32'hbb8969a5),
	.w6(32'hbbcf1e53),
	.w7(32'hbb339d79),
	.w8(32'h3bbbb89e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc46558),
	.w1(32'h393f1166),
	.w2(32'hbc2320ea),
	.w3(32'hbb21b7c2),
	.w4(32'hba6adb0c),
	.w5(32'hb93752e9),
	.w6(32'h3c064ec7),
	.w7(32'h3c52f5ce),
	.w8(32'hbb9b2eea),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf9f3b),
	.w1(32'hbc68706f),
	.w2(32'hbc836bf6),
	.w3(32'hbc165556),
	.w4(32'hbc10c36c),
	.w5(32'h3b27a2c0),
	.w6(32'h3c43cf91),
	.w7(32'h3d1f520f),
	.w8(32'hbb829afb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37d1e4),
	.w1(32'h3b4f1a4e),
	.w2(32'hbc200c89),
	.w3(32'hbaf19f5e),
	.w4(32'hbb175bca),
	.w5(32'h3b632259),
	.w6(32'h3a4ffd74),
	.w7(32'hbc212cfc),
	.w8(32'h3be24ca8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33475a42),
	.w1(32'hbc83cb60),
	.w2(32'h3ce272db),
	.w3(32'h3963d6bf),
	.w4(32'h3d08268f),
	.w5(32'h3bc0c9da),
	.w6(32'h3ab2a33c),
	.w7(32'hbc0b8f24),
	.w8(32'hbb8c7d1e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc250707),
	.w1(32'h3c6c390d),
	.w2(32'hbbf0d9bf),
	.w3(32'hbc020572),
	.w4(32'h3be33f38),
	.w5(32'hbb96d4a7),
	.w6(32'h3c8abb19),
	.w7(32'h3b563b70),
	.w8(32'hbc886a06),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafddf8),
	.w1(32'h3c651505),
	.w2(32'hbbb619d9),
	.w3(32'hba3b558d),
	.w4(32'h3c882f7e),
	.w5(32'h3c1160b8),
	.w6(32'hba6f826c),
	.w7(32'hb975b482),
	.w8(32'h3be7e26d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb57c12),
	.w1(32'h3b5b8c2a),
	.w2(32'h3acaa3ef),
	.w3(32'h3c45dd89),
	.w4(32'hb98fb613),
	.w5(32'hba99cdd0),
	.w6(32'h3b0e3b46),
	.w7(32'hbaf393aa),
	.w8(32'hb9e3d4ff),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc001f31),
	.w1(32'h3b8e0176),
	.w2(32'hbb2bf465),
	.w3(32'hba58fc97),
	.w4(32'hbb702ecc),
	.w5(32'h3a825002),
	.w6(32'hbc18d50a),
	.w7(32'h3c0b0322),
	.w8(32'h35bc66d6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b012b89),
	.w1(32'h3b9f028d),
	.w2(32'hbcb7eb1d),
	.w3(32'hbb883632),
	.w4(32'hbb97ef3f),
	.w5(32'hbb010802),
	.w6(32'hbc0b638b),
	.w7(32'h3c21e55c),
	.w8(32'hbb7e5bdf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba86213),
	.w1(32'hbbcacc75),
	.w2(32'h3c11274b),
	.w3(32'hbc31dcb8),
	.w4(32'hbac0326b),
	.w5(32'hbb98507d),
	.w6(32'h391dafc9),
	.w7(32'h39980e72),
	.w8(32'h39ce0257),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc543e9),
	.w1(32'h39c1bb24),
	.w2(32'hbbe6c58e),
	.w3(32'h3bdaf8f9),
	.w4(32'h3c2dcdf9),
	.w5(32'hbc581090),
	.w6(32'h3b14589b),
	.w7(32'hbbbdbc93),
	.w8(32'h3b8c55c6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf401ee),
	.w1(32'h3a566309),
	.w2(32'hba637d9f),
	.w3(32'hbbbdc26e),
	.w4(32'hbc1853c4),
	.w5(32'h3b0d0372),
	.w6(32'h3c850a4e),
	.w7(32'hbc51bed2),
	.w8(32'hbc600a4a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11afed),
	.w1(32'hbb9dad89),
	.w2(32'hbbff6c9e),
	.w3(32'hbb79f644),
	.w4(32'hbc17ee37),
	.w5(32'hbb538a00),
	.w6(32'hbb51c7dd),
	.w7(32'hba5c83d5),
	.w8(32'h3b81d9f9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d6e81),
	.w1(32'h3c6aa60b),
	.w2(32'h3b71e593),
	.w3(32'hbb6fa0b0),
	.w4(32'hbadf21be),
	.w5(32'hb93895c8),
	.w6(32'hbbc9b4c4),
	.w7(32'hba0400ee),
	.w8(32'hba4554d2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c3c60),
	.w1(32'h395521ad),
	.w2(32'h3c1bded4),
	.w3(32'h3c22015a),
	.w4(32'hba16c99c),
	.w5(32'hbba29da1),
	.w6(32'h3c3c8978),
	.w7(32'hbc040f4e),
	.w8(32'h3babed9a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1a56a),
	.w1(32'hbb783998),
	.w2(32'hbb1b884f),
	.w3(32'hbbd62a67),
	.w4(32'hbbc4cbca),
	.w5(32'hba2fcc1f),
	.w6(32'hbb574263),
	.w7(32'hbc03a6db),
	.w8(32'h39ef18e4),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6e592),
	.w1(32'hbc2bc2cc),
	.w2(32'h3b908048),
	.w3(32'hbb080889),
	.w4(32'hbc36863b),
	.w5(32'h3b3e6d14),
	.w6(32'h3be7b951),
	.w7(32'h3c00a6bb),
	.w8(32'h3be3d7bd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c6b6),
	.w1(32'hbb93bfbf),
	.w2(32'hbb31f8f0),
	.w3(32'h3bfe32a7),
	.w4(32'hbaad8ef0),
	.w5(32'h3b20b573),
	.w6(32'hbb839a9e),
	.w7(32'h3bde4df3),
	.w8(32'h3bd07879),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e7289),
	.w1(32'h3b467f51),
	.w2(32'hbb331b45),
	.w3(32'hba875752),
	.w4(32'h3bc240da),
	.w5(32'hbb850e24),
	.w6(32'h39e2876f),
	.w7(32'hbcb2f95b),
	.w8(32'h3b8a18ac),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1e38),
	.w1(32'h3c1c2767),
	.w2(32'hbcfffb0c),
	.w3(32'hbbc6355b),
	.w4(32'h3c4598fc),
	.w5(32'h3c9412ce),
	.w6(32'hbb8434d9),
	.w7(32'hbba39b7e),
	.w8(32'hbbe4e011),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66bec9),
	.w1(32'hbb9dc231),
	.w2(32'hbb79137a),
	.w3(32'h3af0cfcc),
	.w4(32'h3c388054),
	.w5(32'h3a631971),
	.w6(32'hbb91756a),
	.w7(32'h3c61011f),
	.w8(32'hbbf328f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc832edd),
	.w1(32'hbcc3e704),
	.w2(32'hbb85f414),
	.w3(32'h3c530528),
	.w4(32'h3bdbfb0e),
	.w5(32'hbc6d295e),
	.w6(32'h3cc6d653),
	.w7(32'hbc02582b),
	.w8(32'h3c431f5a),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ae1d7),
	.w1(32'hbc0c7ba4),
	.w2(32'h39bfe0b1),
	.w3(32'hbc227dc6),
	.w4(32'hbbb332cf),
	.w5(32'hbcdd8692),
	.w6(32'hbc80c9ba),
	.w7(32'hbc51101b),
	.w8(32'h3b7e869d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd57d9e),
	.w1(32'hbc88a20e),
	.w2(32'hbbf891d2),
	.w3(32'h383aa962),
	.w4(32'hbc0b01ee),
	.w5(32'hbbd872a3),
	.w6(32'hbc46181c),
	.w7(32'hbba47178),
	.w8(32'h3c7e1a8b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba380aed),
	.w1(32'hbb5063be),
	.w2(32'hbab773ca),
	.w3(32'hba6c7fcd),
	.w4(32'hbc39ea05),
	.w5(32'hbac473ea),
	.w6(32'hbb60b515),
	.w7(32'h3a7a64e4),
	.w8(32'h3c69c322),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b64d9),
	.w1(32'h399a3d21),
	.w2(32'h3a175ac3),
	.w3(32'h3a304281),
	.w4(32'hbca4449b),
	.w5(32'hbbc953eb),
	.w6(32'hbbba5f95),
	.w7(32'hbbe75dd9),
	.w8(32'hbb9ffc92),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c92c5),
	.w1(32'h3c31cccd),
	.w2(32'h3b84e196),
	.w3(32'hbb5ce965),
	.w4(32'hbc849fbe),
	.w5(32'h3b3348c9),
	.w6(32'h3bc1c293),
	.w7(32'hbb3584e4),
	.w8(32'h3c27e702),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc123d17),
	.w1(32'hb9d1268a),
	.w2(32'h3bb87131),
	.w3(32'hbc651491),
	.w4(32'h3cb74a38),
	.w5(32'h3c0222fc),
	.w6(32'h3bfb2d6e),
	.w7(32'h3b9a319c),
	.w8(32'hbbb7640b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95fd5d),
	.w1(32'hbbb9c1c9),
	.w2(32'hbba56ff4),
	.w3(32'h3b391740),
	.w4(32'hbc183b36),
	.w5(32'hba9a4883),
	.w6(32'hbc043de3),
	.w7(32'hba662e9d),
	.w8(32'hbb7ea976),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c735e),
	.w1(32'h3c8654e8),
	.w2(32'h3bd4b196),
	.w3(32'h3907f040),
	.w4(32'hbc3b0f2f),
	.w5(32'hbcce7dde),
	.w6(32'hb99e58cf),
	.w7(32'h3cf1c2ed),
	.w8(32'hbbb6ecfd),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad014c),
	.w1(32'h3a5a15d0),
	.w2(32'hbb8c5654),
	.w3(32'hbb8ec9ff),
	.w4(32'hbba27a79),
	.w5(32'h3c66b6ac),
	.w6(32'hbc226cb9),
	.w7(32'hbc212df3),
	.w8(32'h3a87cde4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42362),
	.w1(32'h3b080525),
	.w2(32'hb9a53750),
	.w3(32'hbbad8ddf),
	.w4(32'hb5adc1ef),
	.w5(32'h3cbbe065),
	.w6(32'hb952c941),
	.w7(32'hbaaad763),
	.w8(32'h3c80ad46),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10d0c5),
	.w1(32'hbbff1363),
	.w2(32'h3ca933ad),
	.w3(32'hbbdb5651),
	.w4(32'hbb9b1731),
	.w5(32'h39f7a84b),
	.w6(32'hbb6d9f5d),
	.w7(32'hbbe8ba1e),
	.w8(32'h3b828628),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83782),
	.w1(32'h3c479562),
	.w2(32'hbc3adae3),
	.w3(32'h3b47c691),
	.w4(32'h3b926e63),
	.w5(32'h391fcde9),
	.w6(32'h391b4359),
	.w7(32'h3ccf1e4b),
	.w8(32'hbbf7c5fd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99fb69),
	.w1(32'hbc3b022a),
	.w2(32'h3c83713b),
	.w3(32'hbc83e8ad),
	.w4(32'h3b446241),
	.w5(32'hba8bc369),
	.w6(32'hbc70b37b),
	.w7(32'hbc416256),
	.w8(32'hbcb1e528),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2918),
	.w1(32'hbc1ec18b),
	.w2(32'hbc05e2d7),
	.w3(32'hbc1d0ece),
	.w4(32'h3c6ab52f),
	.w5(32'hbc246f98),
	.w6(32'hbc7723b4),
	.w7(32'hbbeeafe8),
	.w8(32'hbbbaff74),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3661c6),
	.w1(32'h355251f0),
	.w2(32'hb8cb22fe),
	.w3(32'h3a2059f7),
	.w4(32'hbc8d96b0),
	.w5(32'h3cedc506),
	.w6(32'h3b6549f2),
	.w7(32'h3bd656fd),
	.w8(32'hbc8f5ea6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ab25),
	.w1(32'hbc9c3d27),
	.w2(32'hba331654),
	.w3(32'h3c9943d5),
	.w4(32'h3b96c09d),
	.w5(32'h3a1e3621),
	.w6(32'hbb18febc),
	.w7(32'hbbca4126),
	.w8(32'hbafffa1c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91f140),
	.w1(32'hbcb1e334),
	.w2(32'hbc5f241e),
	.w3(32'hbc1bcf02),
	.w4(32'h3b414564),
	.w5(32'hbc2b992e),
	.w6(32'h3bb8b688),
	.w7(32'hbbe8b9a1),
	.w8(32'hbb3c6426),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2517bf),
	.w1(32'hbcc5871d),
	.w2(32'hbb1a1ca3),
	.w3(32'hbc49eae5),
	.w4(32'hbca040bc),
	.w5(32'hbb20e753),
	.w6(32'hbb3d76be),
	.w7(32'h3c61a336),
	.w8(32'hbbb3ff37),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebc788),
	.w1(32'hbc28151e),
	.w2(32'h3cfc96cb),
	.w3(32'h3c096443),
	.w4(32'h3c15e76e),
	.w5(32'h3aa37919),
	.w6(32'hbbe2f0c4),
	.w7(32'h3bfc55b9),
	.w8(32'hbbb85c83),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb38f2),
	.w1(32'hbb219f2c),
	.w2(32'hbc4bbc14),
	.w3(32'h3be0e241),
	.w4(32'h3a12ad9f),
	.w5(32'hbc512d65),
	.w6(32'h3ca7932f),
	.w7(32'hbc147db6),
	.w8(32'hbcb1a8bc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510978),
	.w1(32'hbbea94cf),
	.w2(32'h3c9b157c),
	.w3(32'h3af21847),
	.w4(32'h3bac3c9b),
	.w5(32'h3c94b3f1),
	.w6(32'hb8ace1ae),
	.w7(32'hbc5e911e),
	.w8(32'hbbf6bdc8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f253),
	.w1(32'hbccb9e23),
	.w2(32'hbbd20918),
	.w3(32'hbc9c22e2),
	.w4(32'hbcabb654),
	.w5(32'hbc1d2760),
	.w6(32'hbc85008d),
	.w7(32'h3cf6af60),
	.w8(32'hbc89cb3c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c6edd),
	.w1(32'hbc12a58d),
	.w2(32'hbc74e379),
	.w3(32'h3bcc1799),
	.w4(32'hbb10eb8d),
	.w5(32'h3b0239a2),
	.w6(32'hbbbcc5c6),
	.w7(32'hbb9ad073),
	.w8(32'h3bf6cc9f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267aad),
	.w1(32'hbc138d24),
	.w2(32'h3c2e1232),
	.w3(32'h391d1e47),
	.w4(32'hba53b8ae),
	.w5(32'h3c33ac45),
	.w6(32'hbcf73c81),
	.w7(32'h3be704b0),
	.w8(32'hbd78bace),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31ccdf),
	.w1(32'h3bd3178b),
	.w2(32'h3bbbb308),
	.w3(32'h3b89e01f),
	.w4(32'hbbebd186),
	.w5(32'hb8eba059),
	.w6(32'hbbc6297a),
	.w7(32'hbb6a02f4),
	.w8(32'hba1d22a3),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bdb1d),
	.w1(32'hbb898624),
	.w2(32'hbc0a1a02),
	.w3(32'h3ba58add),
	.w4(32'hbc386e16),
	.w5(32'hbba27efe),
	.w6(32'hbc5901f3),
	.w7(32'h3b875ed8),
	.w8(32'h3bc8abe0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b9d9b),
	.w1(32'h3a8c61aa),
	.w2(32'h3b7ccf9c),
	.w3(32'hba82ad2a),
	.w4(32'hba371fe5),
	.w5(32'h399cb665),
	.w6(32'h3bcb676a),
	.w7(32'hbc7383a6),
	.w8(32'h3b8c4ce5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bceddcb),
	.w1(32'h3c59e2ba),
	.w2(32'hbc8b7cb6),
	.w3(32'h3c4b6a3d),
	.w4(32'hbc58eac9),
	.w5(32'h3b05b5da),
	.w6(32'h3c8dd081),
	.w7(32'h3c9a394c),
	.w8(32'hbc76a66c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cbe20),
	.w1(32'hbb225a9f),
	.w2(32'h3ba0e6a1),
	.w3(32'hbbc01d75),
	.w4(32'h3ac318cc),
	.w5(32'h39748b63),
	.w6(32'hbb19d77a),
	.w7(32'hbc8336f8),
	.w8(32'h3b3208bd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49289d),
	.w1(32'hbc641141),
	.w2(32'hbbc3a480),
	.w3(32'h3b9b4dbc),
	.w4(32'hbc30b65f),
	.w5(32'hbc1d5685),
	.w6(32'hbbe0dc53),
	.w7(32'hbbcd6847),
	.w8(32'h3c259884),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1edc69),
	.w1(32'hbc3c35b3),
	.w2(32'hbc3ea94f),
	.w3(32'h3bcea094),
	.w4(32'h3af8d3a6),
	.w5(32'hba9566ea),
	.w6(32'hbb3d51db),
	.w7(32'h3c14103d),
	.w8(32'hbb312aa4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133fa5),
	.w1(32'h3c443336),
	.w2(32'h3cb6fec8),
	.w3(32'hba9b181b),
	.w4(32'h3ad5b9a3),
	.w5(32'h39ca68f1),
	.w6(32'h3d29c787),
	.w7(32'h3c7141e9),
	.w8(32'h3b8d2e61),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa377f5),
	.w1(32'h3b144e38),
	.w2(32'hbb7a9b9a),
	.w3(32'h3c1617dd),
	.w4(32'hbc66b1c5),
	.w5(32'h3c7558ac),
	.w6(32'hbc4a5f05),
	.w7(32'hbc38ed48),
	.w8(32'h3bf48472),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1811b6),
	.w1(32'hbb1cbc6b),
	.w2(32'h3bc83e9d),
	.w3(32'hbb89f18b),
	.w4(32'hbc471c67),
	.w5(32'hba1361b8),
	.w6(32'hbc2a60f9),
	.w7(32'hbab636ba),
	.w8(32'hbb91fa0b),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca59427),
	.w1(32'h3ce0f46e),
	.w2(32'h39c9c2d2),
	.w3(32'hbb39b35d),
	.w4(32'h3a44b6b9),
	.w5(32'hbb959910),
	.w6(32'hbc9004cc),
	.w7(32'hbb291b0f),
	.w8(32'h3b639afb),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce9cdc),
	.w1(32'hbc1664a8),
	.w2(32'hb98ff4ba),
	.w3(32'hbb5ae5e1),
	.w4(32'hbba276c0),
	.w5(32'h3b39d962),
	.w6(32'hbbc04601),
	.w7(32'h3bdef17d),
	.w8(32'h3aafe9ed),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c399681),
	.w1(32'hbb6721a9),
	.w2(32'hbb0b448b),
	.w3(32'hbc08e969),
	.w4(32'hbac625a8),
	.w5(32'hb93d7e63),
	.w6(32'h3a45d549),
	.w7(32'h3bbcb7b7),
	.w8(32'hbb2aabde),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8a2b),
	.w1(32'hbbaa475d),
	.w2(32'h3b7daab6),
	.w3(32'h3be10e0e),
	.w4(32'h3c4cb604),
	.w5(32'h3c1dd837),
	.w6(32'hb949cfb6),
	.w7(32'hbb9f7025),
	.w8(32'hb4275416),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4271c2),
	.w1(32'hbc554589),
	.w2(32'hbae13e8c),
	.w3(32'hb9807023),
	.w4(32'h3a1ba0a3),
	.w5(32'hbb19f466),
	.w6(32'h3c756b23),
	.w7(32'h3c4a3688),
	.w8(32'h3a96f83c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c170ee1),
	.w1(32'h3c9220fa),
	.w2(32'h3c653bd7),
	.w3(32'h3cb558cc),
	.w4(32'hbbf7b8ea),
	.w5(32'hba0d2421),
	.w6(32'h3b40c948),
	.w7(32'hbc5e4c39),
	.w8(32'hbaf57c34),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ba7f0),
	.w1(32'h3be7a2fc),
	.w2(32'hba5e5df5),
	.w3(32'hbccc16da),
	.w4(32'hbb836bb2),
	.w5(32'h3c1ce121),
	.w6(32'hbb9e7933),
	.w7(32'hbba7fcf4),
	.w8(32'hbc80a185),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b630756),
	.w1(32'hbbaae2e5),
	.w2(32'hbbcefdae),
	.w3(32'hbbe512cb),
	.w4(32'hbc20fe92),
	.w5(32'h3b8ff24c),
	.w6(32'h3b0c7590),
	.w7(32'hb95793f8),
	.w8(32'hbbc29175),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc302c8f),
	.w1(32'h3b840e22),
	.w2(32'hba88891a),
	.w3(32'hbaaf14b8),
	.w4(32'h3ade1925),
	.w5(32'hb584171b),
	.w6(32'h3cdc3b0c),
	.w7(32'hbbca24cc),
	.w8(32'h3ca340b5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085180),
	.w1(32'h3a97b861),
	.w2(32'hba71c5e2),
	.w3(32'h3b0343ef),
	.w4(32'hbc0245ac),
	.w5(32'h3b8388d0),
	.w6(32'hbbbd955f),
	.w7(32'h3d37c37f),
	.w8(32'h3cf5bb6d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87e941),
	.w1(32'h3c5ccc47),
	.w2(32'hbbecb2a5),
	.w3(32'h3acd737b),
	.w4(32'h3acc2e04),
	.w5(32'h3b800c6f),
	.w6(32'h3c3ad0bd),
	.w7(32'hbb5a793f),
	.w8(32'h3b828b1f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd0526),
	.w1(32'hbc2749cb),
	.w2(32'h39289269),
	.w3(32'hbc51c8de),
	.w4(32'hbbbe222e),
	.w5(32'hbd68ae55),
	.w6(32'h3bcd0bda),
	.w7(32'h3c19e129),
	.w8(32'h3b2aec01),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc033fef),
	.w1(32'h3cab7283),
	.w2(32'hbb95326d),
	.w3(32'hbb2098ad),
	.w4(32'hbc478607),
	.w5(32'hbc32c356),
	.w6(32'hbbe0482c),
	.w7(32'hbbfe8993),
	.w8(32'hbc1f1e59),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd212ee2),
	.w1(32'hbc1dbe81),
	.w2(32'hbb040cf4),
	.w3(32'hbc15bdaa),
	.w4(32'h3b69beec),
	.w5(32'h3af288e5),
	.w6(32'h3ce4852c),
	.w7(32'hbbbb8c71),
	.w8(32'hb9455ae8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10691a),
	.w1(32'h3bbe915c),
	.w2(32'hb9834d88),
	.w3(32'hba88bed0),
	.w4(32'hbb37b179),
	.w5(32'hbae2c6d1),
	.w6(32'h3a4bf1c8),
	.w7(32'h3b9589f6),
	.w8(32'h39e20927),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72fe9),
	.w1(32'hbc13c21d),
	.w2(32'h3cc1b5f4),
	.w3(32'h3c2e5958),
	.w4(32'h3b420ae7),
	.w5(32'hbab2a126),
	.w6(32'hbc885e63),
	.w7(32'h3b8c552f),
	.w8(32'hbbbde866),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc440321),
	.w1(32'h3a6e9ae0),
	.w2(32'hbc760dc9),
	.w3(32'h3b82d8b2),
	.w4(32'hbbef9140),
	.w5(32'hbbc11f08),
	.w6(32'hbb201dd9),
	.w7(32'h3a9ee8cc),
	.w8(32'h3c7862ec),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2b666),
	.w1(32'h3c882a27),
	.w2(32'hbc61a7a9),
	.w3(32'h3c1e3149),
	.w4(32'h3b05213a),
	.w5(32'hbc408d7b),
	.w6(32'h3b890bbf),
	.w7(32'h3a50b23f),
	.w8(32'h3c17f214),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81af10),
	.w1(32'hbb61318d),
	.w2(32'hbbad7019),
	.w3(32'h3b4edb64),
	.w4(32'hbbdd3421),
	.w5(32'h3b9f67e3),
	.w6(32'hba1a675b),
	.w7(32'h3bea9016),
	.w8(32'h3b9e1937),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2a55a6),
	.w1(32'hbf0acf14),
	.w2(32'hbf87581f),
	.w3(32'hbe65369f),
	.w4(32'hbf02f6cc),
	.w5(32'hbf21b9fc),
	.w6(32'hbf04b66f),
	.w7(32'hbe92f13f),
	.w8(32'hbe49b015),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf08c8dd),
	.w1(32'hbddb0af2),
	.w2(32'hbe7b38a8),
	.w3(32'hbeee8101),
	.w4(32'hbed2d143),
	.w5(32'hbf09c315),
	.w6(32'hbf1c6c56),
	.w7(32'h3e81d645),
	.w8(32'hbf3062ae),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef8b97a),
	.w1(32'hbf0c8d48),
	.w2(32'hbdbc3c51),
	.w3(32'hbf16cc95),
	.w4(32'hbf157afa),
	.w5(32'hbf3178c4),
	.w6(32'hbf032891),
	.w7(32'hbe86b1ae),
	.w8(32'h3ee9ac52),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1a36e8),
	.w1(32'hbf131980),
	.w2(32'hbea34e68),
	.w3(32'hbf1ee495),
	.w4(32'hbea45c24),
	.w5(32'hbf07ea6e),
	.w6(32'hbd2e5952),
	.w7(32'hbf09325e),
	.w8(32'hbf303e98),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf336808),
	.w1(32'hbf06cc37),
	.w2(32'hbef4512d),
	.w3(32'hbf470e33),
	.w4(32'hbe3ddac2),
	.w5(32'h3e0867fc),
	.w6(32'hbf05220a),
	.w7(32'hbf2de3c9),
	.w8(32'hbeb3e542),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1d8b98),
	.w1(32'hbd11d036),
	.w2(32'hbdfb71e2),
	.w3(32'hbf06cc80),
	.w4(32'hbf1ecc2e),
	.w5(32'hbf206c9b),
	.w6(32'hbf026a14),
	.w7(32'hbf3148cf),
	.w8(32'hbf183fb7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeee098e),
	.w1(32'hbd0bbec4),
	.w2(32'hbf267bb5),
	.w3(32'hbf160d11),
	.w4(32'hbf0ced19),
	.w5(32'hbf15ecf4),
	.w6(32'hbf3e92b9),
	.w7(32'hbf175662),
	.w8(32'hbd6df867),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb2a1f8),
	.w1(32'hbefe16ca),
	.w2(32'hbefc53eb),
	.w3(32'hbf5bfcf8),
	.w4(32'hbed0bbeb),
	.w5(32'h3d3b7617),
	.w6(32'hbf288a66),
	.w7(32'hbebac4f1),
	.w8(32'hbf26fca4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf12154f),
	.w1(32'hbf178b97),
	.w2(32'hbed8025e),
	.w3(32'hbf014fe5),
	.w4(32'hbe88f2c6),
	.w5(32'hbf1e2cd3),
	.w6(32'hbf834ada),
	.w7(32'hbf107241),
	.w8(32'hbefa4347),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe97a3f4),
	.w1(32'hbf10d817),
	.w2(32'hbf314a1c),
	.w3(32'hbe25a1ec),
	.w4(32'hbf2199ad),
	.w5(32'hbe8e73a8),
	.w6(32'hbf3dea14),
	.w7(32'hbe6f3a7f),
	.w8(32'hbdce4216),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf17256c),
	.w1(32'hbe3a1b2c),
	.w2(32'hbec86746),
	.w3(32'hbede8484),
	.w4(32'hbf157da4),
	.w5(32'hbf0eba56),
	.w6(32'hbec19c12),
	.w7(32'hbef821b3),
	.w8(32'hbee45764),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbee43181),
	.w1(32'hbed593fa),
	.w2(32'hbf13cc1d),
	.w3(32'h3d12243f),
	.w4(32'h3f5634a8),
	.w5(32'hbf0699d7),
	.w6(32'hbf107ed0),
	.w7(32'hbf004b46),
	.w8(32'hbe9d077a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe8d95ec),
	.w1(32'hbebdaab5),
	.w2(32'h3f486e4b),
	.w3(32'hbf36af0b),
	.w4(32'hbf35a21c),
	.w5(32'hbf13094f),
	.w6(32'hbf32e85a),
	.w7(32'hbf6c114b),
	.w8(32'hbf04d817),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2db162),
	.w1(32'hbefd70a7),
	.w2(32'hbe8801c0),
	.w3(32'hbe424662),
	.w4(32'hbf1914b8),
	.w5(32'h3d6150e2),
	.w6(32'hbf9589ad),
	.w7(32'hbec0e6cf),
	.w8(32'hbf0002d9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4b285b),
	.w1(32'hbf179e1f),
	.w2(32'hbf0c49a7),
	.w3(32'hbe888b34),
	.w4(32'hbdb57e3e),
	.w5(32'hbf1b320d),
	.w6(32'hbeb63a2c),
	.w7(32'hbeb271b6),
	.w8(32'hbefab849),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1069e6),
	.w1(32'hbf0856a8),
	.w2(32'hbed828fc),
	.w3(32'hbeb3c186),
	.w4(32'hbf052ac2),
	.w5(32'hbeeee55a),
	.w6(32'hbfa497dc),
	.w7(32'hbef70409),
	.w8(32'hbeabd37b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd40360),
	.w1(32'hbf267b5c),
	.w2(32'hbcf4a295),
	.w3(32'hbeebbda4),
	.w4(32'h3b9d6908),
	.w5(32'hbf141b4f),
	.w6(32'hbf0e9ad1),
	.w7(32'hbecafb00),
	.w8(32'hbf1984c8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe9a140e),
	.w1(32'hbf163cf5),
	.w2(32'hbf424f04),
	.w3(32'hbe38628e),
	.w4(32'hbba784ec),
	.w5(32'hbf0b3fc4),
	.w6(32'hbf12ba8d),
	.w7(32'hbef5e94c),
	.w8(32'hbf28d063),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe83d61c),
	.w1(32'hbede0f88),
	.w2(32'hbf0b26c2),
	.w3(32'hbe3e832a),
	.w4(32'hbef7fa75),
	.w5(32'h3e84ad6e),
	.w6(32'hbf1b7627),
	.w7(32'hbe922ba4),
	.w8(32'hbed1509c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0dff18),
	.w1(32'hbf22fabd),
	.w2(32'hbedd3170),
	.w3(32'hbf58e556),
	.w4(32'hbeedc18d),
	.w5(32'hbefc9a9f),
	.w6(32'h3d3857e1),
	.w7(32'hbea4fab2),
	.w8(32'hbf304c8e),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe73ebdf),
	.w1(32'hbef3755d),
	.w2(32'hbebbfb14),
	.w3(32'hbf1a9b41),
	.w4(32'hbf03d2f6),
	.w5(32'hbf00bf73),
	.w6(32'hbe973292),
	.w7(32'hbf2f9764),
	.w8(32'hbec2aff3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1eeb9f),
	.w1(32'h3cefc137),
	.w2(32'hbf2c8293),
	.w3(32'hbf2d8d2c),
	.w4(32'hbeca6c1c),
	.w5(32'hbf2a974d),
	.w6(32'hbf913184),
	.w7(32'hbd41b732),
	.w8(32'hbed50e54),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe4c1e6f),
	.w1(32'hbefc72a7),
	.w2(32'hbf091bdb),
	.w3(32'hbe0731a1),
	.w4(32'hbf0810bb),
	.w5(32'hbeb51cb1),
	.w6(32'hbf0ec586),
	.w7(32'h3eaff79f),
	.w8(32'hbee76a68),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe5c7f8f),
	.w1(32'hbe5f95fe),
	.w2(32'hbecbcbd3),
	.w3(32'hbf269504),
	.w4(32'hbf2b9931),
	.w5(32'hbf1806ff),
	.w6(32'hbf2b751f),
	.w7(32'hbf043294),
	.w8(32'hbf30d72c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe8e1a2a),
	.w1(32'hbed1a0ce),
	.w2(32'hbf2708c3),
	.w3(32'hbef4f3ea),
	.w4(32'hbefc4972),
	.w5(32'hbf2fb7e6),
	.w6(32'hbe54c4b7),
	.w7(32'hbf1c18a6),
	.w8(32'hbeefbf96),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3de50723),
	.w1(32'hbf0562a4),
	.w2(32'hbee50631),
	.w3(32'hbcb77588),
	.w4(32'hbf0ff7f1),
	.w5(32'hbe284ba2),
	.w6(32'hbe8df6a5),
	.w7(32'hbefeeeb7),
	.w8(32'hbefc4980),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeee9c2f),
	.w1(32'hbef31be8),
	.w2(32'hbeedb46e),
	.w3(32'hbee0cad8),
	.w4(32'hbefe4c39),
	.w5(32'hbe7d8b79),
	.w6(32'hbf1adb69),
	.w7(32'hbf062f52),
	.w8(32'hbf21f232),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec30742),
	.w1(32'hbf6348b6),
	.w2(32'hbe9c937e),
	.w3(32'h3c80cbe1),
	.w4(32'hbcd445fe),
	.w5(32'h3cabc0e2),
	.w6(32'hbf1a5232),
	.w7(32'hbf1a5c46),
	.w8(32'hbed26ac5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef0fea6),
	.w1(32'hbee979b3),
	.w2(32'h3e5237ee),
	.w3(32'hbef3881a),
	.w4(32'h3e6c4e59),
	.w5(32'h3dd7d669),
	.w6(32'hbed9b97e),
	.w7(32'h3e675d96),
	.w8(32'h3eed0de6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e3efc47),
	.w1(32'h36495776),
	.w2(32'h3e80e917),
	.w3(32'h3f964bf9),
	.w4(32'h3a4fe785),
	.w5(32'h3e893b81),
	.w6(32'h3892a7e0),
	.w7(32'h3f2aa0c7),
	.w8(32'h3f521801),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e5e20f9),
	.w1(32'h3e8adc4c),
	.w2(32'h3d8709b6),
	.w3(32'h3e938848),
	.w4(32'h3f2c8dbb),
	.w5(32'h3e566e62),
	.w6(32'h3f0bc7b5),
	.w7(32'hb87bbe3d),
	.w8(32'h3e370825),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dab42c3),
	.w1(32'h3ea21cb8),
	.w2(32'h3f10dc4a),
	.w3(32'h3e9f7906),
	.w4(32'h3e88254c),
	.w5(32'h3f338150),
	.w6(32'h3f4383af),
	.w7(32'h3e617912),
	.w8(32'h3f1a9ff2),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e61d0c2),
	.w1(32'h3fabba2d),
	.w2(32'h3f523167),
	.w3(32'h3ecffadb),
	.w4(32'h3ed61a91),
	.w5(32'h3e3457d1),
	.w6(32'h3e548eaa),
	.w7(32'h3eb3407e),
	.w8(32'h3f6cb859),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e4f01b0),
	.w1(32'h3e89d0ac),
	.w2(32'h3d321ff6),
	.w3(32'h3eb3595a),
	.w4(32'h3f72a5c7),
	.w5(32'h3ea034d6),
	.w6(32'h3f69a784),
	.w7(32'h3f1d0463),
	.w8(32'h3e531a4e),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f025db6),
	.w1(32'h3f08bf9a),
	.w2(32'h3faee9a9),
	.w3(32'h3f148ba7),
	.w4(32'h3f010bc5),
	.w5(32'h3dd5b1e0),
	.w6(32'h3ed13bec),
	.w7(32'hb6385311),
	.w8(32'h3e8d752f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e37dffd),
	.w1(32'h3e2773ea),
	.w2(32'h3eba9fd4),
	.w3(32'h3f28263f),
	.w4(32'hb7540579),
	.w5(32'h3eb512c2),
	.w6(32'h3e0c7536),
	.w7(32'h3f86f8a4),
	.w8(32'h3ea83eef),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f780d43),
	.w1(32'h3f12a616),
	.w2(32'h3f707f7a),
	.w3(32'h3eff7cea),
	.w4(32'h3ef1fce2),
	.w5(32'h3db8b75d),
	.w6(32'h3f0a4dd2),
	.w7(32'h3ea7f95b),
	.w8(32'h3ed63c6b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e237753),
	.w1(32'h3e9aede2),
	.w2(32'h3f80faf7),
	.w3(32'h3d256585),
	.w4(32'h3f415112),
	.w5(32'h3f023170),
	.w6(32'h3dac3877),
	.w7(32'h3ee7e64d),
	.w8(32'h37e7d859),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3ec260),
	.w1(32'h3f15acac),
	.w2(32'h3f2dbbb6),
	.w3(32'h3f6742a3),
	.w4(32'h3903b94b),
	.w5(32'h3eba3500),
	.w6(32'h3d856576),
	.w7(32'h3f2703b0),
	.w8(32'h3d561e9e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ed54e66),
	.w1(32'h3f03ab5d),
	.w2(32'h3e6ffa39),
	.w3(32'h3e9aba3c),
	.w4(32'h3f052ee7),
	.w5(32'h3d3f134c),
	.w6(32'h3eafa1f9),
	.w7(32'h3e191cf3),
	.w8(32'h3f86efe1),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d387fb9),
	.w1(32'h3e6f1e6b),
	.w2(32'h3dc693d6),
	.w3(32'h382b1646),
	.w4(32'h3f4d2e41),
	.w5(32'h3eccf993),
	.w6(32'h3ee72bd0),
	.w7(32'h3f83853d),
	.w8(32'h3ee2b5de),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3ded47),
	.w1(32'h3ede1dc3),
	.w2(32'h3f8edb91),
	.w3(32'h3f8caa6f),
	.w4(32'h3eabf6c1),
	.w5(32'h3e44789d),
	.w6(32'h37dd9e56),
	.w7(32'h3d938143),
	.w8(32'h3e981b1d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1c94dc),
	.w1(32'h3ef8c58c),
	.w2(32'h3eab38ce),
	.w3(32'h3f286520),
	.w4(32'h3f36ff1c),
	.w5(32'h3d1b1938),
	.w6(32'h3f6d36e5),
	.w7(32'h3efc20aa),
	.w8(32'h3f07a1d0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4c1bab),
	.w1(32'h3d7e7ac1),
	.w2(32'h3f8201d4),
	.w3(32'h3efb6927),
	.w4(32'h3e2745aa),
	.w5(32'h37f0d698),
	.w6(32'h3f2a349b),
	.w7(32'h3eefe695),
	.w8(32'h3f692d50),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0a3dbf),
	.w1(32'h3ece079c),
	.w2(32'h3e8d2fa3),
	.w3(32'h3e1c0b3a),
	.w4(32'h3f237821),
	.w5(32'h3e118e2e),
	.w6(32'h3f310c02),
	.w7(32'h3f000f73),
	.w8(32'h3e433da1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e8f5333),
	.w1(32'h37280dca),
	.w2(32'h3edb9bfc),
	.w3(32'h36209509),
	.w4(32'h3c9867cc),
	.w5(32'h3ee01591),
	.w6(32'h3ef1c8ae),
	.w7(32'h3e888ba3),
	.w8(32'h3e14c50c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e6a3de1),
	.w1(32'h3f59539d),
	.w2(32'h3e864f4a),
	.w3(32'h3f4f5496),
	.w4(32'h3dbeb122),
	.w5(32'h3e2992a4),
	.w6(32'h3ec02d5d),
	.w7(32'h3772f36f),
	.w8(32'h36edf456),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e9084a0),
	.w1(32'h3e8446f6),
	.w2(32'h3f224d48),
	.w3(32'h3d38d6a0),
	.w4(32'h3f26343f),
	.w5(32'h3f30840e),
	.w6(32'h3e8b1fb4),
	.w7(32'h3f664d84),
	.w8(32'h3f1c4cc9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ea5e129),
	.w1(32'h3ecbee7a),
	.w2(32'h3ddc6a21),
	.w3(32'h3e937b23),
	.w4(32'h36caee6a),
	.w5(32'h3edde229),
	.w6(32'h3e888815),
	.w7(32'h370c5128),
	.w8(32'h3e987c75),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e603d60),
	.w1(32'h3ee5040d),
	.w2(32'h3f49f11c),
	.w3(32'h3e87a540),
	.w4(32'h3f18eaa1),
	.w5(32'h3e95cd62),
	.w6(32'h3f0b80ac),
	.w7(32'h3e6bd88e),
	.w8(32'h3e945390),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7bed48),
	.w1(32'h3dabe8a5),
	.w2(32'h3eacb6ae),
	.w3(32'h3d90b360),
	.w4(32'h3e768ec4),
	.w5(32'h3d509c77),
	.w6(32'h3f16f3a3),
	.w7(32'h3e88616d),
	.w8(32'h3f1bb839),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e841aa9),
	.w1(32'h3ecdc952),
	.w2(32'h3eaa44b8),
	.w3(32'h3ec4acdd),
	.w4(32'h3f24b81d),
	.w5(32'h3e846480),
	.w6(32'hb79f656f),
	.w7(32'h3eb29846),
	.w8(32'h3eb0de70),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f36f4cf),
	.w1(32'h3ec02092),
	.w2(32'h3e9e0a89),
	.w3(32'h3ec5196b),
	.w4(32'h3e94f196),
	.w5(32'h3f134b4b),
	.w6(32'h3ee81f44),
	.w7(32'h3e21ad5e),
	.w8(32'h3ef4df90),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ecc0fde),
	.w1(32'h3eb51434),
	.w2(32'h3f1040e7),
	.w3(32'h3eb5fd20),
	.w4(32'h3e879b5e),
	.w5(32'h3f4e9b78),
	.w6(32'h3f2277b4),
	.w7(32'h3f25d61d),
	.w8(32'h3ebf3c99),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ec59c7b),
	.w1(32'h3ed33981),
	.w2(32'h3e013501),
	.w3(32'h3e7ff044),
	.w4(32'h3db14b7e),
	.w5(32'h3ec05e43),
	.w6(32'h3edac8a3),
	.w7(32'h3ecea03d),
	.w8(32'h3ee51134),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ead4e22),
	.w1(32'h3e4cdca7),
	.w2(32'h3f5057be),
	.w3(32'h3ebae4b7),
	.w4(32'h3e1c4bab),
	.w5(32'h3fcdbbc6),
	.w6(32'h3e872c97),
	.w7(32'h3f25210c),
	.w8(32'h3f323608),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e943bb0),
	.w1(32'h3eb42276),
	.w2(32'h3dff9481),
	.w3(32'h3e2691b7),
	.w4(32'h3eeecce1),
	.w5(32'h3eca8d8e),
	.w6(32'h3f4ffbe2),
	.w7(32'h3f2acb54),
	.w8(32'hbc7479bf),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb10190),
	.w1(32'hbd21aa6b),
	.w2(32'h3981eed8),
	.w3(32'hbc6eac8b),
	.w4(32'hbb13da63),
	.w5(32'h392f725c),
	.w6(32'h3b3693dd),
	.w7(32'hbdd8246d),
	.w8(32'hba68f27a),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe5565c9),
	.w1(32'hbdb8cbda),
	.w2(32'h3cc444aa),
	.w3(32'h3d8e3c89),
	.w4(32'hbd9edd59),
	.w5(32'h3d43b73a),
	.w6(32'h3d3f6d2d),
	.w7(32'hbd7464cc),
	.w8(32'hbda161ec),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39056c23),
	.w1(32'h3c2d805e),
	.w2(32'hbdc1ae9b),
	.w3(32'hbd1de9bc),
	.w4(32'h3c748d58),
	.w5(32'h3df558d2),
	.w6(32'hbd47f72d),
	.w7(32'hbc2048ec),
	.w8(32'h3d458931),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d344772),
	.w1(32'hbbb406f8),
	.w2(32'hbd2302f3),
	.w3(32'hbe2164b2),
	.w4(32'h3ca71302),
	.w5(32'hbd81534e),
	.w6(32'hbded6596),
	.w7(32'hbd586b7e),
	.w8(32'hbd7cd1ef),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda8d0ca),
	.w1(32'h3b1c239f),
	.w2(32'hbd1d416d),
	.w3(32'h3ad55be8),
	.w4(32'hbd8ee94c),
	.w5(32'hbd04dfc3),
	.w6(32'hbd8c380b),
	.w7(32'hbb891e0c),
	.w8(32'hbe1b3dc0),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd145c16),
	.w1(32'hbd0c1d9f),
	.w2(32'hbd0d5ebb),
	.w3(32'hba9ea517),
	.w4(32'h3cff0cff),
	.w5(32'hbd55e1a2),
	.w6(32'hbdc2a453),
	.w7(32'hbda5d4ec),
	.w8(32'hbde0afcf),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb849a881),
	.w1(32'hbd78a0ee),
	.w2(32'hbc01e995),
	.w3(32'hbdd19315),
	.w4(32'hbcfbfced),
	.w5(32'hbd065a91),
	.w6(32'h3c84b8b0),
	.w7(32'hbdbef07b),
	.w8(32'hb7fa9b4f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd54162),
	.w1(32'h3cc5a542),
	.w2(32'h3d311472),
	.w3(32'h3d1f76a1),
	.w4(32'hbe6000db),
	.w5(32'h3d18053d),
	.w6(32'h3d955312),
	.w7(32'h3db28937),
	.w8(32'h3d910bd4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e4dc249),
	.w1(32'h3d5ee7bf),
	.w2(32'h3c321c54),
	.w3(32'hbd8a7597),
	.w4(32'h3cb549a0),
	.w5(32'hbd544a3a),
	.w6(32'hbd6cc4fd),
	.w7(32'h3c59fa2e),
	.w8(32'h3dae45c5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd910eec),
	.w1(32'h38580829),
	.w2(32'h3b380d96),
	.w3(32'hbc410049),
	.w4(32'hbc18a972),
	.w5(32'hbe2cccd1),
	.w6(32'h3c548531),
	.w7(32'hbd0f2210),
	.w8(32'hb8da06bb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e5cf1d7),
	.w1(32'h3c605d72),
	.w2(32'h3c8b1bb6),
	.w3(32'h3da2bde2),
	.w4(32'h3dcaac84),
	.w5(32'h3c331217),
	.w6(32'hbd890df4),
	.w7(32'h3aad83f6),
	.w8(32'hbe3613d2),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dd2a5e1),
	.w1(32'hbc2b1e82),
	.w2(32'hbce940bc),
	.w3(32'hbd1d3aa5),
	.w4(32'h3bea3606),
	.w5(32'hbdcc5464),
	.w6(32'hbbc7a985),
	.w7(32'h399d6ce0),
	.w8(32'h3c94c46e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd887af5),
	.w1(32'hbc7e95c3),
	.w2(32'h37e976a8),
	.w3(32'hbc7572ce),
	.w4(32'hbd86b117),
	.w5(32'hbd1db1e5),
	.w6(32'h3ca04a43),
	.w7(32'hbe331dbd),
	.w8(32'hbc85fd4a),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6105d),
	.w1(32'hbc99a136),
	.w2(32'h3d60c8f3),
	.w3(32'hbe24869b),
	.w4(32'h3d38f48d),
	.w5(32'h3d01f372),
	.w6(32'hbb7298db),
	.w7(32'hbd1de440),
	.w8(32'hbb51571c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe50654c),
	.w1(32'h3cfd8534),
	.w2(32'hbd94d207),
	.w3(32'h3d4c865f),
	.w4(32'h3d37152e),
	.w5(32'hbc25629b),
	.w6(32'hbcabdb18),
	.w7(32'h3d3ceb6e),
	.w8(32'h3a545ee1),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce29079),
	.w1(32'h3da0a59c),
	.w2(32'hbdfe204f),
	.w3(32'hbc458505),
	.w4(32'hbd4cc102),
	.w5(32'h3e0dffbe),
	.w6(32'hb7e183c0),
	.w7(32'hbc99ca2b),
	.w8(32'h3d3b348b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d116652),
	.w1(32'h3d5f62d0),
	.w2(32'hbc8a660e),
	.w3(32'h3cddaede),
	.w4(32'hbceb9e16),
	.w5(32'h37ce92d1),
	.w6(32'hbc9f78bd),
	.w7(32'h3833735b),
	.w8(32'hbc0e35d7),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42c7d2),
	.w1(32'h37931ba8),
	.w2(32'hbd82bc87),
	.w3(32'h3ca6a279),
	.w4(32'hbcb21839),
	.w5(32'hbe3caa00),
	.w6(32'h3db6e804),
	.w7(32'hbe00282f),
	.w8(32'h3b872533),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b0f84e),
	.w1(32'hb8883fcb),
	.w2(32'hbb6a31a9),
	.w3(32'hbcebf308),
	.w4(32'h3e34d7d5),
	.w5(32'hbda7fd6e),
	.w6(32'hbcd9f6e0),
	.w7(32'hbc799a33),
	.w8(32'h3d3b38b5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc6e791),
	.w1(32'h3ca54a1c),
	.w2(32'h3d50806f),
	.w3(32'hbc4c2198),
	.w4(32'hbc229958),
	.w5(32'h3bba9cad),
	.w6(32'hbdaae75d),
	.w7(32'h3d261171),
	.w8(32'hb580501e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930a953),
	.w1(32'hbd6ed9f5),
	.w2(32'hbd2a081b),
	.w3(32'h37592edb),
	.w4(32'hbc4abc72),
	.w5(32'h3d97d946),
	.w6(32'hbe02c6c8),
	.w7(32'hbc11dace),
	.w8(32'h3cdb4fb0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad5d4),
	.w1(32'h3cd88dde),
	.w2(32'hbdb9674a),
	.w3(32'hbd5a0e7f),
	.w4(32'h3d91dd05),
	.w5(32'hb98fc189),
	.w6(32'h3d2415c7),
	.w7(32'h3c1ea2db),
	.w8(32'h3ded9959),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2bac2c),
	.w1(32'hbe238eb9),
	.w2(32'h379eab07),
	.w3(32'h3d732fcd),
	.w4(32'hbeb2d9f6),
	.w5(32'hbcdddfdc),
	.w6(32'hbc8bef9a),
	.w7(32'hbd8b6460),
	.w8(32'h3d9ead3e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd31caa4),
	.w1(32'h3bdac612),
	.w2(32'h3df2955d),
	.w3(32'hbc3e926e),
	.w4(32'h3de01364),
	.w5(32'hbe09b27b),
	.w6(32'h3cc77354),
	.w7(32'hbd7ceb0d),
	.w8(32'hbd2b2aea),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0e9eb5),
	.w1(32'hbda5e248),
	.w2(32'hbd135447),
	.w3(32'h3db83796),
	.w4(32'hbd9de386),
	.w5(32'h3d997b3f),
	.w6(32'h3dad07e7),
	.w7(32'hbbcdbb67),
	.w8(32'h3d15b755),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc283768),
	.w1(32'hbd9390a5),
	.w2(32'h3abcb20a),
	.w3(32'h3cc9b778),
	.w4(32'hbb9ce5eb),
	.w5(32'hbe032baa),
	.w6(32'hbccff6c3),
	.w7(32'hbd0b9199),
	.w8(32'hbd3585b4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c24e),
	.w1(32'hbdaa3520),
	.w2(32'hbde13dda),
	.w3(32'hbcdb234c),
	.w4(32'hbb4b928b),
	.w5(32'hbc90ff86),
	.w6(32'hbcfb3a8f),
	.w7(32'hbd16cb87),
	.w8(32'hbcb6e62f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3df20732),
	.w1(32'hbda22b0f),
	.w2(32'h3e39bbd2),
	.w3(32'hbe157a20),
	.w4(32'hbd7f31bf),
	.w5(32'h3dc27319),
	.w6(32'hbdb7bd0e),
	.w7(32'hbc79e902),
	.w8(32'hbe3a7842),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd87543c),
	.w1(32'h3bedf00e),
	.w2(32'h3b2327e5),
	.w3(32'hbcd3c3ab),
	.w4(32'h3c37e691),
	.w5(32'h3cea01e5),
	.w6(32'h3d11362d),
	.w7(32'h3c015f1f),
	.w8(32'h3c40a4a1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d9f6487),
	.w1(32'h3702eda7),
	.w2(32'h3d296e74),
	.w3(32'h344e9221),
	.w4(32'h3d600a7b),
	.w5(32'h3d8d6611),
	.w6(32'h3539b9c9),
	.w7(32'h3c0252a1),
	.w8(32'h3d9d8753),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92cabd),
	.w1(32'h3d645497),
	.w2(32'h3b991966),
	.w3(32'h3cd2582f),
	.w4(32'h34341789),
	.w5(32'h3b44371f),
	.w6(32'h3bad5a63),
	.w7(32'h3aa22845),
	.w8(32'h3c1038eb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03792e),
	.w1(32'h3bc44ec1),
	.w2(32'h3d833dfd),
	.w3(32'h3d909648),
	.w4(32'h3bc5bd01),
	.w5(32'h3d32b8ff),
	.w6(32'h3ddb3901),
	.w7(32'h3dcc36f9),
	.w8(32'h3c0aa64f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3feffb),
	.w1(32'h3c9addc2),
	.w2(32'h3b6adc52),
	.w3(32'h3b1e98e7),
	.w4(32'h3c3b1e22),
	.w5(32'h3df7b61c),
	.w6(32'h3dd1cd47),
	.w7(32'h3da7a5e6),
	.w8(32'h3bed7853),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2ea1),
	.w1(32'h3e12c884),
	.w2(32'h3d0806cc),
	.w3(32'h3e189fee),
	.w4(32'h3d80eb34),
	.w5(32'h3bd6bfec),
	.w6(32'h3c7d89f6),
	.w7(32'h3a297829),
	.w8(32'h3c9ac8e5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e029fcb),
	.w1(32'h3ce85216),
	.w2(32'h3c94ea6e),
	.w3(32'h3c241be2),
	.w4(32'hb611d790),
	.w5(32'h3c02a324),
	.w6(32'h3ccc0ce6),
	.w7(32'h3de87264),
	.w8(32'h3bb4442e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5b14ec),
	.w1(32'hb52585a9),
	.w2(32'h3c8dd3be),
	.w3(32'h3b3d4755),
	.w4(32'h3d88f8ef),
	.w5(32'h3c96c88f),
	.w6(32'h3c8a2771),
	.w7(32'h3c8d039f),
	.w8(32'h3e88f52f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc31d14),
	.w1(32'h3cae8a6c),
	.w2(32'h3b7b9782),
	.w3(32'h3d99a14c),
	.w4(32'h3ccddf0a),
	.w5(32'h3cc9884e),
	.w6(32'h3cf8a851),
	.w7(32'h3d72dc32),
	.w8(32'h3abeef36),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacc719),
	.w1(32'h3d9109b1),
	.w2(32'h3ccc2867),
	.w3(32'h3b8417a5),
	.w4(32'h3d7e7d24),
	.w5(32'h34f8fab8),
	.w6(32'h3c812a3b),
	.w7(32'h3d914827),
	.w8(32'h3ad3947a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4b05a5),
	.w1(32'h34cbbb42),
	.w2(32'h3d21a8f2),
	.w3(32'h3ae3c562),
	.w4(32'h3d79dde8),
	.w5(32'h3adc8cc1),
	.w6(32'h3ddd5c06),
	.w7(32'h3d8b1703),
	.w8(32'h3c99a7ac),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc92929),
	.w1(32'h3d0fcc3d),
	.w2(32'h3b016745),
	.w3(32'h3c5bda8e),
	.w4(32'h3c9ae7c1),
	.w5(32'h3e656166),
	.w6(32'h3cba40da),
	.w7(32'h3c106c9d),
	.w8(32'h3a17ba62),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362f1b74),
	.w1(32'h3d6d36c2),
	.w2(32'h3cd315c4),
	.w3(32'h3cd3af8f),
	.w4(32'h3d9a385f),
	.w5(32'h3cf0d9a0),
	.w6(32'h3c9dbba1),
	.w7(32'h3b9628f2),
	.w8(32'h3d345dc6),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e7dc887),
	.w1(32'h3c62e9d2),
	.w2(32'h3c27da2f),
	.w3(32'h33717c84),
	.w4(32'h3b817000),
	.w5(32'h3c21db10),
	.w6(32'h3cb085a6),
	.w7(32'h3d97f73d),
	.w8(32'h3b9ebdb2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d87667a),
	.w1(32'h3d0e22c9),
	.w2(32'h3a6fa0a2),
	.w3(32'h3e2021ca),
	.w4(32'h3d21a694),
	.w5(32'h3d251296),
	.w6(32'h3cf4a4dd),
	.w7(32'h3caf66db),
	.w8(32'h3db16ff9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc21105),
	.w1(32'h3b77c5c5),
	.w2(32'h3599a6a1),
	.w3(32'h3d4ace81),
	.w4(32'h3cf66a1b),
	.w5(32'h3d6aaca0),
	.w6(32'h3acc7e8d),
	.w7(32'h3db3f045),
	.w8(32'h3cdb0583),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90739d),
	.w1(32'h3de16693),
	.w2(32'h3b5eddf4),
	.w3(32'h3d66800a),
	.w4(32'h3cdecd8b),
	.w5(32'h3c93abfc),
	.w6(32'h3d2a6c46),
	.w7(32'h3c1d3822),
	.w8(32'h3c827ac3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4ba4f86),
	.w1(32'h39e07f0c),
	.w2(32'h3cc08805),
	.w3(32'h3d20e335),
	.w4(32'h3d0d8fe4),
	.w5(32'h3c96ef00),
	.w6(32'h362a240e),
	.w7(32'h3ca9e643),
	.w8(32'h3c26edba),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dab1d26),
	.w1(32'h3b2dcb44),
	.w2(32'h3b8820e1),
	.w3(32'h3c9a3943),
	.w4(32'h33845a71),
	.w5(32'hb4725aff),
	.w6(32'h3d56f265),
	.w7(32'h3be82b9a),
	.w8(32'h3cd95b84),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad16351),
	.w1(32'h3d18c330),
	.w2(32'h3d7048da),
	.w3(32'h3d8f496e),
	.w4(32'h3d858b8e),
	.w5(32'h3d7ad866),
	.w6(32'h3bff7beb),
	.w7(32'h3dd2d0e8),
	.w8(32'h3d0da131),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35c6cf),
	.w1(32'h36c3604d),
	.w2(32'h3cdb80dd),
	.w3(32'h3c5658ea),
	.w4(32'h36d22ee7),
	.w5(32'h3c82fc5a),
	.w6(32'h3c6f0a8c),
	.w7(32'h3b91faf5),
	.w8(32'h3bb835a6),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45300d),
	.w1(32'h3cd98101),
	.w2(32'h3d2bb5eb),
	.w3(32'h3d1aebbd),
	.w4(32'h3bc46658),
	.w5(32'h3c5d42a9),
	.w6(32'h3cbc4427),
	.w7(32'h3d71a759),
	.w8(32'h3cf0e790),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af54565),
	.w1(32'h3cefb04b),
	.w2(32'h3ad37739),
	.w3(32'h3d1198dc),
	.w4(32'h3ca9ae88),
	.w5(32'h3d1d180d),
	.w6(32'h3b0ad96e),
	.w7(32'h3cb3c756),
	.w8(32'h3dd4b419),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e3fd3),
	.w1(32'h3d5fefe0),
	.w2(32'h3d25307d),
	.w3(32'h34b0da13),
	.w4(32'h3c4335fe),
	.w5(32'h3c3e36c2),
	.w6(32'h3cf92673),
	.w7(32'h3bd6106b),
	.w8(32'h3d54af64),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb58e29),
	.w1(32'h3cb94b4c),
	.w2(32'h3cc539fe),
	.w3(32'h3d379f30),
	.w4(32'h3b986b6b),
	.w5(32'h3d04a3cd),
	.w6(32'h3c372e1b),
	.w7(32'h3cf2d5ad),
	.w8(32'h3c9333e5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca17bcc),
	.w1(32'h3d115fe8),
	.w2(32'h3d85a681),
	.w3(32'h3cd5dd1d),
	.w4(32'h3dbb0d55),
	.w5(32'h3c509ad1),
	.w6(32'h3cb6eb7c),
	.w7(32'h3d0d2eb3),
	.w8(32'h3cc3d594),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cdab3),
	.w1(32'h3ae393d0),
	.w2(32'h3caf5616),
	.w3(32'h3d201961),
	.w4(32'h3c9eb49a),
	.w5(32'h3cb08349),
	.w6(32'h3cccdbd8),
	.w7(32'h3b074ae8),
	.w8(32'h3c0cc723),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e59e8),
	.w1(32'h3b74d7fe),
	.w2(32'h3e0e42aa),
	.w3(32'h3ca49e2c),
	.w4(32'h3e018686),
	.w5(32'h3de1ca24),
	.w6(32'h3b721699),
	.w7(32'h3e484f0d),
	.w8(32'h3c255e59),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd793f),
	.w1(32'h3d7d082b),
	.w2(32'h3ce192a2),
	.w3(32'h3e3cbb05),
	.w4(32'h3d604600),
	.w5(32'hba2c4395),
	.w6(32'h3cc99292),
	.w7(32'h3babd66d),
	.w8(32'hba02c3e5),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b95a),
	.w1(32'hbae22bc5),
	.w2(32'hba51aedd),
	.w3(32'hbabfaef3),
	.w4(32'hb9e25c5a),
	.w5(32'hbaed7d18),
	.w6(32'hbac8cbb6),
	.w7(32'hb920daf6),
	.w8(32'hbaff4788),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e668b),
	.w1(32'hbabdfd90),
	.w2(32'hbae6799d),
	.w3(32'hba8d20ab),
	.w4(32'hba832982),
	.w5(32'hba4d3842),
	.w6(32'h3a41c3d7),
	.w7(32'hba544551),
	.w8(32'hbb4a15a3),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15fd4b),
	.w1(32'hbad8fad6),
	.w2(32'hbab469bd),
	.w3(32'hba221b41),
	.w4(32'h3988caf1),
	.w5(32'hbadf5e80),
	.w6(32'hbb0bfd49),
	.w7(32'hbafad829),
	.w8(32'hb7940a85),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bef4f),
	.w1(32'h3b1933a0),
	.w2(32'h3a99df0f),
	.w3(32'hbb0658d9),
	.w4(32'hba00f8ed),
	.w5(32'h3ab31e45),
	.w6(32'h3b5754c5),
	.w7(32'h3ae1b8a7),
	.w8(32'hb87b0aca),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba864d1e),
	.w1(32'hba3adf42),
	.w2(32'hb940d7a6),
	.w3(32'hb8d5015d),
	.w4(32'h3988ec41),
	.w5(32'hb86d8f0b),
	.w6(32'hb97eb399),
	.w7(32'h39fee688),
	.w8(32'h3b539b25),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d9a5c),
	.w1(32'h3b19bd17),
	.w2(32'h3acf3e99),
	.w3(32'h3a7d07ea),
	.w4(32'h3a005ad6),
	.w5(32'hba7fab8f),
	.w6(32'h3ab6408b),
	.w7(32'h3aeeec22),
	.w8(32'h37281dab),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0919bb),
	.w1(32'h3a2c9475),
	.w2(32'h3ae59d4d),
	.w3(32'hbacee734),
	.w4(32'hbaf6c3fe),
	.w5(32'hbaaedf25),
	.w6(32'h36d049eb),
	.w7(32'h37253d56),
	.w8(32'hb9b951e0),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8fcb),
	.w1(32'hba9ed3c5),
	.w2(32'hba89bfaf),
	.w3(32'hbaa6f525),
	.w4(32'hbab657e6),
	.w5(32'hbaf64cfd),
	.w6(32'hb983862c),
	.w7(32'hba74d4ea),
	.w8(32'hbb145957),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb459bac),
	.w1(32'h39f30c38),
	.w2(32'h3a94c61f),
	.w3(32'hb95f40e6),
	.w4(32'hb9d10e1d),
	.w5(32'hbabb7291),
	.w6(32'h3a43dcd8),
	.w7(32'h3a296a96),
	.w8(32'hbab8be2e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9adf2),
	.w1(32'h39036dbf),
	.w2(32'hb984b90c),
	.w3(32'hba414bb0),
	.w4(32'hba4ddf9b),
	.w5(32'h39e426d4),
	.w6(32'h3ad4dfb9),
	.w7(32'h3941dd9d),
	.w8(32'h3a123f78),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ab7bc),
	.w1(32'hbaada73d),
	.w2(32'hba9cd850),
	.w3(32'hbab30a56),
	.w4(32'hb8d82fb1),
	.w5(32'hbb1d626d),
	.w6(32'hbacfd6e2),
	.w7(32'hb9f87440),
	.w8(32'hbb2bbe80),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa78812),
	.w1(32'hb83061a2),
	.w2(32'h3a1f6945),
	.w3(32'hbad0b5ec),
	.w4(32'hbaa47e2e),
	.w5(32'h3a68206f),
	.w6(32'hbaa730fe),
	.w7(32'hb9a5f221),
	.w8(32'h3a1e682b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39579f27),
	.w1(32'h388e646d),
	.w2(32'h39137b06),
	.w3(32'hb51d77f0),
	.w4(32'h3a373557),
	.w5(32'hbae1ded9),
	.w6(32'h3a6fdc88),
	.w7(32'hb9eb9b35),
	.w8(32'hbb186266),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0446a7),
	.w1(32'hb89bc061),
	.w2(32'hba33af56),
	.w3(32'hba0f1d13),
	.w4(32'hba1e6fc8),
	.w5(32'hb99c4986),
	.w6(32'hba1e5a87),
	.w7(32'h38bcc5fb),
	.w8(32'hba9ad180),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a490fc2),
	.w1(32'h386b26d1),
	.w2(32'h39b8525e),
	.w3(32'hb71eb542),
	.w4(32'h3a1a50cb),
	.w5(32'h3a9cc067),
	.w6(32'hba6c8e63),
	.w7(32'hba4738a0),
	.w8(32'h3a978305),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b33ae),
	.w1(32'h3acad6dc),
	.w2(32'h3a7f432b),
	.w3(32'h3af6f585),
	.w4(32'h3ae2d3ba),
	.w5(32'h39a532c2),
	.w6(32'h3a2c3e9e),
	.w7(32'h3a63511a),
	.w8(32'h3addfc66),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e967d1),
	.w1(32'h392089b7),
	.w2(32'hbad88b70),
	.w3(32'h398c2193),
	.w4(32'h37e0afec),
	.w5(32'hbb2ac1ba),
	.w6(32'h3a95b33b),
	.w7(32'hb87b2012),
	.w8(32'hbb297a9c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a537f),
	.w1(32'hb9eb6fbf),
	.w2(32'h3a03c807),
	.w3(32'hbb28ebed),
	.w4(32'hba80cc10),
	.w5(32'h3872d043),
	.w6(32'hb8e6d3be),
	.w7(32'h39e8aaaf),
	.w8(32'h39d464b8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928074a),
	.w1(32'hba17b37a),
	.w2(32'hb9fa087b),
	.w3(32'hba0a6f03),
	.w4(32'hb8e69723),
	.w5(32'hba657723),
	.w6(32'hb94a76fb),
	.w7(32'h3a7608d7),
	.w8(32'h39d30cee),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a461cb9),
	.w1(32'hba173545),
	.w2(32'h3a326df1),
	.w3(32'hbac8a9da),
	.w4(32'hb9a967e2),
	.w5(32'hba43bcc0),
	.w6(32'h3ae69bc0),
	.w7(32'h3a9dd46a),
	.w8(32'hba7db5b4),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ea342),
	.w1(32'h38548ac9),
	.w2(32'h3915eda2),
	.w3(32'hba1c7559),
	.w4(32'hbac3ebba),
	.w5(32'hba9196ce),
	.w6(32'hb9cbaa74),
	.w7(32'hba624cb1),
	.w8(32'hbaba42d1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafca473),
	.w1(32'hbb2fe241),
	.w2(32'hba50babb),
	.w3(32'hbb50df97),
	.w4(32'hbadc0987),
	.w5(32'hb95b051d),
	.w6(32'hbb9ba84d),
	.w7(32'hbac72f29),
	.w8(32'h3a2773ac),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4833e6),
	.w1(32'h3b156529),
	.w2(32'h3af6326c),
	.w3(32'h39a8ab4c),
	.w4(32'hb90731a3),
	.w5(32'hb9169f7a),
	.w6(32'h3a4cd09b),
	.w7(32'h3adb4c09),
	.w8(32'hba48568e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899ecc9),
	.w1(32'hba054022),
	.w2(32'hba844f47),
	.w3(32'hb94ee323),
	.w4(32'hbaa924a2),
	.w5(32'h3a3b470a),
	.w6(32'hb9777453),
	.w7(32'hb9fb7959),
	.w8(32'hbb02feb2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f7505),
	.w1(32'h3af06f24),
	.w2(32'h39bd479c),
	.w3(32'h3b4618e2),
	.w4(32'h3afd2f1e),
	.w5(32'h3a575f05),
	.w6(32'h3968d69c),
	.w7(32'hba02b06f),
	.w8(32'hb96dc332),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a656e63),
	.w1(32'h3a92e5cd),
	.w2(32'hb96f0575),
	.w3(32'h3a0ebd6f),
	.w4(32'hba9c9d6c),
	.w5(32'h39908b4f),
	.w6(32'h3ad2b9c0),
	.w7(32'hba9f8ef1),
	.w8(32'hb9f7faa2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac98ba9),
	.w1(32'h3b625389),
	.w2(32'h3b235e5b),
	.w3(32'h3af318a7),
	.w4(32'h3a9bac69),
	.w5(32'h386eb547),
	.w6(32'h3b45ba6f),
	.w7(32'h3adb5647),
	.w8(32'hb998e486),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e1bbb0),
	.w1(32'h39be6d3a),
	.w2(32'h3a77c7a4),
	.w3(32'h3af923cf),
	.w4(32'h3b6f0d1e),
	.w5(32'hbb1f8818),
	.w6(32'h3b1ec01a),
	.w7(32'h3af7d3dc),
	.w8(32'hbb04ad67),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e987),
	.w1(32'hba3cbf4f),
	.w2(32'hba9342b6),
	.w3(32'hbab58348),
	.w4(32'hbb050ec4),
	.w5(32'hba071129),
	.w6(32'h3a96a767),
	.w7(32'hba6b7cb7),
	.w8(32'hb9cee2e7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d373a),
	.w1(32'hba5e3343),
	.w2(32'hba6c485c),
	.w3(32'h3a1859f6),
	.w4(32'hba1cf8c3),
	.w5(32'hbb115a24),
	.w6(32'hb9731237),
	.w7(32'hbab8296f),
	.w8(32'hbafd8476),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule