module layer_10_featuremap_179(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae985d),
	.w1(32'hbc52baca),
	.w2(32'h3ab91a52),
	.w3(32'hbb15d078),
	.w4(32'hbbefecf0),
	.w5(32'h3bd3b4e3),
	.w6(32'hbb01cac8),
	.w7(32'h3b2e8781),
	.w8(32'h3b2004e3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977a9bf),
	.w1(32'hbc2f88be),
	.w2(32'h3b2bff83),
	.w3(32'hbb93b8dc),
	.w4(32'h3a26789f),
	.w5(32'hbb713256),
	.w6(32'h3b19f0d4),
	.w7(32'hbb1d21fc),
	.w8(32'hbc4c9816),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3912ad),
	.w1(32'hbbc6a1e5),
	.w2(32'h3be7d1a5),
	.w3(32'hbc7c263a),
	.w4(32'hbb14bc09),
	.w5(32'hbb275de7),
	.w6(32'h3abfd817),
	.w7(32'h3b6b4e0a),
	.w8(32'hbaede1b8),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0fbc1),
	.w1(32'h3c68e98f),
	.w2(32'h3a2af376),
	.w3(32'hbbc575a7),
	.w4(32'h3bdf29d3),
	.w5(32'hbbc337f6),
	.w6(32'hbb7763b7),
	.w7(32'hbc4c388c),
	.w8(32'hbb3d26b4),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44dcda),
	.w1(32'h3bef371c),
	.w2(32'hbb71b6e5),
	.w3(32'h3a3acd60),
	.w4(32'h38711a38),
	.w5(32'hbbe0ec02),
	.w6(32'hb956b351),
	.w7(32'h396af460),
	.w8(32'h3bf942d3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c156bc3),
	.w1(32'h3d2d4077),
	.w2(32'h3b67e9fe),
	.w3(32'h3b4ec08a),
	.w4(32'h3c5ff62c),
	.w5(32'h3be34276),
	.w6(32'h3c4b7f63),
	.w7(32'h3ba70894),
	.w8(32'hbc73bd94),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f0367),
	.w1(32'hbc8af1ec),
	.w2(32'hbbbf9dca),
	.w3(32'hbc2ed55c),
	.w4(32'hbb523d27),
	.w5(32'hbc5780a1),
	.w6(32'hbb152ddd),
	.w7(32'hbc31dcae),
	.w8(32'hbc95fadb),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9245b5),
	.w1(32'h3d018b44),
	.w2(32'hbc3d8a8e),
	.w3(32'hbcd18e87),
	.w4(32'h3ac60bad),
	.w5(32'h3b19fb00),
	.w6(32'h3b6620ee),
	.w7(32'hbaf4dd7f),
	.w8(32'hbbf71b41),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca928fb),
	.w1(32'h3c61d1f5),
	.w2(32'hbcbb9f53),
	.w3(32'hba246b6d),
	.w4(32'hbb1fa077),
	.w5(32'hbc02ec46),
	.w6(32'hbb3be413),
	.w7(32'hbb8bf255),
	.w8(32'hbb8283a3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fef49),
	.w1(32'hbd24bb6f),
	.w2(32'h3c4784d4),
	.w3(32'hb9aa4aa2),
	.w4(32'hbb3fc8fc),
	.w5(32'hbba6b796),
	.w6(32'hbc2c8648),
	.w7(32'hbbe88b4c),
	.w8(32'h3bef8fcb),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01ad26),
	.w1(32'h3c877d41),
	.w2(32'h3c4c135c),
	.w3(32'h380d241d),
	.w4(32'h3b98d9fe),
	.w5(32'h3bd0f8aa),
	.w6(32'hbb0c6fa9),
	.w7(32'hbb5bec02),
	.w8(32'hbbfe633b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb5614),
	.w1(32'h3b99c5ca),
	.w2(32'hbc97ae6c),
	.w3(32'hbb95ffff),
	.w4(32'hbb2048b4),
	.w5(32'hbb0a2b44),
	.w6(32'h3bc9ff9e),
	.w7(32'hbb35c8de),
	.w8(32'hbbd05eec),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba01152),
	.w1(32'h3bee822a),
	.w2(32'h3bdddb5e),
	.w3(32'h3a21469e),
	.w4(32'h3992188b),
	.w5(32'h3bbdd5de),
	.w6(32'hbb938ca8),
	.w7(32'hba8853de),
	.w8(32'hbb8d90e5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f49f),
	.w1(32'h3cd0ecc8),
	.w2(32'hbc848a2a),
	.w3(32'hbb02b5c3),
	.w4(32'hbbc16689),
	.w5(32'hba89cb98),
	.w6(32'hbb167615),
	.w7(32'hbb277cf2),
	.w8(32'h3b58ee52),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eeba9),
	.w1(32'hbb459a5c),
	.w2(32'h3b73210f),
	.w3(32'h3c2d82ae),
	.w4(32'hbc02d768),
	.w5(32'hba9a2eb4),
	.w6(32'hb8826af6),
	.w7(32'h3b613c78),
	.w8(32'hbadd05a4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c06b7),
	.w1(32'h3cae9928),
	.w2(32'hbc47a8b1),
	.w3(32'hbbe7f7fd),
	.w4(32'hba3ad3fa),
	.w5(32'hbace92ef),
	.w6(32'h3b775adf),
	.w7(32'h3aa52cb2),
	.w8(32'hbb5de38b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c38ca),
	.w1(32'h3bd71261),
	.w2(32'h3bad27df),
	.w3(32'hb98eeffa),
	.w4(32'hba9c1045),
	.w5(32'h3b61ae38),
	.w6(32'h3c2fa5f0),
	.w7(32'h3c0bbca7),
	.w8(32'hbb2a6a62),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d0e26),
	.w1(32'hbd16b8ad),
	.w2(32'h39a681a8),
	.w3(32'hbbd8ee76),
	.w4(32'hbc65c47d),
	.w5(32'hbc31cad5),
	.w6(32'hbc8b8be3),
	.w7(32'hbc301a93),
	.w8(32'hbb48b5ba),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18bceb),
	.w1(32'hbbd301de),
	.w2(32'hbb9c4796),
	.w3(32'hbc2afb7e),
	.w4(32'hba6d8712),
	.w5(32'hbbe0e23c),
	.w6(32'hba8a3ef4),
	.w7(32'hbc0c657d),
	.w8(32'hbc53804c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc372ce3),
	.w1(32'h3c6fd12f),
	.w2(32'hbcacad01),
	.w3(32'hbc48cb1e),
	.w4(32'h3b02f7ba),
	.w5(32'hbbfed1b1),
	.w6(32'h3b438b13),
	.w7(32'hbba189a1),
	.w8(32'hbbcb240a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e93ab),
	.w1(32'h3cd6b5b3),
	.w2(32'hbc9994b3),
	.w3(32'hbb75a23d),
	.w4(32'h3a44409b),
	.w5(32'hbb0226a7),
	.w6(32'h3ad93e40),
	.w7(32'hbb495023),
	.w8(32'hbb4b092d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc734136),
	.w1(32'hbb613e97),
	.w2(32'h3b878df4),
	.w3(32'h3bbe81cd),
	.w4(32'hbbbe59b6),
	.w5(32'hbb9a298a),
	.w6(32'h3987d34a),
	.w7(32'hbbdcd539),
	.w8(32'hbad8fc2f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5b89),
	.w1(32'hbc375987),
	.w2(32'hbc4395ff),
	.w3(32'hbca3a038),
	.w4(32'hbc7a3cf9),
	.w5(32'hbc1aeb69),
	.w6(32'hbc909b8b),
	.w7(32'hbb888f38),
	.w8(32'h3957c638),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b807032),
	.w1(32'h3d15b730),
	.w2(32'hbbfa3ac0),
	.w3(32'h3b5db892),
	.w4(32'h3bf7899e),
	.w5(32'h3bb7187d),
	.w6(32'h3c25b688),
	.w7(32'h3ad806c9),
	.w8(32'hbbecca63),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaf642f),
	.w1(32'hba114306),
	.w2(32'h3b520eb5),
	.w3(32'h3b4494d5),
	.w4(32'hbaa60e57),
	.w5(32'h3ae79e03),
	.w6(32'hbbb5f8f7),
	.w7(32'hba0fa7dd),
	.w8(32'hbb21ea16),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c6760),
	.w1(32'h3c6f4737),
	.w2(32'h3b6bd2a3),
	.w3(32'hba9273b9),
	.w4(32'h3bab08d0),
	.w5(32'h3b83cb9f),
	.w6(32'h3bd371f2),
	.w7(32'hbb914531),
	.w8(32'hbbaff853),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b967c22),
	.w1(32'h3c4f9cf6),
	.w2(32'hbc52f852),
	.w3(32'hbb8ab52b),
	.w4(32'hbb37afee),
	.w5(32'hbb243954),
	.w6(32'h3ae9e8e5),
	.w7(32'hbb872d8c),
	.w8(32'hbbb4e1fd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80d0b4),
	.w1(32'hbc3c8f6c),
	.w2(32'h3bebcdf2),
	.w3(32'h3a94951e),
	.w4(32'hbb3ba0f9),
	.w5(32'h3ae8780d),
	.w6(32'hbc336d50),
	.w7(32'hbbcc3ac6),
	.w8(32'hbb0148ba),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f66ba),
	.w1(32'hbcc707d6),
	.w2(32'hbb633eea),
	.w3(32'hb95f31b5),
	.w4(32'hbd0a729c),
	.w5(32'hbb71e116),
	.w6(32'hbce3cc74),
	.w7(32'hbb213e45),
	.w8(32'h3b640948),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a0eba),
	.w1(32'hba1ab5f4),
	.w2(32'h3aaea70a),
	.w3(32'h3b5e545b),
	.w4(32'h3af22454),
	.w5(32'h3b80af00),
	.w6(32'h3b64a8c7),
	.w7(32'h3ad492c7),
	.w8(32'h398f6fb7),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac169b5),
	.w1(32'h3c7ec063),
	.w2(32'hbbc08b76),
	.w3(32'h3b122d41),
	.w4(32'h3a1186c1),
	.w5(32'h3a891d26),
	.w6(32'h3ac16899),
	.w7(32'hbac3af71),
	.w8(32'hbbb0dd9e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68b5a2),
	.w1(32'h3c951fa9),
	.w2(32'h39a9ac25),
	.w3(32'hba73a2cd),
	.w4(32'h3b3f4052),
	.w5(32'h3bd42cff),
	.w6(32'h3abf40a7),
	.w7(32'h39ea7bb8),
	.w8(32'hbc163e56),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc848ed4),
	.w1(32'hbb18c317),
	.w2(32'hbc2fccf1),
	.w3(32'h3ab8ff78),
	.w4(32'h3a867c8a),
	.w5(32'hbb8a6736),
	.w6(32'h3b4ed067),
	.w7(32'h3966e270),
	.w8(32'hbba892f6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce030e),
	.w1(32'hbbf0cd3b),
	.w2(32'h3ac1754e),
	.w3(32'h3915bea6),
	.w4(32'hba54f157),
	.w5(32'hbc12ef00),
	.w6(32'h3a6ab885),
	.w7(32'h3987430e),
	.w8(32'h3b2bcc9b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab3d31),
	.w1(32'hbcf8eb1b),
	.w2(32'hbb0546bc),
	.w3(32'hbb1ac4a4),
	.w4(32'hbc1f8562),
	.w5(32'hbc13e6c1),
	.w6(32'hbc3888e3),
	.w7(32'hbbcf3be0),
	.w8(32'h3bf9001b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57ae9e),
	.w1(32'h3c84d06a),
	.w2(32'hbb9ce04b),
	.w3(32'hbaaec2c1),
	.w4(32'hbb2da1c2),
	.w5(32'h3b6a5f7a),
	.w6(32'h3b52e927),
	.w7(32'hbb864af5),
	.w8(32'hbc52f0b7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5461b6),
	.w1(32'hbc9f7c57),
	.w2(32'hbc1f9b28),
	.w3(32'h3a9054a7),
	.w4(32'hbb90f555),
	.w5(32'hbc8563ca),
	.w6(32'hbbff6389),
	.w7(32'hbc4b7a19),
	.w8(32'hbc6e2002),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00b47f),
	.w1(32'hbbbcd110),
	.w2(32'h3bc3e0c5),
	.w3(32'hbc11cfca),
	.w4(32'h3c2b5d82),
	.w5(32'h39b546de),
	.w6(32'h3c04f8af),
	.w7(32'h3b9ab8a3),
	.w8(32'hbbf6c459),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b17f5c),
	.w1(32'h3d254f48),
	.w2(32'hba768f9b),
	.w3(32'hbb798d05),
	.w4(32'h3c547aed),
	.w5(32'h3c00905b),
	.w6(32'h3c98d283),
	.w7(32'h3c12392e),
	.w8(32'hbbbd45c2),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab2369),
	.w1(32'hbbae5ccb),
	.w2(32'hbb2b0728),
	.w3(32'hb6d13dd7),
	.w4(32'h3b88b96a),
	.w5(32'hbbe79d25),
	.w6(32'h3b3da6b7),
	.w7(32'hbbab3979),
	.w8(32'hbc2c466a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26735a),
	.w1(32'hbba8298c),
	.w2(32'hba818c76),
	.w3(32'hbc55b59b),
	.w4(32'hbb7a8992),
	.w5(32'h3a887476),
	.w6(32'h3b087b17),
	.w7(32'h3b38a07f),
	.w8(32'h3b24e734),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc178),
	.w1(32'h3aa973a1),
	.w2(32'h3af76761),
	.w3(32'h3ab63ab9),
	.w4(32'h3b8de9b8),
	.w5(32'hbada8d7c),
	.w6(32'h3a129083),
	.w7(32'hb9002f72),
	.w8(32'hbbd8d9d6),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892e98),
	.w1(32'h3c532496),
	.w2(32'hbb851c54),
	.w3(32'hbbfcbdbb),
	.w4(32'h3b5fb3ed),
	.w5(32'hbb102dd2),
	.w6(32'hb92cb7d2),
	.w7(32'hbaf8d4b8),
	.w8(32'hbc2261cd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d18c5),
	.w1(32'hbd644dcc),
	.w2(32'h3c6fee15),
	.w3(32'hbaa05395),
	.w4(32'hbc0e5217),
	.w5(32'hbc215a37),
	.w6(32'hbc5e3c50),
	.w7(32'hbc17653d),
	.w8(32'h3cac0742),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d43b243),
	.w1(32'hbcdd051b),
	.w2(32'h3c1d45fd),
	.w3(32'h3bae06e3),
	.w4(32'hbc0c3a3a),
	.w5(32'h3ac9d9ab),
	.w6(32'hbc13d1c2),
	.w7(32'h3bf15e15),
	.w8(32'h3c51764d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d082e3c),
	.w1(32'hbc9e238c),
	.w2(32'h3be55656),
	.w3(32'h3c0caf0f),
	.w4(32'hbc04bdd3),
	.w5(32'hbb683698),
	.w6(32'hbb1bd1e3),
	.w7(32'hbb409ea8),
	.w8(32'h3b53438e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1643e),
	.w1(32'h3b0255d4),
	.w2(32'hbacd39f0),
	.w3(32'hbb425c4d),
	.w4(32'hbbc58530),
	.w5(32'hbb8e3889),
	.w6(32'h3b113238),
	.w7(32'hbb47e3aa),
	.w8(32'h3b36cd12),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5892eb),
	.w1(32'hbc13722f),
	.w2(32'hbc3123cc),
	.w3(32'hbc2aafb6),
	.w4(32'hbc55db95),
	.w5(32'hbbf4b9a3),
	.w6(32'hbc17b5e2),
	.w7(32'hbc2ef4f2),
	.w8(32'hbbd65f19),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4338aa),
	.w1(32'h3c52ef69),
	.w2(32'hbbde94b5),
	.w3(32'hbad90659),
	.w4(32'h3ba7ea48),
	.w5(32'hba9909dc),
	.w6(32'h3a1b1fb4),
	.w7(32'hbb9aa890),
	.w8(32'hbc1b77c9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9355d8),
	.w1(32'h3ce04ef5),
	.w2(32'hbbc001dc),
	.w3(32'hbb3d76c0),
	.w4(32'h3adcd47c),
	.w5(32'h3b47f73b),
	.w6(32'h3bcf4daa),
	.w7(32'h3b57b5b6),
	.w8(32'hbb1b94d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e1884),
	.w1(32'hbcb5259c),
	.w2(32'h3cd184cc),
	.w3(32'h3b0cd40f),
	.w4(32'hbb8eb845),
	.w5(32'h3ba67ae6),
	.w6(32'hbc411243),
	.w7(32'h3c067328),
	.w8(32'h3c5306f9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce9d4cb),
	.w1(32'hbc2965e3),
	.w2(32'hbd04e728),
	.w3(32'h3b9f3257),
	.w4(32'hbc631670),
	.w5(32'hbc0348a1),
	.w6(32'hba2ee338),
	.w7(32'hbbbcd16e),
	.w8(32'hbbae6ead),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b23470),
	.w1(32'h3d08c527),
	.w2(32'h3bda49ae),
	.w3(32'h3bd6c312),
	.w4(32'h3c077594),
	.w5(32'h3c562eb5),
	.w6(32'h3c2caf74),
	.w7(32'h3c001a69),
	.w8(32'hbc3656ff),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfca283),
	.w1(32'hbbd210c7),
	.w2(32'hbc9de885),
	.w3(32'hbbde642e),
	.w4(32'hbad5ec35),
	.w5(32'hbcbce087),
	.w6(32'hbb27f75c),
	.w7(32'hbc677fc5),
	.w8(32'h3b1d1385),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb3d46),
	.w1(32'hbb2cf8b8),
	.w2(32'h3ae514fe),
	.w3(32'hbba72002),
	.w4(32'h3b4a4d47),
	.w5(32'h39a6d833),
	.w6(32'h3af69031),
	.w7(32'hba9c2398),
	.w8(32'hbb6f60bf),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867faeb),
	.w1(32'hbab33f83),
	.w2(32'h3bad13e8),
	.w3(32'h3a081618),
	.w4(32'hb8ebf3f4),
	.w5(32'h3b47aa9c),
	.w6(32'h3a41f786),
	.w7(32'h3b4516b1),
	.w8(32'h3b78226d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29c206),
	.w1(32'hbbc208bf),
	.w2(32'h3beb2b51),
	.w3(32'hbad20607),
	.w4(32'hbb2ffb41),
	.w5(32'hbac29099),
	.w6(32'h3ad99e1e),
	.w7(32'h3b4d188b),
	.w8(32'h3b9bb837),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6690e),
	.w1(32'hbc1de071),
	.w2(32'h3cc38a05),
	.w3(32'h3ae46bea),
	.w4(32'hbc015787),
	.w5(32'hbb75ee37),
	.w6(32'hbbf56276),
	.w7(32'hb85b5dd1),
	.w8(32'hbb864b8b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ba451),
	.w1(32'hbc296708),
	.w2(32'h3b95e801),
	.w3(32'hbc068418),
	.w4(32'hbaca093c),
	.w5(32'hbb17db84),
	.w6(32'hbb258b43),
	.w7(32'hbb6606c3),
	.w8(32'hbc4386de),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f97d),
	.w1(32'h3d0c095f),
	.w2(32'hbc1e6d21),
	.w3(32'hbc60acb3),
	.w4(32'h3bc53867),
	.w5(32'h3b1114e4),
	.w6(32'h3bf2b9fe),
	.w7(32'h399489cc),
	.w8(32'hbc08f24b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc97bef),
	.w1(32'hbbc9cde2),
	.w2(32'h3b08f6ec),
	.w3(32'hbbba1a49),
	.w4(32'h3b362da6),
	.w5(32'hbb7079fe),
	.w6(32'h3ad4af06),
	.w7(32'hbb16cbee),
	.w8(32'hbc341bf5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf83156),
	.w1(32'h3c151e38),
	.w2(32'hbcb00110),
	.w3(32'hbc884c7e),
	.w4(32'hbb0978f8),
	.w5(32'hbc28c182),
	.w6(32'hbbfd0ce8),
	.w7(32'hbb75dd3a),
	.w8(32'hba1bc13e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c89c0),
	.w1(32'h3b1d578f),
	.w2(32'hbcc087d6),
	.w3(32'hbbe66834),
	.w4(32'hbac1b164),
	.w5(32'hbc1f836c),
	.w6(32'hbbb40444),
	.w7(32'hb990cda7),
	.w8(32'hba60277e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35c9b6),
	.w1(32'hbd1c28b6),
	.w2(32'h3c0b8dde),
	.w3(32'hbbff0236),
	.w4(32'hbba373c1),
	.w5(32'hbc0a7dd2),
	.w6(32'hbc0a99a1),
	.w7(32'hbbe5e07e),
	.w8(32'h3c33d652),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfe49d2),
	.w1(32'hbc036beb),
	.w2(32'hba90ac9b),
	.w3(32'h3abdef89),
	.w4(32'hbb1c89b0),
	.w5(32'hbb716305),
	.w6(32'hbbbe9454),
	.w7(32'hbb6c60d9),
	.w8(32'hbbf5121e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2b78d),
	.w1(32'hbb9e20df),
	.w2(32'h3c844d4b),
	.w3(32'hbb97f81f),
	.w4(32'h3a781926),
	.w5(32'h3bba4e8b),
	.w6(32'hbc535532),
	.w7(32'hbbcf7601),
	.w8(32'h3bbb7282),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19de07),
	.w1(32'hba063a5a),
	.w2(32'h3b63fa7a),
	.w3(32'h3abe5b52),
	.w4(32'h3b3a0c1b),
	.w5(32'h3b903572),
	.w6(32'hba16b4eb),
	.w7(32'h3b3dc998),
	.w8(32'hbb3506e6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6173),
	.w1(32'hbb88225d),
	.w2(32'hba0b7c66),
	.w3(32'hbb61ee7f),
	.w4(32'hba2fa7b6),
	.w5(32'h3ac3fa5e),
	.w6(32'hbb74b2e0),
	.w7(32'hba0c38db),
	.w8(32'hba405d5b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81201),
	.w1(32'h3cc8902e),
	.w2(32'hbc40c892),
	.w3(32'hbb66a167),
	.w4(32'hbbafa423),
	.w5(32'hba58deec),
	.w6(32'h3bc57797),
	.w7(32'h3b25b7df),
	.w8(32'hbbde5e12),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb01bd5),
	.w1(32'hbd004212),
	.w2(32'h3d0c6fe8),
	.w3(32'h3bfad836),
	.w4(32'hbc06654c),
	.w5(32'h3ba7a1d6),
	.w6(32'hbc858178),
	.w7(32'hbac47ce1),
	.w8(32'h3ca01f71),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d25baca),
	.w1(32'hbc9b8912),
	.w2(32'h3b88ef9f),
	.w3(32'h3c93acfa),
	.w4(32'hbb924734),
	.w5(32'hbb34b419),
	.w6(32'hbb9b9e13),
	.w7(32'hbb4f5abf),
	.w8(32'hbb540915),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ead3c),
	.w1(32'h3cc69e5b),
	.w2(32'hbb576cb0),
	.w3(32'hbbb97703),
	.w4(32'h3984e36d),
	.w5(32'h3b5faefd),
	.w6(32'hb7adadf1),
	.w7(32'hb9c1b9c9),
	.w8(32'hbb5e7cc9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95d673),
	.w1(32'h3cf7b817),
	.w2(32'hbbdec8da),
	.w3(32'hb9f2a1d1),
	.w4(32'h3b87fd50),
	.w5(32'h3b322caf),
	.w6(32'h3bdcdab9),
	.w7(32'h3a087e10),
	.w8(32'hbbf112ed),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0043e),
	.w1(32'h3cb84db1),
	.w2(32'hbbbb1db0),
	.w3(32'hbb1696ca),
	.w4(32'hbb7d49d8),
	.w5(32'h3b517e7d),
	.w6(32'h3bd44653),
	.w7(32'hbb3668f9),
	.w8(32'hbc69e0dd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca47c5d),
	.w1(32'hbbbc1185),
	.w2(32'h3b365540),
	.w3(32'h3b29c3a0),
	.w4(32'hbaf60d22),
	.w5(32'hbac4010c),
	.w6(32'hbae7a21a),
	.w7(32'hbb0e0e8e),
	.w8(32'hbc0ed5c8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd31c9),
	.w1(32'hbb1b9131),
	.w2(32'hbc838aa6),
	.w3(32'hbc5c735d),
	.w4(32'hba8edd38),
	.w5(32'hbb5c5834),
	.w6(32'hbc140397),
	.w7(32'hbc0411bd),
	.w8(32'hbb5349fb),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b051567),
	.w1(32'h3cf5d117),
	.w2(32'hbc5ddb60),
	.w3(32'hbb6ad1d4),
	.w4(32'hbbe59c20),
	.w5(32'hbacd941d),
	.w6(32'hbbdaf24c),
	.w7(32'hbbfdc083),
	.w8(32'hba4269e2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bd20c),
	.w1(32'hbbbb0f35),
	.w2(32'h3a77dc4f),
	.w3(32'h3c205dd3),
	.w4(32'h3b962041),
	.w5(32'hbaef23e1),
	.w6(32'h3b1495be),
	.w7(32'hba66ee2b),
	.w8(32'hbc681766),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d678b),
	.w1(32'h3c05b1b1),
	.w2(32'hbb832723),
	.w3(32'hbc8f9dbf),
	.w4(32'h3c1f966a),
	.w5(32'hbbf390e8),
	.w6(32'h3bce6465),
	.w7(32'hbc182059),
	.w8(32'hbc646b51),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc820de0),
	.w1(32'h3c924d46),
	.w2(32'hbc4c3a9b),
	.w3(32'hb9e6e0b4),
	.w4(32'hbbeaf705),
	.w5(32'h3b4c6a29),
	.w6(32'hbb4bd237),
	.w7(32'hbafe0b6d),
	.w8(32'h3a8f7fb3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc303f81),
	.w1(32'hbb58613a),
	.w2(32'hbb33c871),
	.w3(32'h3c1d49f0),
	.w4(32'hbb8c2a37),
	.w5(32'hbb5ac2ae),
	.w6(32'h3b0502b4),
	.w7(32'h3b2e50b4),
	.w8(32'h3b1dc9c7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8354b),
	.w1(32'hbb9dce12),
	.w2(32'h3b871b1e),
	.w3(32'hbbdc3a78),
	.w4(32'h37beb7b6),
	.w5(32'hba224dc1),
	.w6(32'h3a04e01f),
	.w7(32'h39abc59e),
	.w8(32'hbc044fa7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f9a9),
	.w1(32'hbabefd1f),
	.w2(32'hbac1780e),
	.w3(32'hbbf75211),
	.w4(32'hbb81fc80),
	.w5(32'hbaef9281),
	.w6(32'hbbb1cadc),
	.w7(32'hbb5169b6),
	.w8(32'hbba7dc2b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581bc0),
	.w1(32'hbbc74489),
	.w2(32'h38d65950),
	.w3(32'hbabeb600),
	.w4(32'h3a86f660),
	.w5(32'hbb235b88),
	.w6(32'h3a0adcd1),
	.w7(32'hbb420115),
	.w8(32'hbc592f0a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf184a6),
	.w1(32'h3bb05f64),
	.w2(32'h3b9d7851),
	.w3(32'hbc3d79c1),
	.w4(32'h3aaf6c49),
	.w5(32'h3ae78111),
	.w6(32'h3b92be26),
	.w7(32'h3bfb46d9),
	.w8(32'h3b9f7bb2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0896c3),
	.w1(32'hba0d528c),
	.w2(32'h3c5c33ea),
	.w3(32'h386ff88a),
	.w4(32'h3a9229bd),
	.w5(32'h3ba2b744),
	.w6(32'h3b97435f),
	.w7(32'h3c0a797c),
	.w8(32'hbb1b737f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad75209),
	.w1(32'hbc48a6e1),
	.w2(32'h3c8efc61),
	.w3(32'hbb9cc9d0),
	.w4(32'h3b2374ef),
	.w5(32'h3c14f43b),
	.w6(32'hbb14df61),
	.w7(32'h3b6db1cb),
	.w8(32'h3b3e8cd6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c107438),
	.w1(32'h3c88c5a0),
	.w2(32'hbc059370),
	.w3(32'h3bed56ae),
	.w4(32'hbb2f7f37),
	.w5(32'hba3b6e9a),
	.w6(32'h3b25e8f9),
	.w7(32'hba613410),
	.w8(32'hbb824b57),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ba33a),
	.w1(32'hbb03060c),
	.w2(32'h3b614ea3),
	.w3(32'h3b1f5f2a),
	.w4(32'h3b6d62fc),
	.w5(32'h3ab9b90c),
	.w6(32'h3b790446),
	.w7(32'h3a8be80a),
	.w8(32'hbb919f25),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085dd1),
	.w1(32'h3c6db4ee),
	.w2(32'hbc859c49),
	.w3(32'hbc3fd3ae),
	.w4(32'hbc3a9a77),
	.w5(32'hba5137dd),
	.w6(32'hbc206999),
	.w7(32'hbc1872bd),
	.w8(32'hbb80394c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4da403),
	.w1(32'h3cc03536),
	.w2(32'hb9f54f8c),
	.w3(32'h3c2b28f6),
	.w4(32'h3c067c9c),
	.w5(32'h3bb29637),
	.w6(32'h3b9baeb0),
	.w7(32'hbab3b7de),
	.w8(32'hbc579eb5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d13b5),
	.w1(32'hbce6a9bc),
	.w2(32'h3b83f675),
	.w3(32'hbae4b4a8),
	.w4(32'hbc093562),
	.w5(32'hbb9b40b6),
	.w6(32'hbc0eeea3),
	.w7(32'hba81eeaf),
	.w8(32'h3b02abbe),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8575dc),
	.w1(32'hbc07eada),
	.w2(32'hbb194d75),
	.w3(32'hbad8f54d),
	.w4(32'hbb06792e),
	.w5(32'hbad9a9bb),
	.w6(32'h383fbaa6),
	.w7(32'hbaa5f995),
	.w8(32'hbbaf8e70),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd856d1),
	.w1(32'hbbce3c1c),
	.w2(32'hbb3797d6),
	.w3(32'hbb7d9f02),
	.w4(32'hbbfe6413),
	.w5(32'hbad43459),
	.w6(32'hbb1f3582),
	.w7(32'h3aaf19de),
	.w8(32'h3b5a88f5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2723bc),
	.w1(32'hbbb186ae),
	.w2(32'h3befd1e4),
	.w3(32'h398eb5d9),
	.w4(32'h3b457fa4),
	.w5(32'h3b343e6c),
	.w6(32'h3b51008f),
	.w7(32'h3b7ba4bf),
	.w8(32'hbb53b558),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a235fa2),
	.w1(32'h3c2ba18d),
	.w2(32'h3c1c52d9),
	.w3(32'h39f5e1ed),
	.w4(32'h3c492ead),
	.w5(32'h3c61db5a),
	.w6(32'hbac7859e),
	.w7(32'h3a015f85),
	.w8(32'hbbd070e4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfeb787),
	.w1(32'hbbb72796),
	.w2(32'hbb94012c),
	.w3(32'hbac9b4f3),
	.w4(32'hb91d45ea),
	.w5(32'hbb87429a),
	.w6(32'hbb7bded5),
	.w7(32'hbae4deb5),
	.w8(32'h3b4e7e31),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62de2e),
	.w1(32'hbce85621),
	.w2(32'hbbaf36fd),
	.w3(32'hba409513),
	.w4(32'hbc9172ba),
	.w5(32'hbbbcd613),
	.w6(32'hbcbfcebb),
	.w7(32'hbc0f0513),
	.w8(32'h3b593398),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5bfb2),
	.w1(32'hbb3be1d5),
	.w2(32'h3b830b1f),
	.w3(32'h3c1a03f7),
	.w4(32'h3c1f1f80),
	.w5(32'h3a2bf74a),
	.w6(32'h3bd69614),
	.w7(32'h39c82862),
	.w8(32'hbc40aa7e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fcc7b),
	.w1(32'hbc6b6a5a),
	.w2(32'hbc591a14),
	.w3(32'hbca7176b),
	.w4(32'hbc9fbf23),
	.w5(32'hbc1ec75d),
	.w6(32'hbca7e622),
	.w7(32'hbc3f6398),
	.w8(32'hbc03f53d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d4fe2),
	.w1(32'hbc79a002),
	.w2(32'hbca5925b),
	.w3(32'h3b999025),
	.w4(32'h3a76e92c),
	.w5(32'hbce8194a),
	.w6(32'h3bb66e93),
	.w7(32'hbc54811c),
	.w8(32'hbc2d70ed),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc966ed3),
	.w1(32'h3c05378a),
	.w2(32'hbbaeb1d1),
	.w3(32'hbbb62b95),
	.w4(32'hba8324ff),
	.w5(32'hbbd168fd),
	.w6(32'h3c10d151),
	.w7(32'h3c3a2756),
	.w8(32'h3bda9b98),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff48bf),
	.w1(32'h3d489f35),
	.w2(32'hbc7693ba),
	.w3(32'hbb8f7d77),
	.w4(32'h396780be),
	.w5(32'h3b2b128a),
	.w6(32'h3abf7d3e),
	.w7(32'h3a250ac0),
	.w8(32'h3b97a740),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8049d5),
	.w1(32'h3ccff142),
	.w2(32'h3b592766),
	.w3(32'h3c328e84),
	.w4(32'hbb00ec1a),
	.w5(32'h3c1aaa0f),
	.w6(32'h38d2b8f7),
	.w7(32'h3bc4fb72),
	.w8(32'hbb1cc2aa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc8c747),
	.w1(32'h3c90eece),
	.w2(32'hbc9adc92),
	.w3(32'hbbfc5523),
	.w4(32'hbc0cdd30),
	.w5(32'hbbc81121),
	.w6(32'hbc01bb27),
	.w7(32'hbc17817d),
	.w8(32'hbb3d159b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce1e5b),
	.w1(32'h3c3eec26),
	.w2(32'hbc9b9466),
	.w3(32'h3c041f46),
	.w4(32'h3a8864c7),
	.w5(32'hbbe5010b),
	.w6(32'h3bb64ec0),
	.w7(32'hbb9a4444),
	.w8(32'hbbec3467),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84c4fb),
	.w1(32'hbb8bb855),
	.w2(32'h3bd900d8),
	.w3(32'hbb482a09),
	.w4(32'h3a119582),
	.w5(32'h3a2afd2b),
	.w6(32'hba5c01ab),
	.w7(32'h3b1c3d0d),
	.w8(32'hbabc23d9),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034d16),
	.w1(32'h3ce44731),
	.w2(32'hbbe7789a),
	.w3(32'hbbb466a4),
	.w4(32'h3bc898de),
	.w5(32'hba65beeb),
	.w6(32'h3bbc67ed),
	.w7(32'hbb310e54),
	.w8(32'hbc29e0ba),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc985ea6),
	.w1(32'h3ce8c5d8),
	.w2(32'hbb5521cd),
	.w3(32'hba4da777),
	.w4(32'h3b132040),
	.w5(32'h3b4f89b9),
	.w6(32'h3b6fdad5),
	.w7(32'h3ac157f1),
	.w8(32'h3b6ac78c),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc329f),
	.w1(32'hbca7bc81),
	.w2(32'h3c7e824f),
	.w3(32'h3c248646),
	.w4(32'hbada82c0),
	.w5(32'h3bc355ff),
	.w6(32'hbbdbfc7d),
	.w7(32'h3b949250),
	.w8(32'h3ba6b9aa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac6efd),
	.w1(32'h3ce349ac),
	.w2(32'hbca2c495),
	.w3(32'hba688137),
	.w4(32'h3b55a5be),
	.w5(32'hbb14bc00),
	.w6(32'h3c56fb8f),
	.w7(32'hb8ce8494),
	.w8(32'hbc31770b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0c254),
	.w1(32'hbc0e2841),
	.w2(32'hbd73dc12),
	.w3(32'hbb63774e),
	.w4(32'h3b32d8e2),
	.w5(32'hbcd3aac1),
	.w6(32'hbc680611),
	.w7(32'hbc98eeb0),
	.w8(32'h3ad2f6b5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a78b8),
	.w1(32'h3cdab060),
	.w2(32'hbbf8a363),
	.w3(32'hba74d7ff),
	.w4(32'hbb064d33),
	.w5(32'h3b8889eb),
	.w6(32'h3c3afecc),
	.w7(32'h3b980784),
	.w8(32'hbc0cc3e0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaee7f1),
	.w1(32'hbc3c798c),
	.w2(32'h3c385e98),
	.w3(32'hbb226e82),
	.w4(32'hbb2e4de0),
	.w5(32'hbb48fbe8),
	.w6(32'hbbbd8fd0),
	.w7(32'hba4daa09),
	.w8(32'hbbf23a98),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57036b),
	.w1(32'h3c669837),
	.w2(32'hbc1bc1e3),
	.w3(32'hbc4f45bc),
	.w4(32'h3c1409b2),
	.w5(32'h3b694d8f),
	.w6(32'h3bc594b0),
	.w7(32'h3b753d7d),
	.w8(32'h3c11dcb4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e1bd9),
	.w1(32'h3d1c6eb5),
	.w2(32'hbc116bdb),
	.w3(32'h3c0dd6b5),
	.w4(32'h3a9c903d),
	.w5(32'h3b3f2f13),
	.w6(32'h3b3283cd),
	.w7(32'h3a91bd3b),
	.w8(32'h3b80190f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b248b),
	.w1(32'h3d006551),
	.w2(32'hbba8c80e),
	.w3(32'h3c034612),
	.w4(32'h3ba34b84),
	.w5(32'h3b0c7b32),
	.w6(32'h3be6363b),
	.w7(32'h3a89e98a),
	.w8(32'hbbce475b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadd756),
	.w1(32'h3d0b1941),
	.w2(32'hbbba6236),
	.w3(32'hba56254b),
	.w4(32'h3bb486e0),
	.w5(32'h3b577836),
	.w6(32'h3c10c02c),
	.w7(32'h3aef5a29),
	.w8(32'hbbaccc60),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8b14d),
	.w1(32'hba8b94de),
	.w2(32'hba2f0729),
	.w3(32'hb99c6d19),
	.w4(32'h396bd53b),
	.w5(32'hbbabcd63),
	.w6(32'hbc182160),
	.w7(32'hbc1915fd),
	.w8(32'hbbba6b8b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9c31),
	.w1(32'hbc25c78e),
	.w2(32'hbca81dc4),
	.w3(32'hbbb38648),
	.w4(32'hb95e4447),
	.w5(32'hbcdc82d5),
	.w6(32'h3b177299),
	.w7(32'hbcd83d0d),
	.w8(32'hbccab229),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfd6d8c),
	.w1(32'h3cb6b22b),
	.w2(32'h3bc51dc5),
	.w3(32'hbcea136a),
	.w4(32'h3bde9786),
	.w5(32'h3bded0f1),
	.w6(32'h3ba8af34),
	.w7(32'h3b62c178),
	.w8(32'hbc487e5d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca880b1),
	.w1(32'h3c828e8e),
	.w2(32'hbc687bf3),
	.w3(32'hbc276ddf),
	.w4(32'h3bc578e9),
	.w5(32'hbbc1bd41),
	.w6(32'hb954b647),
	.w7(32'hbc0850e6),
	.w8(32'hbc8b7bd1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadf363),
	.w1(32'h3d24da47),
	.w2(32'hbbd4ae50),
	.w3(32'hbc332685),
	.w4(32'h3c288e71),
	.w5(32'h3ba7334e),
	.w6(32'h3c5da606),
	.w7(32'h3b8fee50),
	.w8(32'hbbfbce92),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc13ec4),
	.w1(32'hba83bffa),
	.w2(32'hbbf7ef41),
	.w3(32'hbacdd7a8),
	.w4(32'hb915a0af),
	.w5(32'hbbcb4c3f),
	.w6(32'hbc291db6),
	.w7(32'hbb40dc8d),
	.w8(32'h3abd1c12),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37cce0),
	.w1(32'h3d15218c),
	.w2(32'h3c8d9699),
	.w3(32'hbc08dec3),
	.w4(32'h3c107963),
	.w5(32'h3c8494ca),
	.w6(32'h3bfff339),
	.w7(32'h3c50f3de),
	.w8(32'hbc42752c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0793a2),
	.w1(32'h3cbf2bac),
	.w2(32'hbc6e6268),
	.w3(32'hbc143b2d),
	.w4(32'hbb829a1b),
	.w5(32'hbba1743e),
	.w6(32'h3a1a8c68),
	.w7(32'hbba46752),
	.w8(32'hbc2fc415),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb47f37),
	.w1(32'h399576b5),
	.w2(32'h399db4bb),
	.w3(32'hbaada4c1),
	.w4(32'h3a36428c),
	.w5(32'h394429a4),
	.w6(32'h3a774ca5),
	.w7(32'h3a0be0dc),
	.w8(32'hb9835d7f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4ff3b),
	.w1(32'hb9dbefae),
	.w2(32'hb9616844),
	.w3(32'hbaa7e12a),
	.w4(32'hb9a4bf9c),
	.w5(32'h398e716e),
	.w6(32'hba15e4ab),
	.w7(32'hba638429),
	.w8(32'hb9fffcbe),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c30af),
	.w1(32'hb94b8192),
	.w2(32'h3a77349a),
	.w3(32'hb604bfd0),
	.w4(32'h38296d03),
	.w5(32'h3aa214f0),
	.w6(32'hba8c267a),
	.w7(32'hba2fe7f4),
	.w8(32'h39f7cf97),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fe1e6),
	.w1(32'hba62ae2a),
	.w2(32'hbaae1d2a),
	.w3(32'hba8bcd73),
	.w4(32'hba86858c),
	.w5(32'hba9a1779),
	.w6(32'hba57a850),
	.w7(32'hba87ec4d),
	.w8(32'hba2fac3a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001eeb),
	.w1(32'hbada7817),
	.w2(32'hba841bf2),
	.w3(32'hbad4d48f),
	.w4(32'hb9ea6868),
	.w5(32'h39c30f17),
	.w6(32'hbab529db),
	.w7(32'hba5628e0),
	.w8(32'hb8c390aa),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91c2b29),
	.w1(32'h3905184d),
	.w2(32'hb9558a37),
	.w3(32'h3a318282),
	.w4(32'h3a62868a),
	.w5(32'h3929314f),
	.w6(32'h3a3b604d),
	.w7(32'h39e22a06),
	.w8(32'hb994d6eb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d98d4),
	.w1(32'h395fb7b8),
	.w2(32'h3a4c72ab),
	.w3(32'hb9ae8dab),
	.w4(32'h39e4664e),
	.w5(32'h3a2ec6a2),
	.w6(32'hb9110019),
	.w7(32'h394dc209),
	.w8(32'h3a6c74cb),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911c6cc),
	.w1(32'h3b0b5fc5),
	.w2(32'h3b5d5476),
	.w3(32'h3a4624c5),
	.w4(32'h3b26296e),
	.w5(32'h3b48ec85),
	.w6(32'h39b67c10),
	.w7(32'h3b0ce844),
	.w8(32'h3b208460),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc4887),
	.w1(32'hbb886b34),
	.w2(32'hbb857dbb),
	.w3(32'hbb7dfff9),
	.w4(32'hbb9ae4e2),
	.w5(32'hbb28f1d3),
	.w6(32'hbbcb4129),
	.w7(32'hbbb0dcc1),
	.w8(32'hbae623bf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d3aa5),
	.w1(32'h3a876d40),
	.w2(32'h3ada9a46),
	.w3(32'h3b43c76c),
	.w4(32'h3ad6180b),
	.w5(32'h3a07a242),
	.w6(32'h3b259718),
	.w7(32'h3aaefc66),
	.w8(32'h3a5c8543),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a5983),
	.w1(32'h39c70a21),
	.w2(32'hb73d7a97),
	.w3(32'h3a0b2e72),
	.w4(32'h3aa1f241),
	.w5(32'h3a0df453),
	.w6(32'h38c77af3),
	.w7(32'h3a33477a),
	.w8(32'h388e5894),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbbd7),
	.w1(32'hbb446e42),
	.w2(32'hbb433f6f),
	.w3(32'hbb417d02),
	.w4(32'hbb3b2285),
	.w5(32'hba8a52b8),
	.w6(32'hbb96d47b),
	.w7(32'hbb1e295b),
	.w8(32'hb9cad771),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b64532),
	.w1(32'h3963438a),
	.w2(32'h3ab28be8),
	.w3(32'h3a0e52b6),
	.w4(32'h3a86bfa2),
	.w5(32'h3a30f4cc),
	.w6(32'h39778e4b),
	.w7(32'hb744a274),
	.w8(32'h39e59db5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05843c),
	.w1(32'h38b05a92),
	.w2(32'h3996ba34),
	.w3(32'h38a2ca02),
	.w4(32'h395b1d67),
	.w5(32'hb895ee39),
	.w6(32'h39a57a22),
	.w7(32'h395429a2),
	.w8(32'hb9e33241),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e27c76),
	.w1(32'h381220ea),
	.w2(32'h399d9835),
	.w3(32'hb931fb20),
	.w4(32'h39786f82),
	.w5(32'h396d4a78),
	.w6(32'hb9574882),
	.w7(32'hb96f198b),
	.w8(32'hb8dbf390),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa29df6),
	.w1(32'h3b4e08eb),
	.w2(32'h3b3bce15),
	.w3(32'h3bbc658a),
	.w4(32'h3baa572e),
	.w5(32'h3ad94218),
	.w6(32'h3ba6f9a1),
	.w7(32'h3b8ecd43),
	.w8(32'h3a10d92d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03e330),
	.w1(32'hba31f5a5),
	.w2(32'hba8effc9),
	.w3(32'hb9864b86),
	.w4(32'h3886e0ae),
	.w5(32'hba85a77c),
	.w6(32'hb91020d8),
	.w7(32'h3a617283),
	.w8(32'hb88b1979),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9995ac3),
	.w1(32'hb92b2e08),
	.w2(32'hb71594a6),
	.w3(32'hba52c87e),
	.w4(32'hb94b9258),
	.w5(32'hb7ff2de7),
	.w6(32'hb931ed38),
	.w7(32'h38f6b09d),
	.w8(32'h39418ab3),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f961cb),
	.w1(32'h39c7ca31),
	.w2(32'h393c54e3),
	.w3(32'h39035daa),
	.w4(32'h392e830d),
	.w5(32'h3938d8b8),
	.w6(32'h399a481e),
	.w7(32'h39a9d9d8),
	.w8(32'h397eb14b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac9c53),
	.w1(32'hb8cd5a21),
	.w2(32'h39fcee4a),
	.w3(32'h3a86da50),
	.w4(32'hb9486812),
	.w5(32'hb91cc318),
	.w6(32'h3a47e818),
	.w7(32'hb98fb9aa),
	.w8(32'hb99ccf39),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a54a5),
	.w1(32'h3b04a830),
	.w2(32'h39a2ef6b),
	.w3(32'h3b5a1980),
	.w4(32'h3b1ef1b2),
	.w5(32'hb8af456b),
	.w6(32'h3ad71345),
	.w7(32'h3a901a72),
	.w8(32'hb9d8dc9b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c36cc),
	.w1(32'hba22ecae),
	.w2(32'h3ae8e3a6),
	.w3(32'h3a2c3702),
	.w4(32'hb9c41bb7),
	.w5(32'h3aa31889),
	.w6(32'h3939e421),
	.w7(32'hba850ba7),
	.w8(32'h3a9832ea),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b05456),
	.w1(32'hb9dd8523),
	.w2(32'hb994f05b),
	.w3(32'h38d20d31),
	.w4(32'hb99c6249),
	.w5(32'hb9292ba6),
	.w6(32'hb9b691e8),
	.w7(32'hb8ac4dcc),
	.w8(32'hb97416a6),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ab6ea),
	.w1(32'h3836daf0),
	.w2(32'h3acdca49),
	.w3(32'h3a9a7e7d),
	.w4(32'h3ace6e1e),
	.w5(32'h3b065b4e),
	.w6(32'h397af07d),
	.w7(32'hb9003bb6),
	.w8(32'h399d4d2c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec6907),
	.w1(32'h3acb8412),
	.w2(32'h3b1019a9),
	.w3(32'h3b57e304),
	.w4(32'h3af2d37e),
	.w5(32'h3a9c7590),
	.w6(32'h3b1c65e3),
	.w7(32'h3aa99a5a),
	.w8(32'h39d9a7bf),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c8e7),
	.w1(32'hbb546df5),
	.w2(32'hbb5c4206),
	.w3(32'hbb2393d1),
	.w4(32'hbb81668c),
	.w5(32'hbb2cad50),
	.w6(32'hbb88c338),
	.w7(32'hbb76e57c),
	.w8(32'hbb12c2b9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de682e),
	.w1(32'h3a524f9c),
	.w2(32'h3a5c4ead),
	.w3(32'h3b2b9887),
	.w4(32'h3b4ba24e),
	.w5(32'h3aa99029),
	.w6(32'h3b141fe9),
	.w7(32'h3a93c83f),
	.w8(32'h39c5c038),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac268f9),
	.w1(32'h3b23dcbf),
	.w2(32'h3ab863d1),
	.w3(32'h3b21e8cf),
	.w4(32'h3b3d202e),
	.w5(32'h3aa299a7),
	.w6(32'h3b5748b5),
	.w7(32'h3b0633ff),
	.w8(32'h3a0a88dc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c08c2),
	.w1(32'h3a207e13),
	.w2(32'h39c732c3),
	.w3(32'h3a7bb72c),
	.w4(32'h3adfc097),
	.w5(32'h3a6b2553),
	.w6(32'h3aac2998),
	.w7(32'h3a9aa72a),
	.w8(32'h3a670fc0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baeb17),
	.w1(32'h37bcfaf2),
	.w2(32'hb97772a1),
	.w3(32'h3a892f05),
	.w4(32'h3a193de0),
	.w5(32'hb914263b),
	.w6(32'h3ab6c9d4),
	.w7(32'h397a2099),
	.w8(32'hbaa46e1f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a18eb66),
	.w1(32'h3b05d72e),
	.w2(32'h3abeff95),
	.w3(32'h3b30ac5c),
	.w4(32'h3b7e4991),
	.w5(32'h3b0012d4),
	.w6(32'h3b6bb7b9),
	.w7(32'h3b5a2cc6),
	.w8(32'h3a919423),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6cafd8),
	.w1(32'h3abf3b3d),
	.w2(32'h3a3c786f),
	.w3(32'h3a9cdd4f),
	.w4(32'h3aafc345),
	.w5(32'h3a23581d),
	.w6(32'h3a9bf363),
	.w7(32'h3a7e3913),
	.w8(32'h3a2e9e6a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed0d05),
	.w1(32'hba9a717c),
	.w2(32'hbaa96e2d),
	.w3(32'hba6abab5),
	.w4(32'hbad2e0b0),
	.w5(32'hba6036d3),
	.w6(32'hbb103c58),
	.w7(32'hbacb8a18),
	.w8(32'hb9639c73),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866968c),
	.w1(32'h390b729f),
	.w2(32'h38dec17e),
	.w3(32'h398c5a7d),
	.w4(32'h3974845a),
	.w5(32'h38cf24fc),
	.w6(32'h393b6cde),
	.w7(32'h396b7654),
	.w8(32'h38cae6eb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb969d6cb),
	.w1(32'h397b829b),
	.w2(32'h395f684d),
	.w3(32'hb9fb3fbb),
	.w4(32'h38517334),
	.w5(32'h3a4ecb59),
	.w6(32'hb8c93658),
	.w7(32'hba2f25f2),
	.w8(32'h39070267),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952e427),
	.w1(32'h3a391f43),
	.w2(32'h3a26bd2a),
	.w3(32'h3a09f27e),
	.w4(32'h3a1936cf),
	.w5(32'h3955a2d7),
	.w6(32'h3a182044),
	.w7(32'h39d0674c),
	.w8(32'h3a128c2e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da530e),
	.w1(32'hb8d5edeb),
	.w2(32'h3a0f722c),
	.w3(32'h3a60c91b),
	.w4(32'h3a84e663),
	.w5(32'h39e089bd),
	.w6(32'h3a04ea24),
	.w7(32'h3994a4af),
	.w8(32'hb910a7f1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c868d8),
	.w1(32'h38b26ddb),
	.w2(32'hb78f41fb),
	.w3(32'hb9a7ee21),
	.w4(32'hb5921215),
	.w5(32'h389d9617),
	.w6(32'hb8e36dc3),
	.w7(32'h3987e88e),
	.w8(32'h38b5e45d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0890da),
	.w1(32'h3a8ab897),
	.w2(32'h3ad93274),
	.w3(32'h3a6163f6),
	.w4(32'h3a044da6),
	.w5(32'h3aa57d65),
	.w6(32'h3a137e87),
	.w7(32'hb98495e2),
	.w8(32'h39b4f59b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959c6a5),
	.w1(32'hb97e5e12),
	.w2(32'hb7b94526),
	.w3(32'hb8f23285),
	.w4(32'hb8ad3ba4),
	.w5(32'h38c0c7a5),
	.w6(32'hb906b440),
	.w7(32'h380a2a96),
	.w8(32'h3944db9e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923a34f),
	.w1(32'hb9c80b92),
	.w2(32'hb9ce083e),
	.w3(32'h39893e8e),
	.w4(32'hb94c1f5b),
	.w5(32'hb97fadd0),
	.w6(32'hb8531684),
	.w7(32'hb9013db3),
	.w8(32'hb8fa1184),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08a802),
	.w1(32'h3a20ebe9),
	.w2(32'h38f1d263),
	.w3(32'h3b369d02),
	.w4(32'h3b0967cc),
	.w5(32'h38c66336),
	.w6(32'h3b4252b3),
	.w7(32'h3adee84d),
	.w8(32'h39019d2d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f8b60),
	.w1(32'hbad8920f),
	.w2(32'hbb001ced),
	.w3(32'hbb2fd3da),
	.w4(32'hbb31fe2f),
	.w5(32'hbaa661a9),
	.w6(32'hbb8863b5),
	.w7(32'hbb6166d3),
	.w8(32'hbaeecdf0),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd163),
	.w1(32'h3a4c94fc),
	.w2(32'h395ae1ba),
	.w3(32'h3aa1f3a6),
	.w4(32'h39b54eb8),
	.w5(32'hb967e962),
	.w6(32'h3a7cbe82),
	.w7(32'h3a1d1a64),
	.w8(32'hb8d45622),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c8d0b),
	.w1(32'h3b084ff6),
	.w2(32'h3af668b6),
	.w3(32'h3b45f0ac),
	.w4(32'h3b4363ac),
	.w5(32'h3acf93a2),
	.w6(32'h3b3c0ebf),
	.w7(32'h3a9fff61),
	.w8(32'h3a1b59d4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867e66a),
	.w1(32'hb9371016),
	.w2(32'hb9423b42),
	.w3(32'h396cb970),
	.w4(32'h38d7eaa5),
	.w5(32'h38a7acad),
	.w6(32'h389b4ee1),
	.w7(32'h390f44a6),
	.w8(32'h3a049220),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9788886),
	.w1(32'hba05601b),
	.w2(32'h3a88c0df),
	.w3(32'h3a633b54),
	.w4(32'h36e350ea),
	.w5(32'h3afca749),
	.w6(32'hba0018d4),
	.w7(32'hba9b4a27),
	.w8(32'h3a80239c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926465),
	.w1(32'hba5aceca),
	.w2(32'hb9fd204b),
	.w3(32'hba30b1c7),
	.w4(32'hb9526afd),
	.w5(32'h39a79619),
	.w6(32'hbab3f9e8),
	.w7(32'hba8b1ff3),
	.w8(32'hba30e833),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd968c),
	.w1(32'hbae918b3),
	.w2(32'h39a21787),
	.w3(32'hbb14397b),
	.w4(32'hbb042ea7),
	.w5(32'h39ad2d22),
	.w6(32'hbb59a17b),
	.w7(32'hbb1b59b8),
	.w8(32'h3a13286f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1ef02),
	.w1(32'h391d9353),
	.w2(32'hb81cc4f6),
	.w3(32'h3757e8d9),
	.w4(32'h39e2b74d),
	.w5(32'h396429aa),
	.w6(32'h39311516),
	.w7(32'h3a4788d1),
	.w8(32'h3a380dfd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39879725),
	.w1(32'h37ed81d3),
	.w2(32'hb8a2f494),
	.w3(32'h3a7e5e52),
	.w4(32'h398f4223),
	.w5(32'h3810ab5e),
	.w6(32'h3a43f1d0),
	.w7(32'h388950f6),
	.w8(32'hb9a292a8),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9114515),
	.w1(32'hb9106586),
	.w2(32'hb84007e5),
	.w3(32'hb71c67ea),
	.w4(32'hb92e4cb9),
	.w5(32'hb8c8d5e9),
	.w6(32'hb8dca5b4),
	.w7(32'h382147de),
	.w8(32'h375823db),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed60a7),
	.w1(32'hb9c7d856),
	.w2(32'h399911d9),
	.w3(32'hba28fc05),
	.w4(32'hb9a9f409),
	.w5(32'h39cee094),
	.w6(32'hba69d93e),
	.w7(32'hba0ec568),
	.w8(32'h38868ff1),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab83bb),
	.w1(32'h3836ba77),
	.w2(32'h39a905b0),
	.w3(32'hb9d79c55),
	.w4(32'h37557fd9),
	.w5(32'hb8465180),
	.w6(32'h39b6c74d),
	.w7(32'h39736380),
	.w8(32'hb98beb7d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a1be),
	.w1(32'hb929e0ed),
	.w2(32'h39dba897),
	.w3(32'hb77f170c),
	.w4(32'h39b8e511),
	.w5(32'h3a5aa581),
	.w6(32'hb965ff85),
	.w7(32'hba0c514e),
	.w8(32'hb9416fbe),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ef924),
	.w1(32'h39eaed93),
	.w2(32'h394e870d),
	.w3(32'h3977e337),
	.w4(32'h39ef3e31),
	.w5(32'h3953b5a8),
	.w6(32'h39d26561),
	.w7(32'h38dfaf7d),
	.w8(32'h38c22ddf),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8011be7),
	.w1(32'h39b17958),
	.w2(32'h39097240),
	.w3(32'h37985174),
	.w4(32'h39c2c5dc),
	.w5(32'h3918d14c),
	.w6(32'h39691433),
	.w7(32'h387c2146),
	.w8(32'hb94eb9c9),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983f908),
	.w1(32'hb9c4a01b),
	.w2(32'h39401066),
	.w3(32'h3a38d96d),
	.w4(32'h3a4a5572),
	.w5(32'h39b1d278),
	.w6(32'h3a01e4a6),
	.w7(32'hb948ce69),
	.w8(32'hb986bf75),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79daf9b),
	.w1(32'hbaada0ee),
	.w2(32'hba149b4b),
	.w3(32'h3b13a3ee),
	.w4(32'h3a461175),
	.w5(32'h38c29f27),
	.w6(32'h3aa03944),
	.w7(32'hba2e53f8),
	.w8(32'hba77bf3b),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e538b),
	.w1(32'h391e2cfd),
	.w2(32'hb8dc61a9),
	.w3(32'hbaa8fa2c),
	.w4(32'h395d3b4e),
	.w5(32'h3a1d364d),
	.w6(32'hb9904b56),
	.w7(32'h3814d0e3),
	.w8(32'hb969da23),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2673f),
	.w1(32'hbabd6413),
	.w2(32'hbae0187a),
	.w3(32'hbb0eebe5),
	.w4(32'hbaacfaad),
	.w5(32'hbabfa617),
	.w6(32'hba9fa863),
	.w7(32'hba83b4c5),
	.w8(32'hb9d66329),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45c9ff),
	.w1(32'hbb693788),
	.w2(32'h39cdff25),
	.w3(32'hbb90393c),
	.w4(32'hbbbd2806),
	.w5(32'hb9f6b06a),
	.w6(32'hbbb7cbfe),
	.w7(32'hbbbe1289),
	.w8(32'hbaa76c51),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf02a6),
	.w1(32'h3b73cc04),
	.w2(32'h3b43a7e6),
	.w3(32'h3bc3937e),
	.w4(32'h3bd70eeb),
	.w5(32'h3b096a33),
	.w6(32'h3bae6c59),
	.w7(32'h3b918edc),
	.w8(32'h3a35b7b2),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3875b509),
	.w1(32'h3840e04d),
	.w2(32'hb980ec7f),
	.w3(32'h39539792),
	.w4(32'h3961e634),
	.w5(32'hb9328688),
	.w6(32'h37864bbf),
	.w7(32'h38e24454),
	.w8(32'h36de1b1c),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38877e22),
	.w1(32'h3a873db0),
	.w2(32'h3a2c95fc),
	.w3(32'h3891d044),
	.w4(32'h3a64f5de),
	.w5(32'h3a38d2ae),
	.w6(32'h3a095a65),
	.w7(32'h3a0fc8d2),
	.w8(32'h39ce813d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc9c31),
	.w1(32'hb98bcfdc),
	.w2(32'hb8f35395),
	.w3(32'h39d57fdc),
	.w4(32'hb778be5e),
	.w5(32'h38af57a1),
	.w6(32'h39066767),
	.w7(32'hb82e7b29),
	.w8(32'h3923153c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3972bde4),
	.w1(32'h38407010),
	.w2(32'hb8248410),
	.w3(32'h3992bd84),
	.w4(32'h38eac2d2),
	.w5(32'hb86047bb),
	.w6(32'hb82e7ce1),
	.w7(32'hb8fc7cda),
	.w8(32'hb896ab9f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c649e1),
	.w1(32'h3a98636e),
	.w2(32'h39c32e69),
	.w3(32'h3a0625c7),
	.w4(32'h3a93b535),
	.w5(32'h391d4a86),
	.w6(32'h3a9a1871),
	.w7(32'h3a203033),
	.w8(32'hb9cc1dde),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c61f1),
	.w1(32'h3a1ae12f),
	.w2(32'hb92cf749),
	.w3(32'h3ae96e36),
	.w4(32'h3b1e0244),
	.w5(32'h3a91245d),
	.w6(32'h3a33e2ed),
	.w7(32'h3a2b62df),
	.w8(32'h399b7288),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c053e),
	.w1(32'h39e489f5),
	.w2(32'h3b2f7c27),
	.w3(32'h3b4c1f8d),
	.w4(32'h3a9d9714),
	.w5(32'h3b09ff71),
	.w6(32'h3a7aa54b),
	.w7(32'h3a0b1664),
	.w8(32'h3adebe52),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9172b),
	.w1(32'hba33f5ff),
	.w2(32'h3977046d),
	.w3(32'h3915f508),
	.w4(32'hb84c898c),
	.w5(32'h3980b694),
	.w6(32'hb7d0228a),
	.w7(32'h3908ca65),
	.w8(32'h399557f7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac8b66),
	.w1(32'hb98be2ce),
	.w2(32'h3995c00d),
	.w3(32'h3a53793c),
	.w4(32'h38c4ed8b),
	.w5(32'hb9ddb3c2),
	.w6(32'hb89f56b0),
	.w7(32'hbab9edca),
	.w8(32'hbad82352),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30a215),
	.w1(32'hba459196),
	.w2(32'hb994b970),
	.w3(32'h38e30b4f),
	.w4(32'hba107e23),
	.w5(32'hba436aa5),
	.w6(32'h389b6b33),
	.w7(32'hba3c9862),
	.w8(32'hb9feb3c6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98d3a5a),
	.w1(32'hb925d722),
	.w2(32'h37d08124),
	.w3(32'hb8b155f5),
	.w4(32'hb9015400),
	.w5(32'hb77fa27d),
	.w6(32'hb928be9a),
	.w7(32'h38129959),
	.w8(32'h39024dd8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47c628),
	.w1(32'hbacd1729),
	.w2(32'hba8e8e46),
	.w3(32'hbad20926),
	.w4(32'hbafbe347),
	.w5(32'hba3278f5),
	.w6(32'hba919a89),
	.w7(32'hba302e05),
	.w8(32'hb90c6c73),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700e2a7),
	.w1(32'hb84c8edf),
	.w2(32'hb5be9e77),
	.w3(32'h37cd7f01),
	.w4(32'hb7ff0699),
	.w5(32'h386f4d4d),
	.w6(32'hb800e916),
	.w7(32'h374187ff),
	.w8(32'hb748ee29),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdbdaa),
	.w1(32'hb9ecff15),
	.w2(32'hba5cd123),
	.w3(32'hba8882b3),
	.w4(32'hb99e6e04),
	.w5(32'hb91e196f),
	.w6(32'hba9c346a),
	.w7(32'hba32e70c),
	.w8(32'hba03e2a6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f19d7),
	.w1(32'h3b3121b3),
	.w2(32'h3af61341),
	.w3(32'h3b5421b1),
	.w4(32'h3b72d6ff),
	.w5(32'h3b01dfc3),
	.w6(32'h3b8e1f6b),
	.w7(32'h3b4b3d8c),
	.w8(32'h3a0c1bc7),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391cd159),
	.w1(32'h3a8b3ced),
	.w2(32'h3ab27053),
	.w3(32'h3adbba3b),
	.w4(32'h3b09b603),
	.w5(32'h3a870a56),
	.w6(32'h3b0ad3cf),
	.w7(32'h3a95b0b9),
	.w8(32'h39fe7cdd),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dd156d),
	.w1(32'h3963194e),
	.w2(32'hb86c6ffb),
	.w3(32'h39cf6d1c),
	.w4(32'h38b724d3),
	.w5(32'hb90a37f9),
	.w6(32'h37d10e2e),
	.w7(32'hb7655198),
	.w8(32'hb9ab50c8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acea5e1),
	.w1(32'h3b4c64da),
	.w2(32'h3b252b9c),
	.w3(32'h3b94f67e),
	.w4(32'h3b753ab7),
	.w5(32'h3abcaefc),
	.w6(32'h3b91bd4a),
	.w7(32'h3b3f9769),
	.w8(32'h3a76e5e8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b8314),
	.w1(32'hb9df5a53),
	.w2(32'h3a4bc291),
	.w3(32'hb81d2c41),
	.w4(32'hb88853d0),
	.w5(32'h3a34df35),
	.w6(32'hba0ff9f0),
	.w7(32'hb984d443),
	.w8(32'h39e919e0),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6807e0),
	.w1(32'h390c43a2),
	.w2(32'h3b16f5e1),
	.w3(32'h3a4e3bb3),
	.w4(32'h38fff53f),
	.w5(32'h3afe6e33),
	.w6(32'hb9537b2e),
	.w7(32'hba8cb3b2),
	.w8(32'h3a3359d7),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a5059),
	.w1(32'hb82b358b),
	.w2(32'hb8783cbf),
	.w3(32'h39b11d54),
	.w4(32'hb9287ff8),
	.w5(32'hb91e7760),
	.w6(32'hb867e831),
	.w7(32'hb88052cc),
	.w8(32'hb87a0a92),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fdcdd1),
	.w1(32'hb74b73a2),
	.w2(32'hb8a923a2),
	.w3(32'hb984de61),
	.w4(32'hb9226e28),
	.w5(32'h36a327cf),
	.w6(32'h3884b984),
	.w7(32'h3892110c),
	.w8(32'h373883b9),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983721a),
	.w1(32'h3a6f3700),
	.w2(32'h3a9ce1bb),
	.w3(32'h3b2a6b8a),
	.w4(32'h3a86d46d),
	.w5(32'hb8ff3808),
	.w6(32'h3a072b05),
	.w7(32'hba229cf7),
	.w8(32'hb9568d40),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13bbc6),
	.w1(32'hbbae735e),
	.w2(32'hbb4d35ef),
	.w3(32'hbb4e7411),
	.w4(32'hbb44ddb6),
	.w5(32'hba97797c),
	.w6(32'hbb428008),
	.w7(32'hbb902e38),
	.w8(32'hbb69c0cb),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d6e4c),
	.w1(32'h3a41ddbf),
	.w2(32'h3b03803d),
	.w3(32'h3b16b47d),
	.w4(32'h3af4be6c),
	.w5(32'h3ad0a345),
	.w6(32'h3ab8e4d7),
	.w7(32'hb9181baa),
	.w8(32'h3a07a73b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39958913),
	.w1(32'hb7133602),
	.w2(32'hb95320dc),
	.w3(32'hb97615d3),
	.w4(32'h361fc0f9),
	.w5(32'h3a0d4967),
	.w6(32'hba57ba97),
	.w7(32'hba532d83),
	.w8(32'hb9fb55c3),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c830cb),
	.w1(32'hb9841faf),
	.w2(32'hb867f34f),
	.w3(32'hb9b974ad),
	.w4(32'hb959229e),
	.w5(32'hb8843264),
	.w6(32'hb99f2a4c),
	.w7(32'hb8c0797f),
	.w8(32'hb8978880),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98cbb54),
	.w1(32'h385b3b0c),
	.w2(32'h3874676f),
	.w3(32'hb9c7a065),
	.w4(32'h36342d5e),
	.w5(32'h36852d9a),
	.w6(32'hb974997f),
	.w7(32'hb9564539),
	.w8(32'hb9473594),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb59c4),
	.w1(32'hba1c7082),
	.w2(32'hbab2c7f6),
	.w3(32'hba98804e),
	.w4(32'hbaf16aa2),
	.w5(32'hbac502e7),
	.w6(32'hbb03de9c),
	.w7(32'hbaea359f),
	.w8(32'hba9e7f86),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d4ccf),
	.w1(32'hbba48143),
	.w2(32'hbacdcf3d),
	.w3(32'hbbcfe953),
	.w4(32'hbbaab0be),
	.w5(32'hb8e25747),
	.w6(32'hbbecdbfc),
	.w7(32'hbba41a82),
	.w8(32'hba4dd589),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadeb9ee),
	.w1(32'hbb40ba6b),
	.w2(32'hbb70c129),
	.w3(32'hbb3b0246),
	.w4(32'hbb9df966),
	.w5(32'hbb75d9ee),
	.w6(32'hbb9cf61d),
	.w7(32'hbb95d6ef),
	.w8(32'hbb40765b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21e54e),
	.w1(32'h3aa5661a),
	.w2(32'h3a328c4d),
	.w3(32'h3b0ad2da),
	.w4(32'h3b178c5c),
	.w5(32'h3a28af3a),
	.w6(32'h3b07b938),
	.w7(32'h3ad1df9e),
	.w8(32'h3910e8b9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d5259),
	.w1(32'h3a8c911c),
	.w2(32'h3addaca4),
	.w3(32'h3af0d870),
	.w4(32'h3b1c425f),
	.w5(32'h3acfda98),
	.w6(32'h3a9f0270),
	.w7(32'h3a7e4a48),
	.w8(32'h3a0f2112),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391df172),
	.w1(32'hb795ef93),
	.w2(32'hb92dc361),
	.w3(32'h3987f062),
	.w4(32'h38f8272d),
	.w5(32'h37a2379d),
	.w6(32'h36818fdf),
	.w7(32'hb9016b2a),
	.w8(32'hb90a131e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb28b9),
	.w1(32'h38dcf9de),
	.w2(32'h398fb1ca),
	.w3(32'hb89a7f55),
	.w4(32'hb92b5988),
	.w5(32'hb887e6c1),
	.w6(32'hb858c3dd),
	.w7(32'hb89070a7),
	.w8(32'h377daa91),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9e269),
	.w1(32'h376b761f),
	.w2(32'h3a0fb201),
	.w3(32'hb8e4aeb6),
	.w4(32'hb8db9732),
	.w5(32'h39988080),
	.w6(32'hb9efbbfb),
	.w7(32'h39e40e03),
	.w8(32'hb70b8e9c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39864921),
	.w1(32'h39a8d000),
	.w2(32'h39dffc1b),
	.w3(32'h39bd98dd),
	.w4(32'h398e30f4),
	.w5(32'h39cc8594),
	.w6(32'h39df3520),
	.w7(32'h393efbf5),
	.w8(32'hb9d81952),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8baad3d),
	.w1(32'h395e8736),
	.w2(32'hb997adbb),
	.w3(32'h392696f4),
	.w4(32'h3842e58a),
	.w5(32'hba13297e),
	.w6(32'h3991d4c2),
	.w7(32'hb93112f2),
	.w8(32'hba09fe20),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c4c96),
	.w1(32'hba3c1e2f),
	.w2(32'hba3a0679),
	.w3(32'hba3d4cc3),
	.w4(32'hb94c08c9),
	.w5(32'hba3bb1c6),
	.w6(32'hba12b8d2),
	.w7(32'hb9f83759),
	.w8(32'hbae8e519),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb904b70e),
	.w1(32'h3aff1b0b),
	.w2(32'h3ab6bf0e),
	.w3(32'h3aded6c0),
	.w4(32'h3b1b460f),
	.w5(32'h3aadeff7),
	.w6(32'h3b419620),
	.w7(32'h3a8645f0),
	.w8(32'hba1a44f4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ee614),
	.w1(32'h3a07340b),
	.w2(32'h399e9d25),
	.w3(32'hb917523c),
	.w4(32'h39571285),
	.w5(32'h373b7389),
	.w6(32'h3a08bb79),
	.w7(32'hb8990f22),
	.w8(32'hb90de86c),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31383d),
	.w1(32'hbb9ab342),
	.w2(32'hbb9faa08),
	.w3(32'hbbae6001),
	.w4(32'hbbe058c9),
	.w5(32'hbb7949d1),
	.w6(32'hbbe76d38),
	.w7(32'hbbbe49bb),
	.w8(32'hbb48bf80),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95abaf8),
	.w1(32'hba72c6f8),
	.w2(32'h37a358b0),
	.w3(32'hba5af572),
	.w4(32'hbaaf9ad2),
	.w5(32'hb7901eb5),
	.w6(32'hbaf06a12),
	.w7(32'hbaa11a8d),
	.w8(32'h36efdf2c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80498b5),
	.w1(32'hb6ec29c6),
	.w2(32'h38e3f762),
	.w3(32'h38140493),
	.w4(32'h3890f9b8),
	.w5(32'h39613a60),
	.w6(32'h37b79f3c),
	.w7(32'h396ff676),
	.w8(32'h397bb719),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba907447),
	.w1(32'hbac2ef8b),
	.w2(32'hbaa16781),
	.w3(32'hbafb73b3),
	.w4(32'hbb02a669),
	.w5(32'hba562641),
	.w6(32'hbb266fc3),
	.w7(32'hbb08b030),
	.w8(32'hba6b4a1e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6ecb9),
	.w1(32'hb8105dae),
	.w2(32'hb98b242d),
	.w3(32'h395b2099),
	.w4(32'h398752ed),
	.w5(32'h38968d7a),
	.w6(32'hb907e39f),
	.w7(32'hb901f677),
	.w8(32'hb8a2a29c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f64ef8),
	.w1(32'hba014b1f),
	.w2(32'hb99b0f2a),
	.w3(32'hb9c74889),
	.w4(32'hb9b8bbbf),
	.w5(32'hb8aec99a),
	.w6(32'hba0c102d),
	.w7(32'hb93e611d),
	.w8(32'hb8b12217),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ebe15),
	.w1(32'hb6b5b744),
	.w2(32'h39215b8d),
	.w3(32'hb93fa642),
	.w4(32'h384438ee),
	.w5(32'h39566025),
	.w6(32'h37ec678d),
	.w7(32'h396e9395),
	.w8(32'h397c9353),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3924f2fe),
	.w1(32'hb92ff2ac),
	.w2(32'hb90af3b2),
	.w3(32'h394d9ee5),
	.w4(32'hb82ad231),
	.w5(32'hb8101063),
	.w6(32'hb9853678),
	.w7(32'hb945dce5),
	.w8(32'h3875d557),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86a81fe),
	.w1(32'h3a17b17c),
	.w2(32'h39e0e54b),
	.w3(32'h3a16814c),
	.w4(32'h3a7016af),
	.w5(32'h3a4d336e),
	.w6(32'h3a370dbf),
	.w7(32'h3a58daa1),
	.w8(32'h39fcab43),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9769c),
	.w1(32'h3a2a526c),
	.w2(32'h3a7f6e02),
	.w3(32'h3a43b4a3),
	.w4(32'h3a482a7a),
	.w5(32'h3ab9aefa),
	.w6(32'hba34b180),
	.w7(32'hba3a03d3),
	.w8(32'h3999dc6e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5eca3),
	.w1(32'hbad42655),
	.w2(32'h379d54b9),
	.w3(32'hba754909),
	.w4(32'hba8d1ab0),
	.w5(32'h39b6ebe2),
	.w6(32'hbaa359a7),
	.w7(32'hba4ea3b3),
	.w8(32'h399e6645),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba59d1fa),
	.w1(32'hbac1231b),
	.w2(32'hba001ce6),
	.w3(32'hbabcadc1),
	.w4(32'hbaca59f1),
	.w5(32'hb89d1240),
	.w6(32'hbaf3cd8f),
	.w7(32'hbb1290d9),
	.w8(32'hba084fa5),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8e6e4),
	.w1(32'hb79481f8),
	.w2(32'hb9b5e6d6),
	.w3(32'hb938f462),
	.w4(32'h389a07d2),
	.w5(32'hb9499ccf),
	.w6(32'hb99373d5),
	.w7(32'hb9501374),
	.w8(32'hb9ed7ae8),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aa192),
	.w1(32'h3786610c),
	.w2(32'h39847e8b),
	.w3(32'hba08db60),
	.w4(32'h37e05c60),
	.w5(32'h398c2085),
	.w6(32'hb75f7c13),
	.w7(32'h39972a2e),
	.w8(32'h399ac225),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928a47f),
	.w1(32'h371b5214),
	.w2(32'h391ba95c),
	.w3(32'h3975bfd8),
	.w4(32'h37806a2e),
	.w5(32'h3916d023),
	.w6(32'h37f0bc8b),
	.w7(32'h393316e1),
	.w8(32'h397d17dd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d7520a),
	.w1(32'h380713fd),
	.w2(32'h3910b1a8),
	.w3(32'h392e9ae7),
	.w4(32'h388ee061),
	.w5(32'h39402481),
	.w6(32'h38b64c96),
	.w7(32'h39761924),
	.w8(32'h398abfe8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b9dd4),
	.w1(32'hba0e816c),
	.w2(32'hba5ed959),
	.w3(32'hba6b158d),
	.w4(32'hba1b34be),
	.w5(32'hb9920a41),
	.w6(32'hbab6f453),
	.w7(32'hbab12f07),
	.w8(32'hba4b47fb),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07b5e7),
	.w1(32'h39154586),
	.w2(32'h38d957fa),
	.w3(32'hb991ec9c),
	.w4(32'h3971c82c),
	.w5(32'h385e7499),
	.w6(32'h396129c9),
	.w7(32'hb8ea5891),
	.w8(32'hb9d5f7cf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6db9d),
	.w1(32'h39f0f259),
	.w2(32'h39bbb014),
	.w3(32'h3a15157c),
	.w4(32'h3a4a1eb5),
	.w5(32'h39e91861),
	.w6(32'h39eb1d64),
	.w7(32'h3a05281b),
	.w8(32'h38f8fbf0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3712b8ca),
	.w1(32'h39124bc8),
	.w2(32'h37e64440),
	.w3(32'h38091dfa),
	.w4(32'h3935b6e9),
	.w5(32'h395b6017),
	.w6(32'h38e403ba),
	.w7(32'h39755365),
	.w8(32'h399e1a50),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69029d0),
	.w1(32'hb8a903a7),
	.w2(32'h3826a1ce),
	.w3(32'h3828c218),
	.w4(32'hb900a4e5),
	.w5(32'hb7866777),
	.w6(32'hb89f7460),
	.w7(32'h38d06b08),
	.w8(32'h3910ad5f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb863a12c),
	.w1(32'hb99902b4),
	.w2(32'h38f79d74),
	.w3(32'h399f14d7),
	.w4(32'hb89e6009),
	.w5(32'h39ec8c3b),
	.w6(32'h39d76fca),
	.w7(32'hb99940b9),
	.w8(32'hb92f7de6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d74602),
	.w1(32'h395fc88c),
	.w2(32'h3a281541),
	.w3(32'h39bb1dba),
	.w4(32'h386e755a),
	.w5(32'h39bf04dc),
	.w6(32'hb855ff7b),
	.w7(32'h3993ad88),
	.w8(32'h39aebc3b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa2215),
	.w1(32'hbad50853),
	.w2(32'hbafcb201),
	.w3(32'hbb2a2c58),
	.w4(32'hbaec22cd),
	.w5(32'hba17d84b),
	.w6(32'hbb83df56),
	.w7(32'hbb054b06),
	.w8(32'h38be7056),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8803691),
	.w1(32'hbb25079a),
	.w2(32'hb9b05e1c),
	.w3(32'hb73f5fb9),
	.w4(32'hbb9455d8),
	.w5(32'h3b2c3642),
	.w6(32'hbb9f49d4),
	.w7(32'h3aea6919),
	.w8(32'h3a3092e4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb710dcd),
	.w1(32'hbc6ddd77),
	.w2(32'hbb86d5b0),
	.w3(32'h3a7683c1),
	.w4(32'hbb8d2404),
	.w5(32'h3b58b19a),
	.w6(32'hbbfb1070),
	.w7(32'hbb5133ae),
	.w8(32'h3bb85282),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule