module layer_6_featuremap_32(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf9a641),
	.w1(32'hbcd10e27),
	.w2(32'hbcedbe19),
	.w3(32'hbcaffc24),
	.w4(32'hbcc792ba),
	.w5(32'hbc9f0efd),
	.w6(32'hbce6c807),
	.w7(32'hbd0c6a04),
	.w8(32'hbcc526d5),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbad24a),
	.w1(32'h3a9fd628),
	.w2(32'h38a0c6b1),
	.w3(32'h3bbb7144),
	.w4(32'h3ba996a0),
	.w5(32'h3b5521ea),
	.w6(32'h3ba572f3),
	.w7(32'h3b96e2dc),
	.w8(32'h3bae1ca8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14d8b0),
	.w1(32'hbbfa1e8d),
	.w2(32'hbb3fd0f5),
	.w3(32'hbb9f764a),
	.w4(32'hbb51db7c),
	.w5(32'hbaa1f72c),
	.w6(32'hbc2bb60d),
	.w7(32'hbad92ff2),
	.w8(32'h3b918641),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99195d),
	.w1(32'hbb09e966),
	.w2(32'h3b7610e3),
	.w3(32'hbb1a7af1),
	.w4(32'h3b6e454a),
	.w5(32'h3a380799),
	.w6(32'h3b2e1cf3),
	.w7(32'h3c390edd),
	.w8(32'h3bc9cc73),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb833099a),
	.w1(32'hbaa65964),
	.w2(32'h3b9f3387),
	.w3(32'h3c177cb0),
	.w4(32'h3c5860db),
	.w5(32'h3bf4701a),
	.w6(32'h3c18d638),
	.w7(32'h3c5098dc),
	.w8(32'h3c5dddf1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae52edf),
	.w1(32'h3b832d15),
	.w2(32'hbb6ec22f),
	.w3(32'hbad3833d),
	.w4(32'hbbac1355),
	.w5(32'hba6f42b3),
	.w6(32'hba9089ef),
	.w7(32'hbc1f150e),
	.w8(32'hbbaa1b64),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6a4f6),
	.w1(32'h3c1fb6ad),
	.w2(32'h3cb2c445),
	.w3(32'h3b539bec),
	.w4(32'h3c1c1626),
	.w5(32'h3b999449),
	.w6(32'h3c82b131),
	.w7(32'h3cf82b64),
	.w8(32'h3ca4ee66),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5438f0),
	.w1(32'h396294ab),
	.w2(32'h3b9a4772),
	.w3(32'h3a1cfd85),
	.w4(32'hbb1443e4),
	.w5(32'h398f3112),
	.w6(32'hbb14532b),
	.w7(32'h3b3f61f2),
	.w8(32'hbb132844),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94573c),
	.w1(32'h3c1b5303),
	.w2(32'h3c260f39),
	.w3(32'hbad5d1ef),
	.w4(32'h3b0ab7da),
	.w5(32'h3bb4681e),
	.w6(32'hba326ef4),
	.w7(32'h3b9f9583),
	.w8(32'h3c27b557),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ac92b),
	.w1(32'h3cbe696a),
	.w2(32'h3d222604),
	.w3(32'h3c85462d),
	.w4(32'h3cd72d8f),
	.w5(32'h3c8b88f1),
	.w6(32'h3cfa3bbb),
	.w7(32'h3d401f6a),
	.w8(32'h3d15ad59),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08b787),
	.w1(32'h38e55875),
	.w2(32'hbbbe5e69),
	.w3(32'hbac00207),
	.w4(32'hba8490dc),
	.w5(32'hbb42534a),
	.w6(32'hbbc06b54),
	.w7(32'hbb53d656),
	.w8(32'hbb33c9c9),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d7c2f),
	.w1(32'h3bc2b6d1),
	.w2(32'h3bd6c0eb),
	.w3(32'hbb127a2a),
	.w4(32'h3afd38d8),
	.w5(32'h3bde2309),
	.w6(32'hbb0099d8),
	.w7(32'hb972afe3),
	.w8(32'h3bddd49b),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c312c8b),
	.w1(32'h3b85dd5d),
	.w2(32'h3c4bf453),
	.w3(32'hb9ea6716),
	.w4(32'h3b9fd028),
	.w5(32'hbb14aa9f),
	.w6(32'h3adb129f),
	.w7(32'h3c1707be),
	.w8(32'hba35ba2e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc25b0),
	.w1(32'hbb481c3e),
	.w2(32'hbb8f11a3),
	.w3(32'hbba5bb84),
	.w4(32'hbba1164c),
	.w5(32'hbb361f73),
	.w6(32'hbb1250fe),
	.w7(32'hbab51e9f),
	.w8(32'hbbdeb8f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b7161),
	.w1(32'h3c393b5a),
	.w2(32'h3c471a99),
	.w3(32'h3c35de19),
	.w4(32'h3c5ca9f6),
	.w5(32'h3c46f8de),
	.w6(32'h3c5dde00),
	.w7(32'h3c5d2149),
	.w8(32'h3c6c227d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f917a),
	.w1(32'h3b02f397),
	.w2(32'h3a889b09),
	.w3(32'h39a2b6fa),
	.w4(32'h3a80420c),
	.w5(32'h3a15b5a3),
	.w6(32'h3b843a90),
	.w7(32'h3b6df0c7),
	.w8(32'h3b3ac599),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b8d23),
	.w1(32'hbb0fe9e7),
	.w2(32'hbb8686f1),
	.w3(32'hbb95591a),
	.w4(32'hbb38034c),
	.w5(32'hbabf32ba),
	.w6(32'hbba03c2a),
	.w7(32'hbc18988c),
	.w8(32'hbc0b80cc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1dd8d4),
	.w1(32'h3cf7b9e1),
	.w2(32'h3d1336a8),
	.w3(32'h3d050861),
	.w4(32'h3d1cad1d),
	.w5(32'h3cfaa127),
	.w6(32'h3d201adc),
	.w7(32'h3d393c2b),
	.w8(32'h3d15a696),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdcf631),
	.w1(32'hb9e15c7b),
	.w2(32'h3b69585d),
	.w3(32'h3b3acb0e),
	.w4(32'h3bbf3708),
	.w5(32'hbb0e8196),
	.w6(32'h3c2a72d8),
	.w7(32'h3c88ff6a),
	.w8(32'h3bb48b53),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8869e2),
	.w1(32'h3a80ea51),
	.w2(32'h3a105a7a),
	.w3(32'h3b61db5c),
	.w4(32'h3bd95bff),
	.w5(32'h3afc5ade),
	.w6(32'h396f3566),
	.w7(32'h3be207b8),
	.w8(32'h3a654a33),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d8e53),
	.w1(32'h3b6c5589),
	.w2(32'h3b142a55),
	.w3(32'h3b6c3493),
	.w4(32'h3ab057e9),
	.w5(32'h3b937e73),
	.w6(32'h3b5b5147),
	.w7(32'h3b3d49d7),
	.w8(32'h3b17e898),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19a156),
	.w1(32'h3cceb73f),
	.w2(32'h3ccd237f),
	.w3(32'h3cbca19c),
	.w4(32'h3cef8157),
	.w5(32'h3cb711f5),
	.w6(32'h3ced0769),
	.w7(32'h3cf6202c),
	.w8(32'h3ccb37e8),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca758c6),
	.w1(32'h3ad51088),
	.w2(32'h3b25c5a6),
	.w3(32'h3b11bc8e),
	.w4(32'hba0dddf9),
	.w5(32'hbb255be4),
	.w6(32'h3bd671e1),
	.w7(32'h3b63dc70),
	.w8(32'h3b91c57e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc29e8a),
	.w1(32'hbb5a62cc),
	.w2(32'h3b153540),
	.w3(32'hbb7fb2df),
	.w4(32'hbb089954),
	.w5(32'hba3c1124),
	.w6(32'h3b9adee3),
	.w7(32'h3b51b334),
	.w8(32'h3afe43c7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1235ad),
	.w1(32'hb922d95e),
	.w2(32'h39fe347d),
	.w3(32'h3a6dee29),
	.w4(32'hb9b6254e),
	.w5(32'hb98184e2),
	.w6(32'hbb05fad0),
	.w7(32'h3a533730),
	.w8(32'h398bf09d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07b202),
	.w1(32'hbb9f0c9d),
	.w2(32'hbb517128),
	.w3(32'hbb66b476),
	.w4(32'hba8b9b12),
	.w5(32'h3b6e482c),
	.w6(32'hbad83861),
	.w7(32'hbbcd63f2),
	.w8(32'h3a879f79),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a794e27),
	.w1(32'h3bf04b6d),
	.w2(32'h3c872319),
	.w3(32'h3b9e60d8),
	.w4(32'h3c2d8a4f),
	.w5(32'h3bbec5f9),
	.w6(32'h3c60c725),
	.w7(32'h3d03e72d),
	.w8(32'h3c9fe0e2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6781df),
	.w1(32'h3c3d02c1),
	.w2(32'h3c8dcf84),
	.w3(32'h3c340500),
	.w4(32'h3c372d61),
	.w5(32'h3c11f44e),
	.w6(32'h3c8bfd0b),
	.w7(32'h3cb37883),
	.w8(32'h3c8bac48),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5738b6),
	.w1(32'hbbae767c),
	.w2(32'hbc36f47c),
	.w3(32'hbb85401d),
	.w4(32'hbc04860c),
	.w5(32'hbbcae393),
	.w6(32'hbc0821f9),
	.w7(32'hbc71c766),
	.w8(32'hbc531825),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc204fe1),
	.w1(32'hba7e6e2a),
	.w2(32'hbb9a797b),
	.w3(32'hbb83ea09),
	.w4(32'hbb8977e3),
	.w5(32'hbb70d7a2),
	.w6(32'hbb5305fe),
	.w7(32'hbb4d4f85),
	.w8(32'hbba94a46),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b705c),
	.w1(32'hba88e795),
	.w2(32'h3bfe82bf),
	.w3(32'h3b830cab),
	.w4(32'h3b952278),
	.w5(32'hb9ebc480),
	.w6(32'h3aae544a),
	.w7(32'h3ba828f7),
	.w8(32'h3b9a7b28),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cec5c),
	.w1(32'h3b0c1daf),
	.w2(32'h3b163995),
	.w3(32'h3b9458b8),
	.w4(32'h3bae206a),
	.w5(32'h3b418a08),
	.w6(32'h3b6574cd),
	.w7(32'h3b877ef6),
	.w8(32'h3b121273),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd56627),
	.w1(32'h3b166b7e),
	.w2(32'hb9e78e65),
	.w3(32'hbb623c11),
	.w4(32'hb97a3590),
	.w5(32'hb98e61ba),
	.w6(32'hba288d92),
	.w7(32'h3b6e07a6),
	.w8(32'h3b625df1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c6dca),
	.w1(32'hbb191adf),
	.w2(32'hbbaaea1e),
	.w3(32'h38d5d25c),
	.w4(32'hbb3ae9ec),
	.w5(32'hbb7059b6),
	.w6(32'hbafe281c),
	.w7(32'hbbf7775c),
	.w8(32'hbb5baf77),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c5a1),
	.w1(32'h3c294e70),
	.w2(32'h3c2d87f0),
	.w3(32'h3b8176e1),
	.w4(32'h3b87edd0),
	.w5(32'h3ba43371),
	.w6(32'h3c0f6dab),
	.w7(32'h3c1b5439),
	.w8(32'h3c2a42da),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c310e0f),
	.w1(32'h3bd5fa31),
	.w2(32'h3c16d574),
	.w3(32'h3a92ff9e),
	.w4(32'h3b49fe08),
	.w5(32'h3b854a3f),
	.w6(32'h3bf16056),
	.w7(32'h3c1cbe21),
	.w8(32'h3b28d8b5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5266cd),
	.w1(32'h3cc8cd04),
	.w2(32'h3d0e84eb),
	.w3(32'h3c8ab4c9),
	.w4(32'h3cb72f41),
	.w5(32'h3c74f2c6),
	.w6(32'h3ce12b11),
	.w7(32'h3d0f053f),
	.w8(32'h3d09a4b4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce40563),
	.w1(32'h3b4b8039),
	.w2(32'h3bac4583),
	.w3(32'hba9fe6fd),
	.w4(32'hb928e648),
	.w5(32'hb9ac0d68),
	.w6(32'h3b483214),
	.w7(32'h3b9de8ac),
	.w8(32'h3b7c6112),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b3a06),
	.w1(32'h3b75f8b3),
	.w2(32'hba160c34),
	.w3(32'h3b491d09),
	.w4(32'h3b421cc9),
	.w5(32'h3ab3b2b8),
	.w6(32'hb8e2bd3d),
	.w7(32'hba8a68f6),
	.w8(32'h3afce152),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d9737),
	.w1(32'h3a5b91b5),
	.w2(32'h3bddeffe),
	.w3(32'hbbb107d4),
	.w4(32'h3988995c),
	.w5(32'h3aff3ad5),
	.w6(32'h3b4f972a),
	.w7(32'h3c20d556),
	.w8(32'h3c1c1c76),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11d3cc),
	.w1(32'hbb73971d),
	.w2(32'hba30f033),
	.w3(32'h3aa2712c),
	.w4(32'h3c16c041),
	.w5(32'hb9100987),
	.w6(32'h3ba5898a),
	.w7(32'h3b861528),
	.w8(32'h3bcd1f11),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab06582),
	.w1(32'h3bb17771),
	.w2(32'h3c383450),
	.w3(32'h3ad6be16),
	.w4(32'h3bbb55c3),
	.w5(32'h3bba231c),
	.w6(32'h3beaef5f),
	.w7(32'h3c575c29),
	.w8(32'h3c37881e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f72fc),
	.w1(32'h3bfde0e6),
	.w2(32'h3c7bf2aa),
	.w3(32'h3b1dbbaf),
	.w4(32'h3bb6a315),
	.w5(32'h3b4c4e2b),
	.w6(32'h3bc1417d),
	.w7(32'h3c33bdfe),
	.w8(32'h3c157cff),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c560c19),
	.w1(32'hbaef4b60),
	.w2(32'hbb141d12),
	.w3(32'hba31980b),
	.w4(32'hbaeac145),
	.w5(32'h3ae709d1),
	.w6(32'hb9f5b8f4),
	.w7(32'h3b2957fa),
	.w8(32'hb9b7d3ec),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb764520),
	.w1(32'hbb72d7ef),
	.w2(32'hbc044297),
	.w3(32'hbb424f5f),
	.w4(32'hbba42f99),
	.w5(32'hbb610dfc),
	.w6(32'hbbe392e4),
	.w7(32'hbc21d86b),
	.w8(32'hbbf5deaa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadaa9b),
	.w1(32'hbc2e1abc),
	.w2(32'hbc87325e),
	.w3(32'hbbe9aa31),
	.w4(32'hbc0cc41a),
	.w5(32'hbc293201),
	.w6(32'hbbe3738d),
	.w7(32'hbc45dbb5),
	.w8(32'hbc6333b8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12c62c),
	.w1(32'hbb58f2b8),
	.w2(32'hbb3b2564),
	.w3(32'h3ad1a34b),
	.w4(32'hb9c565ff),
	.w5(32'hbb30d73c),
	.w6(32'hbad09a4d),
	.w7(32'h3a9c2175),
	.w8(32'hba13ba4c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d3d74),
	.w1(32'hbaf98561),
	.w2(32'hbb006e6a),
	.w3(32'hbb45d783),
	.w4(32'hbad1216e),
	.w5(32'h3b94a7bd),
	.w6(32'h39ffeae6),
	.w7(32'hbb4d6182),
	.w8(32'h3a0b5389),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cf422),
	.w1(32'hbc3a7638),
	.w2(32'hbccaa295),
	.w3(32'hbbfb3024),
	.w4(32'hbc7362f8),
	.w5(32'hbbe7e4c1),
	.w6(32'hbc939582),
	.w7(32'hbd0053da),
	.w8(32'hbcb7ad79),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93bda6),
	.w1(32'h3c4e9d47),
	.w2(32'h3c338dfe),
	.w3(32'h3c4229b9),
	.w4(32'h3c738212),
	.w5(32'h3bc5b796),
	.w6(32'h3c9f4fdc),
	.w7(32'h3c908ae6),
	.w8(32'h3c38e6dc),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb2801),
	.w1(32'h3bfe890e),
	.w2(32'h3bf6dba8),
	.w3(32'h3b0e80ce),
	.w4(32'h3ade601e),
	.w5(32'h3b94bcb6),
	.w6(32'h3be73d0a),
	.w7(32'h3c1d3fbb),
	.w8(32'h3c0ef62d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffb708),
	.w1(32'h3c0ba5bf),
	.w2(32'h3c4a83e6),
	.w3(32'h3c04eb11),
	.w4(32'h3c19103f),
	.w5(32'h3bee0e85),
	.w6(32'h3c23a290),
	.w7(32'h3c384ffc),
	.w8(32'h3c2d5427),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c166718),
	.w1(32'hbb6406e7),
	.w2(32'hbc9c6854),
	.w3(32'h3b20311d),
	.w4(32'hbbdc2602),
	.w5(32'h3b3a45ed),
	.w6(32'hbbb6ca51),
	.w7(32'hbc99294f),
	.w8(32'hbc212eef),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc450aeb),
	.w1(32'hbd8dc584),
	.w2(32'hbdd43827),
	.w3(32'hbd836b71),
	.w4(32'hbdb5dc0f),
	.w5(32'hbd78df26),
	.w6(32'hbdc3b3a1),
	.w7(32'hbe0827ba),
	.w8(32'hbdccc722),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda4fb88),
	.w1(32'h3c2bbf02),
	.w2(32'h3c02c3c3),
	.w3(32'h3c204877),
	.w4(32'h3c06d854),
	.w5(32'h3c0d745a),
	.w6(32'h3c2c22bc),
	.w7(32'h3c47b09b),
	.w8(32'h3c071c24),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc5f7a),
	.w1(32'h3c4b3177),
	.w2(32'h3c8971e9),
	.w3(32'h3b06fe06),
	.w4(32'hbae4cc85),
	.w5(32'hbc1a70f5),
	.w6(32'h3b907358),
	.w7(32'hbb188410),
	.w8(32'hbb2929cf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51cecb),
	.w1(32'hbc06837f),
	.w2(32'hbbb08204),
	.w3(32'hbbb88906),
	.w4(32'h3a68868a),
	.w5(32'hba65e400),
	.w6(32'hba74134a),
	.w7(32'h3bc06f5f),
	.w8(32'h3b9af689),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41df47),
	.w1(32'hbb04796a),
	.w2(32'h3c193fb6),
	.w3(32'h3c1f10a7),
	.w4(32'h3bf4826a),
	.w5(32'h3c20b173),
	.w6(32'h3b84ab3e),
	.w7(32'hbc23e767),
	.w8(32'hbacae5ad),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b067864),
	.w1(32'h3bb82bb0),
	.w2(32'h3b38a4fa),
	.w3(32'h3b15f2d9),
	.w4(32'hbb27569f),
	.w5(32'hbb63ca58),
	.w6(32'h3a8913db),
	.w7(32'hbb145418),
	.w8(32'hbb879c60),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ad709),
	.w1(32'hbc1dba46),
	.w2(32'hbbf93de5),
	.w3(32'h3ba2934e),
	.w4(32'h3bfc6a41),
	.w5(32'h3b44f173),
	.w6(32'hbc064fcf),
	.w7(32'h3c532ea4),
	.w8(32'h3c974c35),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc88bf3),
	.w1(32'hbb4635c1),
	.w2(32'hba712391),
	.w3(32'hba58e7df),
	.w4(32'hbbe30285),
	.w5(32'hbc123c4f),
	.w6(32'hbb3c88e6),
	.w7(32'hbc171d28),
	.w8(32'hbc21c2a7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb121c66),
	.w1(32'hbb86205b),
	.w2(32'h3b56f5ec),
	.w3(32'hbb98ee7c),
	.w4(32'h3c1d521d),
	.w5(32'hbb75b821),
	.w6(32'hba5da7b7),
	.w7(32'h3aa848c0),
	.w8(32'hbba57b8a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4df1a),
	.w1(32'h3bd33ae3),
	.w2(32'hbbfe1624),
	.w3(32'h3c242f2d),
	.w4(32'h3cebe938),
	.w5(32'h3cd27b2b),
	.w6(32'hba7b042d),
	.w7(32'h3cc8d789),
	.w8(32'h3d0d859c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4214aa),
	.w1(32'h3c3311c8),
	.w2(32'h3c7b99af),
	.w3(32'hbb2b1a67),
	.w4(32'hbbe8e328),
	.w5(32'hbbbbdd30),
	.w6(32'h3a30129c),
	.w7(32'hbb2807c3),
	.w8(32'hbbaab3cc),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule