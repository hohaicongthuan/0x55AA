module layer_10_featuremap_263(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef49a9),
	.w1(32'hbc1666f5),
	.w2(32'hbc48a67b),
	.w3(32'hbb8b942b),
	.w4(32'hbc7730dc),
	.w5(32'h3aa4b27d),
	.w6(32'hbba50621),
	.w7(32'hbc1ffecb),
	.w8(32'hbba48a62),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bdcc4),
	.w1(32'hbbdce53e),
	.w2(32'hbb30d0bc),
	.w3(32'h3b076b5f),
	.w4(32'hba04fffc),
	.w5(32'hbb40a0d5),
	.w6(32'h3a8dfe1c),
	.w7(32'hbaa58b23),
	.w8(32'hbbe36567),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc1099),
	.w1(32'h3c1075d0),
	.w2(32'h3be96066),
	.w3(32'hbb684162),
	.w4(32'h3ab8c40f),
	.w5(32'h3b4a39ae),
	.w6(32'h3b4a85b4),
	.w7(32'h3b729a5a),
	.w8(32'h3a258b89),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76ad37),
	.w1(32'h3b7af8f1),
	.w2(32'h3b8a9b99),
	.w3(32'h3a78f0b4),
	.w4(32'h3b866b0a),
	.w5(32'hbace5fa0),
	.w6(32'h3abdee33),
	.w7(32'h3b37b390),
	.w8(32'hbb7440f3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb464741),
	.w1(32'hb9d562a4),
	.w2(32'hbbaa513f),
	.w3(32'hbb6e87a4),
	.w4(32'hbc1e81e4),
	.w5(32'h3b651c70),
	.w6(32'hbbf2f1fb),
	.w7(32'hbc58605e),
	.w8(32'h3a0f987b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae05300),
	.w1(32'h3a89864e),
	.w2(32'h3a775f00),
	.w3(32'h3acb36af),
	.w4(32'hb9fa5719),
	.w5(32'hb86e6bf4),
	.w6(32'h3b4f50e1),
	.w7(32'h3b522656),
	.w8(32'hbae5ba02),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba37996),
	.w1(32'h3c20cda1),
	.w2(32'h3b87cad0),
	.w3(32'h3c1c4252),
	.w4(32'h3b7ecdda),
	.w5(32'hbc3f6a86),
	.w6(32'h3b19b70d),
	.w7(32'h3c0df9fc),
	.w8(32'hbc0300b9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2d53a),
	.w1(32'hbc239479),
	.w2(32'hbc48d35d),
	.w3(32'hbc908573),
	.w4(32'hbca8d158),
	.w5(32'hbbef5384),
	.w6(32'hbb0fadd1),
	.w7(32'hbb02c967),
	.w8(32'hbc04eb38),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7a00c),
	.w1(32'hbba92dfb),
	.w2(32'hbb8552b2),
	.w3(32'hbaa36c9d),
	.w4(32'hbb2a10fb),
	.w5(32'h3b8eced0),
	.w6(32'hbba98e76),
	.w7(32'hbab8b4dc),
	.w8(32'h3b0b740b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba886137),
	.w1(32'h3b309db5),
	.w2(32'hbb576769),
	.w3(32'hbb680732),
	.w4(32'hbacb196d),
	.w5(32'hb9aebefa),
	.w6(32'hbb02b667),
	.w7(32'h399d43f2),
	.w8(32'hbba38f65),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab634e),
	.w1(32'h3b7d6546),
	.w2(32'hb933bf4f),
	.w3(32'hba88e984),
	.w4(32'hbae9a68c),
	.w5(32'hbba4f421),
	.w6(32'h3b0a989e),
	.w7(32'h3b839e03),
	.w8(32'hbb576f54),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b240b61),
	.w1(32'h3cc9116b),
	.w2(32'h3c1691a5),
	.w3(32'h3b62028f),
	.w4(32'h3a54577c),
	.w5(32'hbbaed968),
	.w6(32'hbb9a70b5),
	.w7(32'h3c5de9c0),
	.w8(32'h3b53cd47),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99a478),
	.w1(32'h3bcc34e7),
	.w2(32'h3b810bce),
	.w3(32'hbc92f531),
	.w4(32'hbb6a3a20),
	.w5(32'hbb48a6ab),
	.w6(32'h3b2acf18),
	.w7(32'h3b5def16),
	.w8(32'hbaebc9bd),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f883da),
	.w1(32'hbc29ada4),
	.w2(32'hbc6a33fc),
	.w3(32'hbb54035b),
	.w4(32'hbbd12fb9),
	.w5(32'hbaba9ed9),
	.w6(32'h3a480137),
	.w7(32'hbb479a05),
	.w8(32'hbbb77618),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba207c03),
	.w1(32'hbb0450cd),
	.w2(32'h3ac37380),
	.w3(32'h3b049d35),
	.w4(32'h3b41901e),
	.w5(32'h391aef23),
	.w6(32'h3abcdc54),
	.w7(32'h3bb4dcf2),
	.w8(32'h3ad28f5a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af63e76),
	.w1(32'hbc188e3f),
	.w2(32'hbc5d96f0),
	.w3(32'hbab57b97),
	.w4(32'hbb2e98d4),
	.w5(32'hbbc5a2ed),
	.w6(32'hbc9709cc),
	.w7(32'hbb623dca),
	.w8(32'hbbe7504f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce9364),
	.w1(32'hbafbb904),
	.w2(32'hbb0137e9),
	.w3(32'hba92e8c0),
	.w4(32'hbb192cd8),
	.w5(32'hbaf64fe8),
	.w6(32'h393e2416),
	.w7(32'h39cc84a2),
	.w8(32'hbb1d6fc7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd6f7a),
	.w1(32'h3c469381),
	.w2(32'h3bf26ccd),
	.w3(32'hbbf06824),
	.w4(32'hbaffbe86),
	.w5(32'hbbe4ca4e),
	.w6(32'h3bf421ec),
	.w7(32'h3c1a180b),
	.w8(32'h3a9a7416),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102109),
	.w1(32'h3be2baf6),
	.w2(32'h3b3d7900),
	.w3(32'hbc0e9f00),
	.w4(32'hbb1ecfe3),
	.w5(32'hbbcdaec0),
	.w6(32'hba05938e),
	.w7(32'h3ba4cff9),
	.w8(32'h3b1afe29),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49fba0),
	.w1(32'hbb691008),
	.w2(32'hbb69355f),
	.w3(32'h3ad4c113),
	.w4(32'h3b958370),
	.w5(32'h3bd9d362),
	.w6(32'hbaadd067),
	.w7(32'h3b112c42),
	.w8(32'h3c72a246),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a2570),
	.w1(32'hbba8cf8d),
	.w2(32'h398724a3),
	.w3(32'hbc0b8156),
	.w4(32'h3c221fe7),
	.w5(32'h3a35d8b8),
	.w6(32'hbc477bc6),
	.w7(32'h3bc07c20),
	.w8(32'hbb4ca43f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe9cda),
	.w1(32'hbba400c5),
	.w2(32'hbaa7b191),
	.w3(32'hba2b4172),
	.w4(32'h3b28d5c9),
	.w5(32'h39dc470e),
	.w6(32'hbb7d9599),
	.w7(32'h3b111186),
	.w8(32'hb8a201ee),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23432a),
	.w1(32'h3bd7e578),
	.w2(32'hbc6a60ac),
	.w3(32'hbc03e5e0),
	.w4(32'hbc1cc2fd),
	.w5(32'hbc1a361e),
	.w6(32'hbc1a6d2d),
	.w7(32'h3b13dd72),
	.w8(32'hbb0930de),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93f98d),
	.w1(32'hbc38e485),
	.w2(32'hbba21f46),
	.w3(32'hbc3fe3d9),
	.w4(32'hbbb39fe4),
	.w5(32'hba6f5acd),
	.w6(32'hbc9de195),
	.w7(32'h3b98ff0c),
	.w8(32'hbbaf43e5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc564d2b),
	.w1(32'hbc23158f),
	.w2(32'hbab263d8),
	.w3(32'hbbdcbd70),
	.w4(32'hbc06fb67),
	.w5(32'h3b3115c9),
	.w6(32'hbc3cf4f2),
	.w7(32'hbc4ffc64),
	.w8(32'hbb2a53a2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a822b),
	.w1(32'h3956d295),
	.w2(32'hba0ffd41),
	.w3(32'h3bceb25b),
	.w4(32'h3a94fe07),
	.w5(32'hbb958049),
	.w6(32'h3b47385d),
	.w7(32'h3b0ef187),
	.w8(32'hbbe6f269),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb15ce0),
	.w1(32'hbb5619f0),
	.w2(32'hbacec9f2),
	.w3(32'hbadb9c55),
	.w4(32'hb7ee90d7),
	.w5(32'hbbc54a5d),
	.w6(32'hbb965e78),
	.w7(32'hbb22f834),
	.w8(32'hbb871788),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9aac65),
	.w1(32'h3b80d4c1),
	.w2(32'hbbbbdfbd),
	.w3(32'hbc2fcee6),
	.w4(32'h3b84ecae),
	.w5(32'h3b6c1961),
	.w6(32'hbc4eeda0),
	.w7(32'hb9aeb875),
	.w8(32'hbb61e23e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5d383),
	.w1(32'hbb19e57d),
	.w2(32'hbba73366),
	.w3(32'h3bc5c3a0),
	.w4(32'h39f97a92),
	.w5(32'hbb839df5),
	.w6(32'h3b417fe8),
	.w7(32'h3b080582),
	.w8(32'hbbba251a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc838aeb),
	.w1(32'h3b93c84b),
	.w2(32'hbba1ee2a),
	.w3(32'h3c1f9f44),
	.w4(32'h3bba5bdb),
	.w5(32'hbc0d4c23),
	.w6(32'h3bad1107),
	.w7(32'hbb6caccd),
	.w8(32'hbc01de67),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14e9b5),
	.w1(32'hba20b398),
	.w2(32'h3b01edd6),
	.w3(32'hbb96b751),
	.w4(32'hbbd1b524),
	.w5(32'hbb0970fc),
	.w6(32'hbb4a8dac),
	.w7(32'hba9d5693),
	.w8(32'h3bac9dd5),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a295c),
	.w1(32'h3b0b2560),
	.w2(32'hba6379fb),
	.w3(32'hbb8c2ca1),
	.w4(32'hbbbb6b4e),
	.w5(32'hbbab5c85),
	.w6(32'hbb8180bc),
	.w7(32'h3a214dee),
	.w8(32'hba068cb6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92251e),
	.w1(32'h3b64b5fc),
	.w2(32'h3b883077),
	.w3(32'h3b1fb4c9),
	.w4(32'h3b84f988),
	.w5(32'hba6ee92a),
	.w6(32'h3be0917c),
	.w7(32'h3bd7aed1),
	.w8(32'hbb1d9a48),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad904ac),
	.w1(32'h3be6eebe),
	.w2(32'h3b92da82),
	.w3(32'hbab1c3ac),
	.w4(32'h3b0116dc),
	.w5(32'h3a8b5e4a),
	.w6(32'h3b5cd928),
	.w7(32'h3c6b3990),
	.w8(32'hb8a4f463),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5b8c6),
	.w1(32'hbad41188),
	.w2(32'h388ee7b4),
	.w3(32'h3aa5fec1),
	.w4(32'hbafc8c06),
	.w5(32'h3bbe90e6),
	.w6(32'h3b35c906),
	.w7(32'h3b27b0fa),
	.w8(32'h3bb378ca),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13cbb7),
	.w1(32'hbb0f64ca),
	.w2(32'h3b6d3cb0),
	.w3(32'hbc244ec7),
	.w4(32'hbbade116),
	.w5(32'hbc0030cf),
	.w6(32'hbc00e03b),
	.w7(32'h3b424f4c),
	.w8(32'h3b9752a0),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb05bc8),
	.w1(32'hbade219c),
	.w2(32'hbc6b7bce),
	.w3(32'hbc31aa78),
	.w4(32'h3997f414),
	.w5(32'hbc3d699a),
	.w6(32'hbc8af0fb),
	.w7(32'hbc967f95),
	.w8(32'hbc562e34),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc56eb3a),
	.w1(32'hbad9ce15),
	.w2(32'h3ad042f4),
	.w3(32'h3aa793b2),
	.w4(32'h3be246f6),
	.w5(32'h3c690cb2),
	.w6(32'hbb7393ac),
	.w7(32'h3b99db8e),
	.w8(32'h3a1275f6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc776906),
	.w1(32'hbc25e0f0),
	.w2(32'hb9d78326),
	.w3(32'hbb239398),
	.w4(32'hba2570b3),
	.w5(32'h3bff0f7b),
	.w6(32'hbb5adae9),
	.w7(32'hbb43a0d7),
	.w8(32'h3b66a3fc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a689370),
	.w1(32'hbc2bbd0f),
	.w2(32'h3b26be55),
	.w3(32'hbb4de579),
	.w4(32'h3c1ae87e),
	.w5(32'hbbb61fbe),
	.w6(32'hbc21f6ab),
	.w7(32'h3be101a3),
	.w8(32'hbbd1d26b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6ad17),
	.w1(32'h3b9a580f),
	.w2(32'hb96c4ac2),
	.w3(32'hbb32840b),
	.w4(32'hbafda2f7),
	.w5(32'h3bd2776a),
	.w6(32'h3bea0fb2),
	.w7(32'h3be74bc7),
	.w8(32'h3b68a82a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0ebc0),
	.w1(32'h3af6d857),
	.w2(32'h3a494548),
	.w3(32'h3bddd242),
	.w4(32'h3ac4102f),
	.w5(32'hbb8f7ad0),
	.w6(32'h3b91872b),
	.w7(32'h3b0b41e2),
	.w8(32'hbae10c07),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b5ad9),
	.w1(32'hbb8cbb34),
	.w2(32'hbaf45032),
	.w3(32'hb90ba4de),
	.w4(32'hbb8bd4d7),
	.w5(32'h3b89a8b8),
	.w6(32'hbba86742),
	.w7(32'hbb0938d1),
	.w8(32'hbc0263a2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfb12e),
	.w1(32'h3af174d6),
	.w2(32'hbb9d2057),
	.w3(32'hbb2e47f2),
	.w4(32'hbb2ef708),
	.w5(32'hbbc727ec),
	.w6(32'hbb72789a),
	.w7(32'h3a6e78b5),
	.w8(32'hba9f4316),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5bbb39),
	.w1(32'hbb1820fe),
	.w2(32'hbc13a501),
	.w3(32'hbc073995),
	.w4(32'h3ad7e34e),
	.w5(32'h3ba68ea6),
	.w6(32'hbbb32189),
	.w7(32'hba95b643),
	.w8(32'h3b1742dd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ce9df),
	.w1(32'h3adea43c),
	.w2(32'hbb7cee87),
	.w3(32'hbc0e144e),
	.w4(32'hbbda9b0d),
	.w5(32'hbb8d4c48),
	.w6(32'h3ab69310),
	.w7(32'h3b97c858),
	.w8(32'hba8d2dac),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb744a7c),
	.w1(32'h399a2ebe),
	.w2(32'hb98e28fb),
	.w3(32'hbb902eca),
	.w4(32'h3bc2441b),
	.w5(32'h3b463faa),
	.w6(32'hb9ea6792),
	.w7(32'h3b8122a6),
	.w8(32'hbaee138b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf98ad),
	.w1(32'h3b7a433f),
	.w2(32'hbb27c466),
	.w3(32'hbbfefb88),
	.w4(32'hbc0725c2),
	.w5(32'hbc3bf9fe),
	.w6(32'hba8b59bc),
	.w7(32'hbb11c33c),
	.w8(32'hbc1fd52c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96ab14),
	.w1(32'hb9ee86ea),
	.w2(32'hbb9d9b8d),
	.w3(32'hbb84cef1),
	.w4(32'hbb878867),
	.w5(32'h3b458df8),
	.w6(32'hb98c7047),
	.w7(32'hbaeed8f0),
	.w8(32'hbb108201),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1423e4),
	.w1(32'hbba3240b),
	.w2(32'hba59cad3),
	.w3(32'h3b1be8ea),
	.w4(32'h3b8f2454),
	.w5(32'hbbdacf51),
	.w6(32'hbb66c35b),
	.w7(32'h3b34992c),
	.w8(32'hbbe0b5b5),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcca743),
	.w1(32'hbb08759e),
	.w2(32'h3b873418),
	.w3(32'hbb9ba435),
	.w4(32'hbb401d3b),
	.w5(32'hbb816081),
	.w6(32'hbba90f94),
	.w7(32'hb8573f73),
	.w8(32'h3a5a8c89),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4e300),
	.w1(32'hbb80fa6e),
	.w2(32'hbb591ec9),
	.w3(32'hbb68c040),
	.w4(32'hbbd47185),
	.w5(32'hbb9d5b07),
	.w6(32'hbbab8b2c),
	.w7(32'hb9a2480b),
	.w8(32'hbc13f85d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b9c5b),
	.w1(32'h3b9e27fc),
	.w2(32'h3b9a5d45),
	.w3(32'hbba107f9),
	.w4(32'hbbe09f1b),
	.w5(32'hbb688f91),
	.w6(32'h3b4ba300),
	.w7(32'h3c218614),
	.w8(32'hbb685543),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6458b),
	.w1(32'h3c3722d9),
	.w2(32'h39ba0774),
	.w3(32'h3b52bcb2),
	.w4(32'h3b84ad56),
	.w5(32'hbbc2d6fd),
	.w6(32'hba1c4adc),
	.w7(32'h3c490842),
	.w8(32'h3abebcf8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70b7e3),
	.w1(32'hbae886a0),
	.w2(32'hbb9c4b7c),
	.w3(32'hbbdfeb3b),
	.w4(32'hb93672ae),
	.w5(32'h3b2a99ed),
	.w6(32'hbb3d27ae),
	.w7(32'hbaad0217),
	.w8(32'hbaebf6b3),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895787e),
	.w1(32'hbb3210ef),
	.w2(32'hbab2fb49),
	.w3(32'h3bca2114),
	.w4(32'h3a4b3f36),
	.w5(32'hbb4a3de8),
	.w6(32'h3c02b376),
	.w7(32'h3b3fd4b1),
	.w8(32'hbaf81cfe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb441827),
	.w1(32'hbb6e922c),
	.w2(32'hbbdfe555),
	.w3(32'h38a99f93),
	.w4(32'hbb1f2f6e),
	.w5(32'hbba61f9a),
	.w6(32'h3b17e5b9),
	.w7(32'hbaa2e215),
	.w8(32'hbbb73ab7),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0968d8),
	.w1(32'h3b69755a),
	.w2(32'hbb98087a),
	.w3(32'hbac01fec),
	.w4(32'hbaa2781c),
	.w5(32'h3b045c41),
	.w6(32'h39a49ffc),
	.w7(32'h3ae379d1),
	.w8(32'hbae424ef),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57ce25),
	.w1(32'hbb8fd942),
	.w2(32'h3a39b966),
	.w3(32'h3b44f59f),
	.w4(32'h3ba0ffd0),
	.w5(32'hb8ded547),
	.w6(32'hbbf357d0),
	.w7(32'h3b638d50),
	.w8(32'hbb8019cf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd447a6),
	.w1(32'hbbd09d35),
	.w2(32'hbbf77c28),
	.w3(32'hbb479a92),
	.w4(32'hbc138f40),
	.w5(32'h3975e317),
	.w6(32'hbb0a64fd),
	.w7(32'hbc3a5526),
	.w8(32'hbb1131c7),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3c872),
	.w1(32'hbb5541ac),
	.w2(32'hbb592a5d),
	.w3(32'hbafb175f),
	.w4(32'hbafec73c),
	.w5(32'h3acc6536),
	.w6(32'hbb48f646),
	.w7(32'hbb9eaf15),
	.w8(32'h3b93e9ae),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4cd4),
	.w1(32'hbae74c1d),
	.w2(32'hbba134f1),
	.w3(32'hbbdc6e41),
	.w4(32'h3b956d6e),
	.w5(32'hbbb6ed38),
	.w6(32'hbb424063),
	.w7(32'h3a6979d8),
	.w8(32'hbb908e8f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87b072),
	.w1(32'hbaf7b839),
	.w2(32'hba249a59),
	.w3(32'hbbaa8172),
	.w4(32'hbb8321b3),
	.w5(32'hbafaedbc),
	.w6(32'hbba5b42a),
	.w7(32'hbc076077),
	.w8(32'hbb39612c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925698),
	.w1(32'hba88f6aa),
	.w2(32'hbb552fc2),
	.w3(32'hbae8fc03),
	.w4(32'h3a05019b),
	.w5(32'hbb565931),
	.w6(32'h3b7ff027),
	.w7(32'h3b623afa),
	.w8(32'h3a623caf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0c8d6),
	.w1(32'h3ae02657),
	.w2(32'hbadd6e2e),
	.w3(32'h3b9e7894),
	.w4(32'h3accd1e8),
	.w5(32'hbbcbc050),
	.w6(32'h3b0fedcc),
	.w7(32'hbaab1163),
	.w8(32'hbb0f7fb3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ad138),
	.w1(32'h3b536c49),
	.w2(32'hbaafc51f),
	.w3(32'hbb92868a),
	.w4(32'hbbae2186),
	.w5(32'hbae52f07),
	.w6(32'hbb28fb2e),
	.w7(32'hbb3b08d2),
	.w8(32'hbb440bee),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71514e),
	.w1(32'h3c701748),
	.w2(32'hbb96991b),
	.w3(32'h3beef058),
	.w4(32'h3b38a6b3),
	.w5(32'h3c3f1837),
	.w6(32'h393161b3),
	.w7(32'hbb5eeeb0),
	.w8(32'h3afe4ad9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ad9f3),
	.w1(32'h3c374ff8),
	.w2(32'h3b46f3cb),
	.w3(32'h3bee607b),
	.w4(32'h3b5a5390),
	.w5(32'hbc5cbff6),
	.w6(32'h3ce981f1),
	.w7(32'h3c56a3be),
	.w8(32'hb9a9be9a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1db313),
	.w1(32'hbb0c1b94),
	.w2(32'hbb745bd6),
	.w3(32'hbbc4ce9e),
	.w4(32'hbaf20df3),
	.w5(32'hbb603603),
	.w6(32'h3bb5638f),
	.w7(32'h3beca4ac),
	.w8(32'hbb8a31d9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f9805),
	.w1(32'hbb820707),
	.w2(32'hbb0f2a71),
	.w3(32'hbbe275bf),
	.w4(32'h3a8ae195),
	.w5(32'h3a6d0699),
	.w6(32'hbb9ad5d8),
	.w7(32'h3b6b5b9c),
	.w8(32'h39f7c232),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace972d),
	.w1(32'hbb8a5195),
	.w2(32'hbb573c26),
	.w3(32'hbb5cbcb6),
	.w4(32'hbb91a767),
	.w5(32'h3c0d4db6),
	.w6(32'hbb6bf9e4),
	.w7(32'hbb38c7d1),
	.w8(32'h3c258130),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bc411),
	.w1(32'hbc19ab71),
	.w2(32'h3bda12a6),
	.w3(32'h3b0dbdea),
	.w4(32'hbbce27bf),
	.w5(32'hbbb91c5f),
	.w6(32'hbc229e04),
	.w7(32'hbaaf201c),
	.w8(32'h3b84750e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa025c),
	.w1(32'hbae8c274),
	.w2(32'h3ad97114),
	.w3(32'hbb1b7dc7),
	.w4(32'hbaeed25b),
	.w5(32'hbb9b1593),
	.w6(32'hbb24a198),
	.w7(32'hbb8e4fc0),
	.w8(32'hbb64f10a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5bddb),
	.w1(32'hbb0816b8),
	.w2(32'hb9c2827f),
	.w3(32'h3afd4f26),
	.w4(32'h39a64d4d),
	.w5(32'hba139bc0),
	.w6(32'h3b0ea637),
	.w7(32'h3b9b0747),
	.w8(32'hbb162149),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974e2d6),
	.w1(32'h3ab851bb),
	.w2(32'hbb4ddf9c),
	.w3(32'h39140874),
	.w4(32'hbb302d41),
	.w5(32'hbbc89d06),
	.w6(32'h3bd4b1fa),
	.w7(32'h3bb71cfc),
	.w8(32'hbb1284b7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6c7f),
	.w1(32'h3bdbf428),
	.w2(32'h3a47c121),
	.w3(32'hbbfeb745),
	.w4(32'hbb4b11f4),
	.w5(32'h3b23b56b),
	.w6(32'h3b3253a5),
	.w7(32'h39cb0367),
	.w8(32'hbb976bf0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d56a),
	.w1(32'h3c2e7318),
	.w2(32'hbb0d478c),
	.w3(32'hbba7c7f1),
	.w4(32'hbb88e3e7),
	.w5(32'hbbcddc9e),
	.w6(32'h3b21bb60),
	.w7(32'h3c2a69f8),
	.w8(32'hbb4c505f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71d2e6),
	.w1(32'hbbaf592b),
	.w2(32'h3b5129a2),
	.w3(32'hbc887861),
	.w4(32'hbbc755a3),
	.w5(32'hbba90838),
	.w6(32'hbc20665e),
	.w7(32'hbb4a9104),
	.w8(32'h39367eaf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57683a),
	.w1(32'h3887877c),
	.w2(32'h3b3302a1),
	.w3(32'h3aa31f68),
	.w4(32'h396cd2e0),
	.w5(32'hba3e46ca),
	.w6(32'h3b93afde),
	.w7(32'h3b84e60d),
	.w8(32'hbb36f153),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde5404),
	.w1(32'h3bb856b0),
	.w2(32'hbb3ee013),
	.w3(32'h3ad2399b),
	.w4(32'hbad6c6c0),
	.w5(32'hbb5f0118),
	.w6(32'h3b770ba1),
	.w7(32'h3a4310c5),
	.w8(32'hbbc413a3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc320bc1),
	.w1(32'hbc2325a0),
	.w2(32'hbc056930),
	.w3(32'h3b07c690),
	.w4(32'hba67dbc9),
	.w5(32'hbb923d4b),
	.w6(32'hbab466a8),
	.w7(32'hbae00bd3),
	.w8(32'hba76a9d3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277a66),
	.w1(32'h3ba0a430),
	.w2(32'h3b27d581),
	.w3(32'hbbbbf1f0),
	.w4(32'hbac26a7a),
	.w5(32'hbc289d4d),
	.w6(32'hb980e91e),
	.w7(32'h3b9225ec),
	.w8(32'hbc27e007),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804fdf),
	.w1(32'h3b558e39),
	.w2(32'h3af4a33e),
	.w3(32'hbbfcf381),
	.w4(32'hbb39cb04),
	.w5(32'h3c51adb1),
	.w6(32'h3b48a005),
	.w7(32'h3b205c35),
	.w8(32'h3c0b5f96),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb6667),
	.w1(32'h3a8e8b9e),
	.w2(32'h3c086580),
	.w3(32'h3c3f5e31),
	.w4(32'h3c8c77f9),
	.w5(32'hbbb602a6),
	.w6(32'h3be31b69),
	.w7(32'h3bbf6f02),
	.w8(32'hbb78766c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02854a),
	.w1(32'hbb28d620),
	.w2(32'hbb6c5733),
	.w3(32'hbbc2f259),
	.w4(32'hb9da8c04),
	.w5(32'hb7d4d3b8),
	.w6(32'hbb003eb8),
	.w7(32'hbb7390da),
	.w8(32'h3a03868c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34823b),
	.w1(32'hb8a150a0),
	.w2(32'h3a14c49c),
	.w3(32'hbbf17801),
	.w4(32'hbbbb0848),
	.w5(32'h3b522977),
	.w6(32'h39a62d0f),
	.w7(32'h3b1038dd),
	.w8(32'h3bd8d4a6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc44ad),
	.w1(32'h3b2822cd),
	.w2(32'h3a991aee),
	.w3(32'h3aa64e84),
	.w4(32'h3ba768e6),
	.w5(32'hbac7635e),
	.w6(32'hbb883f7a),
	.w7(32'h3b024386),
	.w8(32'h3af05e0e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b837516),
	.w1(32'hbb8f7f09),
	.w2(32'hbbe07bd5),
	.w3(32'hbb559ab2),
	.w4(32'hbbc360b7),
	.w5(32'h3acad178),
	.w6(32'hbb3afe5d),
	.w7(32'hbbb5a830),
	.w8(32'hbac0595d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0748fa),
	.w1(32'hbbb4579a),
	.w2(32'hbacdfe85),
	.w3(32'hba57b1b0),
	.w4(32'hb9d0a4cc),
	.w5(32'hbaf63a01),
	.w6(32'hbb85be84),
	.w7(32'h3ba0f502),
	.w8(32'h3b37a338),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b238f),
	.w1(32'h3c8c29c7),
	.w2(32'hbc45d467),
	.w3(32'h3cae5361),
	.w4(32'hbb2a95ff),
	.w5(32'hbbfa558f),
	.w6(32'h3cf77ebb),
	.w7(32'hbaf03662),
	.w8(32'hbbf50da4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c78f5),
	.w1(32'hbbee7f83),
	.w2(32'h3b95828d),
	.w3(32'h3bf05f07),
	.w4(32'h3c6a173c),
	.w5(32'h3b255123),
	.w6(32'hba7b3187),
	.w7(32'h3c9d4911),
	.w8(32'h3c4be197),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6290f),
	.w1(32'h3d03a9d1),
	.w2(32'hb98677c2),
	.w3(32'h3cf43edc),
	.w4(32'h3ca2aa4e),
	.w5(32'h3a31d736),
	.w6(32'h3cc8f410),
	.w7(32'h3b8ed4e9),
	.w8(32'hbc140035),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd53552),
	.w1(32'hbb2dd18f),
	.w2(32'h39d327eb),
	.w3(32'hba606cf5),
	.w4(32'h3bb25639),
	.w5(32'h3bbf33af),
	.w6(32'hbb4467d0),
	.w7(32'h3bc3fc8c),
	.w8(32'h3be80961),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c674f61),
	.w1(32'h3c0cd956),
	.w2(32'hbc512529),
	.w3(32'h3c85b0b6),
	.w4(32'hbb49dc91),
	.w5(32'hbc06f565),
	.w6(32'h3c783dd3),
	.w7(32'h3b3deb8f),
	.w8(32'hbb942e6f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a477b52),
	.w1(32'hbb0b7bed),
	.w2(32'hbc12fca4),
	.w3(32'h3c0a35fd),
	.w4(32'hbb2cedb0),
	.w5(32'hbbb43429),
	.w6(32'h3b89859a),
	.w7(32'hbb4fa20e),
	.w8(32'hbbf6ec6e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd223e),
	.w1(32'h3ac014f4),
	.w2(32'h3afed9d9),
	.w3(32'hbb97b053),
	.w4(32'h39f625af),
	.w5(32'h3bb021dd),
	.w6(32'hbbeb6b79),
	.w7(32'hbbcd0903),
	.w8(32'h3acfa6e1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9802586),
	.w1(32'hbbcfdcf5),
	.w2(32'h3a31bc84),
	.w3(32'h386ef345),
	.w4(32'h3b96d03f),
	.w5(32'hbaea0db9),
	.w6(32'hbaaa5268),
	.w7(32'h39b1457d),
	.w8(32'hb9bb78bf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86758c),
	.w1(32'h3a0491c4),
	.w2(32'hbbc4633c),
	.w3(32'hba5f05ef),
	.w4(32'hbba81376),
	.w5(32'hbb824b81),
	.w6(32'h3b67df5b),
	.w7(32'h3c051b23),
	.w8(32'hbadf46d2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ef60e),
	.w1(32'h3c24ffa0),
	.w2(32'h3b9ed1cc),
	.w3(32'h3c0ac6ca),
	.w4(32'h3c67d199),
	.w5(32'h3b9919dd),
	.w6(32'h3aa90f86),
	.w7(32'h3ba44292),
	.w8(32'h3a1e493e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e8325),
	.w1(32'hbb408847),
	.w2(32'hbc722f59),
	.w3(32'hbc40b853),
	.w4(32'hbc7b0e30),
	.w5(32'hbc94179d),
	.w6(32'hbbd0c0ce),
	.w7(32'hbc19b437),
	.w8(32'hbbaec135),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef1cec),
	.w1(32'h3c098754),
	.w2(32'h3c032757),
	.w3(32'h3bae6957),
	.w4(32'h3c415d11),
	.w5(32'h3bff5196),
	.w6(32'h3939117a),
	.w7(32'h3c3e046d),
	.w8(32'h3bcc3d0a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0668fc),
	.w1(32'hbb859e72),
	.w2(32'hbb929cf9),
	.w3(32'hbbf8183a),
	.w4(32'hbbb378ee),
	.w5(32'hbb995331),
	.w6(32'hbb62c85c),
	.w7(32'hbb81d2b8),
	.w8(32'hbb9d137c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7cdb0),
	.w1(32'h3c0651a4),
	.w2(32'hbb0dd0a6),
	.w3(32'h3b4bf221),
	.w4(32'h3b74cc6c),
	.w5(32'hb94475d4),
	.w6(32'hb9d357d8),
	.w7(32'hbabcccc2),
	.w8(32'hbba9e968),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baf9fd),
	.w1(32'hba754da9),
	.w2(32'hba32b9b6),
	.w3(32'hb9c242a3),
	.w4(32'hba77254f),
	.w5(32'hba4f2930),
	.w6(32'hb9dcb747),
	.w7(32'hba3d3b6a),
	.w8(32'hba016eed),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04daa5),
	.w1(32'hbc5a4ff5),
	.w2(32'hbb8dea6d),
	.w3(32'hbbaa736f),
	.w4(32'hbb485320),
	.w5(32'hbc1b87bd),
	.w6(32'hbb3ae538),
	.w7(32'hbc0f7c30),
	.w8(32'hbc086bce),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d8d40),
	.w1(32'hb8db8926),
	.w2(32'h3b2cb27c),
	.w3(32'h3b2ffd21),
	.w4(32'h3b181444),
	.w5(32'hbb127adc),
	.w6(32'h3af8691f),
	.w7(32'h3b46b2cd),
	.w8(32'hb9946604),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960b1fb),
	.w1(32'h3819d763),
	.w2(32'h3909b4e1),
	.w3(32'hb960baa4),
	.w4(32'h38c5d314),
	.w5(32'h393e0df6),
	.w6(32'hb94e90e3),
	.w7(32'h38a32623),
	.w8(32'h38eeec29),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa09168),
	.w1(32'hbadef07c),
	.w2(32'hbb967a8f),
	.w3(32'h39847752),
	.w4(32'hbab4e448),
	.w5(32'hbb5fc9f3),
	.w6(32'hba4336c8),
	.w7(32'hba95f9dd),
	.w8(32'hba776811),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3206b4),
	.w1(32'h3aeed263),
	.w2(32'hb9d75838),
	.w3(32'hbbbcd06d),
	.w4(32'hbb82ce0a),
	.w5(32'hbba43dba),
	.w6(32'hbb1f4ba9),
	.w7(32'hbafbe2af),
	.w8(32'hbae1f94b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a630),
	.w1(32'hbb4134f7),
	.w2(32'hbb010711),
	.w3(32'hbb353d9e),
	.w4(32'hbab34446),
	.w5(32'hba3774d1),
	.w6(32'hbadc6474),
	.w7(32'hbac19534),
	.w8(32'hbaeed2f0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace3fb2),
	.w1(32'hbb44f146),
	.w2(32'h39ca89b3),
	.w3(32'h3ad57bda),
	.w4(32'hbabb4c55),
	.w5(32'hb9e6ed2d),
	.w6(32'hba81fe0d),
	.w7(32'hb9af90e4),
	.w8(32'h3a6d0861),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5bbcc),
	.w1(32'hbb0a283f),
	.w2(32'hbabff070),
	.w3(32'hba3963b9),
	.w4(32'hbb08d69f),
	.w5(32'hbb056e1d),
	.w6(32'hbadd8e0f),
	.w7(32'hbb77305e),
	.w8(32'hbb84bbcf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b974b58),
	.w1(32'h3bb96ce7),
	.w2(32'h3b5d26fc),
	.w3(32'hbb5f345b),
	.w4(32'hbb0bdefd),
	.w5(32'hbb94c4c1),
	.w6(32'h3b95aed7),
	.w7(32'h3bcae7c9),
	.w8(32'h3b26046a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04c9e0),
	.w1(32'hbb92d097),
	.w2(32'hbc5b6dd6),
	.w3(32'hbaed0ae8),
	.w4(32'hbba40284),
	.w5(32'hbc0690e6),
	.w6(32'hbbc20996),
	.w7(32'hbbba4fd6),
	.w8(32'hbbfb97a4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca3b7f),
	.w1(32'h3968bfc7),
	.w2(32'hb9857c45),
	.w3(32'hba9d6318),
	.w4(32'hb95c836e),
	.w5(32'hb9ba3561),
	.w6(32'hb954112b),
	.w7(32'h3a38f322),
	.w8(32'hb9d38205),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3857aa7e),
	.w1(32'hb7a9262c),
	.w2(32'hb783c426),
	.w3(32'h38242418),
	.w4(32'h379c217c),
	.w5(32'h37929f09),
	.w6(32'h37c23ffa),
	.w7(32'hb7e05a2b),
	.w8(32'h366c0003),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12d067),
	.w1(32'hbaa58462),
	.w2(32'hbb069368),
	.w3(32'hba3c6075),
	.w4(32'hbaa40928),
	.w5(32'hbabb4169),
	.w6(32'hb9acf2fd),
	.w7(32'hba84e153),
	.w8(32'hba848e71),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66ef807),
	.w1(32'hb92e87a2),
	.w2(32'hb8f142e2),
	.w3(32'hb79deb14),
	.w4(32'hb8aee806),
	.w5(32'hb85a6e0e),
	.w6(32'hb8599bf5),
	.w7(32'h38206fb6),
	.w8(32'hb8936498),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fefe8f),
	.w1(32'hba664042),
	.w2(32'hba5ecc5e),
	.w3(32'hba137c6a),
	.w4(32'hba48bc27),
	.w5(32'hba2acc73),
	.w6(32'hb89c381b),
	.w7(32'hb901bb3a),
	.w8(32'hb99a7127),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ed826),
	.w1(32'hbb127cd4),
	.w2(32'hbb47bb0c),
	.w3(32'hbb52d4ec),
	.w4(32'hba9584d2),
	.w5(32'hbaab24d7),
	.w6(32'hbaab3c3e),
	.w7(32'h3a66417c),
	.w8(32'hba304f6e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba347e),
	.w1(32'h385693ac),
	.w2(32'h3a0d6267),
	.w3(32'hba0b13ff),
	.w4(32'hb9915ee0),
	.w5(32'h39916c6f),
	.w6(32'hba69d21f),
	.w7(32'hb9d625e4),
	.w8(32'hb861e765),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc3129),
	.w1(32'h3b8e714a),
	.w2(32'h3b00bd38),
	.w3(32'hbad2f7ea),
	.w4(32'h3a8f661a),
	.w5(32'h39327243),
	.w6(32'h3b0199bb),
	.w7(32'h3b18dd25),
	.w8(32'h38cc4ae0),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd307db),
	.w1(32'hbbba589b),
	.w2(32'h38718b60),
	.w3(32'hbbaf41a8),
	.w4(32'hbbb02904),
	.w5(32'hba3fc6bb),
	.w6(32'hbbc33be1),
	.w7(32'hbc049fb9),
	.w8(32'hbbca9d87),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78d6743),
	.w1(32'hb8b21fb0),
	.w2(32'hb8638a0b),
	.w3(32'h3724bcc8),
	.w4(32'hb7e64784),
	.w5(32'hb80d6bc2),
	.w6(32'h38287b41),
	.w7(32'h346ccdcb),
	.w8(32'hb73f9e92),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dae4c8),
	.w1(32'h38d0a0a6),
	.w2(32'h3935c7a5),
	.w3(32'hb8dd054e),
	.w4(32'h379caec3),
	.w5(32'h3931a2a2),
	.w6(32'h37905bb4),
	.w7(32'h392cbe38),
	.w8(32'h39465e1b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379d78eb),
	.w1(32'hb694364e),
	.w2(32'h361cb794),
	.w3(32'h380b9af6),
	.w4(32'h37523fe9),
	.w5(32'h378c3a86),
	.w6(32'h37a9d8ea),
	.w7(32'h370b74e1),
	.w8(32'h37612e25),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9926249),
	.w1(32'h39bb366e),
	.w2(32'h3a4a3aa9),
	.w3(32'hbaaa176c),
	.w4(32'hba6e4ced),
	.w5(32'h3967f7c1),
	.w6(32'hba27df94),
	.w7(32'hbac98768),
	.w8(32'hba4017ac),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c395e4a),
	.w1(32'h3bcbb772),
	.w2(32'hbc02e325),
	.w3(32'hb98a33fe),
	.w4(32'hba93796e),
	.w5(32'hbc38b0eb),
	.w6(32'h3c01f087),
	.w7(32'h3c189634),
	.w8(32'hba6b5efa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b735c),
	.w1(32'h3b3b434c),
	.w2(32'hbb3b6366),
	.w3(32'h3a059944),
	.w4(32'h39a148ae),
	.w5(32'hbb56943e),
	.w6(32'h39332b33),
	.w7(32'h3aea512f),
	.w8(32'hbb048879),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade36d3),
	.w1(32'h3a9893cd),
	.w2(32'hb93c71af),
	.w3(32'h3a971655),
	.w4(32'h3a48bd16),
	.w5(32'h3790d442),
	.w6(32'h39a7e367),
	.w7(32'h3a024ca1),
	.w8(32'hb9da4c92),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38592263),
	.w1(32'hbaa22739),
	.w2(32'hbb597695),
	.w3(32'hbb1f5db9),
	.w4(32'hbafaee43),
	.w5(32'hbb31cf04),
	.w6(32'h3ab70939),
	.w7(32'hba53e2a0),
	.w8(32'hbb37e2fa),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112698),
	.w1(32'hba74d301),
	.w2(32'hba8af2f4),
	.w3(32'hbac0e8dc),
	.w4(32'hb98d4906),
	.w5(32'hba7b59d1),
	.w6(32'hba8ba816),
	.w7(32'hba34a03e),
	.w8(32'hba9b6df0),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dbf68),
	.w1(32'hba4642da),
	.w2(32'hbb8a8aec),
	.w3(32'hbb0b5307),
	.w4(32'hbac1f0b0),
	.w5(32'hbb5cbfd9),
	.w6(32'hba3a7f86),
	.w7(32'hbaa38dde),
	.w8(32'hbb2eea32),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb118fa6),
	.w1(32'hbb8582fd),
	.w2(32'hbba53ff7),
	.w3(32'h3985392d),
	.w4(32'hbb33d381),
	.w5(32'hbb8c1241),
	.w6(32'hb8e053e4),
	.w7(32'hbb1f57e0),
	.w8(32'hbbac6719),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c9b4f),
	.w1(32'h3bde9da6),
	.w2(32'hbb148f8e),
	.w3(32'hbafc3d58),
	.w4(32'h3b79c834),
	.w5(32'hba781283),
	.w6(32'hb9977b01),
	.w7(32'h3b00c945),
	.w8(32'hbb64bf56),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada3dd5),
	.w1(32'hba95733e),
	.w2(32'h3a87e961),
	.w3(32'hb8c141cd),
	.w4(32'h39efe8c8),
	.w5(32'h3a2c4820),
	.w6(32'hbae38f8c),
	.w7(32'hba290283),
	.w8(32'hba0e1265),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3f3b8),
	.w1(32'hb9b274d7),
	.w2(32'hbb92eb96),
	.w3(32'h3ab0d32a),
	.w4(32'h38775286),
	.w5(32'hbb1c9f75),
	.w6(32'hba00dc54),
	.w7(32'hba65dada),
	.w8(32'hbb061ade),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c1209),
	.w1(32'h3bb55a1f),
	.w2(32'hba35d785),
	.w3(32'h3b7065bd),
	.w4(32'h3b9cf60c),
	.w5(32'hba1f18f7),
	.w6(32'h3b4caf9f),
	.w7(32'h3ba6ced2),
	.w8(32'hb9bcec56),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2768a6),
	.w1(32'hba259d86),
	.w2(32'hb91ef433),
	.w3(32'hbb28d9d4),
	.w4(32'hb994a644),
	.w5(32'hbac0975b),
	.w6(32'h36c7b848),
	.w7(32'h3b1e8361),
	.w8(32'h3a9d2622),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b95a9),
	.w1(32'h3b1c1063),
	.w2(32'hbb83536a),
	.w3(32'h3aeca0f3),
	.w4(32'h3a4bafc3),
	.w5(32'hbac97f30),
	.w6(32'h3a4c6e29),
	.w7(32'h3a8dc94c),
	.w8(32'hbb311822),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27b06),
	.w1(32'hb9d8f7eb),
	.w2(32'hba536b75),
	.w3(32'hbab40cfc),
	.w4(32'hba00afbf),
	.w5(32'hba185f6a),
	.w6(32'hba6f5675),
	.w7(32'hb9de9a24),
	.w8(32'hb9bfd4ca),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab682e),
	.w1(32'h3ace241b),
	.w2(32'h3b892f1a),
	.w3(32'hbb96ff21),
	.w4(32'h3abb1f55),
	.w5(32'h3ab960bc),
	.w6(32'hbbb09b9e),
	.w7(32'hbaa7f509),
	.w8(32'hb9b10cdb),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa09708),
	.w1(32'h393863c9),
	.w2(32'hbaa4bc35),
	.w3(32'hb98af9a4),
	.w4(32'hb9f50b74),
	.w5(32'hbaabd75e),
	.w6(32'h39e41024),
	.w7(32'hba28b536),
	.w8(32'hb93d0038),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3903b060),
	.w1(32'h38b89ffe),
	.w2(32'h37b31cd5),
	.w3(32'h381c6815),
	.w4(32'h38fefb0a),
	.w5(32'hb8d2be15),
	.w6(32'h39940d29),
	.w7(32'h380e585e),
	.w8(32'hb5e88164),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a789e),
	.w1(32'h391939d9),
	.w2(32'h3855ec37),
	.w3(32'hb906cb6d),
	.w4(32'h38e7db02),
	.w5(32'h394a1826),
	.w6(32'h37eb4a00),
	.w7(32'h3828534e),
	.w8(32'h39202951),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a2bfd6),
	.w1(32'h38494e51),
	.w2(32'h3adc6a42),
	.w3(32'hb9b32bdf),
	.w4(32'hb7e32810),
	.w5(32'h3b0ef645),
	.w6(32'h386fae1f),
	.w7(32'h3a357d8a),
	.w8(32'h3b2a6d1f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a201),
	.w1(32'h39f287e8),
	.w2(32'h3a820e3d),
	.w3(32'h3b44b35a),
	.w4(32'h3b8148cd),
	.w5(32'h3b853968),
	.w6(32'h3aae7fe5),
	.w7(32'h3ac7e3ae),
	.w8(32'h3b1760fb),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f6c14),
	.w1(32'h3acbccf1),
	.w2(32'h3b7bb3d7),
	.w3(32'hbc54e1fd),
	.w4(32'hbc035b60),
	.w5(32'hbb6d2b8b),
	.w6(32'hbba079be),
	.w7(32'hbb208a23),
	.w8(32'h3a3fe1d4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81eabe6),
	.w1(32'hb807617c),
	.w2(32'hb589d1f8),
	.w3(32'hb7d2187a),
	.w4(32'hb7fda5c5),
	.w5(32'hb6ab89ed),
	.w6(32'hb7d15389),
	.w7(32'hb7f3efac),
	.w8(32'hb79f81dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff8edd),
	.w1(32'h3b3b87ea),
	.w2(32'hbacac840),
	.w3(32'hbb4ce816),
	.w4(32'h3a5c7441),
	.w5(32'hbb2df4b6),
	.w6(32'hbb3ca270),
	.w7(32'hbaa0891b),
	.w8(32'hbb23df2b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae74691),
	.w1(32'hb9969502),
	.w2(32'hba3bbf71),
	.w3(32'hbb17c299),
	.w4(32'hbadea34e),
	.w5(32'hbab89b4a),
	.w6(32'hba9b0dfe),
	.w7(32'hbacbcd8a),
	.w8(32'hbab991e3),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b522b2a),
	.w1(32'h3bec0079),
	.w2(32'h3b0dd4ef),
	.w3(32'h3a420f53),
	.w4(32'h3b5c3d32),
	.w5(32'h3a2a6d59),
	.w6(32'h3a734050),
	.w7(32'h38a3a905),
	.w8(32'hbb08c9af),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26c523),
	.w1(32'h3ae82698),
	.w2(32'hba203e5c),
	.w3(32'hbba3da67),
	.w4(32'h3bcafceb),
	.w5(32'h3b6bccf1),
	.w6(32'hbb314eff),
	.w7(32'h3a09ed17),
	.w8(32'hbab529c6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39262974),
	.w1(32'hbad4d892),
	.w2(32'hbb36aebd),
	.w3(32'hb8d86e93),
	.w4(32'hbb07c28e),
	.w5(32'hbb094ed1),
	.w6(32'h39d78574),
	.w7(32'hbb0db151),
	.w8(32'hbb08daf6),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179d1c),
	.w1(32'hb980adb4),
	.w2(32'hb962d87c),
	.w3(32'hb9d3e4d5),
	.w4(32'hb9aa5836),
	.w5(32'hb8890b9a),
	.w6(32'hb9f1d8be),
	.w7(32'hb96829df),
	.w8(32'hb92b89b8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfec19),
	.w1(32'h36a43335),
	.w2(32'h3a72e0a7),
	.w3(32'h3a85d667),
	.w4(32'h3b5c006a),
	.w5(32'h3b832b6b),
	.w6(32'h3adb825c),
	.w7(32'h3bb3c5f7),
	.w8(32'h3b948cb6),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba111971),
	.w1(32'h3a4b683d),
	.w2(32'h3ac10515),
	.w3(32'h3baf82cf),
	.w4(32'h3bd7e5d4),
	.w5(32'h3bacb1dd),
	.w6(32'h3b24194a),
	.w7(32'h3bb95f17),
	.w8(32'h3b8ef24d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55118c),
	.w1(32'hbacea18c),
	.w2(32'h39a60b98),
	.w3(32'hbb082b08),
	.w4(32'hba34d299),
	.w5(32'h3a3983bf),
	.w6(32'hbaf296c3),
	.w7(32'hba99e899),
	.w8(32'hb78e9ee9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaed11c),
	.w1(32'h3ab8852b),
	.w2(32'h38fe47f8),
	.w3(32'h3a20604b),
	.w4(32'h3aa1e0c8),
	.w5(32'h3a01aa5c),
	.w6(32'h3a90c922),
	.w7(32'h3a3cc5d1),
	.w8(32'hba4595f6),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981d9b2),
	.w1(32'hb9de204b),
	.w2(32'hba2fa957),
	.w3(32'hb99c9e44),
	.w4(32'hba30f87b),
	.w5(32'hba3efeba),
	.w6(32'hb9b3e5c3),
	.w7(32'hba2ac074),
	.w8(32'hba53a19b),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56ae30),
	.w1(32'h3b316d04),
	.w2(32'hbb360945),
	.w3(32'h3aa495f1),
	.w4(32'h39e5bfb2),
	.w5(32'hbb81ca7c),
	.w6(32'h39cd7087),
	.w7(32'h3b3a28a0),
	.w8(32'hba576c14),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27fa7b),
	.w1(32'h3b2ca6b0),
	.w2(32'h3afa385c),
	.w3(32'h3b4fa04f),
	.w4(32'h3b34857f),
	.w5(32'h3a6fc9bf),
	.w6(32'h3aeba9e0),
	.w7(32'h3a8a18c5),
	.w8(32'h3975da94),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510aca),
	.w1(32'h38dd849a),
	.w2(32'h3a9f0193),
	.w3(32'hbadb9010),
	.w4(32'hb7f4cbd7),
	.w5(32'h3ab4d4b6),
	.w6(32'hba13c429),
	.w7(32'h3b82b035),
	.w8(32'h3b4c3190),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a3911),
	.w1(32'hb8d5ea72),
	.w2(32'h38bbb285),
	.w3(32'hb919e16c),
	.w4(32'h36ba3cbd),
	.w5(32'h392ac526),
	.w6(32'hb76b42bf),
	.w7(32'h387d5fef),
	.w8(32'h39292868),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62cefa),
	.w1(32'h3ae0bd91),
	.w2(32'hbb643853),
	.w3(32'h3a9310fc),
	.w4(32'hbb22293b),
	.w5(32'hbb91f621),
	.w6(32'h3b8e2215),
	.w7(32'h3b08ea1d),
	.w8(32'h3aa5eb3f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a79454),
	.w1(32'hb893e5b4),
	.w2(32'hb8361099),
	.w3(32'hb904b5d4),
	.w4(32'hb8cf18e4),
	.w5(32'hb8b05d10),
	.w6(32'hb8f39b5f),
	.w7(32'hb8c61807),
	.w8(32'hb88b93c8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bc6b28),
	.w1(32'h3874f292),
	.w2(32'h38a39de8),
	.w3(32'hb774ee20),
	.w4(32'h37e64af8),
	.w5(32'h37b3702c),
	.w6(32'hb86fa940),
	.w7(32'h378cacab),
	.w8(32'h3879744a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985957),
	.w1(32'h3a81ca85),
	.w2(32'h3b0d4719),
	.w3(32'h3b573935),
	.w4(32'h3b4f0117),
	.w5(32'h3b570330),
	.w6(32'h3ae33a5c),
	.w7(32'h3b3a34aa),
	.w8(32'h3b126b93),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba87c51),
	.w1(32'h3b966d06),
	.w2(32'hbb095421),
	.w3(32'h3af667a5),
	.w4(32'h3a0cf6c0),
	.w5(32'hbb7e9655),
	.w6(32'h3be76c59),
	.w7(32'h3bf85552),
	.w8(32'h38aa7666),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad01fbd),
	.w1(32'hba8187d6),
	.w2(32'hb9b2c393),
	.w3(32'hbaa3e170),
	.w4(32'hba1ff59b),
	.w5(32'h391287f9),
	.w6(32'hbb09604c),
	.w7(32'hba7c6623),
	.w8(32'hb9a15992),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23a88b),
	.w1(32'hb94c2252),
	.w2(32'h36cdbc38),
	.w3(32'hbb516d90),
	.w4(32'hbb0b21dd),
	.w5(32'hba04cbc4),
	.w6(32'hbb32d270),
	.w7(32'hbae16c89),
	.w8(32'hba6c3d9e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15c474),
	.w1(32'h3b23813a),
	.w2(32'hba06ddf7),
	.w3(32'h39952839),
	.w4(32'h3b446e1a),
	.w5(32'hba5259fd),
	.w6(32'hba3dbbb1),
	.w7(32'h3a790db2),
	.w8(32'h3966201c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f00d3),
	.w1(32'h3abe7d59),
	.w2(32'hbaa09eaa),
	.w3(32'hbbe4a1bb),
	.w4(32'h3af3680e),
	.w5(32'h3ab95646),
	.w6(32'hbb6d1466),
	.w7(32'h3b83fe68),
	.w8(32'h3b2c3e09),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1230),
	.w1(32'hbab67806),
	.w2(32'hbb0f0b74),
	.w3(32'h3ae2f5f2),
	.w4(32'h39ee4c19),
	.w5(32'hb9f8750c),
	.w6(32'h3a9aca28),
	.w7(32'h3a0ef68a),
	.w8(32'hb8f6633c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafc0f0),
	.w1(32'h3ab0ba10),
	.w2(32'hbb95524e),
	.w3(32'hba02ca3f),
	.w4(32'h393b3fc4),
	.w5(32'hbba89e3d),
	.w6(32'h3a983347),
	.w7(32'h3a9e97d8),
	.w8(32'hbb532f5a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9713d3a),
	.w1(32'hb9a36189),
	.w2(32'hb9a25416),
	.w3(32'hb9672689),
	.w4(32'hb9c5ae86),
	.w5(32'hba01e94a),
	.w6(32'hb9672a35),
	.w7(32'hb99b1155),
	.w8(32'hb9c8a065),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b157291),
	.w1(32'h38ed387d),
	.w2(32'hbb5f9265),
	.w3(32'h3a3dfef4),
	.w4(32'h389c7a14),
	.w5(32'hbb2fba75),
	.w6(32'hba27f592),
	.w7(32'hba42f6e0),
	.w8(32'hbb3a7865),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb656c95e),
	.w1(32'h369cc673),
	.w2(32'h379a58ed),
	.w3(32'h37005d73),
	.w4(32'h35c89609),
	.w5(32'h37883ad8),
	.w6(32'hb7015986),
	.w7(32'hb759c708),
	.w8(32'h37c5b97d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d4baf),
	.w1(32'h3a7973f6),
	.w2(32'h39d28237),
	.w3(32'h390f523c),
	.w4(32'h37bea366),
	.w5(32'hb917ffae),
	.w6(32'hb959b4b6),
	.w7(32'hba1d42ee),
	.w8(32'hba73a6ab),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7685571),
	.w1(32'hb9a8ec28),
	.w2(32'hb9819294),
	.w3(32'h39866867),
	.w4(32'h38e79618),
	.w5(32'hb9a49792),
	.w6(32'h397a7806),
	.w7(32'hba002da9),
	.w8(32'hba97b471),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddf930),
	.w1(32'hbb7d444e),
	.w2(32'hbbcbb3a0),
	.w3(32'hbb820119),
	.w4(32'hbbae8b43),
	.w5(32'hbbc31aef),
	.w6(32'hbbe91f7d),
	.w7(32'hbbfd1ec2),
	.w8(32'hbbe1c605),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c741d1),
	.w1(32'hb70d4216),
	.w2(32'h3559bb26),
	.w3(32'hb81c0f48),
	.w4(32'hb60fadd2),
	.w5(32'hb6a8c716),
	.w6(32'hb7c65880),
	.w7(32'hb76bd6f0),
	.w8(32'hb6328749),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39270e93),
	.w1(32'h38c2d629),
	.w2(32'h37d6f0e3),
	.w3(32'h37fe4c25),
	.w4(32'h36641f09),
	.w5(32'hb792c12d),
	.w6(32'h390e8150),
	.w7(32'h38c082be),
	.w8(32'h3856f385),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4207f8),
	.w1(32'hba5d42ee),
	.w2(32'hba69a96d),
	.w3(32'hba757b15),
	.w4(32'hbae54c0c),
	.w5(32'hbaa5f9fc),
	.w6(32'h3adc8f87),
	.w7(32'h3a599d39),
	.w8(32'hb9ee8c7c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae54c7b),
	.w1(32'hba490d0c),
	.w2(32'hbbf475ea),
	.w3(32'hbab93262),
	.w4(32'h3988796c),
	.w5(32'hbb3b4818),
	.w6(32'h3a5df037),
	.w7(32'h3a825a6a),
	.w8(32'hbb57e592),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40e07f),
	.w1(32'hbb013fa9),
	.w2(32'hbb2fc0fa),
	.w3(32'hbb3fc7ad),
	.w4(32'hba872d2c),
	.w5(32'hbb46059c),
	.w6(32'hbb9aa811),
	.w7(32'hbbc06200),
	.w8(32'hbb15d9d1),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39697ae2),
	.w1(32'h3905d7ee),
	.w2(32'h37b38847),
	.w3(32'h392286ed),
	.w4(32'hb99cb216),
	.w5(32'hb997c61f),
	.w6(32'h3850b0e1),
	.w7(32'hb731c39f),
	.w8(32'hb937b6a6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc2017),
	.w1(32'h3b45f625),
	.w2(32'h3bcfde76),
	.w3(32'hbb7f8d6f),
	.w4(32'h3b30290d),
	.w5(32'h3baaa0c7),
	.w6(32'h3c2212a3),
	.w7(32'h3cc30678),
	.w8(32'h3ca16249),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d7946),
	.w1(32'h3bd2f4a4),
	.w2(32'h3b809b5b),
	.w3(32'h3bb0e5e7),
	.w4(32'h3c25f947),
	.w5(32'h3be72358),
	.w6(32'hba8f4d5f),
	.w7(32'h3b91a093),
	.w8(32'h3a6876eb),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68e24c),
	.w1(32'h3b6b6ed2),
	.w2(32'h3acf75d2),
	.w3(32'h3b32c5ee),
	.w4(32'h3b0d94b1),
	.w5(32'h3a409d64),
	.w6(32'h3ad2cc43),
	.w7(32'hb9ab6391),
	.w8(32'hbb0262fd),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba46fc),
	.w1(32'hb89f7a85),
	.w2(32'h36fa3fe6),
	.w3(32'hb8271ac6),
	.w4(32'hb939737f),
	.w5(32'hb8fc1a76),
	.w6(32'h3739aa0a),
	.w7(32'hb71e26b6),
	.w8(32'h36b0fd99),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f44991),
	.w1(32'hb7e54770),
	.w2(32'h3919c903),
	.w3(32'h383297db),
	.w4(32'h37e03f2e),
	.w5(32'h392b1d9c),
	.w6(32'h394c10dd),
	.w7(32'h3911adf9),
	.w8(32'h395f30e0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e95584),
	.w1(32'h370fb1fc),
	.w2(32'h373a9f82),
	.w3(32'h37646460),
	.w4(32'h3660f0c3),
	.w5(32'h37084380),
	.w6(32'h3642d551),
	.w7(32'hb691a007),
	.w8(32'hb59f0f92),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9b24),
	.w1(32'h3bbd267a),
	.w2(32'hba0c9f6b),
	.w3(32'h3b42acff),
	.w4(32'h3b08e69a),
	.w5(32'hbb412554),
	.w6(32'h3b36637c),
	.w7(32'h3b3d035a),
	.w8(32'hba896e5c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3f8d2),
	.w1(32'h3a810ff2),
	.w2(32'hb6910ffa),
	.w3(32'h3afdfdc3),
	.w4(32'h3abce511),
	.w5(32'h3a931b27),
	.w6(32'h3a8bc7c7),
	.w7(32'h3b013c8b),
	.w8(32'h3a170920),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b6de8),
	.w1(32'hbbab3f00),
	.w2(32'hbb81f7ab),
	.w3(32'hbc2e084a),
	.w4(32'hbbd32f99),
	.w5(32'hbb84a3d4),
	.w6(32'hbc039241),
	.w7(32'hbbfcdce1),
	.w8(32'hba88e461),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5e8ad),
	.w1(32'hbaadbb5d),
	.w2(32'hbad65337),
	.w3(32'hba87487f),
	.w4(32'hba7ac66b),
	.w5(32'hba2514ab),
	.w6(32'hba1e8d6a),
	.w7(32'h39e76171),
	.w8(32'h3a0df30f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbd096),
	.w1(32'h3b978a51),
	.w2(32'h3b699a24),
	.w3(32'hbb1008a2),
	.w4(32'h3aaeffb4),
	.w5(32'h3adb76a7),
	.w6(32'h39869c6a),
	.w7(32'h3b677731),
	.w8(32'h3a56b6e0),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a8ae),
	.w1(32'hbb043630),
	.w2(32'hba1c2119),
	.w3(32'hbb6778d7),
	.w4(32'hbb1c595b),
	.w5(32'hbacf00ef),
	.w6(32'hba753ea2),
	.w7(32'h3918c1db),
	.w8(32'h39cdf584),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7725da1),
	.w1(32'hb767f3d5),
	.w2(32'hb7644d77),
	.w3(32'h365cc7f5),
	.w4(32'h35ffde2f),
	.w5(32'hb70eb882),
	.w6(32'h3727818a),
	.w7(32'h36180540),
	.w8(32'h364e3079),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6334b4),
	.w1(32'hbba290e8),
	.w2(32'hbb8a08b3),
	.w3(32'hbb060fcd),
	.w4(32'hbb6d86f4),
	.w5(32'hbb38c9bb),
	.w6(32'hba86320b),
	.w7(32'hbb9c9f30),
	.w8(32'hbb2d884c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37913fc4),
	.w1(32'hb7cf4600),
	.w2(32'h37c978c1),
	.w3(32'h382e27ee),
	.w4(32'h37f78589),
	.w5(32'h385b9169),
	.w6(32'hb6eaa737),
	.w7(32'hb4a4caad),
	.w8(32'h3830dbad),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae914f4),
	.w1(32'h39491bd8),
	.w2(32'hbb085148),
	.w3(32'hbb8216f5),
	.w4(32'hba4b6cd4),
	.w5(32'hbacaeccf),
	.w6(32'hbaa234dc),
	.w7(32'h3a293d40),
	.w8(32'hbb20f1d2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb397f5d),
	.w1(32'hbaccb404),
	.w2(32'hbad9f9c1),
	.w3(32'h3b10ccfa),
	.w4(32'h3ae13587),
	.w5(32'h3aeefafc),
	.w6(32'h39c504f7),
	.w7(32'h3abbd9eb),
	.w8(32'h3a7642cc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb24c777),
	.w1(32'hb9af3350),
	.w2(32'hba2a2a0d),
	.w3(32'hbac50abf),
	.w4(32'h3a2d126c),
	.w5(32'h3a80db84),
	.w6(32'hbabc85a5),
	.w7(32'h3a4e71ee),
	.w8(32'h3a398628),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9722df9),
	.w1(32'hb99965e4),
	.w2(32'h3a15824b),
	.w3(32'hb803d931),
	.w4(32'h3a179d4c),
	.w5(32'h3a775439),
	.w6(32'hba7e951e),
	.w7(32'h37f62aa3),
	.w8(32'h3a08955a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac7795),
	.w1(32'hbb32e83d),
	.w2(32'hba22c904),
	.w3(32'hbb81b434),
	.w4(32'hbb17900c),
	.w5(32'h39f74ac6),
	.w6(32'hbb54cffe),
	.w7(32'hbafa12a0),
	.w8(32'hba3b3c3b),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393736c0),
	.w1(32'h3a354028),
	.w2(32'hbb68cfe7),
	.w3(32'hba850c9c),
	.w4(32'hbaf11b4c),
	.w5(32'hbb52585c),
	.w6(32'hba677bab),
	.w7(32'hba1dbc4b),
	.w8(32'hbb5a9b1a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f2dbf),
	.w1(32'hba736088),
	.w2(32'hb9c71fde),
	.w3(32'hbc711f3d),
	.w4(32'hbc05757e),
	.w5(32'hbb86b221),
	.w6(32'hbbdee425),
	.w7(32'hbb49a99a),
	.w8(32'h3a85bd95),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c602a6),
	.w1(32'h370a2910),
	.w2(32'h3382c199),
	.w3(32'h37cd068c),
	.w4(32'h37a0a364),
	.w5(32'hb7015320),
	.w6(32'h361ca04c),
	.w7(32'h372885d4),
	.w8(32'h3644dfab),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377f9e79),
	.w1(32'h37a83ec0),
	.w2(32'hb8c72f69),
	.w3(32'hb860f3a3),
	.w4(32'h367fedeb),
	.w5(32'h37bf4000),
	.w6(32'h391c0bab),
	.w7(32'h37e18b37),
	.w8(32'h3868e381),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517ce3),
	.w1(32'h3b430e13),
	.w2(32'hba03fc98),
	.w3(32'h3ad711f3),
	.w4(32'hbb58c940),
	.w5(32'hbbe28d31),
	.w6(32'h3bff24bf),
	.w7(32'h3c0871bd),
	.w8(32'h3aec6c95),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24adf8),
	.w1(32'h3b03a19c),
	.w2(32'hbb547b43),
	.w3(32'h3ad0bf31),
	.w4(32'h3a18ea58),
	.w5(32'hbb2f268e),
	.w6(32'h3bc84c67),
	.w7(32'h3bf351b3),
	.w8(32'h3a7902be),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fe383),
	.w1(32'hbb4b95cf),
	.w2(32'hbb6cfd96),
	.w3(32'hbba09ca7),
	.w4(32'hbb1faa34),
	.w5(32'hbb1b5538),
	.w6(32'hbb2608aa),
	.w7(32'hba1ae209),
	.w8(32'hba9e0eb0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ac9a0),
	.w1(32'h3c47bbb2),
	.w2(32'hba45cb60),
	.w3(32'h3bba0b47),
	.w4(32'h3bf14fd5),
	.w5(32'hb9d89c7e),
	.w6(32'hbaee09ca),
	.w7(32'hb8a0eda2),
	.w8(32'hbb936e92),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4860ff),
	.w1(32'h39f4f7f7),
	.w2(32'h38a65344),
	.w3(32'h3a16fbc0),
	.w4(32'hba22577b),
	.w5(32'hb9bfcdc2),
	.w6(32'h3a0a23ee),
	.w7(32'hb9f25a66),
	.w8(32'hba02edcc),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad08ca8),
	.w1(32'hbaf06ecd),
	.w2(32'hbb690a34),
	.w3(32'h38c398e1),
	.w4(32'h38f7cb0d),
	.w5(32'hbb2bc86e),
	.w6(32'h3a0cebae),
	.w7(32'hba941ec5),
	.w8(32'hbade3632),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea2a7a),
	.w1(32'h3c9eca5f),
	.w2(32'hbb1252cf),
	.w3(32'h3956c47c),
	.w4(32'h3bd5fcd0),
	.w5(32'hbc0e54ca),
	.w6(32'h3ab6a556),
	.w7(32'h3c16be04),
	.w8(32'h3af3d34e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb765df8),
	.w1(32'h3b7a01bf),
	.w2(32'hbaf8b24e),
	.w3(32'hbbb96468),
	.w4(32'h3a4c9372),
	.w5(32'hb9b42292),
	.w6(32'h3bb51d22),
	.w7(32'h3c272ec4),
	.w8(32'h3bc99e98),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace58f2),
	.w1(32'h3b9cdf91),
	.w2(32'h3af70989),
	.w3(32'hbaf75e55),
	.w4(32'hbb2e1d10),
	.w5(32'hbb32380a),
	.w6(32'h398da00b),
	.w7(32'hbb534d97),
	.w8(32'hbb9a60a5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c47d),
	.w1(32'hb920c1fe),
	.w2(32'h39d4b118),
	.w3(32'hbaf31c54),
	.w4(32'h398b7748),
	.w5(32'h3a8b9c9e),
	.w6(32'hba9a4884),
	.w7(32'h3a21d9a6),
	.w8(32'h3979cddf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef9b0a),
	.w1(32'hbbbedc37),
	.w2(32'hbb54c198),
	.w3(32'hbabec6cd),
	.w4(32'hba882f48),
	.w5(32'h3a47ab5f),
	.w6(32'h3993e0a8),
	.w7(32'hb9f31f08),
	.w8(32'hbada0159),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7870fac),
	.w1(32'hb6d199e0),
	.w2(32'h36c82eb7),
	.w3(32'hb71e3da6),
	.w4(32'h3702ab0f),
	.w5(32'h3756b2ca),
	.w6(32'hb65e37f2),
	.w7(32'h373916c6),
	.w8(32'h37a24fda),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6daae4f),
	.w1(32'hb77753b7),
	.w2(32'hb6f315b1),
	.w3(32'h37a0a321),
	.w4(32'h370914d3),
	.w5(32'h347c8b34),
	.w6(32'h37e4286d),
	.w7(32'h37e0c8a0),
	.w8(32'h37c0bc3b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29aaa1),
	.w1(32'h3b8291e8),
	.w2(32'h3aef7c00),
	.w3(32'h3acee7c9),
	.w4(32'hb8108cf1),
	.w5(32'hba8f949c),
	.w6(32'h3b042a83),
	.w7(32'h3afa84bd),
	.w8(32'h3a8e8963),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37147b6c),
	.w1(32'h36983231),
	.w2(32'h37a7a6fe),
	.w3(32'h36776f42),
	.w4(32'hb788932b),
	.w5(32'hbc3d2a32),
	.w6(32'h36894374),
	.w7(32'hb755605a),
	.w8(32'h3b448614),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7bdf),
	.w1(32'h3cee192b),
	.w2(32'hbace5bd4),
	.w3(32'hbc1c1552),
	.w4(32'hbc807ca2),
	.w5(32'hbc1a09e0),
	.w6(32'h3beea64b),
	.w7(32'hbb307016),
	.w8(32'hbb162374),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb122cc),
	.w1(32'h3cf08e76),
	.w2(32'hbbd89255),
	.w3(32'hbc82e97e),
	.w4(32'hba556d42),
	.w5(32'hbc154982),
	.w6(32'h3b48a6f1),
	.w7(32'h3b7d654b),
	.w8(32'h3b71ebdd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4211d4),
	.w1(32'h3cae5be8),
	.w2(32'h3c3d3c92),
	.w3(32'hbcb3934b),
	.w4(32'hbc7f6156),
	.w5(32'h3b3e5140),
	.w6(32'h3b01dd83),
	.w7(32'hbb1fdfaa),
	.w8(32'hbbccef97),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa484ed),
	.w1(32'hb9ab73ff),
	.w2(32'h3b29a136),
	.w3(32'h3bcd5db4),
	.w4(32'h3b448f2c),
	.w5(32'hb9db3864),
	.w6(32'hba97609b),
	.w7(32'hbc1ca138),
	.w8(32'h3a0fab67),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a159414),
	.w1(32'h3b8a8769),
	.w2(32'hbbb49c0d),
	.w3(32'hbb394f00),
	.w4(32'hbbe650c9),
	.w5(32'hbc94aa41),
	.w6(32'h3b22f780),
	.w7(32'h3af926f8),
	.w8(32'h3c3b76a9),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1e3134),
	.w1(32'h3dc214f0),
	.w2(32'h3cb8b1e6),
	.w3(32'hbd9f4559),
	.w4(32'hbd25dacb),
	.w5(32'h3b2e3a54),
	.w6(32'hbba51158),
	.w7(32'hbcd064ad),
	.w8(32'hbb195dbd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb065b1),
	.w1(32'hbbb4fd64),
	.w2(32'hbb5f0a2f),
	.w3(32'hbb01abfc),
	.w4(32'hbac8af0c),
	.w5(32'hbb23f6f4),
	.w6(32'hbc53d0dd),
	.w7(32'h3b2d15b7),
	.w8(32'h3b9a4b8a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2567ac),
	.w1(32'h3c61ad96),
	.w2(32'h3c46d162),
	.w3(32'hbb1c87f5),
	.w4(32'hbbe33fda),
	.w5(32'hbb278b6b),
	.w6(32'h3c1140d0),
	.w7(32'h3bddda31),
	.w8(32'hbbba8265),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe24469),
	.w1(32'h3c9e38ee),
	.w2(32'h3c944853),
	.w3(32'h3c03b08e),
	.w4(32'hbbfbd640),
	.w5(32'h3c0bef00),
	.w6(32'hbc090521),
	.w7(32'hbc3e58ec),
	.w8(32'h3c1974fc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb34f5a),
	.w1(32'hbbb36256),
	.w2(32'h3b3f73f7),
	.w3(32'h3c36492e),
	.w4(32'h3b99045c),
	.w5(32'hbc4a6fb3),
	.w6(32'h3bac57af),
	.w7(32'h3bbf9d3b),
	.w8(32'h3baf1990),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c744),
	.w1(32'h3d22c677),
	.w2(32'h3c338fdf),
	.w3(32'hbb64fc18),
	.w4(32'hbc81586a),
	.w5(32'hbb029e40),
	.w6(32'h3c436788),
	.w7(32'hbb7a13cd),
	.w8(32'hbbfa82ee),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc891e7e),
	.w1(32'hbcc5f02f),
	.w2(32'hbc8ab6fe),
	.w3(32'h3c194792),
	.w4(32'hbb825b8e),
	.w5(32'h3b61087f),
	.w6(32'hba9e6831),
	.w7(32'hbb1e0c9f),
	.w8(32'h3ba264a7),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74f90),
	.w1(32'h3aca7669),
	.w2(32'h3b48aaed),
	.w3(32'h3c0897c1),
	.w4(32'h3b2e6617),
	.w5(32'h3be448a4),
	.w6(32'h3c0bbac2),
	.w7(32'hba93e1b8),
	.w8(32'h3b522808),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345a8a),
	.w1(32'hb9848210),
	.w2(32'hbbc90b6d),
	.w3(32'h3be8d939),
	.w4(32'h3ba3d642),
	.w5(32'h3b574426),
	.w6(32'hbbcb8687),
	.w7(32'h3b573aa6),
	.w8(32'hbc88961d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca4e214),
	.w1(32'hbcfbcc49),
	.w2(32'hbcae4f7b),
	.w3(32'h3d31af3f),
	.w4(32'h3c6512f4),
	.w5(32'h3ae6a0a6),
	.w6(32'h3bd007f4),
	.w7(32'h3b217b93),
	.w8(32'h3a2be637),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ff38c),
	.w1(32'h3b3c029a),
	.w2(32'hbb89701a),
	.w3(32'hbbe935be),
	.w4(32'h3be0f5f6),
	.w5(32'hbb8333a2),
	.w6(32'h3c5877c7),
	.w7(32'h3ba55146),
	.w8(32'h3b256e13),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd12570),
	.w1(32'h3c8272f8),
	.w2(32'h3c1fb0a5),
	.w3(32'hbc9aaf28),
	.w4(32'hba172a9b),
	.w5(32'h3b7551a7),
	.w6(32'hbaa5c4d8),
	.w7(32'hbac34912),
	.w8(32'h3b5e7a75),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d767e),
	.w1(32'hbb72e637),
	.w2(32'h3b6c3f8f),
	.w3(32'hbb3fa283),
	.w4(32'hbb9ab6b4),
	.w5(32'hba2a3e76),
	.w6(32'hbbb2ac9f),
	.w7(32'h3a1b53e0),
	.w8(32'hbb451bca),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc318dfd),
	.w1(32'hbc30639f),
	.w2(32'hbc10d42b),
	.w3(32'h3ac96cd9),
	.w4(32'hba9248f4),
	.w5(32'hbb026d9a),
	.w6(32'hbb4675d0),
	.w7(32'hbb088e6f),
	.w8(32'hbbebd705),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7068df),
	.w1(32'h3be59369),
	.w2(32'hbb00d564),
	.w3(32'hbc0ece82),
	.w4(32'h3c0e3bed),
	.w5(32'hbc792f5b),
	.w6(32'hbca3dd38),
	.w7(32'hbb74b119),
	.w8(32'hbb9f9461),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30c2dd),
	.w1(32'h3c3b50ef),
	.w2(32'hbc77dc9c),
	.w3(32'hbc9ddf49),
	.w4(32'hbc293464),
	.w5(32'hbce259f5),
	.w6(32'hbaf6e33a),
	.w7(32'hbc0d3065),
	.w8(32'hba543a1d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c612415),
	.w1(32'h3d5287e9),
	.w2(32'h3c49219b),
	.w3(32'hbd84111e),
	.w4(32'hbcfeb3fa),
	.w5(32'h3b78e216),
	.w6(32'hbc38bc2a),
	.w7(32'hbc8ba52e),
	.w8(32'h3878053e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc39d),
	.w1(32'hbb419dac),
	.w2(32'h3b5410c5),
	.w3(32'hbbc2f270),
	.w4(32'hbc11624c),
	.w5(32'hba4a8097),
	.w6(32'hbbf5b21d),
	.w7(32'hbbada7ab),
	.w8(32'h3be253df),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1a2a2),
	.w1(32'hbc9aae23),
	.w2(32'hbc40daab),
	.w3(32'h3c85a405),
	.w4(32'h3cac39ee),
	.w5(32'h3b3c620d),
	.w6(32'h3b8cb80a),
	.w7(32'h3c159b05),
	.w8(32'hbc47b2ee),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2a740),
	.w1(32'hbb732f26),
	.w2(32'hbb93e4d9),
	.w3(32'h3ccd532a),
	.w4(32'h3bcf68dd),
	.w5(32'h3c6c9e9b),
	.w6(32'h387c6eca),
	.w7(32'h3ba8038c),
	.w8(32'hb5d896d2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5311fd),
	.w1(32'hbc937d86),
	.w2(32'hbc1688d4),
	.w3(32'h3c97a24a),
	.w4(32'h3984d263),
	.w5(32'h3bfb4f6c),
	.w6(32'hb96f51e5),
	.w7(32'h3a6cda80),
	.w8(32'hbc186c74),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07ad44),
	.w1(32'hbca57617),
	.w2(32'hbc3373cc),
	.w3(32'h3c5b98ae),
	.w4(32'hba83e778),
	.w5(32'hbba01aad),
	.w6(32'h3c3da9da),
	.w7(32'h3c1b01e1),
	.w8(32'hbb13b31f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc24ca2),
	.w1(32'hbaffd3cf),
	.w2(32'hbc702eac),
	.w3(32'hbc6a8781),
	.w4(32'hbb57b3b0),
	.w5(32'hbbe58a5b),
	.w6(32'h3c30d6ea),
	.w7(32'hbc0f309a),
	.w8(32'hbc0a9b0c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baad508),
	.w1(32'hbb3433f5),
	.w2(32'hbb69dc2f),
	.w3(32'h3c38a923),
	.w4(32'hbc312b98),
	.w5(32'h3bc84b9c),
	.w6(32'hbbdf38da),
	.w7(32'hbb439cff),
	.w8(32'h3a0bb2f6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eecab),
	.w1(32'h3a9db2ce),
	.w2(32'h3ba8371a),
	.w3(32'h3a5c6cb0),
	.w4(32'h399437b7),
	.w5(32'hbb5a15a2),
	.w6(32'h3c0736b5),
	.w7(32'h3c561188),
	.w8(32'h395e05a0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule