module layer_8_featuremap_146(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90a716),
	.w1(32'h3b943a4d),
	.w2(32'hbc2e54b6),
	.w3(32'hbb8c1e5f),
	.w4(32'hbae90a67),
	.w5(32'h3bdfbf24),
	.w6(32'h3ba98b3b),
	.w7(32'hbba505b0),
	.w8(32'hbaebb5f6),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f5bf8),
	.w1(32'h3c00626b),
	.w2(32'hbb4f9138),
	.w3(32'hbbb7362b),
	.w4(32'hbb38bcdb),
	.w5(32'h3c779b8e),
	.w6(32'hbc4afff5),
	.w7(32'h3c7da999),
	.w8(32'h3caae936),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd00a2a7),
	.w1(32'hbcab2c07),
	.w2(32'hbb4f4bba),
	.w3(32'h3b4fd7bf),
	.w4(32'h3bbc2d64),
	.w5(32'h3b470161),
	.w6(32'hbc4cea5e),
	.w7(32'h3c6cb07e),
	.w8(32'h3cc683a9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e7e4e),
	.w1(32'hbbc40c13),
	.w2(32'hbc8894eb),
	.w3(32'hbbf40be0),
	.w4(32'h3b6d375a),
	.w5(32'h3b8483e4),
	.w6(32'hbc3a3717),
	.w7(32'hbc859a30),
	.w8(32'hbc0c3095),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc97c05),
	.w1(32'h3c499852),
	.w2(32'hbbcc6c0c),
	.w3(32'hbc356ca3),
	.w4(32'hbb831fdb),
	.w5(32'h3adf9e7c),
	.w6(32'h3a87e248),
	.w7(32'hbbb5aae9),
	.w8(32'hbc41b2ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d481516),
	.w1(32'h3d1fe9f1),
	.w2(32'hbcc6ae74),
	.w3(32'hbb2161f9),
	.w4(32'h3bde43ea),
	.w5(32'hbc3265e5),
	.w6(32'h3b1f85f1),
	.w7(32'hba020337),
	.w8(32'hbbc34618),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a768a81),
	.w1(32'h3cc6d01d),
	.w2(32'hbc9d1368),
	.w3(32'h3c08932d),
	.w4(32'h3ab73869),
	.w5(32'h3c7e7b65),
	.w6(32'h3c4c44df),
	.w7(32'h3ad4d0aa),
	.w8(32'hbc2c5234),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00234e),
	.w1(32'hbd065b94),
	.w2(32'hbbe422b6),
	.w3(32'hbcc9579b),
	.w4(32'hbb4e1453),
	.w5(32'hbc4e6be1),
	.w6(32'hbc54b671),
	.w7(32'h3b195004),
	.w8(32'hbc33784a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3760f3),
	.w1(32'hbba69003),
	.w2(32'hbc37b785),
	.w3(32'h3be50451),
	.w4(32'hb9610d2d),
	.w5(32'h3c2a589c),
	.w6(32'hbba1e175),
	.w7(32'hbbafc24e),
	.w8(32'hbba1bc16),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfb7d7),
	.w1(32'hbbf77fbe),
	.w2(32'h3adece49),
	.w3(32'hbc1f5578),
	.w4(32'hbc47938c),
	.w5(32'hbb97b796),
	.w6(32'hbbe8fa45),
	.w7(32'hbb9b1a2d),
	.w8(32'hbc24fd2c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2aa0b),
	.w1(32'h3c621250),
	.w2(32'h39b7d568),
	.w3(32'hbbdb5b0b),
	.w4(32'h3aef0167),
	.w5(32'h3b04e17e),
	.w6(32'h3c589155),
	.w7(32'hbc913218),
	.w8(32'hbc33e7a1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc74a202),
	.w1(32'h3b6902d6),
	.w2(32'hbc592742),
	.w3(32'h3b34cab4),
	.w4(32'hbb9d20f3),
	.w5(32'hbc5ef7a5),
	.w6(32'h3a5df258),
	.w7(32'hbc536342),
	.w8(32'hbc31c90f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1db09),
	.w1(32'h392612d6),
	.w2(32'h3b506279),
	.w3(32'hbc6a0046),
	.w4(32'h3b768105),
	.w5(32'h3c1563b1),
	.w6(32'hbc4397f3),
	.w7(32'h3b97295b),
	.w8(32'h3c020785),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b753816),
	.w1(32'h3ae95be4),
	.w2(32'h3ba42c27),
	.w3(32'h3c59e4d7),
	.w4(32'h3b908402),
	.w5(32'hba3e3487),
	.w6(32'h3ab09df8),
	.w7(32'h3c4c4bdb),
	.w8(32'h3abc4e2d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b212566),
	.w1(32'hba3ff79c),
	.w2(32'h3c143d18),
	.w3(32'h3a80013d),
	.w4(32'h3beabb92),
	.w5(32'hbb5c6b0f),
	.w6(32'hbbaef0a9),
	.w7(32'h3c3c917f),
	.w8(32'hbb0e496d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2ba6d),
	.w1(32'hba15434e),
	.w2(32'h3c45fc1b),
	.w3(32'h3a16387e),
	.w4(32'hbca65862),
	.w5(32'h3c088d5b),
	.w6(32'hbac8f2b0),
	.w7(32'hbba25406),
	.w8(32'h3cdc1079),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff46a6),
	.w1(32'h3ca75e57),
	.w2(32'hbc50368b),
	.w3(32'h3b87d11f),
	.w4(32'hbca0c350),
	.w5(32'hbd5d5710),
	.w6(32'h3c953d94),
	.w7(32'hbc05dd2e),
	.w8(32'hbd3b1376),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd72bb5a),
	.w1(32'h3ba1ed38),
	.w2(32'h3c8f60ca),
	.w3(32'hbc778468),
	.w4(32'h3c35ba57),
	.w5(32'hbc8ca024),
	.w6(32'h3cca4f33),
	.w7(32'h3c564520),
	.w8(32'hbcc01698),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c56b9c9),
	.w1(32'h3b9fc8b1),
	.w2(32'hbb0b9920),
	.w3(32'h3c166af5),
	.w4(32'hbcfb6707),
	.w5(32'hbc85a53d),
	.w6(32'h3d131c93),
	.w7(32'hbc14505f),
	.w8(32'hbb2a07f6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e1894),
	.w1(32'h3c0f2a9e),
	.w2(32'hbc10a4c4),
	.w3(32'hbc22e1df),
	.w4(32'h3b8ed1d2),
	.w5(32'h3b383ba9),
	.w6(32'h3c372e57),
	.w7(32'h3bc6ef33),
	.w8(32'hbaba8a2b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c454db5),
	.w1(32'hbc8f3a3f),
	.w2(32'hbc776896),
	.w3(32'h3caaed77),
	.w4(32'hbca2510a),
	.w5(32'h3ade9263),
	.w6(32'hbd199664),
	.w7(32'hbc4b74e5),
	.w8(32'h3d279171),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf90417),
	.w1(32'hbcbee4ea),
	.w2(32'h3a814020),
	.w3(32'hbcdfd17e),
	.w4(32'hbbbf0871),
	.w5(32'h3c474595),
	.w6(32'hbd71df0e),
	.w7(32'hbb600c15),
	.w8(32'h3c441e9e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdef450),
	.w1(32'h3cb003c1),
	.w2(32'h3c25c2f8),
	.w3(32'h3c23d1c6),
	.w4(32'hbcdbeb5d),
	.w5(32'h3cbed0e5),
	.w6(32'h3c00e482),
	.w7(32'h3c4f4446),
	.w8(32'h3d925760),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c890ae9),
	.w1(32'hbccd09e2),
	.w2(32'h3b8d7baf),
	.w3(32'hbc726f94),
	.w4(32'h3b0534b1),
	.w5(32'h3b5cd826),
	.w6(32'hbd13bebd),
	.w7(32'h3b5e13d0),
	.w8(32'h3beb53cc),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7581e9),
	.w1(32'hba7bfda3),
	.w2(32'h3b721058),
	.w3(32'h3becb8f3),
	.w4(32'hbc0b89ba),
	.w5(32'h3b08b0dd),
	.w6(32'h3c8ffd79),
	.w7(32'h3b4ebd3d),
	.w8(32'h3c2f9cd7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58f57e),
	.w1(32'hbc2c3bb3),
	.w2(32'hbb71ca56),
	.w3(32'h38c1eb62),
	.w4(32'hbc07df37),
	.w5(32'h3bee8f66),
	.w6(32'h3ac51840),
	.w7(32'h3b15aaeb),
	.w8(32'h3d0a9284),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad54a43),
	.w1(32'hbb674f40),
	.w2(32'hb7db2094),
	.w3(32'hbc4b9c15),
	.w4(32'hb9e951a4),
	.w5(32'hbc34962f),
	.w6(32'h3b650a82),
	.w7(32'hbb27c2df),
	.w8(32'hbc996cda),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d071545),
	.w1(32'hbce5cac0),
	.w2(32'hbc3f4d67),
	.w3(32'h3cb88a98),
	.w4(32'hbd3b78d3),
	.w5(32'hbd053b53),
	.w6(32'hbc7df628),
	.w7(32'hbd6e1c4d),
	.w8(32'hbd2c6954),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3a03f),
	.w1(32'hbb0f6b9b),
	.w2(32'hbbb69ca8),
	.w3(32'h3c12c59a),
	.w4(32'h3b2a678c),
	.w5(32'h3ca894d0),
	.w6(32'hbccebc3b),
	.w7(32'hba98f1c5),
	.w8(32'h3c59057c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7543ed),
	.w1(32'hbbd7c689),
	.w2(32'hbb11a891),
	.w3(32'hbbcab2ed),
	.w4(32'hbb2b1bbf),
	.w5(32'hbb7ca52d),
	.w6(32'hbc587dd2),
	.w7(32'h3a9e2c09),
	.w8(32'h3bbde294),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd65c2),
	.w1(32'hbaea254f),
	.w2(32'h3b8034c2),
	.w3(32'hbb17b217),
	.w4(32'h3a99769f),
	.w5(32'h3a9083f1),
	.w6(32'h3c47ad60),
	.w7(32'h3baa95d5),
	.w8(32'h3bc2f1e1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8db2b8),
	.w1(32'hb9883393),
	.w2(32'hbc1e2808),
	.w3(32'h3b251e07),
	.w4(32'hbb8357c3),
	.w5(32'h3bbb7080),
	.w6(32'h3a79d35e),
	.w7(32'hbc47e5d4),
	.w8(32'hbc8d1245),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32c6f6),
	.w1(32'h3c63bf7e),
	.w2(32'hbbbbb564),
	.w3(32'h3bee976b),
	.w4(32'hbac22283),
	.w5(32'hbc25d652),
	.w6(32'hbcb755e5),
	.w7(32'hbc3d6b28),
	.w8(32'h3bb3b08f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb565f7a),
	.w1(32'hbb750143),
	.w2(32'hbb56503f),
	.w3(32'h3bcea86d),
	.w4(32'h3b331f9d),
	.w5(32'hbce1d0a4),
	.w6(32'h3c3ca22e),
	.w7(32'h3bcab53b),
	.w8(32'hbd2727a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd505059),
	.w1(32'h3c62f855),
	.w2(32'h3bc350a9),
	.w3(32'h3ca0262d),
	.w4(32'h3bec27a6),
	.w5(32'h3ca9b416),
	.w6(32'h3d93e02f),
	.w7(32'h3b98cfa0),
	.w8(32'h3cc5ccf1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83df43),
	.w1(32'hbbf5f213),
	.w2(32'hbb876d5a),
	.w3(32'hbc07de17),
	.w4(32'h3a55e7f8),
	.w5(32'h3bde6d66),
	.w6(32'hbcb2ce73),
	.w7(32'hbb9ea479),
	.w8(32'hbbdbbfaf),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b657372),
	.w1(32'hbc11d991),
	.w2(32'h3be6de57),
	.w3(32'h3b59aa5b),
	.w4(32'hbc3dbc80),
	.w5(32'h3b8d5990),
	.w6(32'hbd04e718),
	.w7(32'hbb96a145),
	.w8(32'h3b340e95),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996917e),
	.w1(32'hbc62119a),
	.w2(32'hbc05d47a),
	.w3(32'hbc72df25),
	.w4(32'hbc3c2dfc),
	.w5(32'hbcaec0d3),
	.w6(32'hbd098471),
	.w7(32'h39961ddb),
	.w8(32'hbc05e409),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe6f14),
	.w1(32'h3c86bc99),
	.w2(32'hbc15e630),
	.w3(32'h3b2a7c2b),
	.w4(32'hba252dcf),
	.w5(32'hbc70b422),
	.w6(32'h3d3114d8),
	.w7(32'hbb67e7e6),
	.w8(32'hbce773a8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c47a4),
	.w1(32'hba7c925d),
	.w2(32'hbc270f94),
	.w3(32'h3bc2330e),
	.w4(32'hbc08495e),
	.w5(32'hbbad3460),
	.w6(32'hbb57eee6),
	.w7(32'h39aeead2),
	.w8(32'h3c24eb0b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cf5aa),
	.w1(32'hbc945434),
	.w2(32'h3b38ac30),
	.w3(32'hbc3efc15),
	.w4(32'hbca233b2),
	.w5(32'h3c333025),
	.w6(32'hbca5abd5),
	.w7(32'hbcb04c14),
	.w8(32'hbccf67e2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb655c78),
	.w1(32'h3c6f24e0),
	.w2(32'h3c7c849f),
	.w3(32'h3b27f9f4),
	.w4(32'hbc0e64c9),
	.w5(32'h3d155f09),
	.w6(32'h3c1a6ae4),
	.w7(32'hbc49ac66),
	.w8(32'h3d1dae27),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d42a12b),
	.w1(32'hbc92f508),
	.w2(32'hbbb811fb),
	.w3(32'hbcc8c534),
	.w4(32'hbb134f7d),
	.w5(32'hbc828c13),
	.w6(32'hbd5c25c3),
	.w7(32'h3b36058e),
	.w8(32'h3ca408a5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe77cd5),
	.w1(32'hbbbed196),
	.w2(32'h3ad0c54e),
	.w3(32'hbc08f75c),
	.w4(32'hbb220004),
	.w5(32'hbb68f310),
	.w6(32'h3c08ae87),
	.w7(32'hba846dca),
	.w8(32'h38eeb798),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5983),
	.w1(32'h39f42eb5),
	.w2(32'h3bc552eb),
	.w3(32'h3bcbf174),
	.w4(32'hbb83ddee),
	.w5(32'h3bdad634),
	.w6(32'hbafed6e8),
	.w7(32'hba9bf2c8),
	.w8(32'hbbef382e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3b6c6),
	.w1(32'h3c355f48),
	.w2(32'hbc5491d5),
	.w3(32'hbc1d7af7),
	.w4(32'hbc848530),
	.w5(32'h3ca79bb3),
	.w6(32'hbb746b76),
	.w7(32'hbc4826a0),
	.w8(32'h3d2cbd27),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caae37c),
	.w1(32'hbc7ef212),
	.w2(32'h3a54e954),
	.w3(32'hbc043f9a),
	.w4(32'h3b37a306),
	.w5(32'h3cd052f9),
	.w6(32'hbd0f4804),
	.w7(32'hbaf274b6),
	.w8(32'h3c893c08),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5089f6),
	.w1(32'hbc31ce42),
	.w2(32'h3c6c4ce7),
	.w3(32'h3b9bf261),
	.w4(32'h3a93db1f),
	.w5(32'hba7345dc),
	.w6(32'hbcdb3d05),
	.w7(32'h3bb8b02a),
	.w8(32'hbc5d2d7e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd05c13c),
	.w1(32'h3aa93672),
	.w2(32'hbc46fe72),
	.w3(32'hbc89c98b),
	.w4(32'hbc322914),
	.w5(32'hbc45c62b),
	.w6(32'h3bf2f3b0),
	.w7(32'hbc9f1189),
	.w8(32'hbcaab3eb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c320630),
	.w1(32'hbbf0fd9e),
	.w2(32'hbcb906f0),
	.w3(32'h3c863840),
	.w4(32'hbcfad43e),
	.w5(32'hbd13e17c),
	.w6(32'hbc4d3fa6),
	.w7(32'hbc4e932d),
	.w8(32'hbd05e10e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd37c97b),
	.w1(32'hbc661f10),
	.w2(32'hbc48d6ac),
	.w3(32'hbc829f43),
	.w4(32'hbb9c4369),
	.w5(32'hbc834059),
	.w6(32'h3c5df7be),
	.w7(32'h3b467e2f),
	.w8(32'h3ce29486),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc150247),
	.w1(32'h3c246a8d),
	.w2(32'hbbbb408c),
	.w3(32'hbc81d30f),
	.w4(32'hbcf887bc),
	.w5(32'h3bcd9327),
	.w6(32'h3d50e65b),
	.w7(32'hbcb76fb7),
	.w8(32'h3d5d4939),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1a6704),
	.w1(32'hbc3a265c),
	.w2(32'h3c952d76),
	.w3(32'hbb6b076c),
	.w4(32'h3b54caf0),
	.w5(32'hbc927b2c),
	.w6(32'hbca622f3),
	.w7(32'h3c935b63),
	.w8(32'hbd18cbcd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae3aca),
	.w1(32'hbbff3d8e),
	.w2(32'hbbce57a9),
	.w3(32'hba893e0f),
	.w4(32'hbb97455a),
	.w5(32'hbae3f0a9),
	.w6(32'h3cd59088),
	.w7(32'h3b4408e7),
	.w8(32'h3b8d6f26),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa119d),
	.w1(32'hbb892e81),
	.w2(32'hbc0929e8),
	.w3(32'h3b612fea),
	.w4(32'hba2a03b3),
	.w5(32'h3c74804b),
	.w6(32'hbb7e6ce9),
	.w7(32'h3a6a68cd),
	.w8(32'h3c9570bc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86af18),
	.w1(32'hbc2659ca),
	.w2(32'hbc1f0b59),
	.w3(32'h3c094b29),
	.w4(32'hbc41a960),
	.w5(32'hbd026b87),
	.w6(32'hbcdaa98c),
	.w7(32'hbbbcd7ea),
	.w8(32'hbceb592c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfaa84d),
	.w1(32'h3c380f21),
	.w2(32'h3ba87e5f),
	.w3(32'h3c43d8eb),
	.w4(32'hba81ce21),
	.w5(32'hba4e8492),
	.w6(32'h3d040a87),
	.w7(32'h3c636e7e),
	.w8(32'hbbbd940c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd32097),
	.w1(32'hbbf5415c),
	.w2(32'hbaa89f29),
	.w3(32'hbc1ebb7f),
	.w4(32'hbc961a1d),
	.w5(32'hbb036d7c),
	.w6(32'hbc87b254),
	.w7(32'hbc033e58),
	.w8(32'h3c72de3a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0705),
	.w1(32'h3aee180f),
	.w2(32'h3af71d9d),
	.w3(32'hbbb1d66a),
	.w4(32'hb9e62b32),
	.w5(32'hbb2eaf9b),
	.w6(32'h3b7c61ae),
	.w7(32'h3b8aad36),
	.w8(32'h3ba6301d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d83a2),
	.w1(32'hb9a1f3ea),
	.w2(32'hbb458481),
	.w3(32'h3bcf3892),
	.w4(32'hba91dd27),
	.w5(32'hbc34a1ab),
	.w6(32'hbabc0431),
	.w7(32'hbb05bbaa),
	.w8(32'h3c81ab2c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c065f02),
	.w1(32'hbc7b74b1),
	.w2(32'hb99b23a5),
	.w3(32'h3b42dad6),
	.w4(32'h3bba9094),
	.w5(32'hbcea98a7),
	.w6(32'hbc85a234),
	.w7(32'h3c456c6a),
	.w8(32'hbd1423b4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8894ec),
	.w1(32'hbaf42747),
	.w2(32'hbaa37d4a),
	.w3(32'h3c72e4c5),
	.w4(32'hb9bb78aa),
	.w5(32'hbc23f735),
	.w6(32'h3c79be07),
	.w7(32'h3bcfd38d),
	.w8(32'h3b5194fe),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1769d1),
	.w1(32'hbcb754e2),
	.w2(32'hba5b37ec),
	.w3(32'hbc76b075),
	.w4(32'hbb6dff8d),
	.w5(32'hbc6c901d),
	.w6(32'hbb846ba4),
	.w7(32'h3cdf60ae),
	.w8(32'hbcefa064),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92d3e8),
	.w1(32'h3b78f0e4),
	.w2(32'hbc424022),
	.w3(32'hbb6d937f),
	.w4(32'h3c10b32e),
	.w5(32'h3c76db7b),
	.w6(32'h3c215ddf),
	.w7(32'hbb0bd1f7),
	.w8(32'h3b44152f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801e82),
	.w1(32'h3c3ed17f),
	.w2(32'hbc96c372),
	.w3(32'h3cae3f5a),
	.w4(32'hbb5a4057),
	.w5(32'h3d1a9102),
	.w6(32'h3c6eacf0),
	.w7(32'h3bff0d9e),
	.w8(32'h3d6c322e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc767b6),
	.w1(32'hbc708fe1),
	.w2(32'h3ad77a7a),
	.w3(32'hbc21ccc5),
	.w4(32'hbc4567a7),
	.w5(32'hbc5dfe79),
	.w6(32'hbce95448),
	.w7(32'h3a5a9fed),
	.w8(32'h3c0616ad),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaef511),
	.w1(32'hbcdf502b),
	.w2(32'h3b09f825),
	.w3(32'hbc8bfa4e),
	.w4(32'h3b9ac1c1),
	.w5(32'hbc2148cb),
	.w6(32'h3c2cb0b3),
	.w7(32'h3bd2970f),
	.w8(32'hbba7bbcc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38c0c6),
	.w1(32'h3ce15c8b),
	.w2(32'hba6adc2b),
	.w3(32'h3c2ba82f),
	.w4(32'hbc2e053a),
	.w5(32'h3c563e14),
	.w6(32'h3d8f16c9),
	.w7(32'hbba98469),
	.w8(32'h3c27fef4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9294f),
	.w1(32'h3bc39be8),
	.w2(32'hbb837a21),
	.w3(32'hbbf039d7),
	.w4(32'hbc75210c),
	.w5(32'hbb1e642d),
	.w6(32'hbca105c7),
	.w7(32'hbc1e1162),
	.w8(32'hbbc32dc3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d326477),
	.w1(32'h3c3386e5),
	.w2(32'h3c1c6b6c),
	.w3(32'h3c088f0f),
	.w4(32'h3baacbbd),
	.w5(32'hbd214194),
	.w6(32'hbacc4192),
	.w7(32'h3b441aa0),
	.w8(32'hbcbf4520),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c539c),
	.w1(32'hbbf52763),
	.w2(32'h3c6b4519),
	.w3(32'hbc0e6898),
	.w4(32'hbc0024f9),
	.w5(32'h3cb41556),
	.w6(32'h3cbdbd4d),
	.w7(32'h3c2e4db1),
	.w8(32'h3c395c9e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceab2ce),
	.w1(32'hbc2db1e5),
	.w2(32'h3b11ceb2),
	.w3(32'hbc61c62a),
	.w4(32'hbb38b0d2),
	.w5(32'hbc0a33c3),
	.w6(32'hbbf6ca69),
	.w7(32'hbb01cbd7),
	.w8(32'hbcd8b384),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b035303),
	.w1(32'h3beaf842),
	.w2(32'hb9d82025),
	.w3(32'h3ce239c3),
	.w4(32'hbbcbe82e),
	.w5(32'h3c9847ad),
	.w6(32'h3ce92172),
	.w7(32'h3ac16d60),
	.w8(32'h3cc73c41),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27e608),
	.w1(32'hbb553f58),
	.w2(32'hbb8fd4fd),
	.w3(32'hbcabb041),
	.w4(32'hbbbf1911),
	.w5(32'hb98223dd),
	.w6(32'hbc9763df),
	.w7(32'h3b6ee17b),
	.w8(32'h3c116a96),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a42564f),
	.w1(32'hbbfe0e82),
	.w2(32'h3c034f4b),
	.w3(32'hbb4b08e9),
	.w4(32'hbba85f0d),
	.w5(32'hbcb5ea12),
	.w6(32'h3b4aa31f),
	.w7(32'hbc1766c0),
	.w8(32'hbd05b54e),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e584d),
	.w1(32'h3ba6c010),
	.w2(32'hbb09bffe),
	.w3(32'h3c78c433),
	.w4(32'h3ba3690f),
	.w5(32'hbcae4f04),
	.w6(32'h3c5f1b0f),
	.w7(32'h3be98208),
	.w8(32'hbaa48ec3),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90489e),
	.w1(32'hbcc5065c),
	.w2(32'hb7de8e00),
	.w3(32'h3b47b090),
	.w4(32'hb8bd8e5b),
	.w5(32'hb82f5672),
	.w6(32'hb9e7c776),
	.w7(32'hb88b0c2b),
	.w8(32'hb852f163),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c331ae7),
	.w1(32'h39a88985),
	.w2(32'hbae0032f),
	.w3(32'h390506b1),
	.w4(32'hbc02ecb5),
	.w5(32'hbc018d9f),
	.w6(32'h376254c9),
	.w7(32'hbbba10b3),
	.w8(32'hbb6db7bc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba171ef7),
	.w1(32'hbafce1ff),
	.w2(32'h3b40c50e),
	.w3(32'hbbb45898),
	.w4(32'hbbad2144),
	.w5(32'h3a29a044),
	.w6(32'hbbe16eef),
	.w7(32'hbbe66f08),
	.w8(32'h385e5a96),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba3402),
	.w1(32'h3987f27d),
	.w2(32'hb6a67247),
	.w3(32'hb9108826),
	.w4(32'h3994bae6),
	.w5(32'h38315f26),
	.w6(32'hb969cd29),
	.w7(32'h3902b59e),
	.w8(32'hb8ca4d8d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b702b2),
	.w1(32'h389a700f),
	.w2(32'h3919ee72),
	.w3(32'h38a69b42),
	.w4(32'h38b3756b),
	.w5(32'h39194a88),
	.w6(32'hb84a5c8d),
	.w7(32'h3819a8b8),
	.w8(32'h38c2757d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ec237),
	.w1(32'h3b0f01b5),
	.w2(32'h39a2d0ce),
	.w3(32'h3bccff86),
	.w4(32'h3b596675),
	.w5(32'h3a78e28a),
	.w6(32'hba08c75a),
	.w7(32'hbb402dae),
	.w8(32'hbbca4337),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6abb5),
	.w1(32'hbab5bdb6),
	.w2(32'hba6a77c8),
	.w3(32'hbba6cdfb),
	.w4(32'hbc1a18ae),
	.w5(32'hbbd4d81a),
	.w6(32'hbb765e1e),
	.w7(32'hbbd4d478),
	.w8(32'hbb55b9c1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf64aae),
	.w1(32'hbc0bb637),
	.w2(32'hbc5b323a),
	.w3(32'hbc84bc04),
	.w4(32'hbc76ff0c),
	.w5(32'hbc24dd77),
	.w6(32'hbb87fa23),
	.w7(32'hbbbb80e1),
	.w8(32'hbbf30fff),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a9be4),
	.w1(32'hba14749f),
	.w2(32'h3ae23a01),
	.w3(32'hbb8fa437),
	.w4(32'hbc5d712d),
	.w5(32'hbbc40ffc),
	.w6(32'hbb9c7a11),
	.w7(32'hbbe73ad7),
	.w8(32'h3a5341ea),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21fb18),
	.w1(32'h3c0fb535),
	.w2(32'h3b95bf4d),
	.w3(32'h3c635691),
	.w4(32'h3bc63c05),
	.w5(32'h3af495d4),
	.w6(32'h3c151b1c),
	.w7(32'h3bac3269),
	.w8(32'h39e44e0f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a84d10),
	.w1(32'hb9adf863),
	.w2(32'hb80017ae),
	.w3(32'hb83b2f1f),
	.w4(32'hb8d8ca1c),
	.w5(32'h3937b780),
	.w6(32'h380f7b17),
	.w7(32'hb9052efe),
	.w8(32'h383bfcac),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb722f012),
	.w1(32'hb86f8816),
	.w2(32'h38499001),
	.w3(32'h37bd00ed),
	.w4(32'hb6bed935),
	.w5(32'hb70ad3a2),
	.w6(32'h38217d2a),
	.w7(32'h379c675e),
	.w8(32'h37a491ec),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378857f5),
	.w1(32'h38bfdc62),
	.w2(32'hb7e4f5fb),
	.w3(32'h386ccdad),
	.w4(32'h38b614c0),
	.w5(32'h37de2cd6),
	.w6(32'hb83345b6),
	.w7(32'hb890aa5e),
	.w8(32'hb89166ee),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7e1c0),
	.w1(32'h3a61a598),
	.w2(32'h3a1b6581),
	.w3(32'h3a954d79),
	.w4(32'hba58f7d3),
	.w5(32'hba6c5b32),
	.w6(32'h3afc3a33),
	.w7(32'h39d933da),
	.w8(32'h3a85042c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3989f942),
	.w1(32'hb9de2504),
	.w2(32'hb9da9eda),
	.w3(32'h3b3a161b),
	.w4(32'h3a9925ad),
	.w5(32'h398086e0),
	.w6(32'h3b58a1c8),
	.w7(32'h3b0fbc7c),
	.w8(32'hb99192b0),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ab4ea),
	.w1(32'h39f376ed),
	.w2(32'h3a5d18ed),
	.w3(32'h3a865a2f),
	.w4(32'h3a212b7c),
	.w5(32'h3aab71e5),
	.w6(32'h39a69b67),
	.w7(32'h3a0eb2e1),
	.w8(32'h3a17264e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23db14),
	.w1(32'h3ba3a2e0),
	.w2(32'h3aa126bb),
	.w3(32'h3ae16953),
	.w4(32'h3b1fa9c2),
	.w5(32'h399cb472),
	.w6(32'h3a4c3580),
	.w7(32'h39c36352),
	.w8(32'hbb1aa01d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3f79f),
	.w1(32'hba6e0097),
	.w2(32'hb9c55d7d),
	.w3(32'hbb2e8430),
	.w4(32'hbb49c52e),
	.w5(32'hbab51daa),
	.w6(32'hbafd1884),
	.w7(32'hba5e0a83),
	.w8(32'h398753ef),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99244e0),
	.w1(32'h3a2cfc68),
	.w2(32'h3aa142d3),
	.w3(32'hbad647f7),
	.w4(32'h3a4a429f),
	.w5(32'h3ab74bca),
	.w6(32'hbaaa7d58),
	.w7(32'h3a22daa6),
	.w8(32'h3b183adb),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be23ace),
	.w1(32'h3ac2a6e6),
	.w2(32'hbae288d7),
	.w3(32'h3b0967ad),
	.w4(32'hbbae6c37),
	.w5(32'hbba4d93e),
	.w6(32'h3ab06b1e),
	.w7(32'hbb8bf54e),
	.w8(32'hbb6261df),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cfd2f),
	.w1(32'h3b420a85),
	.w2(32'h3b92f031),
	.w3(32'h3adf1778),
	.w4(32'h3aa384d3),
	.w5(32'h3b5adaa1),
	.w6(32'h3ba674ae),
	.w7(32'h3b8ec8cb),
	.w8(32'h3b9f1341),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb853953b),
	.w1(32'h37bd6a78),
	.w2(32'h375d4a9a),
	.w3(32'hb85814c8),
	.w4(32'h381184f5),
	.w5(32'h38ba6bf8),
	.w6(32'h382cc083),
	.w7(32'h3897bcbc),
	.w8(32'h381f4438),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d24d7),
	.w1(32'h3916c23c),
	.w2(32'h39828284),
	.w3(32'h395955f8),
	.w4(32'h390f9937),
	.w5(32'h3987de24),
	.w6(32'h396ef032),
	.w7(32'h38dcf41b),
	.w8(32'h396b341f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82158ff),
	.w1(32'hb87b0fbb),
	.w2(32'hb7f56127),
	.w3(32'h365540c2),
	.w4(32'hb8705ac4),
	.w5(32'h383508d7),
	.w6(32'hb857f5fe),
	.w7(32'hb92c4ab1),
	.w8(32'h36412f70),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7778546),
	.w1(32'hb9030775),
	.w2(32'hb8d22ce8),
	.w3(32'hb9489328),
	.w4(32'hb9a4b53b),
	.w5(32'hb9709a1a),
	.w6(32'hb95f60b2),
	.w7(32'hb991b002),
	.w8(32'hb99c8d38),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafed322),
	.w1(32'hb93e6f7e),
	.w2(32'h3a2a2c40),
	.w3(32'hbb57a01b),
	.w4(32'hba8b2ee2),
	.w5(32'h39877067),
	.w6(32'hbb6d24f2),
	.w7(32'hbaa5bffe),
	.w8(32'h3aa913d6),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5328f),
	.w1(32'h3ac06393),
	.w2(32'h3ad7dcf2),
	.w3(32'h3a6e02d3),
	.w4(32'h3a6d2a56),
	.w5(32'h3ab9a83d),
	.w6(32'h39c6cf74),
	.w7(32'h3a37cc35),
	.w8(32'h3aa06eef),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bd391),
	.w1(32'h3b60f89e),
	.w2(32'h3ae6cd97),
	.w3(32'h391c74de),
	.w4(32'h3b7d0b3a),
	.w5(32'h3b52d143),
	.w6(32'hbb1cc090),
	.w7(32'hba984cc4),
	.w8(32'hbb6335a4),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ef10f4),
	.w1(32'h3abb81ba),
	.w2(32'hb922558f),
	.w3(32'h3991debc),
	.w4(32'h3ab3be62),
	.w5(32'hb98a3cba),
	.w6(32'h397d9d0a),
	.w7(32'h3a77b79f),
	.w8(32'hba14c5a9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c871bb4),
	.w1(32'h3bca28ad),
	.w2(32'h3b696c88),
	.w3(32'h3b777230),
	.w4(32'hbb48c141),
	.w5(32'hbb91e6e5),
	.w6(32'hba9685f7),
	.w7(32'hbbaa9808),
	.w8(32'hbb832c35),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ea63e),
	.w1(32'h3b67fb0d),
	.w2(32'h3b133296),
	.w3(32'h3b336f97),
	.w4(32'h3b2096e2),
	.w5(32'h3af03b3c),
	.w6(32'h3ac29165),
	.w7(32'h3ae2fdfb),
	.w8(32'h3ac3d310),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa284f4),
	.w1(32'h3b58e020),
	.w2(32'h3ac1f307),
	.w3(32'h3acd62ff),
	.w4(32'h3b2250ad),
	.w5(32'h3a978f69),
	.w6(32'h3b1b058b),
	.w7(32'h3b3a50f9),
	.w8(32'h3a77a545),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b172504),
	.w1(32'h3b2b2e38),
	.w2(32'h39de904b),
	.w3(32'h3ae96b72),
	.w4(32'h3af3d14c),
	.w5(32'h38ab0c39),
	.w6(32'h3aaefb4d),
	.w7(32'h3aaa85fd),
	.w8(32'hb9f9aec1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8107d),
	.w1(32'hba2813ba),
	.w2(32'h3b92a9a0),
	.w3(32'hbb203894),
	.w4(32'h3b3f2297),
	.w5(32'h3bd3e32b),
	.w6(32'hbb1ba3ea),
	.w7(32'h3ae408ce),
	.w8(32'h3b92c37c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf244e),
	.w1(32'hbac69d4a),
	.w2(32'hbb3f7c89),
	.w3(32'hbb444084),
	.w4(32'hba94855f),
	.w5(32'hbaf93051),
	.w6(32'h3b4b562b),
	.w7(32'h3b0d1a98),
	.w8(32'h39211978),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a544a2b),
	.w1(32'h3aacced6),
	.w2(32'hbaedcc4d),
	.w3(32'hba7df69f),
	.w4(32'hb9649ce1),
	.w5(32'hbb1144d1),
	.w6(32'h373d93fd),
	.w7(32'h3a8494c3),
	.w8(32'hb9c9e0fd),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae52139),
	.w1(32'h3b9c81e7),
	.w2(32'h3b9407bb),
	.w3(32'h3aa04a14),
	.w4(32'h3b70db68),
	.w5(32'h3b5747df),
	.w6(32'h3a67a41a),
	.w7(32'h3b4fb8e0),
	.w8(32'h3b280464),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ecf9bb),
	.w1(32'hb9c94e73),
	.w2(32'hb880dfd8),
	.w3(32'hb832e066),
	.w4(32'hb9673d7a),
	.w5(32'hb8c40567),
	.w6(32'h39041b60),
	.w7(32'hb8ca385f),
	.w8(32'hb90fc81c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb812ebb0),
	.w1(32'hba0c0eea),
	.w2(32'h388a892d),
	.w3(32'hba8aa89a),
	.w4(32'hbae44aa9),
	.w5(32'hb9d281fb),
	.w6(32'hba1488e2),
	.w7(32'hba799f0e),
	.w8(32'hb9b88e61),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9947c6),
	.w1(32'h3ad9469d),
	.w2(32'h3a75972f),
	.w3(32'h3ae524e7),
	.w4(32'h3b0f0075),
	.w5(32'h3abc96b4),
	.w6(32'hb986d7d3),
	.w7(32'h39d92d9a),
	.w8(32'h3a7f94eb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a649d21),
	.w1(32'h3a83cec0),
	.w2(32'hba939327),
	.w3(32'h3ae1a9b9),
	.w4(32'h38baba9c),
	.w5(32'hbb1c2d71),
	.w6(32'h3a8396dd),
	.w7(32'hba124305),
	.w8(32'hbb585514),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b5122),
	.w1(32'hbad5dd7e),
	.w2(32'hbac36244),
	.w3(32'hba9773e6),
	.w4(32'hbb8878f0),
	.w5(32'hbb886c61),
	.w6(32'hba088a4f),
	.w7(32'hbb4a0d67),
	.w8(32'hbadb43b6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a468e1),
	.w1(32'h381ce5f8),
	.w2(32'h3824dd54),
	.w3(32'h37c0eb7c),
	.w4(32'h37064068),
	.w5(32'h380361b1),
	.w6(32'h377038a2),
	.w7(32'hb8999db4),
	.w8(32'h372defd3),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2538d),
	.w1(32'hb93f63d5),
	.w2(32'h3977a219),
	.w3(32'hb9926ca4),
	.w4(32'hb9e3e774),
	.w5(32'h395ce208),
	.w6(32'hb816dd4f),
	.w7(32'hb993c53e),
	.w8(32'h39c70924),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf7ae7),
	.w1(32'h3b58fa59),
	.w2(32'h3b89e3d1),
	.w3(32'h3b468b8b),
	.w4(32'h3ad6e8a1),
	.w5(32'h3ad2ba08),
	.w6(32'h3b5e18dd),
	.w7(32'h3a4eea69),
	.w8(32'hba2b381b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b5c5),
	.w1(32'h3ab36689),
	.w2(32'h3999be3b),
	.w3(32'h3b9deda9),
	.w4(32'h3b860a97),
	.w5(32'h3b801a06),
	.w6(32'h3b7e462b),
	.w7(32'h3b2a9abd),
	.w8(32'h3ae1d74d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b2a40),
	.w1(32'hba92ce80),
	.w2(32'hba2d4e35),
	.w3(32'hba3b6176),
	.w4(32'hba6b22b3),
	.w5(32'hba351a6b),
	.w6(32'hba25f145),
	.w7(32'hbac980a1),
	.w8(32'hbadd8d49),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa4f30),
	.w1(32'h39ec43cf),
	.w2(32'hb9bd42d3),
	.w3(32'h3b0f15a8),
	.w4(32'hba9a3419),
	.w5(32'hbb0038ac),
	.w6(32'h3aa6c9a0),
	.w7(32'hbaad72d3),
	.w8(32'hbaf4af85),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8283ef),
	.w1(32'hba4b1ce7),
	.w2(32'h3afab8e2),
	.w3(32'hbb691667),
	.w4(32'h3a5ca66b),
	.w5(32'h3b5dfb22),
	.w6(32'hbb2af39e),
	.w7(32'h3aceadae),
	.w8(32'h3b806ca5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a84a5e),
	.w1(32'h35182660),
	.w2(32'hb9c073a7),
	.w3(32'hbb31fd04),
	.w4(32'hba38ccca),
	.w5(32'hbb1d0b5f),
	.w6(32'hbad26793),
	.w7(32'hb98c4f49),
	.w8(32'h3a4a9d7e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e7dcc),
	.w1(32'hbaa4c7b7),
	.w2(32'h3a8d518f),
	.w3(32'hbab53ad6),
	.w4(32'h39b58b85),
	.w5(32'h3b1ebaf0),
	.w6(32'h39426a1b),
	.w7(32'h3aafe1a0),
	.w8(32'h3b22251b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77dcf1),
	.w1(32'hb9b02266),
	.w2(32'hbb09dabc),
	.w3(32'hb9e6d91e),
	.w4(32'hbb76f1aa),
	.w5(32'hbb72d456),
	.w6(32'hbb2a4a6f),
	.w7(32'hbb8c0893),
	.w8(32'hbb0f9821),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule