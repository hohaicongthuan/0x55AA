module layer_8_featuremap_101(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27dcb2),
	.w1(32'hbb5ea8d4),
	.w2(32'hbbd8aac0),
	.w3(32'h3b2ada4a),
	.w4(32'hbc3aadcc),
	.w5(32'h3c194fec),
	.w6(32'hbc7a4849),
	.w7(32'hbc98d44a),
	.w8(32'h3c44c25b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb679a),
	.w1(32'hbc4cb264),
	.w2(32'hbb1922dd),
	.w3(32'h3bb84146),
	.w4(32'h3c1f3b98),
	.w5(32'hb713e98c),
	.w6(32'hbbbd2499),
	.w7(32'h3a1d77a2),
	.w8(32'hbb3b3c6e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b20c),
	.w1(32'h3b9d95ea),
	.w2(32'h3c2fe1cc),
	.w3(32'hba5734d0),
	.w4(32'hbaa95228),
	.w5(32'hbc7448fe),
	.w6(32'hbbbe4d0b),
	.w7(32'hbbeab11b),
	.w8(32'h3c5b969f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccd69f0),
	.w1(32'hba291297),
	.w2(32'hbc77c7b5),
	.w3(32'h3c040649),
	.w4(32'hbbb7554f),
	.w5(32'hbcc1cda6),
	.w6(32'hbc5e8596),
	.w7(32'h3cc7ac31),
	.w8(32'h3c65cc52),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14f60e),
	.w1(32'h3b96ccc3),
	.w2(32'h3b22c465),
	.w3(32'hbc3a3b89),
	.w4(32'hb9ec5227),
	.w5(32'hbb813e19),
	.w6(32'h3a87ee63),
	.w7(32'hbc9e7fe2),
	.w8(32'hbccf9a8a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f2e1d),
	.w1(32'h3c467744),
	.w2(32'h3bf6134e),
	.w3(32'hbc1ed863),
	.w4(32'h3c27fb0e),
	.w5(32'hbbef9428),
	.w6(32'hbc1d6496),
	.w7(32'h3c510aba),
	.w8(32'h3d235931),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5699),
	.w1(32'h3c0e8400),
	.w2(32'h3c13a3f4),
	.w3(32'hbc55741f),
	.w4(32'h3c13a833),
	.w5(32'hba9eb904),
	.w6(32'hbc973f38),
	.w7(32'h3c3e069d),
	.w8(32'hbb720f09),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcb586),
	.w1(32'hbb80432c),
	.w2(32'h3b9884f4),
	.w3(32'hbb7a3c16),
	.w4(32'hbad19ae3),
	.w5(32'hbb000b17),
	.w6(32'h3bb0cc4b),
	.w7(32'hbbd626c8),
	.w8(32'hba21959d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01fb2a),
	.w1(32'h3b160aec),
	.w2(32'hbc57db96),
	.w3(32'h39e22e35),
	.w4(32'hbc0159bd),
	.w5(32'hba77b7ad),
	.w6(32'hbc486f4d),
	.w7(32'h3c3c44b4),
	.w8(32'h3c6e776a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99bc02),
	.w1(32'hbba2c3b8),
	.w2(32'h3caf17ad),
	.w3(32'hbb076de1),
	.w4(32'hbb236e6e),
	.w5(32'h3c877e8f),
	.w6(32'hbc79a089),
	.w7(32'hbc4f5418),
	.w8(32'hbdafbf12),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f447a),
	.w1(32'h3bb1f7fb),
	.w2(32'h3a9b314e),
	.w3(32'h3c11be9d),
	.w4(32'hbcddd3f7),
	.w5(32'hbcfed275),
	.w6(32'hbd19c09e),
	.w7(32'h3ba36c08),
	.w8(32'h3d1185e0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14ad4),
	.w1(32'hbc13e069),
	.w2(32'hbbecb526),
	.w3(32'hbc42eb3f),
	.w4(32'hbb133f68),
	.w5(32'hbb89d227),
	.w6(32'hbcfa25e3),
	.w7(32'hbbdd8d52),
	.w8(32'hbca519c1),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec010e),
	.w1(32'hbbab0ae2),
	.w2(32'h3b4471d9),
	.w3(32'hbb3f6f3a),
	.w4(32'h395f7959),
	.w5(32'h3b309a7f),
	.w6(32'hbbec4207),
	.w7(32'hbb7f91b0),
	.w8(32'hba91ddd4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ee945),
	.w1(32'hba20a562),
	.w2(32'hba8a5faa),
	.w3(32'hba93f2c6),
	.w4(32'hba172b7b),
	.w5(32'hba7d13c2),
	.w6(32'hbab2bcd9),
	.w7(32'hba40ac1e),
	.w8(32'hbac9d5d6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879c3fa),
	.w1(32'h3814b037),
	.w2(32'hb880ecb8),
	.w3(32'hb8883a9b),
	.w4(32'hb8aa9803),
	.w5(32'hb8a86010),
	.w6(32'hb877dd64),
	.w7(32'hb8baa1aa),
	.w8(32'hb8e4462f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6d9dd),
	.w1(32'hbad3d508),
	.w2(32'hbb0b2038),
	.w3(32'hbb2fb815),
	.w4(32'hbae53a81),
	.w5(32'hbab41349),
	.w6(32'hba631c55),
	.w7(32'hba4ee0b2),
	.w8(32'hba7c99bb),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6aec61),
	.w1(32'hbb0a4643),
	.w2(32'hbb16683d),
	.w3(32'hbb8eeb17),
	.w4(32'hbb4677f0),
	.w5(32'hbb7018b7),
	.w6(32'hbb4650cb),
	.w7(32'hbb13a486),
	.w8(32'hbb29790d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39396193),
	.w1(32'h3a378b2a),
	.w2(32'h3a100928),
	.w3(32'hbbb8c036),
	.w4(32'hbb5a9f61),
	.w5(32'hb95909f5),
	.w6(32'hbb812d54),
	.w7(32'hbb9f9944),
	.w8(32'h3aee0b74),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2f124),
	.w1(32'hbcdf634b),
	.w2(32'hbcbaa390),
	.w3(32'hbc9b4c60),
	.w4(32'hbca06d12),
	.w5(32'hbc44f974),
	.w6(32'hbbeeb3d5),
	.w7(32'hbbf7eec4),
	.w8(32'hbb269613),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc120652),
	.w1(32'hbc81601d),
	.w2(32'hbc6ded6f),
	.w3(32'hbc4049e9),
	.w4(32'hbc927037),
	.w5(32'hbc72b96f),
	.w6(32'h3b484597),
	.w7(32'h3ad29de1),
	.w8(32'h3a0b021e),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf00c9d),
	.w1(32'h3ac42f9c),
	.w2(32'hbb4657e9),
	.w3(32'h3b134faa),
	.w4(32'h3bd71157),
	.w5(32'h3b4d9872),
	.w6(32'hbb109610),
	.w7(32'h3b1e55cc),
	.w8(32'h3ada5657),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00cd34),
	.w1(32'h3c45a026),
	.w2(32'h3ba0c872),
	.w3(32'h3af2df52),
	.w4(32'h3bf9966d),
	.w5(32'h3b786fb7),
	.w6(32'h3a889046),
	.w7(32'h3b8af313),
	.w8(32'h3a13013e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95680a),
	.w1(32'hbc72b20f),
	.w2(32'hbc9cb776),
	.w3(32'h3a85d28e),
	.w4(32'hbc9dc506),
	.w5(32'hbc8b1e95),
	.w6(32'h3c538c4e),
	.w7(32'h3a95d6a6),
	.w8(32'hba8936aa),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636f9e),
	.w1(32'h3a1113cb),
	.w2(32'h3a2ce9d2),
	.w3(32'hbb075e43),
	.w4(32'hbbb09dfd),
	.w5(32'hbb803484),
	.w6(32'hbb2dacb1),
	.w7(32'hbb984aac),
	.w8(32'hbb2965c0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb461f6),
	.w1(32'hbba5214f),
	.w2(32'hbc0299df),
	.w3(32'hbb68e0e4),
	.w4(32'hbb469bf7),
	.w5(32'hbbfc46fc),
	.w6(32'hbc17c4a9),
	.w7(32'hbb9aa8bd),
	.w8(32'hbc25f883),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c750c),
	.w1(32'hbb2b9eb6),
	.w2(32'hbb55e70a),
	.w3(32'h3aefb543),
	.w4(32'hbb80ab87),
	.w5(32'hbb674e4a),
	.w6(32'h3c0f2829),
	.w7(32'h3b76928f),
	.w8(32'h3b7ab95e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2bf9b),
	.w1(32'h3960dae8),
	.w2(32'h38b11c08),
	.w3(32'h3b2a6228),
	.w4(32'h39e3a5a5),
	.w5(32'hb965a5b9),
	.w6(32'h3b3f6045),
	.w7(32'h3aa1cb7f),
	.w8(32'h39d0f95c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5bad19),
	.w1(32'hbd2951e2),
	.w2(32'hbd8a2e87),
	.w3(32'hbd7aa383),
	.w4(32'hbd5bcfea),
	.w5(32'hbd36278d),
	.w6(32'hbc17bfa0),
	.w7(32'h3d192d54),
	.w8(32'h3beb1ab6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb406f21),
	.w1(32'hbb8e8d09),
	.w2(32'hbba5e7a0),
	.w3(32'hbb447917),
	.w4(32'hbb7c3ed0),
	.w5(32'hbb82a1fd),
	.w6(32'h3a28d6b7),
	.w7(32'h3989cbe2),
	.w8(32'hb9c553b0),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba430060),
	.w1(32'hb8399249),
	.w2(32'hbb0c5558),
	.w3(32'hba1652ef),
	.w4(32'hb9e9e380),
	.w5(32'hbb026405),
	.w6(32'hbacd891e),
	.w7(32'hbacce31e),
	.w8(32'hbb268f9d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2081bb),
	.w1(32'h3c304d5e),
	.w2(32'h3bd3cf69),
	.w3(32'h3c11d3eb),
	.w4(32'h3c2323c5),
	.w5(32'h3bb20845),
	.w6(32'h3bcccc13),
	.w7(32'h3bafce97),
	.w8(32'h3b040db7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9598cb0),
	.w1(32'hbabfd559),
	.w2(32'hba8bb047),
	.w3(32'hba7e2d81),
	.w4(32'h395d593d),
	.w5(32'h3a7ffe82),
	.w6(32'h3a9e15b8),
	.w7(32'h3a84f419),
	.w8(32'h3b0b6804),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d7c509),
	.w1(32'hb943983b),
	.w2(32'hb84ea60c),
	.w3(32'hb823da84),
	.w4(32'hb924f605),
	.w5(32'h3693a1d1),
	.w6(32'hb8ce83eb),
	.w7(32'hb9966918),
	.w8(32'hb8881eb6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb719f895),
	.w1(32'hb90b0331),
	.w2(32'h38d00942),
	.w3(32'hb7f7452d),
	.w4(32'hb945923a),
	.w5(32'hb67c29b2),
	.w6(32'h362b8b0d),
	.w7(32'hb8bf22dd),
	.w8(32'h38ee5c4f),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c61f4),
	.w1(32'h3babfaf2),
	.w2(32'h3b3ddad9),
	.w3(32'h3aac472c),
	.w4(32'h3a541d4d),
	.w5(32'hbaa33baa),
	.w6(32'h39c3ce45),
	.w7(32'h3a65099d),
	.w8(32'hba5e133e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba222cbd),
	.w1(32'hbbdf3009),
	.w2(32'hbbeb32ea),
	.w3(32'hbaf662d5),
	.w4(32'hbbb233e6),
	.w5(32'hbb697962),
	.w6(32'h38944390),
	.w7(32'hbb7a307e),
	.w8(32'hbb2a659f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7d8c6),
	.w1(32'hbab11cbd),
	.w2(32'hbaa0784b),
	.w3(32'hba1a4ae0),
	.w4(32'hba8468cb),
	.w5(32'hbab4a5da),
	.w6(32'h38fa47f8),
	.w7(32'h39676a06),
	.w8(32'hba44f6f9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8da3bf),
	.w1(32'h3b20303c),
	.w2(32'h39fbd59c),
	.w3(32'h3b8a78d8),
	.w4(32'h3b8e9a7a),
	.w5(32'h3b7aa0ed),
	.w6(32'h3bcd53b8),
	.w7(32'h3be26afa),
	.w8(32'h3b9eb4b3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916b55a),
	.w1(32'hb9b5d426),
	.w2(32'h39212e68),
	.w3(32'hb8e61a47),
	.w4(32'hba2d90fc),
	.w5(32'hb91e35b5),
	.w6(32'hb6a32325),
	.w7(32'hb9d8312f),
	.w8(32'h3908b40d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39060a88),
	.w1(32'h3a480193),
	.w2(32'h39e2790c),
	.w3(32'hb9c08c8e),
	.w4(32'hb9a9d61b),
	.w5(32'hb9a90f92),
	.w6(32'h39f307af),
	.w7(32'hba1d6647),
	.w8(32'hba4fa6b3),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc100d76),
	.w1(32'hbbdaee4a),
	.w2(32'hbc32c295),
	.w3(32'hbbd15ae9),
	.w4(32'hbb8b85be),
	.w5(32'hbc0b3967),
	.w6(32'hbb7de727),
	.w7(32'hbb588eb3),
	.w8(32'hbc0a76bb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa915ee),
	.w1(32'h3ab737e4),
	.w2(32'h3b725387),
	.w3(32'h397c1dbc),
	.w4(32'h3a2ccad8),
	.w5(32'h3b6e0c63),
	.w6(32'h38a7f968),
	.w7(32'h3afb5f19),
	.w8(32'h3b846323),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f811),
	.w1(32'hba130eb6),
	.w2(32'hb93f5866),
	.w3(32'hb9f82587),
	.w4(32'hb989617d),
	.w5(32'hb93ee719),
	.w6(32'hba0fa668),
	.w7(32'hb9cf00b3),
	.w8(32'h398cdf03),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570194),
	.w1(32'hbb8bb910),
	.w2(32'hbbbdbece),
	.w3(32'hbb591007),
	.w4(32'hbb40782a),
	.w5(32'hbb89a559),
	.w6(32'hbb3a9818),
	.w7(32'hbb41befe),
	.w8(32'hbb49f2ca),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15c6d0),
	.w1(32'hb93577ab),
	.w2(32'hbb2c3997),
	.w3(32'hba86d2b1),
	.w4(32'hbb5ffa4b),
	.w5(32'hba0ed893),
	.w6(32'h3b284ee8),
	.w7(32'h3b0a3475),
	.w8(32'h3b7c81a0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6d415),
	.w1(32'h3a04de44),
	.w2(32'h3a8f13fd),
	.w3(32'hbb0d704a),
	.w4(32'h39e82006),
	.w5(32'h3a32d410),
	.w6(32'hbb1f5bb2),
	.w7(32'hb9182b1e),
	.w8(32'hba5bdc14),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39241bfa),
	.w1(32'h368e6d0b),
	.w2(32'h38233289),
	.w3(32'hb8812c6b),
	.w4(32'hb72852e8),
	.w5(32'h38c92260),
	.w6(32'h3872cb0e),
	.w7(32'hb826d7b0),
	.w8(32'hb87fd766),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79fa04),
	.w1(32'hbc461087),
	.w2(32'hbc540de5),
	.w3(32'hbc1fcfde),
	.w4(32'hbc7165ff),
	.w5(32'hbc084ebb),
	.w6(32'hbb01af4d),
	.w7(32'hbb2c2efe),
	.w8(32'h3ab0a817),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87ef50),
	.w1(32'hbb1a37d5),
	.w2(32'hbaa8971a),
	.w3(32'hbba315cf),
	.w4(32'hbb4399f5),
	.w5(32'hbb066d98),
	.w6(32'hbb803f24),
	.w7(32'hbacdeba1),
	.w8(32'hba0494b1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d820d),
	.w1(32'hba9ef7b0),
	.w2(32'h39ca7e12),
	.w3(32'h3a89fb6a),
	.w4(32'hba8be8d9),
	.w5(32'h3aa21f83),
	.w6(32'h3b637c74),
	.w7(32'h3a430aa8),
	.w8(32'h3ae30f1e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1c021),
	.w1(32'h3c324d1a),
	.w2(32'h3babb687),
	.w3(32'h3be945c2),
	.w4(32'h3c539890),
	.w5(32'h3c0767d7),
	.w6(32'h3c074701),
	.w7(32'h3c3d29b5),
	.w8(32'h3c0bf032),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31aed2),
	.w1(32'hbc94080a),
	.w2(32'hbcc00af9),
	.w3(32'hbca785c2),
	.w4(32'hbcd567c7),
	.w5(32'hbcd40e83),
	.w6(32'h3ab2db3f),
	.w7(32'hbb27ece1),
	.w8(32'h3aa3e8b0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85289f),
	.w1(32'hbbb67340),
	.w2(32'hbb8176de),
	.w3(32'hbc39ac26),
	.w4(32'hbc5b37ce),
	.w5(32'hbc2c4c2e),
	.w6(32'hba0ea13a),
	.w7(32'hbaa94a89),
	.w8(32'hba84d3e3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82d6e8),
	.w1(32'hbb9d3893),
	.w2(32'hbb350f9d),
	.w3(32'hbb91ca18),
	.w4(32'hbbaf6539),
	.w5(32'hbad399c8),
	.w6(32'hbb980f49),
	.w7(32'hbb97a867),
	.w8(32'hbafe2c98),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dab67f),
	.w1(32'hb9224b08),
	.w2(32'hb92fceeb),
	.w3(32'hb7f0a7ee),
	.w4(32'hb9787fcd),
	.w5(32'hb92b0be6),
	.w6(32'h3632b495),
	.w7(32'hb8cd3f2f),
	.w8(32'hb93ad13e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c9adb),
	.w1(32'hbbbb0611),
	.w2(32'hbbc61c5e),
	.w3(32'hbb8e88b6),
	.w4(32'hbb94fe48),
	.w5(32'h386cbd36),
	.w6(32'hb97e067d),
	.w7(32'h39798f3e),
	.w8(32'h3b883dcb),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f3bb),
	.w1(32'h3b80d042),
	.w2(32'h3b2ce3cc),
	.w3(32'hbb0ed713),
	.w4(32'hba8dd052),
	.w5(32'hbae78b24),
	.w6(32'h3aa7243d),
	.w7(32'h3ba5d28d),
	.w8(32'h3b696e62),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856048),
	.w1(32'hba3064a3),
	.w2(32'hbadd59b8),
	.w3(32'hbbc6d9f9),
	.w4(32'hbbe1f879),
	.w5(32'hbbda8a1e),
	.w6(32'hbbaf4544),
	.w7(32'hbb86e065),
	.w8(32'hba7174db),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c9e09),
	.w1(32'hbb6fc1a0),
	.w2(32'hbba09740),
	.w3(32'hbbc5be0c),
	.w4(32'hbba3537c),
	.w5(32'hbbaa9d33),
	.w6(32'hbb73109d),
	.w7(32'hbabf355b),
	.w8(32'hba689df6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c182c),
	.w1(32'hbab7d2fd),
	.w2(32'hbb281403),
	.w3(32'hbb1afa4b),
	.w4(32'hba917c93),
	.w5(32'hbb3521db),
	.w6(32'hbae8b15f),
	.w7(32'hb9f0c796),
	.w8(32'hbae4a708),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73086b),
	.w1(32'hbb36b28e),
	.w2(32'hbb3d6a47),
	.w3(32'hbb5d7a25),
	.w4(32'hbb4bbc2a),
	.w5(32'hbb84f6b0),
	.w6(32'hbb4fc82d),
	.w7(32'hbb0c13b7),
	.w8(32'hbb408368),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08c8c9),
	.w1(32'h39ee9a41),
	.w2(32'hb8271a7e),
	.w3(32'hba25d5bd),
	.w4(32'hba5f1d2b),
	.w5(32'hba6a618f),
	.w6(32'h3a3e1b07),
	.w7(32'h39e105f7),
	.w8(32'hb81f8f73),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f4c27),
	.w1(32'hbb4dcb2d),
	.w2(32'hbbce6537),
	.w3(32'hbb87d728),
	.w4(32'hbb521e0a),
	.w5(32'hbbae8b58),
	.w6(32'h3a4c5aec),
	.w7(32'h3b4822e2),
	.w8(32'h39b7062e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e273ca),
	.w1(32'hbb3f9bf2),
	.w2(32'hbb5f1e14),
	.w3(32'hbb209150),
	.w4(32'hbbe739b5),
	.w5(32'hbbf32f52),
	.w6(32'hbb7c32e2),
	.w7(32'hbbfabdbf),
	.w8(32'hbb888005),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b8b4b),
	.w1(32'h3a90b622),
	.w2(32'h3a1f5a10),
	.w3(32'h3b1b9f50),
	.w4(32'hb9a4b8a8),
	.w5(32'hba20ca07),
	.w6(32'h3af660b2),
	.w7(32'hb9b061d4),
	.w8(32'h39cb8716),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8937fd),
	.w1(32'hba197423),
	.w2(32'hb9ca4ab9),
	.w3(32'hba32d568),
	.w4(32'hbb4becec),
	.w5(32'hbb2e0d75),
	.w6(32'h3a8e30a8),
	.w7(32'hba9ca270),
	.w8(32'hb95a9e2b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d408b),
	.w1(32'hbb1e10b8),
	.w2(32'hbb718985),
	.w3(32'hb9f0f83e),
	.w4(32'hbb06ecc8),
	.w5(32'hbb138778),
	.w6(32'hbb968ae1),
	.w7(32'hbb3312c1),
	.w8(32'hb986d769),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3810a0),
	.w1(32'hb9d42198),
	.w2(32'hbabd84e0),
	.w3(32'h398a5949),
	.w4(32'h393c2c20),
	.w5(32'hba533827),
	.w6(32'h3af6ff95),
	.w7(32'h3a54d401),
	.w8(32'hb9f75e86),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba857ab9),
	.w1(32'hba147258),
	.w2(32'hba98f4eb),
	.w3(32'h38383ea9),
	.w4(32'hb99d0fcd),
	.w5(32'hb9bd827e),
	.w6(32'h3ad1d827),
	.w7(32'h3aeeb80b),
	.w8(32'h3ab532cf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56471f),
	.w1(32'hbc28fbb9),
	.w2(32'hbca967ab),
	.w3(32'hbbc45aef),
	.w4(32'hbc90b406),
	.w5(32'hbcb92b01),
	.w6(32'hb861a181),
	.w7(32'hbb82697b),
	.w8(32'hbb771e4f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4509a),
	.w1(32'h3ac8ad5b),
	.w2(32'h3a9739dd),
	.w3(32'h3ad0026c),
	.w4(32'h3abf658f),
	.w5(32'h3a69aa54),
	.w6(32'h3ab764d9),
	.w7(32'h3a96bf24),
	.w8(32'h3a3e802e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb566d4f),
	.w1(32'hbb856925),
	.w2(32'hbb225c26),
	.w3(32'hbbf270b0),
	.w4(32'hbbf167e4),
	.w5(32'hbb893af5),
	.w6(32'hbb6a3851),
	.w7(32'hba9632f0),
	.w8(32'h3af5e2cb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a905806),
	.w1(32'h3a6c5701),
	.w2(32'h3a2b3dae),
	.w3(32'h3ab1972b),
	.w4(32'h3a42ad6f),
	.w5(32'h3a3f3e72),
	.w6(32'h3ad67f3d),
	.w7(32'h3a7ed11a),
	.w8(32'h3a397cc9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab8a0),
	.w1(32'hb987cb25),
	.w2(32'hbb88b9b1),
	.w3(32'hbad36da4),
	.w4(32'h3b2d861c),
	.w5(32'hba980819),
	.w6(32'hbaa50656),
	.w7(32'h3b11b096),
	.w8(32'h3a6ea6c5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b9fbcd),
	.w1(32'hb7389b26),
	.w2(32'hb84e7858),
	.w3(32'h39521855),
	.w4(32'hb8c6c9aa),
	.w5(32'h380b8d4e),
	.w6(32'hb823e7aa),
	.w7(32'h381cc4b6),
	.w8(32'hb8b60715),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada16cb),
	.w1(32'hbb85a0e6),
	.w2(32'hbb5082fb),
	.w3(32'h3a9ccb36),
	.w4(32'hb98a57a4),
	.w5(32'hbabdfa32),
	.w6(32'h3bd335f3),
	.w7(32'h3b8f7de6),
	.w8(32'h39cccfd4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c35294),
	.w1(32'hb9ac678d),
	.w2(32'hb8c78485),
	.w3(32'hb83453c7),
	.w4(32'hba0cd4c3),
	.w5(32'h3b9be1c3),
	.w6(32'h39551626),
	.w7(32'h3a154f20),
	.w8(32'h3ba41a70),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9065a9),
	.w1(32'hbc49eb22),
	.w2(32'hbc881ad3),
	.w3(32'hbb570cb5),
	.w4(32'hbc447ad4),
	.w5(32'hbc012e79),
	.w6(32'h3a1cc391),
	.w7(32'hbbcf9b39),
	.w8(32'h3ade5682),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d069b),
	.w1(32'hbad63088),
	.w2(32'hbbe5fd20),
	.w3(32'hbb50610d),
	.w4(32'hbbee0f7d),
	.w5(32'hbc4dce61),
	.w6(32'hbb2ecdf1),
	.w7(32'hbb8cec33),
	.w8(32'hbc064ccd),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36da9c),
	.w1(32'hbb72c9f1),
	.w2(32'h3c3186df),
	.w3(32'hbbb7a06e),
	.w4(32'hbc4dbdd7),
	.w5(32'h3b4f4add),
	.w6(32'hbbaa3e9c),
	.w7(32'hbc087ceb),
	.w8(32'hbc36ecc8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7915cd),
	.w1(32'hbc823333),
	.w2(32'hbc612032),
	.w3(32'hba1e00f1),
	.w4(32'hbbf72f4a),
	.w5(32'hbb29c70d),
	.w6(32'hbca00af0),
	.w7(32'hbb6e3470),
	.w8(32'hbb730edd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a7cb6),
	.w1(32'h3c6b622a),
	.w2(32'hbc8a8c32),
	.w3(32'hbb3e41b3),
	.w4(32'hbca1574e),
	.w5(32'hbccac4d7),
	.w6(32'h3c86ded6),
	.w7(32'hbc0111d8),
	.w8(32'hbc95be9f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7409b6),
	.w1(32'hbb84a0b2),
	.w2(32'hbbe4e27f),
	.w3(32'hbc366264),
	.w4(32'hbab158e0),
	.w5(32'hbb375636),
	.w6(32'hbb358773),
	.w7(32'h3bbef01e),
	.w8(32'h3c289f98),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc663c10),
	.w1(32'h3bda2ff7),
	.w2(32'hbb287b47),
	.w3(32'hbcad012a),
	.w4(32'hba48b3f5),
	.w5(32'hbc832ce7),
	.w6(32'hbbc3cbfa),
	.w7(32'h3c5d6b6f),
	.w8(32'hbc1015ab),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ac8ce),
	.w1(32'hbc531fb2),
	.w2(32'hbc933591),
	.w3(32'hbd1952aa),
	.w4(32'hbc927afb),
	.w5(32'hbbe02b71),
	.w6(32'hbcf5d060),
	.w7(32'h3c386865),
	.w8(32'h3c6f329b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ecc9f),
	.w1(32'hbcb17a24),
	.w2(32'h3a822060),
	.w3(32'hbb8794b6),
	.w4(32'h3ab3b467),
	.w5(32'hbc366b2d),
	.w6(32'hbaa7cec3),
	.w7(32'h3c6f62b0),
	.w8(32'h3c0d9786),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8577fa),
	.w1(32'hbc124984),
	.w2(32'h3c870ea9),
	.w3(32'h3b083ca6),
	.w4(32'hbb5e7df8),
	.w5(32'hbb83a621),
	.w6(32'hbbad1b76),
	.w7(32'h3c815ea3),
	.w8(32'h3bcb2015),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c404571),
	.w1(32'hbc18af00),
	.w2(32'hbbca478f),
	.w3(32'hbc9a84ea),
	.w4(32'hbc05d98c),
	.w5(32'hbc3b5305),
	.w6(32'hbcb8d94e),
	.w7(32'hbc229186),
	.w8(32'hbc19db5b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc33b897),
	.w1(32'h3b30db39),
	.w2(32'h3c3d8385),
	.w3(32'hbb551ecc),
	.w4(32'h3b02a1e7),
	.w5(32'hbbbfaf00),
	.w6(32'h3bcba163),
	.w7(32'h3badc201),
	.w8(32'hbc07ddde),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf4b465),
	.w1(32'hba51f0cb),
	.w2(32'hbc2a285e),
	.w3(32'hbbb2ebfe),
	.w4(32'hbc33939d),
	.w5(32'h3c66c982),
	.w6(32'hbb4b659b),
	.w7(32'hbc73d15a),
	.w8(32'hbc52813a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bb2b2),
	.w1(32'h3cb5bed5),
	.w2(32'hba4caf30),
	.w3(32'h3be04097),
	.w4(32'h3b7679d3),
	.w5(32'hbbe79e7d),
	.w6(32'h3c63e3d4),
	.w7(32'h3c27265c),
	.w8(32'h3b31a8bb),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dbdc0),
	.w1(32'hbb7ababe),
	.w2(32'h3bdfcfd2),
	.w3(32'hbc32106a),
	.w4(32'h3cca0cef),
	.w5(32'h3ae98115),
	.w6(32'hbc9495f9),
	.w7(32'h3cde6a59),
	.w8(32'h3c51672d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7c0f),
	.w1(32'hbcadc1aa),
	.w2(32'hbc123426),
	.w3(32'hbc9f7dbb),
	.w4(32'h3b6a8978),
	.w5(32'h3c05a5a2),
	.w6(32'hbcd70ae7),
	.w7(32'h3ae1fe36),
	.w8(32'h3be165f6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b567f),
	.w1(32'hbaed5563),
	.w2(32'h3c10fe2e),
	.w3(32'h3ad29844),
	.w4(32'hbbb839c7),
	.w5(32'h3a227927),
	.w6(32'h3b60869e),
	.w7(32'h3b99b64f),
	.w8(32'h3b053c8c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb95752),
	.w1(32'h3c18ab35),
	.w2(32'h3a2dd47a),
	.w3(32'h379c5762),
	.w4(32'hbb09b03a),
	.w5(32'h3b92fd3c),
	.w6(32'h3b68e4d4),
	.w7(32'hbaf27f80),
	.w8(32'h3ba05761),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed92e),
	.w1(32'h3c691de6),
	.w2(32'h3d3688fb),
	.w3(32'h3c1bd8e1),
	.w4(32'h3c083b25),
	.w5(32'hbc037721),
	.w6(32'h3c484f5a),
	.w7(32'h3d29fd56),
	.w8(32'h3c8d728e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c806d43),
	.w1(32'hbd99c627),
	.w2(32'hbceb3464),
	.w3(32'hbd3b7305),
	.w4(32'hbc06949c),
	.w5(32'h3bdc5208),
	.w6(32'hbd3d31bf),
	.w7(32'hbc1f6be4),
	.w8(32'h39bb3e33),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc785421),
	.w1(32'h3d11ddb3),
	.w2(32'hbb9a2da8),
	.w3(32'h3cf35d82),
	.w4(32'hba933c98),
	.w5(32'hb9a21652),
	.w6(32'h3d0f32d7),
	.w7(32'h3ad7e9b0),
	.w8(32'hbbfb9d87),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8134e8),
	.w1(32'h3ce2cb21),
	.w2(32'hbc015b66),
	.w3(32'h3c95b24b),
	.w4(32'hbb9156e3),
	.w5(32'h3bf774c2),
	.w6(32'h3d262a88),
	.w7(32'hbc49d612),
	.w8(32'hba89d75a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b671d50),
	.w1(32'h3c85d380),
	.w2(32'hba9f9b04),
	.w3(32'h3cacc766),
	.w4(32'hbc3a175d),
	.w5(32'h3b3a3293),
	.w6(32'h3cac19c3),
	.w7(32'hbbee28e4),
	.w8(32'h3c8805bd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b855d49),
	.w1(32'hbc78bbc9),
	.w2(32'h3cf8c448),
	.w3(32'h3a864ddf),
	.w4(32'h3c08443d),
	.w5(32'hbb904be8),
	.w6(32'h3ba0e871),
	.w7(32'h3cd84928),
	.w8(32'hbbf89d6c),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb431c5),
	.w1(32'hbce4a1cf),
	.w2(32'hbc023227),
	.w3(32'hbbec6b10),
	.w4(32'hbc59b7dc),
	.w5(32'hbc31560d),
	.w6(32'hbcecb1c1),
	.w7(32'hbb630f44),
	.w8(32'hbc0719ee),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bec4e),
	.w1(32'h3bbdc290),
	.w2(32'h3c9092f4),
	.w3(32'hbbf99e79),
	.w4(32'h3bfc6745),
	.w5(32'h3b4eaaba),
	.w6(32'h3b9ec54f),
	.w7(32'h3cbc5c87),
	.w8(32'hbc0a1d32),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6bcadb),
	.w1(32'hbc8b13e6),
	.w2(32'h3b0af55c),
	.w3(32'hbcbc9e68),
	.w4(32'hb7d6bf24),
	.w5(32'hb9ad6538),
	.w6(32'hbcde6317),
	.w7(32'h3b8efbbc),
	.w8(32'hbbca2649),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffe0b2),
	.w1(32'hbc254d5b),
	.w2(32'h3bd83fbf),
	.w3(32'hbb499b08),
	.w4(32'h399f4728),
	.w5(32'hbba6f7ac),
	.w6(32'hbc9b3767),
	.w7(32'hbb308763),
	.w8(32'hbc5bd1b9),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb954296),
	.w1(32'hbc620586),
	.w2(32'hbb756c17),
	.w3(32'hbcc57563),
	.w4(32'hbc6924cd),
	.w5(32'hbce5f9b3),
	.w6(32'hbc8e14ec),
	.w7(32'h3c334516),
	.w8(32'hbbab89d6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e85f2),
	.w1(32'hbc8c9236),
	.w2(32'hbcca6055),
	.w3(32'hbb60f884),
	.w4(32'h3a6b649d),
	.w5(32'h3ba221bc),
	.w6(32'hbc87e444),
	.w7(32'hbae29236),
	.w8(32'hba41f4b3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6d412),
	.w1(32'h3cc8c711),
	.w2(32'hb9b666ea),
	.w3(32'h3c2d06bb),
	.w4(32'hbb845a1f),
	.w5(32'h3b76952c),
	.w6(32'h3d134b9b),
	.w7(32'h3a1f7c4e),
	.w8(32'h3bed91de),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc07be6),
	.w1(32'h3bda8d13),
	.w2(32'h3c15db8b),
	.w3(32'h3bce2c7e),
	.w4(32'h3bf64d18),
	.w5(32'h3bcb51b4),
	.w6(32'h3be7b0d1),
	.w7(32'h3bf05243),
	.w8(32'h3adf0816),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc194b91),
	.w1(32'hba96ca32),
	.w2(32'h3bfbbccc),
	.w3(32'hbc4e9490),
	.w4(32'h3bca60c6),
	.w5(32'h3bda8df1),
	.w6(32'hbc0066e5),
	.w7(32'h3c48f4cf),
	.w8(32'h3c056064),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e670f),
	.w1(32'hbbe24689),
	.w2(32'hbc3a14d1),
	.w3(32'h3c432ab2),
	.w4(32'h3ce01b9d),
	.w5(32'h3cb8f95e),
	.w6(32'hbc0d1c7d),
	.w7(32'h3c4ea6bf),
	.w8(32'h3c771d0d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5a77f),
	.w1(32'hbca62951),
	.w2(32'h3b4a19fb),
	.w3(32'hbc47e3ad),
	.w4(32'hbb0b6eb6),
	.w5(32'h3c9881b0),
	.w6(32'hbc35ec1b),
	.w7(32'hbc06b736),
	.w8(32'h3c29e2ec),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48f73c),
	.w1(32'h3d0a9e89),
	.w2(32'h3ce348db),
	.w3(32'h3be5382a),
	.w4(32'h3c659d23),
	.w5(32'hbb998842),
	.w6(32'h3cec6c83),
	.w7(32'h3cf33da2),
	.w8(32'h3c0e5a93),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb535c0),
	.w1(32'hbd2b7cf6),
	.w2(32'h3d45c466),
	.w3(32'hbce238ab),
	.w4(32'h3cacc9da),
	.w5(32'hbcb4af43),
	.w6(32'hbd3c4540),
	.w7(32'h3d436969),
	.w8(32'h3abe41da),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce560a),
	.w1(32'hbd52e21c),
	.w2(32'hbbe0ded8),
	.w3(32'hbd904701),
	.w4(32'hbc1b602d),
	.w5(32'hbc8623b7),
	.w6(32'hbd91aa9e),
	.w7(32'hbcaffac0),
	.w8(32'hbc24f292),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c496f59),
	.w1(32'h3cf88cba),
	.w2(32'hbb396f82),
	.w3(32'h3c1677ed),
	.w4(32'hbbaf9418),
	.w5(32'hba5e0ad3),
	.w6(32'h3d17f381),
	.w7(32'h3973e60b),
	.w8(32'h3bdc1885),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbe182),
	.w1(32'hbcc54bf4),
	.w2(32'hbc7c1c8f),
	.w3(32'h3ac48be7),
	.w4(32'hbb7337c4),
	.w5(32'hbcaab6f4),
	.w6(32'hbba56579),
	.w7(32'hbc163b6c),
	.w8(32'h3ba17ec2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c097109),
	.w1(32'hbbced44e),
	.w2(32'hbb9fec0a),
	.w3(32'hbc821bf1),
	.w4(32'hbb1a54c9),
	.w5(32'h3ab373f2),
	.w6(32'hbbcc16f0),
	.w7(32'h394f1cbe),
	.w8(32'h3bd9ed2b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc46a19),
	.w1(32'h3b92ee74),
	.w2(32'h3b5cfe30),
	.w3(32'h3b55ed75),
	.w4(32'h3bd8afc0),
	.w5(32'hbc1083ed),
	.w6(32'h3bc336af),
	.w7(32'h3c31e11c),
	.w8(32'hbb04bb81),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7adaf1),
	.w1(32'hbc656140),
	.w2(32'h3c4651ab),
	.w3(32'hbca741bf),
	.w4(32'h3baa23f1),
	.w5(32'hbbb02fc4),
	.w6(32'hbc9f11b6),
	.w7(32'h3ba69c0c),
	.w8(32'hba7d07b5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8328f),
	.w1(32'hbb1f1300),
	.w2(32'h3b7d796f),
	.w3(32'hbc36ca12),
	.w4(32'hbba26a14),
	.w5(32'hbc2047f1),
	.w6(32'hbc076215),
	.w7(32'h3c0905da),
	.w8(32'hbb18511e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb867bc66),
	.w1(32'hbbfe3197),
	.w2(32'hbcf3c480),
	.w3(32'hbbb43682),
	.w4(32'hbcaafadb),
	.w5(32'hbbfd409e),
	.w6(32'h3ac345d4),
	.w7(32'hbce22821),
	.w8(32'hbc9983b7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3407f3),
	.w1(32'h3d1ff446),
	.w2(32'hba844765),
	.w3(32'h3c47c420),
	.w4(32'hbb184253),
	.w5(32'h3b2d2ec5),
	.w6(32'h3cfca37f),
	.w7(32'hb83297f6),
	.w8(32'h3bdfd471),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7479a),
	.w1(32'h3c1dc58d),
	.w2(32'h3c862128),
	.w3(32'h3bd792b0),
	.w4(32'h3cae7a1e),
	.w5(32'h3c23f5ba),
	.w6(32'h3bcd2ad8),
	.w7(32'h3bc1fe05),
	.w8(32'h3beaa7fb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55a26a),
	.w1(32'hba91e552),
	.w2(32'hbc26c813),
	.w3(32'hbb2bc202),
	.w4(32'h3c0e3b67),
	.w5(32'hbba0991c),
	.w6(32'hbb863eb3),
	.w7(32'h3bc2eaf4),
	.w8(32'h3c2a68f6),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c274eff),
	.w1(32'h3c56db7e),
	.w2(32'hb9e111e7),
	.w3(32'h3bacdae9),
	.w4(32'hbb596c69),
	.w5(32'hbb966ee8),
	.w6(32'h3c8854b8),
	.w7(32'h3b3d0e01),
	.w8(32'hbb8c5194),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc177aa5),
	.w1(32'hbbc0a5a7),
	.w2(32'h3a3cbf5a),
	.w3(32'hbb9095b9),
	.w4(32'h3c2be1e7),
	.w5(32'h3c0e4293),
	.w6(32'hba2dcf62),
	.w7(32'hba98f027),
	.w8(32'hbb553bd7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37850a),
	.w1(32'h3b210f4d),
	.w2(32'hba48b6b1),
	.w3(32'hbbfc1f69),
	.w4(32'hba468708),
	.w5(32'hba9e18b2),
	.w6(32'hbbc03422),
	.w7(32'h3b0bd36e),
	.w8(32'hbc409dfb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule