module layer_8_featuremap_178(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb663f52),
	.w1(32'hbb4c5230),
	.w2(32'hbc01fc71),
	.w3(32'hbb3e1cfb),
	.w4(32'hbbd3681b),
	.w5(32'hbc17248c),
	.w6(32'h3b9ce56e),
	.w7(32'hbb9cc9ef),
	.w8(32'hbb9209f2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6a1ad),
	.w1(32'h3b1b2ec6),
	.w2(32'hbb1f8fe4),
	.w3(32'hbc4b9bb1),
	.w4(32'h3b1dc3d4),
	.w5(32'hbb6587b6),
	.w6(32'h3b26c0a2),
	.w7(32'hbab17e7f),
	.w8(32'hbb4113e2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f131a),
	.w1(32'hbbda4b99),
	.w2(32'hbcbaf919),
	.w3(32'hbbba2f79),
	.w4(32'hba972918),
	.w5(32'hbc92e986),
	.w6(32'h3be1612e),
	.w7(32'hbbe3f62d),
	.w8(32'hbc3d84f2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9efc03),
	.w1(32'hbc5dd871),
	.w2(32'hbccaa3a6),
	.w3(32'hbc908e14),
	.w4(32'hbc83086d),
	.w5(32'hbcc3ad91),
	.w6(32'h3b0b5880),
	.w7(32'hbbff2fa7),
	.w8(32'hbbea5afc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc54e668),
	.w1(32'h3aaaeca9),
	.w2(32'h39f5e17a),
	.w3(32'hbbe02145),
	.w4(32'h39eb8c09),
	.w5(32'h38f85f65),
	.w6(32'h3ade2d6b),
	.w7(32'h3b7aac70),
	.w8(32'h3b32b03f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a972896),
	.w1(32'hb9956922),
	.w2(32'h3bd3ab4d),
	.w3(32'h3a90532d),
	.w4(32'h3b9ef43c),
	.w5(32'h3c2c201f),
	.w6(32'hbb51c4f3),
	.w7(32'h3bb9c6bf),
	.w8(32'hbaabb3e8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea6236),
	.w1(32'hb9f51c45),
	.w2(32'hbb17f376),
	.w3(32'h3b83e476),
	.w4(32'hbb1e0f48),
	.w5(32'hb96ddf68),
	.w6(32'hbb5ff5f1),
	.w7(32'hb811a0a3),
	.w8(32'hbb540b25),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b976b30),
	.w1(32'h3c285f8c),
	.w2(32'h3c2a3f9d),
	.w3(32'h3b5ab5f3),
	.w4(32'h3a177da5),
	.w5(32'hbc05fd0e),
	.w6(32'h3c0a2275),
	.w7(32'h3c2e9322),
	.w8(32'hbc0afe63),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc349cb7),
	.w1(32'h3bd87202),
	.w2(32'h3993bff8),
	.w3(32'hbc37786b),
	.w4(32'h3bae8391),
	.w5(32'hba938c27),
	.w6(32'h3baab14f),
	.w7(32'hb942f250),
	.w8(32'hb98f6d9f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b291aa7),
	.w1(32'hba6b45f7),
	.w2(32'hbcaeea6c),
	.w3(32'h3a147bf9),
	.w4(32'h3bccaa9c),
	.w5(32'hbc872cc8),
	.w6(32'h379b3c81),
	.w7(32'hbc72379f),
	.w8(32'hbc6579bd),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b2847),
	.w1(32'h3b8b73b4),
	.w2(32'hbb857b9f),
	.w3(32'hbb2bc564),
	.w4(32'hbbda35ec),
	.w5(32'hbc57b49d),
	.w6(32'h3c0a0021),
	.w7(32'h3b64d888),
	.w8(32'hbb8e6e6f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104856),
	.w1(32'hb9af219a),
	.w2(32'h3abaa380),
	.w3(32'hbc47f6d3),
	.w4(32'h3b3bac00),
	.w5(32'h3a8d94e5),
	.w6(32'hbb136c5f),
	.w7(32'hb963a183),
	.w8(32'hb9246aad),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bcfdc),
	.w1(32'hbb97ee64),
	.w2(32'hbd0289e3),
	.w3(32'h3aaf5145),
	.w4(32'hbbad0217),
	.w5(32'hbcc9ee8c),
	.w6(32'h3bd4c952),
	.w7(32'hbc4d309e),
	.w8(32'hbc3a5715),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcea7917),
	.w1(32'hbc91c388),
	.w2(32'hbca0347c),
	.w3(32'hbc282f4c),
	.w4(32'hbc27c917),
	.w5(32'hbc7e016a),
	.w6(32'hbc2a0015),
	.w7(32'hbc8c6ba6),
	.w8(32'hbc88965b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9ee913),
	.w1(32'h3adc3d2b),
	.w2(32'hbab95d0d),
	.w3(32'hbc6bb328),
	.w4(32'h3addf6de),
	.w5(32'h37add036),
	.w6(32'h3a38ed88),
	.w7(32'hbaf00849),
	.w8(32'hba8e1c09),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0294d1),
	.w1(32'hbb1df17b),
	.w2(32'h3bdc4291),
	.w3(32'h39e05b64),
	.w4(32'hba44a8e1),
	.w5(32'h3bef9d44),
	.w6(32'h3bd3753c),
	.w7(32'h3b011f81),
	.w8(32'h3bfa6df7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c75268e),
	.w1(32'h3a189e80),
	.w2(32'h3c552290),
	.w3(32'h3c765985),
	.w4(32'h3b609219),
	.w5(32'h3bbf18d5),
	.w6(32'h3bc36760),
	.w7(32'hbb9b9612),
	.w8(32'hb9fffe0c),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26f42f),
	.w1(32'hbb89d2bc),
	.w2(32'hbc86ef59),
	.w3(32'h3c09acb8),
	.w4(32'h3a51c49c),
	.w5(32'hbc5ad0f3),
	.w6(32'hbc1b4fd2),
	.w7(32'hbbdc1535),
	.w8(32'h3b313564),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc092688),
	.w1(32'hbc074321),
	.w2(32'h3bf961fc),
	.w3(32'hbbb03f83),
	.w4(32'h3a0b106e),
	.w5(32'h3c34a0ca),
	.w6(32'hbbbc15d1),
	.w7(32'hbb1c3a7a),
	.w8(32'hbb0f7ae8),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d7b5e),
	.w1(32'hbabf8b5f),
	.w2(32'hba1e23db),
	.w3(32'hba1896b3),
	.w4(32'hbb409e29),
	.w5(32'hba8a93ec),
	.w6(32'hb9167eb8),
	.w7(32'hbb164561),
	.w8(32'h39eb28bb),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034c86),
	.w1(32'hbbf8bdc7),
	.w2(32'hbc742305),
	.w3(32'hb9b09353),
	.w4(32'hbae62864),
	.w5(32'hbc50ee19),
	.w6(32'hbc229506),
	.w7(32'h3aee63db),
	.w8(32'h3adf301e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76270d),
	.w1(32'h3c28f8c9),
	.w2(32'h3b3b6ca8),
	.w3(32'hbbf43613),
	.w4(32'h3bf44e3b),
	.w5(32'h3bacc921),
	.w6(32'h3bbd62e0),
	.w7(32'h3b8caa48),
	.w8(32'hbbc2cac0),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e911a),
	.w1(32'h3c8de86f),
	.w2(32'h3c8ad69d),
	.w3(32'h3a99e2bf),
	.w4(32'h3c8eb2e5),
	.w5(32'h3c89fdfe),
	.w6(32'h3b64b281),
	.w7(32'h3c67d0b2),
	.w8(32'h3bcaf1ca),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968cdd4),
	.w1(32'h3bb13264),
	.w2(32'h3a99b992),
	.w3(32'h3b761458),
	.w4(32'h3acc0989),
	.w5(32'hbb0b0e49),
	.w6(32'h3bd8a4c7),
	.w7(32'hbbbe74c4),
	.w8(32'hbb4d2269),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea139),
	.w1(32'h3b871a06),
	.w2(32'h3b439c7f),
	.w3(32'h3b5ccd5b),
	.w4(32'h3bfe4218),
	.w5(32'h3bc23542),
	.w6(32'h3bd7e5bf),
	.w7(32'h3bfbaed0),
	.w8(32'h3c0425e3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7967bfe),
	.w1(32'h3be3d6e7),
	.w2(32'hbac34832),
	.w3(32'h3c0882f2),
	.w4(32'h3b5b1058),
	.w5(32'hbb224315),
	.w6(32'h3c331954),
	.w7(32'h3afa4ff6),
	.w8(32'hbc27966b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f8be9),
	.w1(32'h3bbc0698),
	.w2(32'hbc2e1301),
	.w3(32'hbc0e78d0),
	.w4(32'hbbd85efc),
	.w5(32'hbb993767),
	.w6(32'h3b60f4f0),
	.w7(32'hbab49941),
	.w8(32'hba806093),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17641b),
	.w1(32'hbc7d5d47),
	.w2(32'hbd130a53),
	.w3(32'h3ba3f0f9),
	.w4(32'hbc4b2a5d),
	.w5(32'hbcdfb0a0),
	.w6(32'h3ca0509b),
	.w7(32'h3b1ab16c),
	.w8(32'hbaf88a7f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac90f7),
	.w1(32'h3ba08e93),
	.w2(32'h3b47d506),
	.w3(32'hbbea79ad),
	.w4(32'h3bc9eb84),
	.w5(32'hbb35d334),
	.w6(32'h3c393108),
	.w7(32'h3bb995f8),
	.w8(32'h39eda273),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ee3e8),
	.w1(32'h3c021f34),
	.w2(32'h3b99ba5c),
	.w3(32'hb8fbc1b2),
	.w4(32'h3ab5ab2c),
	.w5(32'h3b229c52),
	.w6(32'h3b95a3cb),
	.w7(32'h3bd76b4b),
	.w8(32'hba80c5c9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba5096),
	.w1(32'h3badc416),
	.w2(32'hba297264),
	.w3(32'hbb994206),
	.w4(32'h3baa1d9a),
	.w5(32'hbb130af6),
	.w6(32'h3bb5d86f),
	.w7(32'h3bb8e5a9),
	.w8(32'h3bf968b1),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39841ee5),
	.w1(32'h3ae672ff),
	.w2(32'h39781ed8),
	.w3(32'h3b0abd6f),
	.w4(32'h3c2b6029),
	.w5(32'hbb78c15f),
	.w6(32'hba648840),
	.w7(32'h3be95c24),
	.w8(32'hbb1bb90a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf06c3c),
	.w1(32'hbc219249),
	.w2(32'hbc9295fa),
	.w3(32'hbc1e1aca),
	.w4(32'hbc285ee2),
	.w5(32'hbc0cbc7c),
	.w6(32'hbb981d66),
	.w7(32'hbc1ae2a6),
	.w8(32'hbbed7681),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfcdb95),
	.w1(32'h3c4c9865),
	.w2(32'h3cacbc3e),
	.w3(32'hbc06b592),
	.w4(32'h3c57c145),
	.w5(32'h3c8a83d7),
	.w6(32'hb9c9b766),
	.w7(32'h3c40413f),
	.w8(32'h3c5b122a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b408),
	.w1(32'hbb251659),
	.w2(32'hbb525e22),
	.w3(32'h3c44e330),
	.w4(32'h3aae1b80),
	.w5(32'h3ba981c4),
	.w6(32'h3a305ec9),
	.w7(32'h3ac1b7a3),
	.w8(32'h3b0620f3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b8ca2),
	.w1(32'h3c8d101f),
	.w2(32'h3cdec4e0),
	.w3(32'h3bded54d),
	.w4(32'h3c5e8669),
	.w5(32'h3c842dc0),
	.w6(32'h3c497c94),
	.w7(32'h3ccd32d6),
	.w8(32'h3c4df5ee),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce3a6b0),
	.w1(32'hbac03cf1),
	.w2(32'hbb723186),
	.w3(32'h3cab12d0),
	.w4(32'hbb801f93),
	.w5(32'hbb85ef16),
	.w6(32'h3b4d4d12),
	.w7(32'h3a4e81b0),
	.w8(32'h3a8a5db4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaed56),
	.w1(32'h399d258b),
	.w2(32'hbb9019f3),
	.w3(32'h3b22d225),
	.w4(32'h3b515e04),
	.w5(32'hba832742),
	.w6(32'hbaccbe97),
	.w7(32'hbbc0f174),
	.w8(32'h3a48f30c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d8fb1),
	.w1(32'h3c3858e2),
	.w2(32'h3d028733),
	.w3(32'h3b91bd0a),
	.w4(32'h3b6d87dd),
	.w5(32'h3c99e425),
	.w6(32'h3b8385f9),
	.w7(32'h3c6b48fe),
	.w8(32'h3c7922dd),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0778b),
	.w1(32'hbc4e6ea5),
	.w2(32'hbcc62ae5),
	.w3(32'h3c9d92b4),
	.w4(32'hbc4ac3e7),
	.w5(32'hbc48b299),
	.w6(32'h3b6edb32),
	.w7(32'hbb89e6d0),
	.w8(32'hbc049f80),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2457),
	.w1(32'h3b274b0c),
	.w2(32'hbba1f22f),
	.w3(32'h3a618fed),
	.w4(32'h3af92e43),
	.w5(32'hbba113c7),
	.w6(32'h3b8c3953),
	.w7(32'hbb72aa8f),
	.w8(32'hbac392c5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92ba5b),
	.w1(32'hbaff6f19),
	.w2(32'hbb88a4e5),
	.w3(32'hbae53239),
	.w4(32'hbb9bedf0),
	.w5(32'hbbbd348a),
	.w6(32'hbc1523e3),
	.w7(32'h3a9a5c80),
	.w8(32'h3bc7568c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394874f2),
	.w1(32'h398eede9),
	.w2(32'h3b42d579),
	.w3(32'hbbe61d03),
	.w4(32'h3a83a100),
	.w5(32'h3ae8ad12),
	.w6(32'h3a4e4ffe),
	.w7(32'h3bd5f325),
	.w8(32'hbb6d08df),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b1751),
	.w1(32'hbc23c000),
	.w2(32'hbcb71b49),
	.w3(32'hbb334418),
	.w4(32'hbc253a12),
	.w5(32'hbc95aa7f),
	.w6(32'hbbf11dae),
	.w7(32'hbc505aea),
	.w8(32'hbc21cfcc),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc432220),
	.w1(32'hbae2908b),
	.w2(32'h3c5b9e81),
	.w3(32'hbbeead47),
	.w4(32'hbc59a718),
	.w5(32'h3c0b4e63),
	.w6(32'hbb91b8f9),
	.w7(32'h3b3af1af),
	.w8(32'hbae143db),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ddd59),
	.w1(32'hbad8a98b),
	.w2(32'hbb1f22bd),
	.w3(32'h3b88440c),
	.w4(32'hbb18ba87),
	.w5(32'hbb375e03),
	.w6(32'h3b4a54da),
	.w7(32'h3a365e84),
	.w8(32'hbbc5b701),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ca3c9),
	.w1(32'hbb00c4d7),
	.w2(32'hbc008ba7),
	.w3(32'hbbd3f468),
	.w4(32'hbac08a58),
	.w5(32'hbc1b0c89),
	.w6(32'hbae082a8),
	.w7(32'hbb1f8ff3),
	.w8(32'hbbf56ec1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc257340),
	.w1(32'h3b535cd3),
	.w2(32'hbc150adc),
	.w3(32'hbc8090a4),
	.w4(32'h3b412ee2),
	.w5(32'hbc014244),
	.w6(32'h3c59fe7f),
	.w7(32'hbb1a5d2b),
	.w8(32'hbaab32b0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11eb9b),
	.w1(32'hbc040896),
	.w2(32'hbc9daa61),
	.w3(32'h3ac4c209),
	.w4(32'hbc0ecfe5),
	.w5(32'hbcc450a8),
	.w6(32'h3ba8a8e9),
	.w7(32'hbc5d9701),
	.w8(32'hbc002eb2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc966d00),
	.w1(32'hbbf927b7),
	.w2(32'hbc1e61c7),
	.w3(32'hbaab1504),
	.w4(32'hbab0314a),
	.w5(32'hbc1f89ba),
	.w6(32'hbbcf9115),
	.w7(32'hbb460771),
	.w8(32'hbc2aa740),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0686e),
	.w1(32'h3aaeffdc),
	.w2(32'hbbc96fed),
	.w3(32'hbc88e985),
	.w4(32'h3b11c00f),
	.w5(32'hbb6a2369),
	.w6(32'h39fc6c71),
	.w7(32'hbb740033),
	.w8(32'h3b28a010),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8b5fb),
	.w1(32'h3bcb1e7e),
	.w2(32'h3b909a68),
	.w3(32'h3a38aa96),
	.w4(32'h3b39e7af),
	.w5(32'h3a69a720),
	.w6(32'hbb538ba5),
	.w7(32'h39af16dc),
	.w8(32'hbbe0639f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e887dc),
	.w1(32'h3aebbab4),
	.w2(32'hbb673635),
	.w3(32'hbb6b4034),
	.w4(32'h3b617541),
	.w5(32'hbb3099dc),
	.w6(32'hb940cb16),
	.w7(32'hbba1ecd5),
	.w8(32'hbb4fd78c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13f9b7),
	.w1(32'h3bcc65b3),
	.w2(32'h3c33270a),
	.w3(32'h39869b3c),
	.w4(32'h3aaf4bb8),
	.w5(32'h3b82219a),
	.w6(32'h3bc433ad),
	.w7(32'h3c5cf9d3),
	.w8(32'hbc1d8918),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2e95f),
	.w1(32'hb7c92a1b),
	.w2(32'hbc88941f),
	.w3(32'h3beef54b),
	.w4(32'hbc117a0c),
	.w5(32'hbbba2c46),
	.w6(32'hbbd92fcf),
	.w7(32'hbc768b8e),
	.w8(32'hbc01b21c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a758d6b),
	.w1(32'h3bf74810),
	.w2(32'hbc9c97d8),
	.w3(32'h3b7bc1ef),
	.w4(32'h3c3491a8),
	.w5(32'hbc0a4f60),
	.w6(32'h3c7596ba),
	.w7(32'h3b2c1a71),
	.w8(32'h3b1e6e5e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb947f7f),
	.w1(32'h3c4a6f04),
	.w2(32'h3c86b07f),
	.w3(32'hbb26a908),
	.w4(32'h3ba4a591),
	.w5(32'h3cb03ad7),
	.w6(32'h3c04dbcc),
	.w7(32'h3ba98a17),
	.w8(32'h3be8d269),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43d5ab),
	.w1(32'hbb39cc03),
	.w2(32'hbb9c9e1e),
	.w3(32'h3baa9c5e),
	.w4(32'hbb58f277),
	.w5(32'hbb875158),
	.w6(32'h3b0f1010),
	.w7(32'hbb2e0941),
	.w8(32'hbb84d422),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ba419),
	.w1(32'hba2a34d3),
	.w2(32'hbb520310),
	.w3(32'h3b01fe5a),
	.w4(32'hba791e7f),
	.w5(32'hbb038732),
	.w6(32'hbb336b80),
	.w7(32'hbb7ebad7),
	.w8(32'hbb4c10c9),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec6d2f),
	.w1(32'h3c51ea90),
	.w2(32'h3c5e62d0),
	.w3(32'hbb0a8f42),
	.w4(32'h3c69e2c1),
	.w5(32'h3c7a690b),
	.w6(32'h3aafb72f),
	.w7(32'h3bbd8add),
	.w8(32'h3bafbe17),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c702702),
	.w1(32'hbaafb7bf),
	.w2(32'hbbf33ea8),
	.w3(32'h3bb2bc0b),
	.w4(32'hbaf0bc30),
	.w5(32'hbc160673),
	.w6(32'h3c458fc3),
	.w7(32'h3b7f4e53),
	.w8(32'hbb011845),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689d77),
	.w1(32'h3b387af7),
	.w2(32'h3abe40aa),
	.w3(32'hbc627e05),
	.w4(32'h3af89e75),
	.w5(32'hbac7f335),
	.w6(32'hbb9a7731),
	.w7(32'h3b7ff731),
	.w8(32'h3bb8d693),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc761b3),
	.w1(32'h3b47b7ea),
	.w2(32'h3c443d55),
	.w3(32'hbb649a98),
	.w4(32'hb7b84db0),
	.w5(32'h3c35daa9),
	.w6(32'hbb61b56a),
	.w7(32'h3ad62838),
	.w8(32'h3b3683b9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5243b3),
	.w1(32'hbc08b069),
	.w2(32'hbc26b7e4),
	.w3(32'h3c154206),
	.w4(32'hbbceb636),
	.w5(32'hbc257cb9),
	.w6(32'hbc08acf8),
	.w7(32'hbc33b7ca),
	.w8(32'hbc082aff),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e6c1),
	.w1(32'h3b905ce9),
	.w2(32'h3b3e4508),
	.w3(32'hbc221ed9),
	.w4(32'h3b842ecb),
	.w5(32'h384eda82),
	.w6(32'h3ac2985b),
	.w7(32'hb9371b66),
	.w8(32'hba2608d6),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b362761),
	.w1(32'hbbff9902),
	.w2(32'hbcaff543),
	.w3(32'h3a5f43a6),
	.w4(32'hbc17a3b8),
	.w5(32'hbcca0250),
	.w6(32'h3b6ac73c),
	.w7(32'hbc5b163f),
	.w8(32'hbc4beae2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82635f),
	.w1(32'hbc868c6c),
	.w2(32'hbc8359a2),
	.w3(32'hbb81eb97),
	.w4(32'hbc183428),
	.w5(32'hbabf2e4b),
	.w6(32'hbb2e440e),
	.w7(32'hbc34f8c0),
	.w8(32'hbba61243),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f1057),
	.w1(32'h3c37a207),
	.w2(32'hbb184792),
	.w3(32'hbb311f6f),
	.w4(32'h3c2f02fa),
	.w5(32'h3aea0b64),
	.w6(32'h3b59fd06),
	.w7(32'h3bbbeee1),
	.w8(32'h3ac4e96d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c0b07),
	.w1(32'h3c4e5f05),
	.w2(32'h3c4cd7fd),
	.w3(32'hbc087c26),
	.w4(32'h3c729331),
	.w5(32'h3b4ab3ea),
	.w6(32'h3c412083),
	.w7(32'h3c6c95e8),
	.w8(32'h3c575016),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba890240),
	.w1(32'h3bcc1dcf),
	.w2(32'h3b8ecd0d),
	.w3(32'hbb5272c8),
	.w4(32'h3b971dd8),
	.w5(32'h3caeb254),
	.w6(32'h3a2ff07c),
	.w7(32'h3bcd0eb1),
	.w8(32'h3ae70a1a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b230751),
	.w1(32'hbacbbf8b),
	.w2(32'hbb2589fe),
	.w3(32'h3c01e4b3),
	.w4(32'hbb6bddad),
	.w5(32'hbb62f15b),
	.w6(32'hbbd93f6c),
	.w7(32'hbbef52a6),
	.w8(32'hbc0c56f5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf29e85),
	.w1(32'h3abb6d37),
	.w2(32'h3c1b5ff8),
	.w3(32'hbbaeeb7c),
	.w4(32'hbb8dda98),
	.w5(32'h3ae7047d),
	.w6(32'hba21ee3c),
	.w7(32'hb991b489),
	.w8(32'h3b026edd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70470c),
	.w1(32'h3ac8639c),
	.w2(32'h3b92a12b),
	.w3(32'hbb32aa53),
	.w4(32'h3b1b1022),
	.w5(32'h3b5413fb),
	.w6(32'h3c1db57f),
	.w7(32'h3be85e1d),
	.w8(32'h3c1d63cb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b9e44),
	.w1(32'hbc2eae65),
	.w2(32'hbc48f827),
	.w3(32'h3bd92b0a),
	.w4(32'hbbd28ffe),
	.w5(32'hbc2bf157),
	.w6(32'hbc32c5d1),
	.w7(32'hbc390fc9),
	.w8(32'hbc00f4d2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a49b1),
	.w1(32'hbc101dd6),
	.w2(32'hbba379b6),
	.w3(32'hbbd14400),
	.w4(32'hbc0a23d1),
	.w5(32'hbbe8bedd),
	.w6(32'hbc2aca4b),
	.w7(32'hba92dcba),
	.w8(32'hbb958d6b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec62a),
	.w1(32'h3cca9ccf),
	.w2(32'h3d0f0e6d),
	.w3(32'hbc40766c),
	.w4(32'h3cb789cf),
	.w5(32'h3cc75a6c),
	.w6(32'h3c4f814f),
	.w7(32'h3cb78316),
	.w8(32'h3c0d8194),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3a6dd),
	.w1(32'h38d628e7),
	.w2(32'hbb7e7257),
	.w3(32'h3c0eb3e4),
	.w4(32'hb9d47d83),
	.w5(32'hbb7cb1ca),
	.w6(32'hbb9dc089),
	.w7(32'hb9fe584a),
	.w8(32'hbc0043e0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13e0c7),
	.w1(32'hb9cbceeb),
	.w2(32'hbb060d06),
	.w3(32'hbbe4b392),
	.w4(32'h3ab044e2),
	.w5(32'hbbf674f7),
	.w6(32'h3a4e0cb8),
	.w7(32'hba6bdf5c),
	.w8(32'hbb3190b1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61357d),
	.w1(32'hbb582851),
	.w2(32'hbbb0350c),
	.w3(32'hbb92bda7),
	.w4(32'h3b1f9ed1),
	.w5(32'hbb1663bc),
	.w6(32'h3b7127ed),
	.w7(32'h3ad20376),
	.w8(32'hbaefad8c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde2e66),
	.w1(32'hbb645860),
	.w2(32'hbbac2ba5),
	.w3(32'hbaa8f7cc),
	.w4(32'h3ba6e4aa),
	.w5(32'hb9fc49c0),
	.w6(32'h3b82d012),
	.w7(32'hb8b733a2),
	.w8(32'h3bda587e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6626d1),
	.w1(32'hbc3a977c),
	.w2(32'hbc972b82),
	.w3(32'hbaa0a031),
	.w4(32'hba6d4748),
	.w5(32'hbc3d4558),
	.w6(32'h3b316f73),
	.w7(32'hbc05fe11),
	.w8(32'hbba91c07),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30b778),
	.w1(32'h3b009aee),
	.w2(32'h3b8b37a7),
	.w3(32'hbc6cb3cd),
	.w4(32'h3c215692),
	.w5(32'h3b542729),
	.w6(32'h399b78e2),
	.w7(32'h3b1ab873),
	.w8(32'h3abbc706),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b937228),
	.w1(32'h3bbcb330),
	.w2(32'h3d0ad3fd),
	.w3(32'hb98f6b02),
	.w4(32'h3c4d39a2),
	.w5(32'h3c6d5455),
	.w6(32'h396b4e70),
	.w7(32'h3ca46fa9),
	.w8(32'h3c4c401b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a50e1),
	.w1(32'h3bf0f76b),
	.w2(32'h3c36e0be),
	.w3(32'h3b98c76b),
	.w4(32'h3bd18a4c),
	.w5(32'h3c5a0763),
	.w6(32'h3bef4bd5),
	.w7(32'h3c1ad9c6),
	.w8(32'h3c09fddd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1ea0c),
	.w1(32'hbc44eafe),
	.w2(32'hbcee4b63),
	.w3(32'h3c735695),
	.w4(32'hbc860afd),
	.w5(32'hbca940f4),
	.w6(32'hb784d852),
	.w7(32'hbc673a98),
	.w8(32'hbbdad427),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc632d07),
	.w1(32'h3bef377f),
	.w2(32'hb9a0dfc1),
	.w3(32'hbc872eb6),
	.w4(32'hba060d24),
	.w5(32'h386dc44c),
	.w6(32'h3c89713d),
	.w7(32'h3b244ea5),
	.w8(32'h3b56e0fa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38e88),
	.w1(32'h3afd3e0b),
	.w2(32'h3b9244b4),
	.w3(32'h3b7672c5),
	.w4(32'h3bef28fd),
	.w5(32'h3c1381c1),
	.w6(32'hb9a41538),
	.w7(32'h3a95f632),
	.w8(32'h3ad33afd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79cb75),
	.w1(32'h3b8a4fc3),
	.w2(32'hbaa75fdb),
	.w3(32'h3c0aef20),
	.w4(32'h3b9b32ca),
	.w5(32'h3b41fbce),
	.w6(32'h3b38ebbc),
	.w7(32'h3bb94ff2),
	.w8(32'hbab86a85),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb290410),
	.w1(32'hbb806c64),
	.w2(32'hbbd70f75),
	.w3(32'h3aca9f94),
	.w4(32'h3b8c6a1e),
	.w5(32'h3a8debfb),
	.w6(32'h3bea2efc),
	.w7(32'h3b09b8a7),
	.w8(32'h3b8f426f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29263a),
	.w1(32'hbbaac6e0),
	.w2(32'hbca7f26e),
	.w3(32'h3b2d8a55),
	.w4(32'hbbc8dfd5),
	.w5(32'hbc3fe6e4),
	.w6(32'h39e8f338),
	.w7(32'hbc716ba0),
	.w8(32'hbc5018f2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c5916),
	.w1(32'hbad783cd),
	.w2(32'h3c67999b),
	.w3(32'hbc38899a),
	.w4(32'h3a0cab98),
	.w5(32'h3c8e4a6e),
	.w6(32'h3b0b700d),
	.w7(32'h3c040268),
	.w8(32'h3bf569e8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c975f04),
	.w1(32'h3bb07b55),
	.w2(32'h3c9e484b),
	.w3(32'h3c70744f),
	.w4(32'h3bc9ee6f),
	.w5(32'h3cc8676d),
	.w6(32'hbb6b8485),
	.w7(32'h3bc44758),
	.w8(32'h3c345d59),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4363bc),
	.w1(32'h3aaf4e97),
	.w2(32'hba98ae43),
	.w3(32'h3beb964e),
	.w4(32'hb96272fd),
	.w5(32'h386b95ff),
	.w6(32'hb9b60986),
	.w7(32'hba2a6d3c),
	.w8(32'hba3bd525),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc4a1f),
	.w1(32'hbb0c4725),
	.w2(32'hbb7e7f9a),
	.w3(32'h3a9ae280),
	.w4(32'hbaa300ef),
	.w5(32'hbb9d9ee2),
	.w6(32'hbade37d3),
	.w7(32'hbb272025),
	.w8(32'hbbb5b8a9),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49ee5e),
	.w1(32'h3b5a85a4),
	.w2(32'h3c26b1a5),
	.w3(32'hbb723c55),
	.w4(32'h3c48071d),
	.w5(32'h3c0e2309),
	.w6(32'hbb2ea61f),
	.w7(32'h3aa0a11c),
	.w8(32'h3a4a083a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1adbd8),
	.w1(32'h3b216a37),
	.w2(32'hbb234bd4),
	.w3(32'h3c018ecb),
	.w4(32'h3b8da7fa),
	.w5(32'hbab9072a),
	.w6(32'h3b8e8336),
	.w7(32'hba670e89),
	.w8(32'hb9c852cf),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b381034),
	.w1(32'h3cde8796),
	.w2(32'h3d6d5454),
	.w3(32'h3b238918),
	.w4(32'h3d0c3a72),
	.w5(32'h3d4e5bb7),
	.w6(32'h3babcc0a),
	.w7(32'h3cc94ffe),
	.w8(32'h3cf8bc38),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d19f40e),
	.w1(32'h3c5961a4),
	.w2(32'h3cf4d020),
	.w3(32'h3cd1e7da),
	.w4(32'h3b68f093),
	.w5(32'h3cd4a917),
	.w6(32'h3af899df),
	.w7(32'h3cabcaab),
	.w8(32'h3c608c47),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd22108),
	.w1(32'h3c0ad448),
	.w2(32'h3c3e5204),
	.w3(32'h3c9378a0),
	.w4(32'h3c4aaf24),
	.w5(32'h3c1910db),
	.w6(32'hbb33e309),
	.w7(32'h3bf7d3b5),
	.w8(32'h3c0ccec0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b082d),
	.w1(32'hbc83abd0),
	.w2(32'hbc6d8358),
	.w3(32'h3b0a0560),
	.w4(32'hbc8b27d4),
	.w5(32'hbc801bae),
	.w6(32'hbb80787b),
	.w7(32'hbb7dc811),
	.w8(32'h3afd40fd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb979d88),
	.w1(32'hbb1ddac9),
	.w2(32'hbbfc8eb5),
	.w3(32'hbaf5c7b6),
	.w4(32'hbb15cbdc),
	.w5(32'hbc077248),
	.w6(32'h3bb7f097),
	.w7(32'hba0239da),
	.w8(32'h3b7e3150),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ac87a),
	.w1(32'hbb5b132e),
	.w2(32'hbc82040d),
	.w3(32'hbba20ac8),
	.w4(32'hbba52a86),
	.w5(32'hbba1e3c8),
	.w6(32'hbb125320),
	.w7(32'hbc657913),
	.w8(32'hbc56e05a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18503a),
	.w1(32'h3a0fe90e),
	.w2(32'h3b856712),
	.w3(32'hbb0b9c4d),
	.w4(32'h3b282209),
	.w5(32'h3a92e707),
	.w6(32'hbb3ab5af),
	.w7(32'hb6c9f6fc),
	.w8(32'h3b3a2f2f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be4c0),
	.w1(32'hbc151a4e),
	.w2(32'hbbfd2d9e),
	.w3(32'h3af2223d),
	.w4(32'hbb84a9a6),
	.w5(32'hbb97513d),
	.w6(32'hbbee7f42),
	.w7(32'hbc5bb4a7),
	.w8(32'hbc2008fc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a316a),
	.w1(32'hbbe2964a),
	.w2(32'hbb416a6c),
	.w3(32'h3c56c010),
	.w4(32'hbc2c9270),
	.w5(32'hb9d7c7e5),
	.w6(32'h3b8c76f6),
	.w7(32'hbc179fa2),
	.w8(32'h3b42727d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b719),
	.w1(32'h3b37e0b9),
	.w2(32'hb874eab1),
	.w3(32'hbb226a95),
	.w4(32'h3b6dd6a0),
	.w5(32'h3b015c7d),
	.w6(32'h3b02faa1),
	.w7(32'h38b690ca),
	.w8(32'hbb210d1f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf036e1),
	.w1(32'h3a8104b6),
	.w2(32'hbaed2a72),
	.w3(32'hba4b8646),
	.w4(32'h3c063b92),
	.w5(32'h3b8e4845),
	.w6(32'hb79739c8),
	.w7(32'hbab77492),
	.w8(32'h3b39ec95),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895d1f),
	.w1(32'hbba29c58),
	.w2(32'hbb918e53),
	.w3(32'h3b4e91dc),
	.w4(32'hbbd8c115),
	.w5(32'hbc205710),
	.w6(32'h3b814578),
	.w7(32'h3b218a8a),
	.w8(32'h3b9ccd7c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07bde5),
	.w1(32'h3c0682a1),
	.w2(32'h3c806325),
	.w3(32'hbbd5c17e),
	.w4(32'h3bdf24b5),
	.w5(32'h3c26dd36),
	.w6(32'hb8fba9f9),
	.w7(32'h3b81bcd6),
	.w8(32'h3bf0b1ce),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e5f64),
	.w1(32'h3be29e37),
	.w2(32'h3bb80add),
	.w3(32'h3c665a1e),
	.w4(32'h3bff2828),
	.w5(32'h3b931a2d),
	.w6(32'h3b55c9e2),
	.w7(32'h3b1ec4ef),
	.w8(32'h3b83badd),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb33759),
	.w1(32'hbbbe9bbb),
	.w2(32'h3bd8c844),
	.w3(32'h3b9ff5f3),
	.w4(32'h3b2a35bb),
	.w5(32'h37d2d294),
	.w6(32'hbc1574d3),
	.w7(32'h3917d93d),
	.w8(32'h3a93bd2d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53c758),
	.w1(32'hbb20a873),
	.w2(32'hbb5d6879),
	.w3(32'h3ae616f2),
	.w4(32'hbb08f3d9),
	.w5(32'hbb8fe9f9),
	.w6(32'hb8bd2310),
	.w7(32'hbacab333),
	.w8(32'hbbbeb22d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdfe0d),
	.w1(32'h3b83848c),
	.w2(32'hb9ab62c2),
	.w3(32'hbbb4a8a7),
	.w4(32'h3b1883e4),
	.w5(32'h3b7ff421),
	.w6(32'hbaf5dbc7),
	.w7(32'hba11e6d4),
	.w8(32'h3b80e77a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995e887),
	.w1(32'hbc0a642a),
	.w2(32'hbc235395),
	.w3(32'h3a602a0d),
	.w4(32'h399d1239),
	.w5(32'hbb7ee2bc),
	.w6(32'hbb8dd385),
	.w7(32'hbc861fda),
	.w8(32'hbc496e9a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc119f5d),
	.w1(32'hbb5ab52e),
	.w2(32'hbb51736a),
	.w3(32'h3b9841ac),
	.w4(32'h3b4b12fc),
	.w5(32'hbaebd9fa),
	.w6(32'h3b9595fd),
	.w7(32'h3b9705b3),
	.w8(32'h3bdcad27),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3962d689),
	.w1(32'h3b5445c4),
	.w2(32'hb9a009be),
	.w3(32'h3ad1b22d),
	.w4(32'h3b24a0cb),
	.w5(32'hba36d798),
	.w6(32'h3a819e47),
	.w7(32'hba35aa75),
	.w8(32'hba0b7c09),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f6da8),
	.w1(32'h3b7098ec),
	.w2(32'h3bddb154),
	.w3(32'h39e61697),
	.w4(32'h3b513133),
	.w5(32'hba13078c),
	.w6(32'h3aeb0da0),
	.w7(32'h3bec38b3),
	.w8(32'h3c27c602),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc02702),
	.w1(32'h3b9a93ab),
	.w2(32'h3bf9228c),
	.w3(32'hbac4507e),
	.w4(32'h3c05a2b7),
	.w5(32'h3bc621cc),
	.w6(32'h3bb8edc2),
	.w7(32'h3b8b2534),
	.w8(32'hb98be5f7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b995a24),
	.w1(32'hbc5186cf),
	.w2(32'hbd1022b6),
	.w3(32'h3af15b6d),
	.w4(32'hbb5cb8ff),
	.w5(32'hbc9414b5),
	.w6(32'hbbdf79c8),
	.w7(32'hbca1367c),
	.w8(32'hbc8dbf9d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cbc29),
	.w1(32'hba86e837),
	.w2(32'h3b0dc0b9),
	.w3(32'hbc205420),
	.w4(32'hbb151386),
	.w5(32'hbb1df323),
	.w6(32'hbb0721b0),
	.w7(32'h3ba524b0),
	.w8(32'h3a02c1de),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb274f9c),
	.w1(32'h3cf6041a),
	.w2(32'h3c82a994),
	.w3(32'hbba7d5db),
	.w4(32'h3ccf374a),
	.w5(32'h3cad9c34),
	.w6(32'h3c6050db),
	.w7(32'h3c66c27f),
	.w8(32'h3c80174f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f06cb),
	.w1(32'hbc6544b2),
	.w2(32'hbc929041),
	.w3(32'h3c7cde01),
	.w4(32'hbc60e99e),
	.w5(32'hbc8519e5),
	.w6(32'hbbc7036d),
	.w7(32'hbbfe4521),
	.w8(32'hbc89cd9f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ebfb8),
	.w1(32'hbbb14eb7),
	.w2(32'hbb81cb6a),
	.w3(32'hbc9f9711),
	.w4(32'hbbb27a17),
	.w5(32'hbbc6f4cb),
	.w6(32'hbb8c0434),
	.w7(32'hbb99cf85),
	.w8(32'hbba30fb0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadb4ab),
	.w1(32'h39824c00),
	.w2(32'hbc0c44c3),
	.w3(32'hbbc7387b),
	.w4(32'hbbe40421),
	.w5(32'hbbb41aed),
	.w6(32'h3b2f1703),
	.w7(32'hbb2f327b),
	.w8(32'hbbcaa3cd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c179b),
	.w1(32'hbc3265ee),
	.w2(32'hbc7e094f),
	.w3(32'h3a25d26c),
	.w4(32'h3732ef38),
	.w5(32'hbb2d168d),
	.w6(32'hbc74f624),
	.w7(32'hbc71a053),
	.w8(32'hbc0adace),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76c640),
	.w1(32'hbc294a8f),
	.w2(32'hbce8c331),
	.w3(32'hbc6a8e9c),
	.w4(32'hbc63878c),
	.w5(32'hbc83f495),
	.w6(32'h3b58faeb),
	.w7(32'hbc402f6a),
	.w8(32'hbc70d99d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9865cf),
	.w1(32'h37f80534),
	.w2(32'hbb5317e6),
	.w3(32'h3b36a45d),
	.w4(32'h3b09f431),
	.w5(32'h3aa67f01),
	.w6(32'h3ab17434),
	.w7(32'h3a9b3400),
	.w8(32'h3af92817),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e5030),
	.w1(32'hbbe1be48),
	.w2(32'hbc37b8d2),
	.w3(32'h3ac2fbd2),
	.w4(32'hb9ec62d7),
	.w5(32'h3b974196),
	.w6(32'hbbe53ff2),
	.w7(32'hbb65e4fc),
	.w8(32'h3c1d7958),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule