module layer_10_featuremap_74(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf16ed9),
	.w1(32'h3c30aee2),
	.w2(32'h3b649983),
	.w3(32'hbbf386ea),
	.w4(32'h3b6b9849),
	.w5(32'hbc1d2fec),
	.w6(32'hbc283b90),
	.w7(32'hba69e2df),
	.w8(32'hbc4a3bdf),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c189c1a),
	.w1(32'h3b45719d),
	.w2(32'hbb37bfdc),
	.w3(32'hbc2098d5),
	.w4(32'hb97157ea),
	.w5(32'h3c5ff2fa),
	.w6(32'hbbf4da5f),
	.w7(32'hbb6ab8a8),
	.w8(32'h3bf5bd94),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36f235),
	.w1(32'hb9d93491),
	.w2(32'h38ac10c6),
	.w3(32'h3c5b1542),
	.w4(32'hbae1ec0b),
	.w5(32'h3a3683d5),
	.w6(32'h3b829f33),
	.w7(32'hbb3dc7f1),
	.w8(32'h3c05109d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04f3f4),
	.w1(32'h392727f7),
	.w2(32'hbbd4bef1),
	.w3(32'hba728475),
	.w4(32'h3b9c7af8),
	.w5(32'hbc3cc1e3),
	.w6(32'h3bbd4641),
	.w7(32'h3bfb9329),
	.w8(32'h3b6286a9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc045d01),
	.w1(32'hbadfd5ee),
	.w2(32'h3b72deae),
	.w3(32'hb864f4fc),
	.w4(32'h3b1c0009),
	.w5(32'hbb303bce),
	.w6(32'hbaed644e),
	.w7(32'h3ba926b4),
	.w8(32'h3b84033b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396803d2),
	.w1(32'h3b302614),
	.w2(32'hbbb13554),
	.w3(32'hbb0f8512),
	.w4(32'h3b698f1e),
	.w5(32'hbb484c2b),
	.w6(32'h3baf3683),
	.w7(32'h3c20dd31),
	.w8(32'hbb253b49),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b29ac),
	.w1(32'hbb380294),
	.w2(32'hbbbb2582),
	.w3(32'h3c3bdb3a),
	.w4(32'h3b950597),
	.w5(32'hbaee31e9),
	.w6(32'h3c3eb4bc),
	.w7(32'h3b3226aa),
	.w8(32'hbc13d54a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc5f12),
	.w1(32'hbb9a310c),
	.w2(32'hbbcd3ac6),
	.w3(32'hbb998d3a),
	.w4(32'hbbdde363),
	.w5(32'hbc1a3404),
	.w6(32'hbbc06879),
	.w7(32'hbb9af0fb),
	.w8(32'hbba6165d),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08facf),
	.w1(32'h3ab11013),
	.w2(32'h3b9bec2b),
	.w3(32'hbba0abb2),
	.w4(32'hbbe271ea),
	.w5(32'h3cb79fdb),
	.w6(32'hbbbafbce),
	.w7(32'hbb9444de),
	.w8(32'h3c8081f8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2d46b),
	.w1(32'h3c5f639c),
	.w2(32'h3b7080a1),
	.w3(32'h3d0e5ace),
	.w4(32'h3ccf9667),
	.w5(32'h3b9e4587),
	.w6(32'h3cdd9800),
	.w7(32'h3cb2a65e),
	.w8(32'h3b91f070),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b929f98),
	.w1(32'h3b3dedc3),
	.w2(32'h3be142fa),
	.w3(32'h3be89808),
	.w4(32'h3bea2c8a),
	.w5(32'hbb0adcfc),
	.w6(32'h3c01844f),
	.w7(32'h3bd3ac1b),
	.w8(32'hbb38b73e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b695dc5),
	.w1(32'h3b58a55c),
	.w2(32'hbb249342),
	.w3(32'h3b7759e4),
	.w4(32'h3c0b7ea1),
	.w5(32'hbb4a6fbf),
	.w6(32'h3be82423),
	.w7(32'h3b16b171),
	.w8(32'h39c98897),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38140b8d),
	.w1(32'hbaa23170),
	.w2(32'h3c166d12),
	.w3(32'h3ab6cd24),
	.w4(32'hba6afedf),
	.w5(32'h3c236a7e),
	.w6(32'h3b503130),
	.w7(32'h3b1f9df7),
	.w8(32'h3c0fd458),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b465d94),
	.w1(32'h3b56aeb6),
	.w2(32'hbb21a0b8),
	.w3(32'hbae92457),
	.w4(32'hbaf6222a),
	.w5(32'hbbefaf8c),
	.w6(32'h3b4c98b3),
	.w7(32'hbb8c02a4),
	.w8(32'h3b91e3fb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01dd8d),
	.w1(32'h3adb9c11),
	.w2(32'hbb15e5eb),
	.w3(32'hbb98446a),
	.w4(32'h3b5d8003),
	.w5(32'h3b9f912c),
	.w6(32'h3c0ecaa3),
	.w7(32'h3bab2f4e),
	.w8(32'hb994bb78),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1020f),
	.w1(32'h3bb70c12),
	.w2(32'h3ae9af54),
	.w3(32'h3bdbcace),
	.w4(32'h3bc9e129),
	.w5(32'h3abd15fa),
	.w6(32'hbb002145),
	.w7(32'hbb02b06b),
	.w8(32'h3b33b9de),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c6363),
	.w1(32'h3b166bb0),
	.w2(32'hbae9ccad),
	.w3(32'h3b81d799),
	.w4(32'h3b962486),
	.w5(32'h3befe274),
	.w6(32'h3bc79aa8),
	.w7(32'h3b8b7006),
	.w8(32'hbbeae196),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15fc1),
	.w1(32'h39c75f3e),
	.w2(32'h3b87fccb),
	.w3(32'h3c4481c6),
	.w4(32'h3b73a46e),
	.w5(32'h3b6f565d),
	.w6(32'hb8e14142),
	.w7(32'hbbd67fbb),
	.w8(32'h3b1d2af8),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d98b),
	.w1(32'h3b3ad077),
	.w2(32'hbc229798),
	.w3(32'h3c02bab1),
	.w4(32'h3b0bf388),
	.w5(32'hbc46535f),
	.w6(32'h3aa030d0),
	.w7(32'hbaabbaa5),
	.w8(32'h3c2e9e92),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbec760),
	.w1(32'hbc56dcb6),
	.w2(32'h3a978a6a),
	.w3(32'hbca64420),
	.w4(32'hbca0fa67),
	.w5(32'hbb26b0f4),
	.w6(32'hba82230b),
	.w7(32'hbc3d2a35),
	.w8(32'hbbc5fd6b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7505e1),
	.w1(32'hbb11e4b9),
	.w2(32'hbbb13611),
	.w3(32'hbc0095bd),
	.w4(32'hbb939134),
	.w5(32'hbbe72647),
	.w6(32'hbbafa636),
	.w7(32'hb714f106),
	.w8(32'h3b0b1f8f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7987bf),
	.w1(32'hbb959ec3),
	.w2(32'hbc230483),
	.w3(32'hbc1700bc),
	.w4(32'hbb9758a1),
	.w5(32'hbc8eb76b),
	.w6(32'h3ac97160),
	.w7(32'h3ae050aa),
	.w8(32'hbbc40585),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96601c),
	.w1(32'hbb53208c),
	.w2(32'h3b920469),
	.w3(32'hbc7b3d4e),
	.w4(32'hbb3e3460),
	.w5(32'h3c19d7c9),
	.w6(32'hbbcba9b6),
	.w7(32'h3b4cd697),
	.w8(32'h3bbfcaf0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb10422),
	.w1(32'h3a6005df),
	.w2(32'h3ba08b07),
	.w3(32'h3c26a26a),
	.w4(32'h3c023924),
	.w5(32'hbad185b7),
	.w6(32'h3be27fa1),
	.w7(32'h3b81dcc2),
	.w8(32'hbabcc68b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2e8c1),
	.w1(32'h3b24d5e9),
	.w2(32'hbc336063),
	.w3(32'h3aaf6e53),
	.w4(32'h3a6f225d),
	.w5(32'hbc1b439d),
	.w6(32'hbb16507c),
	.w7(32'hbb434404),
	.w8(32'h3c39b9ff),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34e738),
	.w1(32'h3a752027),
	.w2(32'h3c3cd617),
	.w3(32'hbc375399),
	.w4(32'hbc03f732),
	.w5(32'h3bf62ec0),
	.w6(32'h3c2f5301),
	.w7(32'h3bcfea62),
	.w8(32'h3ae6cdf4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb483d),
	.w1(32'h3b6a7071),
	.w2(32'hb9b67a8b),
	.w3(32'hbcb030bb),
	.w4(32'hbc2a5c7e),
	.w5(32'hbac5b155),
	.w6(32'hbbaa62f8),
	.w7(32'hbb599f36),
	.w8(32'hba3cae09),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e18b4),
	.w1(32'hb6a692fe),
	.w2(32'h3b82edcc),
	.w3(32'hbaa380c5),
	.w4(32'hba7868d0),
	.w5(32'hb91a0ee3),
	.w6(32'hb89efa2e),
	.w7(32'hb6b80db5),
	.w8(32'h3b28b310),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b041ea7),
	.w1(32'h3a09c2be),
	.w2(32'hbab03114),
	.w3(32'h3b9305d8),
	.w4(32'hbb64bfec),
	.w5(32'hbb98fbcc),
	.w6(32'h3b14c3e9),
	.w7(32'hbb856478),
	.w8(32'hbb3aa823),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91b3c4),
	.w1(32'h3ab261d6),
	.w2(32'hba7cbd78),
	.w3(32'hbc25b0d5),
	.w4(32'h3abe427b),
	.w5(32'hbac2e6ba),
	.w6(32'hbc809e05),
	.w7(32'hbc3166a1),
	.w8(32'h3a27cc0a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205c8a),
	.w1(32'h3a619748),
	.w2(32'hbaf40669),
	.w3(32'hbb72a656),
	.w4(32'h3ab77ec5),
	.w5(32'hbacdef1b),
	.w6(32'h36fc1689),
	.w7(32'h3b855f40),
	.w8(32'h3b04bc41),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b1c51),
	.w1(32'hbc0b27bb),
	.w2(32'hbc22fa64),
	.w3(32'hbc1713c9),
	.w4(32'hbba1aa40),
	.w5(32'hbc4dd782),
	.w6(32'hbbe3846e),
	.w7(32'h3b1c6cfb),
	.w8(32'hbc78737b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f4941),
	.w1(32'hbc14c538),
	.w2(32'hbaac4e98),
	.w3(32'hbc8ce6c8),
	.w4(32'hbc3d21fa),
	.w5(32'h3acdb307),
	.w6(32'hbc897ce5),
	.w7(32'hbc0faf89),
	.w8(32'h3b5c921a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52d45),
	.w1(32'hba029bcc),
	.w2(32'hbb8b5880),
	.w3(32'h3b36866d),
	.w4(32'h3b9f1345),
	.w5(32'hbc2bcb6c),
	.w6(32'h3bb0d977),
	.w7(32'h3b585844),
	.w8(32'hbc53b6f5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba00e4b),
	.w1(32'hbb53bcd0),
	.w2(32'h3b3528fa),
	.w3(32'hbcd38097),
	.w4(32'hbc4be94a),
	.w5(32'h3b433219),
	.w6(32'hbcb02bd1),
	.w7(32'hbb7eabb8),
	.w8(32'h3a9f9d86),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a5412),
	.w1(32'h396ffbe4),
	.w2(32'hbbc37547),
	.w3(32'h3af5f09d),
	.w4(32'hbad11beb),
	.w5(32'hbb81145f),
	.w6(32'hbaa484b7),
	.w7(32'hbb43902d),
	.w8(32'h3c0cac2f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5993e0),
	.w1(32'hbc5cff04),
	.w2(32'hba9ed21c),
	.w3(32'h3be167cc),
	.w4(32'h3b7a0518),
	.w5(32'h3b33671d),
	.w6(32'hbb217500),
	.w7(32'hbb6810f2),
	.w8(32'h3b37299d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba584f4),
	.w1(32'hbba38cff),
	.w2(32'hbc45af86),
	.w3(32'hbaed8121),
	.w4(32'hbb98e633),
	.w5(32'hbc007649),
	.w6(32'hbaf2dee9),
	.w7(32'hbba3b5c8),
	.w8(32'h3bc50adc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79dbd6),
	.w1(32'hba9f984b),
	.w2(32'h3b949159),
	.w3(32'hbbdb2814),
	.w4(32'h3b1ad518),
	.w5(32'h3c2bf8dd),
	.w6(32'h3bc452d7),
	.w7(32'h3c0b2243),
	.w8(32'h3c9d6ab6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7c52f),
	.w1(32'h3b837b5b),
	.w2(32'h3b11951b),
	.w3(32'hbb2cbfcd),
	.w4(32'hbc11ecc7),
	.w5(32'h3aa88d58),
	.w6(32'h3bb72f2e),
	.w7(32'hbb483087),
	.w8(32'hbb496313),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b831ee2),
	.w1(32'h3b9382de),
	.w2(32'hbbc346db),
	.w3(32'h3b5deef7),
	.w4(32'h3b377781),
	.w5(32'hbc3cdfbb),
	.w6(32'hbb1e52c6),
	.w7(32'h3b8f4173),
	.w8(32'h399667ea),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5031f0),
	.w1(32'hbc2504f2),
	.w2(32'hbcd3c15a),
	.w3(32'hbc29846f),
	.w4(32'hbba48208),
	.w5(32'hbd03a577),
	.w6(32'h3b314cd6),
	.w7(32'h3b6c48b6),
	.w8(32'hbb84faa9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf94263),
	.w1(32'hbc9bc56d),
	.w2(32'hbac34f1c),
	.w3(32'hbd25deea),
	.w4(32'hbc8896a5),
	.w5(32'h3a0edb12),
	.w6(32'hbcb640a2),
	.w7(32'hbc1c3067),
	.w8(32'h38c69962),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b05460),
	.w1(32'h3b5ccf87),
	.w2(32'hb96865c3),
	.w3(32'h3a6a304c),
	.w4(32'hba673c32),
	.w5(32'h3ba6c51d),
	.w6(32'hb9d3303f),
	.w7(32'h395ac629),
	.w8(32'hbab3ee8c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33220c),
	.w1(32'h3c29207f),
	.w2(32'hbbf66d8e),
	.w3(32'hbae062d2),
	.w4(32'h3bc2b130),
	.w5(32'hbc3820b9),
	.w6(32'hbbe04285),
	.w7(32'hbb80d654),
	.w8(32'hbb747118),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31274e),
	.w1(32'hbb86afc2),
	.w2(32'h3c5852da),
	.w3(32'hbb42d6e7),
	.w4(32'h3bf6b472),
	.w5(32'h3c9f45d0),
	.w6(32'hb90160f6),
	.w7(32'h3bae132b),
	.w8(32'h3c6f8b6e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c214258),
	.w1(32'hbb31780b),
	.w2(32'h3bced23d),
	.w3(32'h3c22c5b2),
	.w4(32'hb9f108e6),
	.w5(32'hbbc89018),
	.w6(32'h3c8862a6),
	.w7(32'h3b82d287),
	.w8(32'h3af57602),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfff21),
	.w1(32'h39813254),
	.w2(32'h3b4b4903),
	.w3(32'h3a9ad877),
	.w4(32'h3c0d5b99),
	.w5(32'hba85d613),
	.w6(32'h3c26e073),
	.w7(32'h3c24956b),
	.w8(32'hbad41267),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abacc6a),
	.w1(32'hba08aa54),
	.w2(32'h3c104784),
	.w3(32'hba8da741),
	.w4(32'hbb94fa1e),
	.w5(32'h3aa39809),
	.w6(32'hbb1df5c5),
	.w7(32'hbbb72137),
	.w8(32'h3b0eaac9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b4ec0),
	.w1(32'hbad38c71),
	.w2(32'hbcbdbbb8),
	.w3(32'hb9f8ba5e),
	.w4(32'h3b3478c0),
	.w5(32'hbce15312),
	.w6(32'hbb9ba36a),
	.w7(32'h3b5bf60e),
	.w8(32'hbcee76d3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1375cb),
	.w1(32'hbc89c255),
	.w2(32'hbc3a0385),
	.w3(32'hbd4c938e),
	.w4(32'hbcb677c3),
	.w5(32'hbc13c4f7),
	.w6(32'hbd11f3bb),
	.w7(32'hbc70d296),
	.w8(32'hbb218760),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87d129),
	.w1(32'h3a92c41b),
	.w2(32'hbc19b335),
	.w3(32'hbb4c6514),
	.w4(32'h3b509518),
	.w5(32'hbd157ad7),
	.w6(32'h3bd2c51a),
	.w7(32'h3c3537f8),
	.w8(32'hbd0d533a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf11900),
	.w1(32'hbcb6e30d),
	.w2(32'h38c2a219),
	.w3(32'hbd2861ea),
	.w4(32'hbc9a1ff7),
	.w5(32'h3b88486c),
	.w6(32'hbd100a23),
	.w7(32'hbbed0fe0),
	.w8(32'h3ba9a208),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7df56f),
	.w1(32'h3c83df1e),
	.w2(32'hbc38ab33),
	.w3(32'h3c0f3736),
	.w4(32'h3c3afbe2),
	.w5(32'hbad1699e),
	.w6(32'h3afb8127),
	.w7(32'h3b23fb75),
	.w8(32'h3b87561d),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3fd9a),
	.w1(32'h3b665f3d),
	.w2(32'hbb14f87b),
	.w3(32'hba50a95a),
	.w4(32'hba60d90c),
	.w5(32'h3a8247f9),
	.w6(32'hbc33cb79),
	.w7(32'hbba3ac4c),
	.w8(32'hbb8a65db),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63e91e),
	.w1(32'h3bc1bba8),
	.w2(32'h3c39b7cd),
	.w3(32'hbb00a4f0),
	.w4(32'hbc0fe6a3),
	.w5(32'h3a30f31d),
	.w6(32'hbb9a9bd0),
	.w7(32'hbc2c7df4),
	.w8(32'h3c0823dd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52ba9e),
	.w1(32'h3a44e096),
	.w2(32'h3b9ea5d1),
	.w3(32'hbbd0d0dd),
	.w4(32'hbb23ccd6),
	.w5(32'h3bafd9cd),
	.w6(32'h3b95c852),
	.w7(32'h3b20a084),
	.w8(32'h3bcc2ccc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a253e3),
	.w1(32'hb7ec83ed),
	.w2(32'hbb5f45f2),
	.w3(32'hbb4d2c49),
	.w4(32'hbae09bf4),
	.w5(32'hb94e520d),
	.w6(32'hbab94899),
	.w7(32'hbaa8afa8),
	.w8(32'h39a45edb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd338),
	.w1(32'h3a7eb6ff),
	.w2(32'hbb11784b),
	.w3(32'h3b996482),
	.w4(32'h3b2b1756),
	.w5(32'hba8c1d9f),
	.w6(32'h3afabea1),
	.w7(32'hba44a615),
	.w8(32'h3b827a55),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4af013),
	.w1(32'h3b8ed658),
	.w2(32'h3b8a14bd),
	.w3(32'h3b3404ea),
	.w4(32'h3bafa948),
	.w5(32'hbbd3109f),
	.w6(32'h3b70a961),
	.w7(32'h3b0fea38),
	.w8(32'hbb32379e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c233204),
	.w1(32'h3b47171e),
	.w2(32'hbab1424a),
	.w3(32'hbc0c5259),
	.w4(32'hba855fb1),
	.w5(32'hbb0b924d),
	.w6(32'h3781868d),
	.w7(32'h3c0bee3a),
	.w8(32'h3bcaae00),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd87d),
	.w1(32'hbc110781),
	.w2(32'hbb07f2aa),
	.w3(32'hbc98d98b),
	.w4(32'hbc3843f6),
	.w5(32'h3a38618a),
	.w6(32'h3b69331a),
	.w7(32'h3a7bd091),
	.w8(32'h3c30ae40),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3709f),
	.w1(32'h3b28be03),
	.w2(32'h3afb4d61),
	.w3(32'hbb3e1308),
	.w4(32'hb9b575ab),
	.w5(32'h3b718edf),
	.w6(32'h3c36b581),
	.w7(32'h3c3ed2e4),
	.w8(32'h3becd465),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfafc92),
	.w1(32'h3c3a2d13),
	.w2(32'h3c7525a7),
	.w3(32'h3c0a5e7d),
	.w4(32'h3c1d4a50),
	.w5(32'h3ccb15cd),
	.w6(32'h3c65fa58),
	.w7(32'h3c861c92),
	.w8(32'h3ca9131f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbaaca2),
	.w1(32'h3cabc973),
	.w2(32'hb93a95eb),
	.w3(32'h3d1b7216),
	.w4(32'h3ca2cbba),
	.w5(32'h3b20567b),
	.w6(32'h3cb21811),
	.w7(32'h3c51390d),
	.w8(32'h3b6bab56),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e30d5),
	.w1(32'h3ac968f6),
	.w2(32'hbbaedbdd),
	.w3(32'h3adc2dd7),
	.w4(32'h3b52e33f),
	.w5(32'hbb3349f3),
	.w6(32'h3a838d80),
	.w7(32'h3a9aa267),
	.w8(32'hbb5b3929),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70673b),
	.w1(32'hbaca29ef),
	.w2(32'hbc6698fa),
	.w3(32'hba8b2211),
	.w4(32'hbaafb1de),
	.w5(32'hbc788cbf),
	.w6(32'hbacbed6a),
	.w7(32'hbb7b72b0),
	.w8(32'hbc65008b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64a549),
	.w1(32'h3aeb858f),
	.w2(32'h3a34d449),
	.w3(32'hbcc31d4a),
	.w4(32'hbb96c66b),
	.w5(32'hbb9c3212),
	.w6(32'hbca94d74),
	.w7(32'h3919b280),
	.w8(32'hbb45bca0),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1492cf),
	.w1(32'hbba60bce),
	.w2(32'h3b3d925a),
	.w3(32'hbbea5921),
	.w4(32'hbbd87d23),
	.w5(32'h3b934b4c),
	.w6(32'hbc119597),
	.w7(32'h38beb4cf),
	.w8(32'h3b9ad2f3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ffc39),
	.w1(32'h3b7a8fad),
	.w2(32'h3bbac817),
	.w3(32'h3a43664d),
	.w4(32'h3b7a700d),
	.w5(32'h3bcb87cb),
	.w6(32'h37882760),
	.w7(32'h3b0a929b),
	.w8(32'h3b8f03da),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af349c2),
	.w1(32'h3c22240c),
	.w2(32'h3b2db943),
	.w3(32'hbb14d070),
	.w4(32'h3b77ece0),
	.w5(32'h3b2a85b2),
	.w6(32'hb9f2ff80),
	.w7(32'h3b1987a9),
	.w8(32'h3c14b863),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adc8c0),
	.w1(32'h38265123),
	.w2(32'h3c867ef0),
	.w3(32'h3ab68f40),
	.w4(32'h3bc19cb0),
	.w5(32'h3c8a0832),
	.w6(32'h3c68a7a0),
	.w7(32'h3c1d7bc5),
	.w8(32'h3c303cdb),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb11353),
	.w1(32'h3c42ee86),
	.w2(32'hbc3a3d71),
	.w3(32'h3ce042fe),
	.w4(32'h3c6fd0f2),
	.w5(32'hbc1730d2),
	.w6(32'h3cb2461c),
	.w7(32'h3c1a2661),
	.w8(32'hbaae9175),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc043da7),
	.w1(32'h3b03e57b),
	.w2(32'h3c3a7686),
	.w3(32'hbc940ff5),
	.w4(32'h39c7dc38),
	.w5(32'h3b909a68),
	.w6(32'hbc4ac627),
	.w7(32'h3b9e9354),
	.w8(32'h3ba46b79),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca8f0d),
	.w1(32'h3bea2f71),
	.w2(32'hb9f21f40),
	.w3(32'hbb04d10b),
	.w4(32'h385d3d91),
	.w5(32'hbb9cc8fd),
	.w6(32'hb8987cdd),
	.w7(32'hb9c9ddfa),
	.w8(32'hbac64c9b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3847d3),
	.w1(32'h3adf8028),
	.w2(32'h3c8313b8),
	.w3(32'hbc311f6f),
	.w4(32'hba9bcc61),
	.w5(32'h3cce3c17),
	.w6(32'hbb11b25c),
	.w7(32'h3bb84056),
	.w8(32'h3c6d27ff),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdc0bb5),
	.w1(32'h3cb69d7e),
	.w2(32'h3a1fcb06),
	.w3(32'h3d0caacd),
	.w4(32'h3cbd4979),
	.w5(32'h3c94953c),
	.w6(32'h3d009421),
	.w7(32'h3c241244),
	.w8(32'h3c8f94d7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830a5f),
	.w1(32'h3cbf0e46),
	.w2(32'h3a9c16af),
	.w3(32'h3c98090e),
	.w4(32'h3c856c4c),
	.w5(32'h3b04df99),
	.w6(32'h3c864de1),
	.w7(32'h3bf91f3d),
	.w8(32'hbab68d08),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27f59e),
	.w1(32'hbb906a0a),
	.w2(32'hba7795c4),
	.w3(32'hbc3c0faf),
	.w4(32'hbb4b97d7),
	.w5(32'h3af0629b),
	.w6(32'hba8bc38a),
	.w7(32'h3a643cef),
	.w8(32'h3a6611a3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae4a8f),
	.w1(32'hba579aa5),
	.w2(32'h3ba0ff96),
	.w3(32'hbbb33fc7),
	.w4(32'h3ac942d2),
	.w5(32'h3b5877e6),
	.w6(32'hbb933fe6),
	.w7(32'h39f3d7e5),
	.w8(32'hba96f628),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e31b61),
	.w1(32'h3ba7ab89),
	.w2(32'hbabfc0ed),
	.w3(32'hb8fd9b92),
	.w4(32'h3a86ad89),
	.w5(32'hbb335c2a),
	.w6(32'hb9b8b2de),
	.w7(32'h3ba2d6f4),
	.w8(32'h3ad60fc8),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae53781),
	.w1(32'h3ac06135),
	.w2(32'h3b950c69),
	.w3(32'hbaeff59e),
	.w4(32'h3aedbe5f),
	.w5(32'h3b25d56b),
	.w6(32'h3b1f6c87),
	.w7(32'h3bc60255),
	.w8(32'hba5a9331),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b873e1e),
	.w1(32'hbbc30b0e),
	.w2(32'h3bcef28b),
	.w3(32'h3b4cc2c2),
	.w4(32'hbbd07459),
	.w5(32'h3c02efd1),
	.w6(32'hbc17df14),
	.w7(32'hbbc1ad49),
	.w8(32'h3c2c4a91),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35b7eb),
	.w1(32'hbb969980),
	.w2(32'h3c503545),
	.w3(32'h3af02d85),
	.w4(32'hbbf15bfc),
	.w5(32'h3c8728ed),
	.w6(32'h3c79a0f9),
	.w7(32'h3bb30b45),
	.w8(32'h3c43ee71),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25fc13),
	.w1(32'hbba98232),
	.w2(32'hbaf355f9),
	.w3(32'h3c249efa),
	.w4(32'hbc05558e),
	.w5(32'h3a7c8fca),
	.w6(32'h3c558959),
	.w7(32'h3ad48367),
	.w8(32'hbbe58dcd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb939777),
	.w1(32'hbb5d06b2),
	.w2(32'h3b6eff25),
	.w3(32'h3b969e28),
	.w4(32'h3bf21a60),
	.w5(32'h3bcd885a),
	.w6(32'h3b4ce46f),
	.w7(32'h3bc213fe),
	.w8(32'h3c28a50b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f7ec2),
	.w1(32'h39cd58b2),
	.w2(32'h3a88b62e),
	.w3(32'h3a9f3efd),
	.w4(32'h3b78a9fc),
	.w5(32'h380945b5),
	.w6(32'h3bbe7cab),
	.w7(32'h3c02d2be),
	.w8(32'hba8662c0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390270c8),
	.w1(32'h3a825565),
	.w2(32'hbc88fa3e),
	.w3(32'hba9a2d26),
	.w4(32'hbb0ab00b),
	.w5(32'hbd05938f),
	.w6(32'hba9263e5),
	.w7(32'hb95b2d1b),
	.w8(32'hbcf681fc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd047388),
	.w1(32'hbcac8158),
	.w2(32'hba96450a),
	.w3(32'hbd4c4845),
	.w4(32'hbcb976bc),
	.w5(32'h3acfd7ce),
	.w6(32'hbcf3ca82),
	.w7(32'hbbc626ab),
	.w8(32'h3a353d93),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a256af5),
	.w1(32'h3b8c5f3b),
	.w2(32'hbb09e406),
	.w3(32'hbab0db78),
	.w4(32'hbb3d08c4),
	.w5(32'h3c0b4ab2),
	.w6(32'hbba0311a),
	.w7(32'h3a8677f2),
	.w8(32'h3bcf48a5),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83304b),
	.w1(32'hbb6d8df5),
	.w2(32'h3c277940),
	.w3(32'h3bc6c2b4),
	.w4(32'h39ed3e8d),
	.w5(32'h3c4bca95),
	.w6(32'hbb22285b),
	.w7(32'h3a3ca798),
	.w8(32'h3a7b8200),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d9197),
	.w1(32'h3c3120d2),
	.w2(32'h3b306e61),
	.w3(32'h3c9016b8),
	.w4(32'h3bea21ba),
	.w5(32'h3aef5401),
	.w6(32'h3c0408e5),
	.w7(32'hbaec795f),
	.w8(32'hb9a94958),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0dae1e),
	.w1(32'h3b2442ff),
	.w2(32'h3b09c2f7),
	.w3(32'h3b3d3e7b),
	.w4(32'h38444c52),
	.w5(32'h3b0a28c8),
	.w6(32'hb886c0ad),
	.w7(32'hbb003c1b),
	.w8(32'hba9dc9dc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72716b),
	.w1(32'h3b6d8067),
	.w2(32'h39f2033a),
	.w3(32'h3b19fa0d),
	.w4(32'h3b53a7d0),
	.w5(32'hbb9fd02c),
	.w6(32'hbaa25c31),
	.w7(32'h39052060),
	.w8(32'hbb974b52),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad61a00),
	.w1(32'h3b6f604c),
	.w2(32'h3c4d3d50),
	.w3(32'hbc295d50),
	.w4(32'hbb4c7efa),
	.w5(32'h3b6cd71e),
	.w6(32'hbb7bffef),
	.w7(32'hbb89dedd),
	.w8(32'hbbdbf53b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c567a26),
	.w1(32'h39c18209),
	.w2(32'h3af8e482),
	.w3(32'hbc1231f1),
	.w4(32'hbc24be30),
	.w5(32'hbc0757c3),
	.w6(32'hbca676ed),
	.w7(32'hbc621b85),
	.w8(32'hbaa0db1c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392e722e),
	.w1(32'hbb9a307d),
	.w2(32'hbb021a50),
	.w3(32'hbc56c1c3),
	.w4(32'hbbbf79bb),
	.w5(32'hbb7f73c3),
	.w6(32'hbbb066ce),
	.w7(32'hbb492a5a),
	.w8(32'h3bf636e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc801904),
	.w1(32'hbc577541),
	.w2(32'h3b9e306c),
	.w3(32'hbc88962a),
	.w4(32'hbc22a735),
	.w5(32'h3c897989),
	.w6(32'h3b25f605),
	.w7(32'h3addcefd),
	.w8(32'h3c909e92),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b2097),
	.w1(32'h3c38dad1),
	.w2(32'h3b7fb052),
	.w3(32'h3ca63417),
	.w4(32'h3ccc108a),
	.w5(32'h3a5bec70),
	.w6(32'h3c4ff54d),
	.w7(32'h3c0f2ea7),
	.w8(32'hbaf46a6e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980632c),
	.w1(32'h3b4b43f1),
	.w2(32'hbc2c791e),
	.w3(32'hbb8416c7),
	.w4(32'hbbd8eb0e),
	.w5(32'hbc62d0f9),
	.w6(32'hbbac2bb1),
	.w7(32'hbbfd52e7),
	.w8(32'hbb74e87c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7eae49),
	.w1(32'hbc372327),
	.w2(32'h3c108823),
	.w3(32'hbc8fdefd),
	.w4(32'hbb96ba7a),
	.w5(32'h3b06423b),
	.w6(32'hbbf7bc3e),
	.w7(32'h3c133b2f),
	.w8(32'h3be3ebfb),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb55396),
	.w1(32'h3b4d96ee),
	.w2(32'hbc20cbdc),
	.w3(32'h3ba02548),
	.w4(32'h3a4d2067),
	.w5(32'hbc092a75),
	.w6(32'hb9b70f41),
	.w7(32'h3a1b5c56),
	.w8(32'hbb0bd198),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f81b1),
	.w1(32'hbb5a3cbc),
	.w2(32'h3ab282f3),
	.w3(32'hbaedead3),
	.w4(32'hba8b0336),
	.w5(32'h3c10e679),
	.w6(32'h3ae3f675),
	.w7(32'hbb5dab10),
	.w8(32'h3baee158),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03b77),
	.w1(32'h3b567350),
	.w2(32'hbb58cd37),
	.w3(32'hbb1fc449),
	.w4(32'hbb855687),
	.w5(32'h3aaf823f),
	.w6(32'hbb790d78),
	.w7(32'hba8450de),
	.w8(32'h3c01a458),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010ff2),
	.w1(32'h3a710a92),
	.w2(32'hba439b4d),
	.w3(32'h3be04be2),
	.w4(32'h3c3f3d98),
	.w5(32'h3b688221),
	.w6(32'h3c780ec1),
	.w7(32'h3c41f636),
	.w8(32'h3abe45d8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d9fe6),
	.w1(32'h3bf16e54),
	.w2(32'hbba8460a),
	.w3(32'h3bed0918),
	.w4(32'h3c144da8),
	.w5(32'hbb2a33dc),
	.w6(32'h3c12a0c9),
	.w7(32'h3c0ce9ac),
	.w8(32'h3b4966a5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72bdb5),
	.w1(32'hba95a4d4),
	.w2(32'hbadbc8b3),
	.w3(32'h3ae6079d),
	.w4(32'h3af7d316),
	.w5(32'h3b149adb),
	.w6(32'h3bdcccc9),
	.w7(32'h3bd1949a),
	.w8(32'h3c08c8c8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ad083),
	.w1(32'hb93a4fbb),
	.w2(32'h3c25d9cd),
	.w3(32'hbc0b68c3),
	.w4(32'hba4c7205),
	.w5(32'h3c3a28e7),
	.w6(32'h3b0022ae),
	.w7(32'h3b4c749b),
	.w8(32'h3cafb80f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e172f),
	.w1(32'h3b05dbd6),
	.w2(32'hbc05ae14),
	.w3(32'hbadbeacd),
	.w4(32'hbb143d8d),
	.w5(32'hbbd755e1),
	.w6(32'h3c3c23de),
	.w7(32'hbb574e2a),
	.w8(32'h38a1c05d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0922ac),
	.w1(32'hbc1e8a4b),
	.w2(32'hbc0a8269),
	.w3(32'hbc9a25a4),
	.w4(32'hbb8ec7b1),
	.w5(32'hbc081056),
	.w6(32'h399a1b45),
	.w7(32'h3a8a40c7),
	.w8(32'h3b2750f0),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0384de),
	.w1(32'hbc45bf08),
	.w2(32'h3b73cffc),
	.w3(32'hbc9b2750),
	.w4(32'hbc060dc5),
	.w5(32'h3ae4ad34),
	.w6(32'hbc2a8a4e),
	.w7(32'h3b179071),
	.w8(32'h3bf06282),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc64130),
	.w1(32'h3bdd6b42),
	.w2(32'hbb8fd152),
	.w3(32'h3b85748d),
	.w4(32'h3b88d492),
	.w5(32'hbbd4add0),
	.w6(32'h3c36db2f),
	.w7(32'h3c299290),
	.w8(32'hba57d60e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadee9b),
	.w1(32'hbc09280b),
	.w2(32'hbc32f64c),
	.w3(32'hbc3c29dc),
	.w4(32'hbc153e51),
	.w5(32'hbc9ed6e2),
	.w6(32'hbb583f5b),
	.w7(32'h3ac2d9ff),
	.w8(32'hbad150b3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0dc81),
	.w1(32'hbc9e1565),
	.w2(32'h3c0e43e4),
	.w3(32'hbd05838a),
	.w4(32'hbc9b41db),
	.w5(32'h3b557add),
	.w6(32'hbc360a74),
	.w7(32'hbbc7f971),
	.w8(32'h3bc28a14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae0d2f),
	.w1(32'h3c01235f),
	.w2(32'h3b7d6aa0),
	.w3(32'hbb6ec84b),
	.w4(32'h3ba35066),
	.w5(32'h3b8e01fc),
	.w6(32'h3a9bf539),
	.w7(32'h3b04ef29),
	.w8(32'h3b9c4b40),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba02fe1),
	.w1(32'h3b688b50),
	.w2(32'h3a2e0a9d),
	.w3(32'h3ba36321),
	.w4(32'h3bb021bb),
	.w5(32'h3b8391d5),
	.w6(32'h3b355818),
	.w7(32'h392b800e),
	.w8(32'h3a86df6d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976ea7),
	.w1(32'h3b501013),
	.w2(32'hb9d07a47),
	.w3(32'hba1a19cf),
	.w4(32'hbb6a2ef9),
	.w5(32'hbb047a4f),
	.w6(32'hbbdef1bc),
	.w7(32'hbc15e1b5),
	.w8(32'hba3871c6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7aab8),
	.w1(32'h3b382202),
	.w2(32'h39b636d6),
	.w3(32'hba82c5a8),
	.w4(32'h3aadbd6d),
	.w5(32'h3c80e70e),
	.w6(32'h3ad008e5),
	.w7(32'h3bcb2cc2),
	.w8(32'h3c069550),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b4b8),
	.w1(32'h3c304b71),
	.w2(32'h3ad449c6),
	.w3(32'h3c7694d5),
	.w4(32'h3c69300a),
	.w5(32'hbb42be92),
	.w6(32'h3bd3f101),
	.w7(32'h3a846b4e),
	.w8(32'hb9e76605),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb1810),
	.w1(32'hbb4cdac7),
	.w2(32'hba49950b),
	.w3(32'h3be70955),
	.w4(32'hbad666e5),
	.w5(32'h3b7722e2),
	.w6(32'h3a123fdd),
	.w7(32'h3baa2afb),
	.w8(32'h3c127f7a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97ee73),
	.w1(32'hb9a94f2c),
	.w2(32'h3b05aba6),
	.w3(32'hbb11d5dd),
	.w4(32'hbb27d97e),
	.w5(32'h3982a07d),
	.w6(32'h3c1cfc39),
	.w7(32'h3b91a2f6),
	.w8(32'hbabd9c54),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b248eb6),
	.w1(32'h3b2352b3),
	.w2(32'hbb09eb14),
	.w3(32'hba1900e1),
	.w4(32'h39e4e245),
	.w5(32'hbba04a1b),
	.w6(32'h3a5485b3),
	.w7(32'hbaa2d360),
	.w8(32'hbba9b39f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb402c03),
	.w1(32'hbb223ded),
	.w2(32'hbc93e490),
	.w3(32'hbbe7ad36),
	.w4(32'hbb069b6d),
	.w5(32'hbbe924cb),
	.w6(32'hbb8898d6),
	.w7(32'hba6f5625),
	.w8(32'h3bd4043f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc243563),
	.w1(32'hbae00c5f),
	.w2(32'hbaaca76f),
	.w3(32'h3b9ec9d8),
	.w4(32'h3c046ac8),
	.w5(32'h3a992829),
	.w6(32'h3c5c702f),
	.w7(32'h3c977bb1),
	.w8(32'h3bfc4901),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829755d),
	.w1(32'h3a54fa12),
	.w2(32'hb92f1394),
	.w3(32'h3b685677),
	.w4(32'h3b601712),
	.w5(32'hbb21d8f6),
	.w6(32'h3ba55ac4),
	.w7(32'h3bafd39d),
	.w8(32'h3bc74145),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aa21d),
	.w1(32'h3bc2cb06),
	.w2(32'h3b6c9373),
	.w3(32'h3a374e9e),
	.w4(32'h3c8551c4),
	.w5(32'hba3585de),
	.w6(32'h3c1cde44),
	.w7(32'h3c5f1199),
	.w8(32'hbbc4bc89),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb548ba3),
	.w1(32'hba58630d),
	.w2(32'h3bc4fedc),
	.w3(32'hba9d77d3),
	.w4(32'h3b5a7e42),
	.w5(32'hb97f4926),
	.w6(32'h3b4d2bd4),
	.w7(32'h3b44b568),
	.w8(32'hba2516e7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd55b23),
	.w1(32'hbb23f1eb),
	.w2(32'h3b246b6a),
	.w3(32'hbb1b3590),
	.w4(32'h3a4c7edc),
	.w5(32'hbc525ab2),
	.w6(32'hbc33d47e),
	.w7(32'hba948135),
	.w8(32'h3af50995),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6f760),
	.w1(32'hbba641a0),
	.w2(32'h3c0e20c9),
	.w3(32'hbc5f68a5),
	.w4(32'hbc83f53c),
	.w5(32'h3cb809cc),
	.w6(32'hbab2dbcc),
	.w7(32'h3b9f31a9),
	.w8(32'h3c884b9d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add969a),
	.w1(32'hbbcb0864),
	.w2(32'hbb5c58f8),
	.w3(32'h3c9bb6cf),
	.w4(32'hba16ad76),
	.w5(32'hbbc2aa4d),
	.w6(32'h3cc5a625),
	.w7(32'h3c159ae2),
	.w8(32'h3b9e090b),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9242),
	.w1(32'h3aadf0b0),
	.w2(32'hbc4fded3),
	.w3(32'hbbfa9f82),
	.w4(32'hbb87a192),
	.w5(32'hbc94c6e4),
	.w6(32'hbbe0d38f),
	.w7(32'h390a19b8),
	.w8(32'hbb6dd4a8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca81a89),
	.w1(32'hbba07682),
	.w2(32'hbc3d0048),
	.w3(32'hbce058c2),
	.w4(32'hbc3284d4),
	.w5(32'hb88e6ad3),
	.w6(32'hbb6a08a8),
	.w7(32'hbb4ce808),
	.w8(32'h3b5afb10),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38531cbc),
	.w1(32'h3bb8e58e),
	.w2(32'hbbcfcfe0),
	.w3(32'h3c0e7c1b),
	.w4(32'h3b613d01),
	.w5(32'hbb1744a5),
	.w6(32'h3b2d8683),
	.w7(32'hbb98ebb9),
	.w8(32'hbb88929b),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf55eda),
	.w1(32'hbaaf88b5),
	.w2(32'h3bd2aa2f),
	.w3(32'hbbb186ff),
	.w4(32'h3b834e12),
	.w5(32'h3afc114b),
	.w6(32'hbbb7f80d),
	.w7(32'hbbd10812),
	.w8(32'h3b339993),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1698b7),
	.w1(32'h3b8c11e6),
	.w2(32'hbbcde645),
	.w3(32'hbb35adaa),
	.w4(32'hbaca5c46),
	.w5(32'h3a0a7967),
	.w6(32'hbae90cba),
	.w7(32'h398f70d2),
	.w8(32'h3a7bacda),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fd1f4),
	.w1(32'h3bb073c4),
	.w2(32'hb98438fe),
	.w3(32'h3bdb9335),
	.w4(32'h3b5ee470),
	.w5(32'hb73afc0c),
	.w6(32'h3ab6fd7a),
	.w7(32'h39bdfd7f),
	.w8(32'h3c1f6b2e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce383),
	.w1(32'hbbdf2c4d),
	.w2(32'h3c24f42d),
	.w3(32'h3b26228f),
	.w4(32'h3b2444c4),
	.w5(32'h3c8cb689),
	.w6(32'h3c2d7832),
	.w7(32'h3c1c3b74),
	.w8(32'h3bea4991),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dfe59),
	.w1(32'h3c56d2db),
	.w2(32'h3a409bfa),
	.w3(32'h3c8e4efb),
	.w4(32'h3c194652),
	.w5(32'h3ab0efe1),
	.w6(32'h3b2e5187),
	.w7(32'h3a482f66),
	.w8(32'h3abe3f9a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a412a1f),
	.w1(32'h38ec0ddc),
	.w2(32'hbc3f6e09),
	.w3(32'h3aa8da9c),
	.w4(32'h3b7e91fc),
	.w5(32'hbcca9863),
	.w6(32'h3b3200ba),
	.w7(32'h3af49f2b),
	.w8(32'hbb916efa),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87d244),
	.w1(32'hbc4aa351),
	.w2(32'hbb07111a),
	.w3(32'hbcdfdea8),
	.w4(32'hbc826f8c),
	.w5(32'hbb7f715b),
	.w6(32'hbc7f37a0),
	.w7(32'hb920862e),
	.w8(32'hbc01d70d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d41a4),
	.w1(32'hbbb35745),
	.w2(32'h3c07ad99),
	.w3(32'hbbf03db9),
	.w4(32'hbbb8c042),
	.w5(32'h3c1f392e),
	.w6(32'hbc176769),
	.w7(32'hbc13278f),
	.w8(32'h3c03923d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36e05f),
	.w1(32'h3be196dd),
	.w2(32'hba7c1c0d),
	.w3(32'h3bd07bb1),
	.w4(32'h3c19870e),
	.w5(32'hb9cb37f1),
	.w6(32'h3bff2020),
	.w7(32'h3c5b48a9),
	.w8(32'h3bf29f48),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b9cd4),
	.w1(32'hbbf42412),
	.w2(32'h3b681287),
	.w3(32'hba2e0404),
	.w4(32'hbb8f7e31),
	.w5(32'h3a0cc9ea),
	.w6(32'hb9f98a67),
	.w7(32'hbbaadabc),
	.w8(32'h3b734a68),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9091b3b),
	.w1(32'h3a859f1f),
	.w2(32'hbb0d6fce),
	.w3(32'hbb7777ac),
	.w4(32'hba66939d),
	.w5(32'hba6bf8da),
	.w6(32'h38e34c19),
	.w7(32'h3b063074),
	.w8(32'hbaab3e14),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba35bf8b),
	.w1(32'hbacb3326),
	.w2(32'h3be3f21f),
	.w3(32'h391ef9b1),
	.w4(32'h3ad7d97a),
	.w5(32'h3c5068b1),
	.w6(32'h3a5cbcb1),
	.w7(32'h3ab648dc),
	.w8(32'h3c6f89ec),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1145e4),
	.w1(32'h3c187167),
	.w2(32'hbac6b0b1),
	.w3(32'h3c132924),
	.w4(32'h3ba06e60),
	.w5(32'h3b26093a),
	.w6(32'h3aff2ac1),
	.w7(32'hbbbd1f99),
	.w8(32'h3b867d61),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00493a),
	.w1(32'h3b4cfb0f),
	.w2(32'hbc6ee1fb),
	.w3(32'h3c33a31a),
	.w4(32'h3c0ced76),
	.w5(32'hbc4e0960),
	.w6(32'h3c0981be),
	.w7(32'h3bddf301),
	.w8(32'h3afde93b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc42497),
	.w1(32'hbcb73f9a),
	.w2(32'h3abd4fbb),
	.w3(32'hbcb8e80f),
	.w4(32'hbc96d87c),
	.w5(32'h3b55901b),
	.w6(32'hbc2062e4),
	.w7(32'hba519e69),
	.w8(32'hba230ca5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad75786),
	.w1(32'h3ae85c35),
	.w2(32'h3bb0bf08),
	.w3(32'hbb48fb93),
	.w4(32'hbbe11d9a),
	.w5(32'h3b0748e7),
	.w6(32'hbbd3bba2),
	.w7(32'hbb9896ae),
	.w8(32'h3c2808f8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc544885),
	.w1(32'hbb675725),
	.w2(32'hbba64eb5),
	.w3(32'hbbebaac2),
	.w4(32'hbc31e028),
	.w5(32'hbc2f0ba7),
	.w6(32'h3bd4c986),
	.w7(32'hbb742727),
	.w8(32'h3aa6bdb7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedd9c5),
	.w1(32'hbc309287),
	.w2(32'h3af3815b),
	.w3(32'hbbd23cb9),
	.w4(32'hbb18dfb5),
	.w5(32'h3b4f0200),
	.w6(32'h3b335d55),
	.w7(32'h3bc8ef3e),
	.w8(32'h3b340ba8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e3566b),
	.w1(32'h3b0293b9),
	.w2(32'h3b9013f7),
	.w3(32'h3a3f55ca),
	.w4(32'h3b76f767),
	.w5(32'h3ab15560),
	.w6(32'h3b820115),
	.w7(32'h3b69d1c5),
	.w8(32'h3912af1f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1ee17),
	.w1(32'h3be4fadd),
	.w2(32'hbc6d8ef3),
	.w3(32'h3b88c183),
	.w4(32'h3afd3214),
	.w5(32'hbb9f97b2),
	.w6(32'h3ba3c7a0),
	.w7(32'hba4785cb),
	.w8(32'h3b746232),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca71856),
	.w1(32'hbc4484c4),
	.w2(32'h3c1aa956),
	.w3(32'hbc3b2885),
	.w4(32'hba3a264e),
	.w5(32'h3c4ae457),
	.w6(32'h3b9f807c),
	.w7(32'h3c3842c1),
	.w8(32'h3c86bb1d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830daa),
	.w1(32'h3c40a1e8),
	.w2(32'h388962ba),
	.w3(32'h3cbabead),
	.w4(32'h3c185eca),
	.w5(32'h3b056b5c),
	.w6(32'h3bf6aca3),
	.w7(32'h3b426ed8),
	.w8(32'h3a957815),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114957),
	.w1(32'h3a5cab42),
	.w2(32'h3b9017e8),
	.w3(32'h3b1826c1),
	.w4(32'h3b42c196),
	.w5(32'hba35a334),
	.w6(32'h38c9c8d3),
	.w7(32'h3a64711c),
	.w8(32'h3b9bbb61),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ba82),
	.w1(32'h3b09e710),
	.w2(32'h3c27563f),
	.w3(32'hbc1a52d9),
	.w4(32'h3c19b6a8),
	.w5(32'hbbd31393),
	.w6(32'hbbfb021d),
	.w7(32'h3b87119b),
	.w8(32'hbccff6c8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a22ad),
	.w1(32'h38a845c7),
	.w2(32'h3b497ced),
	.w3(32'h3d0a22ca),
	.w4(32'hbcc1a68d),
	.w5(32'h3b89816c),
	.w6(32'h3c8dce5c),
	.w7(32'h3c2acb67),
	.w8(32'h3b98f475),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff1c3),
	.w1(32'h39ee2d25),
	.w2(32'h3a62ad45),
	.w3(32'h3930f3ca),
	.w4(32'hba5d4cd2),
	.w5(32'h3c4946d2),
	.w6(32'h3b84da3a),
	.w7(32'hbb85cc48),
	.w8(32'h3c3f40a4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb701dc6),
	.w1(32'h3bea0c49),
	.w2(32'h3c27f55b),
	.w3(32'hbb8964fc),
	.w4(32'h3b06b61f),
	.w5(32'h3baa72a9),
	.w6(32'h3b58cc41),
	.w7(32'hbc142ee4),
	.w8(32'h3a7732e3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42fa13),
	.w1(32'h3b3f8641),
	.w2(32'hba850d59),
	.w3(32'h3c2bada2),
	.w4(32'h3ba4a661),
	.w5(32'hba8afc1a),
	.w6(32'h3ba2b3e2),
	.w7(32'h3b085ab3),
	.w8(32'h3af87983),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319966),
	.w1(32'hbb8a81b7),
	.w2(32'hbb420221),
	.w3(32'hbb9be958),
	.w4(32'hbb362dbe),
	.w5(32'h3b03b7d6),
	.w6(32'hbb56e438),
	.w7(32'hbac453e9),
	.w8(32'h3afaeaf7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46c37d),
	.w1(32'hba7db7b6),
	.w2(32'hbb332521),
	.w3(32'hbcba856d),
	.w4(32'hbc4f9867),
	.w5(32'hbaa08428),
	.w6(32'hbc85c523),
	.w7(32'hbc3a1522),
	.w8(32'hbb0d78da),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae39ccd),
	.w1(32'hbb46eaa9),
	.w2(32'hbb900c45),
	.w3(32'h3acbb1c0),
	.w4(32'hb9594d75),
	.w5(32'hba916c7f),
	.w6(32'hbaa3a1d2),
	.w7(32'h3b2f61f8),
	.w8(32'hbbf7e6f2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5ed2c),
	.w1(32'h3bf6356a),
	.w2(32'h3affa1a5),
	.w3(32'hbb97bd9a),
	.w4(32'h3c165f2c),
	.w5(32'h3af71608),
	.w6(32'hbc39cee8),
	.w7(32'h3c36ed53),
	.w8(32'h3b4ecf62),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e624),
	.w1(32'h3a3e9200),
	.w2(32'h3b248fdc),
	.w3(32'hba0edf48),
	.w4(32'h3bc35771),
	.w5(32'hbbddeb25),
	.w6(32'hbb4c6eec),
	.w7(32'h3bba65e1),
	.w8(32'hbc407105),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab051ff),
	.w1(32'hbb019705),
	.w2(32'h3cd34615),
	.w3(32'h3c312a3e),
	.w4(32'hbb96a0d5),
	.w5(32'h3cfe4b95),
	.w6(32'hba73f4bb),
	.w7(32'h3b202091),
	.w8(32'h3c4813c6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc677fa),
	.w1(32'h3bb09c8a),
	.w2(32'hba932951),
	.w3(32'h3ad0eb2a),
	.w4(32'hbc25d797),
	.w5(32'h3b03da5e),
	.w6(32'h3d0d01b6),
	.w7(32'hbcc5cd3f),
	.w8(32'h3affff4d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390214b0),
	.w1(32'h3a1d8d3f),
	.w2(32'hbb4edc2c),
	.w3(32'h3b655458),
	.w4(32'hbb73528f),
	.w5(32'hbbc4d111),
	.w6(32'h3b5626e3),
	.w7(32'hbc0a5326),
	.w8(32'hba897291),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a948eae),
	.w1(32'hba96d904),
	.w2(32'h3c030be7),
	.w3(32'h3bb2c689),
	.w4(32'hbc1e3e04),
	.w5(32'h3b808345),
	.w6(32'h3be599ea),
	.w7(32'hbb9adf88),
	.w8(32'hbb1d8e9f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad5ad5),
	.w1(32'h3a82c734),
	.w2(32'hbb91841c),
	.w3(32'h3be0edaa),
	.w4(32'hbc04e30c),
	.w5(32'hbb1ee6c5),
	.w6(32'h3a0c05e4),
	.w7(32'h3a644772),
	.w8(32'hbb4e0861),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07aaab),
	.w1(32'hba8c61c9),
	.w2(32'hba8eaac3),
	.w3(32'h3a968731),
	.w4(32'h3b8c3f36),
	.w5(32'hbc8be642),
	.w6(32'h3977c73b),
	.w7(32'h3bc31b63),
	.w8(32'hbc9418f7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487fb7),
	.w1(32'hbc6054f8),
	.w2(32'h3c792144),
	.w3(32'h3ca84714),
	.w4(32'hbcc681bc),
	.w5(32'h3cb4a6f6),
	.w6(32'h3c612fab),
	.w7(32'hbba11645),
	.w8(32'h3c0b36dd),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b1677),
	.w1(32'h3c91493f),
	.w2(32'hbc76f4b6),
	.w3(32'hbb917b4f),
	.w4(32'h3c9192c8),
	.w5(32'hbc061df2),
	.w6(32'h3c239e87),
	.w7(32'hbc5cd6ac),
	.w8(32'hbb69ffd3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce82c21),
	.w1(32'h3aa6fc5e),
	.w2(32'hbc68a7dd),
	.w3(32'h3d1ea53f),
	.w4(32'h3d1237a1),
	.w5(32'hbc504c5f),
	.w6(32'h3c020624),
	.w7(32'h3d1226cc),
	.w8(32'hbc0aaac9),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86eca2),
	.w1(32'h3bfad668),
	.w2(32'hba4bb50a),
	.w3(32'hbc147f6a),
	.w4(32'h3b9ba4ea),
	.w5(32'hba52c010),
	.w6(32'hbc3b4eb1),
	.w7(32'h3af10a7e),
	.w8(32'hbb0ddfa2),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c497d),
	.w1(32'h3af015f0),
	.w2(32'hba8fa02c),
	.w3(32'h3b7aac70),
	.w4(32'h3b38c0b3),
	.w5(32'h3a89ecc9),
	.w6(32'h3aba891f),
	.w7(32'h3aa3f45f),
	.w8(32'h3b21a8f6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca79323),
	.w1(32'h3bd817c7),
	.w2(32'h3c48995e),
	.w3(32'hbcca4057),
	.w4(32'hbc05475d),
	.w5(32'h3c444f0e),
	.w6(32'hbc25d78b),
	.w7(32'hbc4dede5),
	.w8(32'hbb2f31f6),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab55b6c),
	.w1(32'hb9fd8967),
	.w2(32'hbb83f210),
	.w3(32'hbbf7fbda),
	.w4(32'hbbc96d80),
	.w5(32'hbbf54d74),
	.w6(32'hb87d7d85),
	.w7(32'hbbc8bb6c),
	.w8(32'hbc616327),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3563ea),
	.w1(32'hbc00f750),
	.w2(32'h3ca6ff52),
	.w3(32'hbbb6bd9e),
	.w4(32'hbc9e6334),
	.w5(32'h3bd975a5),
	.w6(32'h3bc3891a),
	.w7(32'hbbdb7477),
	.w8(32'h3bc00d1b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde43ae),
	.w1(32'h3c898080),
	.w2(32'h3c0a394f),
	.w3(32'h3b51bcf8),
	.w4(32'h3bcccdbc),
	.w5(32'h3b980e87),
	.w6(32'h3c019256),
	.w7(32'h3b40e269),
	.w8(32'h3c2cff60),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58322e),
	.w1(32'h3b80e6bc),
	.w2(32'hbc7b3dff),
	.w3(32'hbba3e7c5),
	.w4(32'hba3309f0),
	.w5(32'hbc33f7cb),
	.w6(32'h3af0e481),
	.w7(32'hbbd41017),
	.w8(32'hbbf77f32),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cd379),
	.w1(32'hbc17814f),
	.w2(32'h3ad94270),
	.w3(32'hbca52dc7),
	.w4(32'hbc684a99),
	.w5(32'hbb98fe0f),
	.w6(32'hbcc04250),
	.w7(32'h3bf17da0),
	.w8(32'hb95f3bd6),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb527815),
	.w1(32'h3aa7a8d1),
	.w2(32'h3c41f195),
	.w3(32'hbc9b8e27),
	.w4(32'hbc2a5558),
	.w5(32'hbc2c1c2b),
	.w6(32'hbb062cca),
	.w7(32'hbc58df2e),
	.w8(32'hbca10b78),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba997da0),
	.w1(32'hba032595),
	.w2(32'hbb18438b),
	.w3(32'h3cdd97c7),
	.w4(32'hbc18d485),
	.w5(32'h38a5f1a7),
	.w6(32'h3cb0d427),
	.w7(32'hbc15f30f),
	.w8(32'hbab378a2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d6b10),
	.w1(32'hbb4b18cf),
	.w2(32'hba9fb0e9),
	.w3(32'h3b0988d4),
	.w4(32'h3b44498e),
	.w5(32'hbb000d95),
	.w6(32'hba975fd0),
	.w7(32'hba077c24),
	.w8(32'h3affed10),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae62e15),
	.w1(32'hbb666d32),
	.w2(32'h39ff50a4),
	.w3(32'hb9dcbed8),
	.w4(32'hbae90fe9),
	.w5(32'hbac52876),
	.w6(32'hb9ecf327),
	.w7(32'hb8c6aee4),
	.w8(32'hbb030c9b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d00c8),
	.w1(32'h3b47ac48),
	.w2(32'hba7b2832),
	.w3(32'hbae3b765),
	.w4(32'hbb862d6b),
	.w5(32'hbb13fa56),
	.w6(32'hbaa92316),
	.w7(32'hbb8e4e64),
	.w8(32'hba5fbd6a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6dfcab),
	.w1(32'h3c3899f1),
	.w2(32'hbc0e0fc1),
	.w3(32'hbc7c2082),
	.w4(32'h3c26b795),
	.w5(32'hba94f2f5),
	.w6(32'hbc1cf836),
	.w7(32'h3addfbce),
	.w8(32'hbc0f0c1c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97592b),
	.w1(32'hbb998bea),
	.w2(32'h3b959821),
	.w3(32'hbba1d15f),
	.w4(32'hbc75d32a),
	.w5(32'hbc430c40),
	.w6(32'h3b7d05e0),
	.w7(32'hbbe3f0f7),
	.w8(32'hba5ee985),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdff0b),
	.w1(32'hbc81bb90),
	.w2(32'h3a516917),
	.w3(32'hba21cde9),
	.w4(32'h3c08848f),
	.w5(32'h3b14cb16),
	.w6(32'hbcb1e1d7),
	.w7(32'h3c80e19e),
	.w8(32'h3c0078c6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38d7b5),
	.w1(32'hbba944b4),
	.w2(32'hbb747f44),
	.w3(32'hbb72224a),
	.w4(32'h3b21033e),
	.w5(32'hbb43fa12),
	.w6(32'hbba6822e),
	.w7(32'hbbd875a7),
	.w8(32'h3b073aaf),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60e82d),
	.w1(32'h3b8938e7),
	.w2(32'h3b11ee78),
	.w3(32'h3aac0185),
	.w4(32'h3c3d496d),
	.w5(32'h39bf1dce),
	.w6(32'h3a7c1c14),
	.w7(32'h3b38936e),
	.w8(32'h3a4375d0),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306569),
	.w1(32'h3b9f6304),
	.w2(32'hbb9b6cd9),
	.w3(32'hbb4ec814),
	.w4(32'h3ad0fa7f),
	.w5(32'hbb43321b),
	.w6(32'hbaca3868),
	.w7(32'h3a428d67),
	.w8(32'h3a0d8a60),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ee12e),
	.w1(32'hbb4824f4),
	.w2(32'h389834e9),
	.w3(32'hbad3588e),
	.w4(32'h3ae20aa4),
	.w5(32'hbb6ebc81),
	.w6(32'hbb49cdb6),
	.w7(32'h3b541384),
	.w8(32'hbb23ccfb),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc651e30),
	.w1(32'hbc8b8d05),
	.w2(32'h3bd4248a),
	.w3(32'hbb975034),
	.w4(32'hbcede640),
	.w5(32'hbb57c05e),
	.w6(32'h3b53eaad),
	.w7(32'hbcaec1b9),
	.w8(32'hbbcf80ca),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5521c4),
	.w1(32'hbb3fcb58),
	.w2(32'h3a940ac7),
	.w3(32'hbbb02ec8),
	.w4(32'hb9da254f),
	.w5(32'hba34553a),
	.w6(32'hbb5a0d70),
	.w7(32'hbbf2dc21),
	.w8(32'hbaa730e7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcada99),
	.w1(32'h3a4611af),
	.w2(32'h3ac3d625),
	.w3(32'hbbe84f6c),
	.w4(32'hbb0a8330),
	.w5(32'hbad61cfd),
	.w6(32'hbba9cd32),
	.w7(32'hbb593c31),
	.w8(32'hbbf0a14e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8c21b),
	.w1(32'hbbec79eb),
	.w2(32'h3a679e8b),
	.w3(32'h3c15b294),
	.w4(32'hbc88b43c),
	.w5(32'h3a63253f),
	.w6(32'h3beee03f),
	.w7(32'hbc144ebd),
	.w8(32'h3b22e2d6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24c1f2),
	.w1(32'h3a6adfc5),
	.w2(32'hbcd4db2f),
	.w3(32'h3bb4be19),
	.w4(32'h3b2fac8d),
	.w5(32'hbc566ec1),
	.w6(32'h3bf18f16),
	.w7(32'h3b648e23),
	.w8(32'hbadb5b3c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6bafa),
	.w1(32'hbc07bf80),
	.w2(32'h3c07c36a),
	.w3(32'h3b7f2f82),
	.w4(32'hb964ddf5),
	.w5(32'h3c13a819),
	.w6(32'hbc34580a),
	.w7(32'h3bccf364),
	.w8(32'h3a2debbe),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf97536),
	.w1(32'h3b854c88),
	.w2(32'hbb77d303),
	.w3(32'hbc3e5015),
	.w4(32'hbcc19784),
	.w5(32'hbb41985b),
	.w6(32'h3bb5dde4),
	.w7(32'hbd114453),
	.w8(32'hbb66e171),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebe12f),
	.w1(32'h3aeee7f1),
	.w2(32'hbabde930),
	.w3(32'h3b12456e),
	.w4(32'h3ab1e8bb),
	.w5(32'hbb843fb0),
	.w6(32'h3b4af1d9),
	.w7(32'h39373087),
	.w8(32'hbb950d99),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d9a3fc),
	.w1(32'hbb85b45e),
	.w2(32'hba70a79e),
	.w3(32'h3b76d914),
	.w4(32'hbab6304f),
	.w5(32'hbc0852b6),
	.w6(32'h3915c5ba),
	.w7(32'h3ade2f9d),
	.w8(32'h362ebd30),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b773f1),
	.w1(32'hba080b3a),
	.w2(32'hb97d7e94),
	.w3(32'h3a09ff57),
	.w4(32'h3b889015),
	.w5(32'hbb309340),
	.w6(32'hbb553895),
	.w7(32'hbb478ce2),
	.w8(32'hbbf91915),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc151660),
	.w1(32'h3c0eb049),
	.w2(32'hbb8ddc60),
	.w3(32'hbba3f19a),
	.w4(32'hbb274b06),
	.w5(32'hbc41fb14),
	.w6(32'h3b27702e),
	.w7(32'hbc2be386),
	.w8(32'hbb7f633d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc357ec),
	.w1(32'hba3338a0),
	.w2(32'h392860f3),
	.w3(32'h3ca3bc9b),
	.w4(32'h3c39a9e6),
	.w5(32'h3afb821e),
	.w6(32'hbc09a21b),
	.w7(32'h3c345c29),
	.w8(32'h3ae8e81c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9913070),
	.w1(32'hb9f7bc4e),
	.w2(32'hbb2dc877),
	.w3(32'h3a7ca5a6),
	.w4(32'hbacdaeb2),
	.w5(32'hbb72e74e),
	.w6(32'h3b639620),
	.w7(32'h3a8ac5f6),
	.w8(32'hba125f1d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b846125),
	.w1(32'hbb9abd13),
	.w2(32'h39e52602),
	.w3(32'h3be882a1),
	.w4(32'hbbe7f67b),
	.w5(32'h3b77bca9),
	.w6(32'h3aeb3365),
	.w7(32'h3ba45cd0),
	.w8(32'h3bd3b1da),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a299f),
	.w1(32'h39f74546),
	.w2(32'hbbb8e09b),
	.w3(32'h3b2269f2),
	.w4(32'h3b965ef0),
	.w5(32'hbbd9a68d),
	.w6(32'h3bad46df),
	.w7(32'h3b2bf3aa),
	.w8(32'h3b9cbd9f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6fb4a5),
	.w1(32'h3c20b2cd),
	.w2(32'hbc3c34a1),
	.w3(32'hbc490f75),
	.w4(32'h3c96af7e),
	.w5(32'hbb90a541),
	.w6(32'hbcb35590),
	.w7(32'h3c622e22),
	.w8(32'h3b3103b7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc87544),
	.w1(32'hbbf22b00),
	.w2(32'h39860a1d),
	.w3(32'h3cb84ba3),
	.w4(32'h3cea44dd),
	.w5(32'hbc6415c3),
	.w6(32'hbbc5336f),
	.w7(32'h3d16de74),
	.w8(32'hbbcef441),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb4024e),
	.w1(32'hbb9d992a),
	.w2(32'hbbaa9b46),
	.w3(32'h3cc53ba7),
	.w4(32'h3c53ca4b),
	.w5(32'hbc8d4b11),
	.w6(32'hbc423e83),
	.w7(32'h3cddf035),
	.w8(32'hbc88ecf5),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71263),
	.w1(32'hbc86ddb0),
	.w2(32'h3b88d2ef),
	.w3(32'hbc87a3f4),
	.w4(32'hbc548caf),
	.w5(32'h3b69f86e),
	.w6(32'hbc030cf7),
	.w7(32'hbc01693c),
	.w8(32'h3b8a6ca0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf74f1f),
	.w1(32'hbbca0246),
	.w2(32'hb9ce78a5),
	.w3(32'hbc07fc4a),
	.w4(32'hbb930a14),
	.w5(32'hbb5e1dc9),
	.w6(32'hbc2929d6),
	.w7(32'hbbbe1e0a),
	.w8(32'hbb09e41a),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de360),
	.w1(32'hbc00433d),
	.w2(32'h3c3cd72f),
	.w3(32'hbbb27117),
	.w4(32'hbc17fbab),
	.w5(32'h3cc98720),
	.w6(32'hbb224c57),
	.w7(32'hbbfcb564),
	.w8(32'h3be7bb19),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc01259),
	.w1(32'h3c7a14b9),
	.w2(32'hbba6dd5f),
	.w3(32'hb9aeb03f),
	.w4(32'h3c14bf3a),
	.w5(32'h3b785fa8),
	.w6(32'h3c264067),
	.w7(32'h3c1c3c72),
	.w8(32'hbbafafb6),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0462e5),
	.w1(32'h3b9c0a25),
	.w2(32'h3a53c859),
	.w3(32'hbc043938),
	.w4(32'h3b80be70),
	.w5(32'h3ab2b1d6),
	.w6(32'h3bd161ae),
	.w7(32'hbb0b2de5),
	.w8(32'hbb046bf2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a6b3f3),
	.w1(32'h3b90e926),
	.w2(32'h3ac75993),
	.w3(32'h3badb0d6),
	.w4(32'h3c3be1c4),
	.w5(32'h3b6de3a4),
	.w6(32'h3bb0c29e),
	.w7(32'h3b916008),
	.w8(32'h3b9cafe7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90559c),
	.w1(32'h3c47a93f),
	.w2(32'hbb2457d4),
	.w3(32'hbbd706f7),
	.w4(32'h3c5d2d68),
	.w5(32'hbbb12517),
	.w6(32'hbbf97134),
	.w7(32'h3bbb350b),
	.w8(32'hbbf1ccce),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc29c8),
	.w1(32'hbc256291),
	.w2(32'hba9dca0e),
	.w3(32'hbc08d48d),
	.w4(32'hbc24695e),
	.w5(32'h3a091e5d),
	.w6(32'hbc2a3f99),
	.w7(32'hbc26176c),
	.w8(32'h3b15beff),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb436bc1),
	.w1(32'hbadd37cd),
	.w2(32'hbb04afbb),
	.w3(32'hbaaec1bd),
	.w4(32'hbb00ea06),
	.w5(32'h3a3f3e24),
	.w6(32'h3b7e9148),
	.w7(32'hbb24f9e9),
	.w8(32'hbb17deb8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc9a5),
	.w1(32'h3a90d9a3),
	.w2(32'hbbd427fd),
	.w3(32'hbb4626cb),
	.w4(32'hbb8855b8),
	.w5(32'h3bd0a74b),
	.w6(32'hbbbf5893),
	.w7(32'hbc0ba04d),
	.w8(32'h39866fdb),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6a83a),
	.w1(32'hbb0e78d1),
	.w2(32'hbb9ffc77),
	.w3(32'h3bac2ed7),
	.w4(32'h3ba36d18),
	.w5(32'hbc3072f1),
	.w6(32'hbb42a4ce),
	.w7(32'h3a627702),
	.w8(32'hbba55191),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9740f6),
	.w1(32'hbb3cfa21),
	.w2(32'h3b75517d),
	.w3(32'hbc7c8af0),
	.w4(32'hbc7798b6),
	.w5(32'hbc3a2b8a),
	.w6(32'hbb19d9c9),
	.w7(32'h3a80e1a5),
	.w8(32'h3b0d8ba5),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cedad6b),
	.w1(32'hbc17df78),
	.w2(32'h3b0eab2e),
	.w3(32'h3cc76ff7),
	.w4(32'h3bcbb1b3),
	.w5(32'h3c0c9636),
	.w6(32'hbc9c7750),
	.w7(32'h3d049c04),
	.w8(32'h3b6fb71e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1055e1),
	.w1(32'h3aa73911),
	.w2(32'hbba0124d),
	.w3(32'hbc54059c),
	.w4(32'hbb244381),
	.w5(32'hbc0dbfe2),
	.w6(32'h3bc5001b),
	.w7(32'hbb803ed6),
	.w8(32'hbbdee4f8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a143def),
	.w1(32'hbb648cba),
	.w2(32'h3c145629),
	.w3(32'h3abfeaa5),
	.w4(32'hbbe8f40d),
	.w5(32'h3c1cdeea),
	.w6(32'hb8dc2d13),
	.w7(32'hbb702b0a),
	.w8(32'h3b09caeb),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba05f20),
	.w1(32'h3b3d6326),
	.w2(32'hbacbc0c5),
	.w3(32'hbb51109d),
	.w4(32'hb7f2205e),
	.w5(32'h3bafb89a),
	.w6(32'h3c8206a9),
	.w7(32'hbc54e535),
	.w8(32'hbbbc51d4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b9016),
	.w1(32'h3c13974d),
	.w2(32'hb889cef4),
	.w3(32'hbb00c98a),
	.w4(32'hba8d7615),
	.w5(32'h3b5e6176),
	.w6(32'h3c16ffa1),
	.w7(32'h3bd4b2c5),
	.w8(32'h3bf80128),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0daaed),
	.w1(32'hb76d6c49),
	.w2(32'h3b1ce86c),
	.w3(32'hbbbb5bbe),
	.w4(32'hbaa99540),
	.w5(32'hb903efcf),
	.w6(32'h390af7aa),
	.w7(32'hbbbeef0e),
	.w8(32'h3b185050),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a236e),
	.w1(32'hbc592687),
	.w2(32'hbc1b2229),
	.w3(32'hb99206f0),
	.w4(32'hbc17701f),
	.w5(32'hbc21d357),
	.w6(32'h3b2ddb52),
	.w7(32'hbab1a5d2),
	.w8(32'hbc804938),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c3e4c),
	.w1(32'hbc87b8cc),
	.w2(32'hbb7237d0),
	.w3(32'hbbb2a6fd),
	.w4(32'hbbf3ad92),
	.w5(32'hbb7c5cee),
	.w6(32'hbb84c4dd),
	.w7(32'hbbd613da),
	.w8(32'hb949fd96),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26f0b2),
	.w1(32'hbb1b8593),
	.w2(32'hbbb50b19),
	.w3(32'hbb99725a),
	.w4(32'hbaffad57),
	.w5(32'hbbd7b824),
	.w6(32'hbb408233),
	.w7(32'h3b5b153a),
	.w8(32'hbb4b03a8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb906613),
	.w1(32'hbb8d053c),
	.w2(32'hbc225686),
	.w3(32'h399d8f22),
	.w4(32'h39e32be5),
	.w5(32'hbc43ab2e),
	.w6(32'hbbfc371a),
	.w7(32'h3bfaa16e),
	.w8(32'hbc1e82b5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c385dd7),
	.w1(32'hbc6200bb),
	.w2(32'hbb83211d),
	.w3(32'h3c389a0a),
	.w4(32'hbc1179f8),
	.w5(32'hbc594566),
	.w6(32'h3b99c6df),
	.w7(32'h3ba177e7),
	.w8(32'hbcb13747),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6be3b7),
	.w1(32'hbc2fa6f6),
	.w2(32'hbbf48494),
	.w3(32'h3d0d3fd6),
	.w4(32'hbc696255),
	.w5(32'hbc557a34),
	.w6(32'h3d08b960),
	.w7(32'h3b86500c),
	.w8(32'hba824858),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc950dec),
	.w1(32'hbb7dab38),
	.w2(32'h3b1938c1),
	.w3(32'hbc3f004a),
	.w4(32'hbc7e2f57),
	.w5(32'hbc5d7f09),
	.w6(32'hbbc0720e),
	.w7(32'hbc8203b5),
	.w8(32'hbc552129),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b17fe),
	.w1(32'hbc6c5c04),
	.w2(32'hbbd7bcf4),
	.w3(32'h3bfae1c1),
	.w4(32'hbc309095),
	.w5(32'hbc4b7444),
	.w6(32'hbc227f11),
	.w7(32'h3bd8cd49),
	.w8(32'hbc7b4697),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf305ee),
	.w1(32'hbbe060eb),
	.w2(32'hbae99c88),
	.w3(32'h3aaad9e3),
	.w4(32'hbc30db5f),
	.w5(32'hbada2b34),
	.w6(32'hbb07f8ea),
	.w7(32'hba862727),
	.w8(32'h3b9fb636),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05d23a),
	.w1(32'h3a3327cc),
	.w2(32'hb9e5f320),
	.w3(32'h3ae1edec),
	.w4(32'h3bd14c16),
	.w5(32'h3a46baaa),
	.w6(32'hbb05b583),
	.w7(32'h3b5a9e79),
	.w8(32'hbb035b50),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8e449),
	.w1(32'hba0de3bb),
	.w2(32'h3c025800),
	.w3(32'hbb72f6f2),
	.w4(32'h3b7b6b2d),
	.w5(32'hb9823cc1),
	.w6(32'h3b1e53d3),
	.w7(32'h39c032bd),
	.w8(32'hbb289e21),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11ce2c),
	.w1(32'hbb9ccba5),
	.w2(32'h3c0ef68f),
	.w3(32'h3c741e4a),
	.w4(32'hbbcb4e8c),
	.w5(32'h3bed67f2),
	.w6(32'h3c807536),
	.w7(32'hbbb350ef),
	.w8(32'h3a3cc271),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054749),
	.w1(32'h3a5f5197),
	.w2(32'h3ad2f23a),
	.w3(32'h3c2fee46),
	.w4(32'hbb70804e),
	.w5(32'h3ae734c8),
	.w6(32'h3c220e31),
	.w7(32'hbae1270c),
	.w8(32'h3b58ffe1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98417bb),
	.w1(32'h3b151079),
	.w2(32'h3b2eef53),
	.w3(32'hbb8d6e47),
	.w4(32'hb993e768),
	.w5(32'hbb7bffcc),
	.w6(32'h3b80b629),
	.w7(32'h3b945ea4),
	.w8(32'hbaa12f41),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d2ad),
	.w1(32'h3b82509a),
	.w2(32'h3bfa65b6),
	.w3(32'h3aa2255e),
	.w4(32'hba199f3a),
	.w5(32'h3c7d7176),
	.w6(32'h3b37b53a),
	.w7(32'hbb75ff3a),
	.w8(32'h3b92f145),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5b8eb),
	.w1(32'h3c862dfb),
	.w2(32'h3b0c9968),
	.w3(32'h3b904b88),
	.w4(32'hba78a4d8),
	.w5(32'h3c17ddfb),
	.w6(32'h3cbe9ae5),
	.w7(32'h3b561842),
	.w8(32'h3be98a15),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68859b),
	.w1(32'h3c61b0ab),
	.w2(32'hbafa5698),
	.w3(32'h3ad6e846),
	.w4(32'h3bac030f),
	.w5(32'hbbdd18a7),
	.w6(32'h3c23b67d),
	.w7(32'h3bdca65f),
	.w8(32'hbb340e77),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2287d7),
	.w1(32'hbbfe9915),
	.w2(32'hbad9b0cc),
	.w3(32'hbc5f6c83),
	.w4(32'hbc4da9bf),
	.w5(32'hb95442f2),
	.w6(32'hbcbaadab),
	.w7(32'hb9a1f4a0),
	.w8(32'hbaa8c1a3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39ebf1),
	.w1(32'hbbd01bad),
	.w2(32'h3ae43829),
	.w3(32'hbb0b5b8e),
	.w4(32'hbba3a3d2),
	.w5(32'h3b26df79),
	.w6(32'hbae4b5b2),
	.w7(32'hbbd668c6),
	.w8(32'h3b1964c5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce1c11),
	.w1(32'h389a19fc),
	.w2(32'hbbaf745c),
	.w3(32'h3aa5d8aa),
	.w4(32'hbb31b04f),
	.w5(32'h3c813b86),
	.w6(32'h3b4b9f8b),
	.w7(32'hbb46e7f2),
	.w8(32'h3d00ba31),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b84ed),
	.w1(32'h3ca81d5a),
	.w2(32'h3bc04785),
	.w3(32'hbd001b39),
	.w4(32'h3d142869),
	.w5(32'h3bc7e2f7),
	.w6(32'hbcfc7dd5),
	.w7(32'h3c8a9bfa),
	.w8(32'h3bd40917),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384455a8),
	.w1(32'h3bfd8392),
	.w2(32'hba10649c),
	.w3(32'hbb513f98),
	.w4(32'h3bc3314c),
	.w5(32'hbb31d0e4),
	.w6(32'hbb4059c5),
	.w7(32'h3af34589),
	.w8(32'h39927e0e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4d8e4),
	.w1(32'hbb9f6551),
	.w2(32'hbcad0870),
	.w3(32'hbbc42b76),
	.w4(32'hbc089bce),
	.w5(32'hbc3054c1),
	.w6(32'h3b2ae703),
	.w7(32'hbbeaebca),
	.w8(32'hbbd1752f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0da5e9),
	.w1(32'hbccba179),
	.w2(32'hbc932211),
	.w3(32'h3c04e361),
	.w4(32'hbcc5f911),
	.w5(32'hbc3247a8),
	.w6(32'h3bde43a9),
	.w7(32'hbc854f14),
	.w8(32'h3ab71adc),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e3e66),
	.w1(32'hbc8c28b1),
	.w2(32'h3be1232e),
	.w3(32'hbc2c04d3),
	.w4(32'hbca3b48c),
	.w5(32'hbb7dc87d),
	.w6(32'h399946f8),
	.w7(32'hbbc15c90),
	.w8(32'hbbeaf9d7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule