module layer_10_featuremap_254(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7334b8),
	.w1(32'h3b9d3bc3),
	.w2(32'h3b95fe19),
	.w3(32'hbb364cf4),
	.w4(32'hbac22116),
	.w5(32'hba01c208),
	.w6(32'hbb4eb982),
	.w7(32'hbafa1ea4),
	.w8(32'h3b53f4e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28af97),
	.w1(32'h3b7e15af),
	.w2(32'hb9b53843),
	.w3(32'hba9e3d8a),
	.w4(32'hbb42f3c1),
	.w5(32'h3b6f0609),
	.w6(32'hba122f61),
	.w7(32'hbb00a350),
	.w8(32'hbb1464a7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ab4b9),
	.w1(32'hbbe5faeb),
	.w2(32'hbaaac7e7),
	.w3(32'h3a9e448a),
	.w4(32'h3be7996e),
	.w5(32'hbaa89dee),
	.w6(32'hbba50fcc),
	.w7(32'hbc0e8263),
	.w8(32'hba8eb7cd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ef5e80),
	.w1(32'hba1e9f92),
	.w2(32'h3a724245),
	.w3(32'hb9cc3377),
	.w4(32'hb9c25725),
	.w5(32'hb95d5780),
	.w6(32'h3b05c735),
	.w7(32'h393e5e09),
	.w8(32'h3be52e7a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd97dd1),
	.w1(32'h3acaf1a7),
	.w2(32'hbb489cac),
	.w3(32'hbb4ca258),
	.w4(32'hbb3bc912),
	.w5(32'hbba31070),
	.w6(32'h3c200499),
	.w7(32'h3bec6db0),
	.w8(32'h3a5aa614),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0845b),
	.w1(32'h3b170061),
	.w2(32'h3aee370c),
	.w3(32'hbb4ba90b),
	.w4(32'hbb21267d),
	.w5(32'hbb516655),
	.w6(32'h3ae1a48a),
	.w7(32'h3acf60a2),
	.w8(32'hb9908827),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9881),
	.w1(32'hbb62a434),
	.w2(32'hbb5e8f9c),
	.w3(32'hbb2f3426),
	.w4(32'hbb8aa32b),
	.w5(32'hbc101548),
	.w6(32'h3952db30),
	.w7(32'hbbb33b0e),
	.w8(32'hbc12bec3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc97bc09),
	.w1(32'hbb03d90e),
	.w2(32'h3b4c5862),
	.w3(32'hbc841048),
	.w4(32'hbc02c0b4),
	.w5(32'hbb1fc449),
	.w6(32'hbc51d531),
	.w7(32'hbb0a1fb7),
	.w8(32'h3b162007),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b027288),
	.w1(32'h3b67ead9),
	.w2(32'h3b793adb),
	.w3(32'hbabb62fd),
	.w4(32'hba6a8fe6),
	.w5(32'hbb77dd47),
	.w6(32'h3adb71dd),
	.w7(32'h3aa27d50),
	.w8(32'h3ad9adcf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b5cc),
	.w1(32'h3b96db28),
	.w2(32'h3ab3e9da),
	.w3(32'hbb20f8b3),
	.w4(32'hbae6cb78),
	.w5(32'hbbb1026e),
	.w6(32'h3b5c72b6),
	.w7(32'h3a147c93),
	.w8(32'h3b32ccf9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5dcee),
	.w1(32'h3b7311b3),
	.w2(32'h3ba68c29),
	.w3(32'hbb5702d0),
	.w4(32'hbb211b73),
	.w5(32'hbb821448),
	.w6(32'h3bbbd750),
	.w7(32'h3b53f9ff),
	.w8(32'h3b3e8675),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b5d0),
	.w1(32'h3a7acd6f),
	.w2(32'h3b03f8ed),
	.w3(32'hbb0d0019),
	.w4(32'hbaac2844),
	.w5(32'hbbc54bdd),
	.w6(32'h3c19680f),
	.w7(32'h3bb68b12),
	.w8(32'hbb9efbd7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c7502),
	.w1(32'hba451f29),
	.w2(32'hbb9ecf95),
	.w3(32'hbb2d6254),
	.w4(32'hbb93d124),
	.w5(32'h39f36fbd),
	.w6(32'hba6cfe1d),
	.w7(32'hbb3e1bde),
	.w8(32'hb9b42d89),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1910),
	.w1(32'hbbb66374),
	.w2(32'hbba9d4cb),
	.w3(32'hbb88645c),
	.w4(32'hbbf2b451),
	.w5(32'hbb06f949),
	.w6(32'hbb36a359),
	.w7(32'hbbf38628),
	.w8(32'hba8da9d8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c5df7),
	.w1(32'h3a2753ea),
	.w2(32'h3a9011ee),
	.w3(32'h398ff4a2),
	.w4(32'hb93d347d),
	.w5(32'hbb90f260),
	.w6(32'hb9ca8b85),
	.w7(32'hb9a2c804),
	.w8(32'hb79db638),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfc0d),
	.w1(32'h3b88e0fe),
	.w2(32'h3a23daec),
	.w3(32'hbb8a191c),
	.w4(32'h397ee332),
	.w5(32'h3a3fd056),
	.w6(32'hbb89ae39),
	.w7(32'hbb5f2e89),
	.w8(32'h3ad582ff),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be05456),
	.w1(32'h3b8c399c),
	.w2(32'h3b703ab1),
	.w3(32'h3a373862),
	.w4(32'h3ae2c7ca),
	.w5(32'hba88a581),
	.w6(32'h3b88b446),
	.w7(32'h3baaa988),
	.w8(32'hba1e5c39),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07c86),
	.w1(32'hbb708ac4),
	.w2(32'hbb7c1685),
	.w3(32'hbc1010f8),
	.w4(32'hbbbc05ac),
	.w5(32'hbb19d09f),
	.w6(32'hbbb5ab17),
	.w7(32'hbac84664),
	.w8(32'h39a89104),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0527e),
	.w1(32'hbb741705),
	.w2(32'hbaccb160),
	.w3(32'hbb1ff563),
	.w4(32'hb795b3c1),
	.w5(32'hbaed3a38),
	.w6(32'h396b6081),
	.w7(32'h3aa6ce00),
	.w8(32'h3b7cd771),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88b3f2),
	.w1(32'hb9365fca),
	.w2(32'hba6a3ea7),
	.w3(32'h391692cc),
	.w4(32'hbb23a934),
	.w5(32'hba77347e),
	.w6(32'h3ba34101),
	.w7(32'h3beb02f1),
	.w8(32'h3b8fb66a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39c616),
	.w1(32'h395bd288),
	.w2(32'hba844016),
	.w3(32'h3ac3b994),
	.w4(32'h3aca6673),
	.w5(32'hb9c9bc08),
	.w6(32'h3a9b39c7),
	.w7(32'h3ac0441b),
	.w8(32'hb87a8db4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a241756),
	.w1(32'h3a612c25),
	.w2(32'h3af864b5),
	.w3(32'hba3cefe4),
	.w4(32'h398e092e),
	.w5(32'hba998752),
	.w6(32'h38918068),
	.w7(32'h3a277aca),
	.w8(32'h3a8b2a2b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f3da4),
	.w1(32'hbb8cd054),
	.w2(32'h3b358543),
	.w3(32'hbc36e387),
	.w4(32'hbb3ce97e),
	.w5(32'hbaf3f41a),
	.w6(32'hba36ef26),
	.w7(32'h39b31602),
	.w8(32'h3b7996af),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ea2c),
	.w1(32'h3b06cf5f),
	.w2(32'hba4018b1),
	.w3(32'h3bccd672),
	.w4(32'h3a3c4327),
	.w5(32'h3bccb362),
	.w6(32'h3bd2dc94),
	.w7(32'h3b2f8ab8),
	.w8(32'hbbd73e85),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0285d1),
	.w1(32'h3bdb8358),
	.w2(32'h3b9323dc),
	.w3(32'h3c5ce5e7),
	.w4(32'h3c367166),
	.w5(32'hbaa844ff),
	.w6(32'hbaaa8a46),
	.w7(32'hbc2ba5ee),
	.w8(32'h39848f62),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57bd7a),
	.w1(32'h3b23a70c),
	.w2(32'h3b77b210),
	.w3(32'hbaba3aa1),
	.w4(32'h3a949ba8),
	.w5(32'h3b2c82a4),
	.w6(32'h3aec1b33),
	.w7(32'h3b5dc478),
	.w8(32'hbb040b0d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb915968),
	.w1(32'hbb1bdd24),
	.w2(32'hbb212e5e),
	.w3(32'h3b2f4b90),
	.w4(32'h3b7e8706),
	.w5(32'h38b0013b),
	.w6(32'h3b347feb),
	.w7(32'h3a9db1eb),
	.w8(32'h3b44a2fd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cef7b),
	.w1(32'h3bc09ef5),
	.w2(32'h3a39cbd4),
	.w3(32'h3b86920b),
	.w4(32'h3a82cb82),
	.w5(32'hbb649035),
	.w6(32'hba713f5e),
	.w7(32'hba33ebc1),
	.w8(32'hbbae48d8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bbc3e),
	.w1(32'hbb4159d9),
	.w2(32'hbb784721),
	.w3(32'hbb8e17e2),
	.w4(32'hbb6b4d90),
	.w5(32'hbaec8249),
	.w6(32'hbbd19e06),
	.w7(32'hbbeeb4f7),
	.w8(32'hb97cdc49),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59a9fe),
	.w1(32'h3ae89f0e),
	.w2(32'h3b26b18b),
	.w3(32'h3b922a09),
	.w4(32'h3aef2480),
	.w5(32'hbb1f7219),
	.w6(32'h3b24cb6a),
	.w7(32'h3b49c732),
	.w8(32'h3b984a90),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4512b),
	.w1(32'hbb5f8d76),
	.w2(32'hbb3a98fa),
	.w3(32'hbb7e9152),
	.w4(32'hbb34c4ab),
	.w5(32'h3ac09aad),
	.w6(32'h3b0f58ee),
	.w7(32'h3a0a02fa),
	.w8(32'hbb8cfe7b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e5399),
	.w1(32'hbae3cdb6),
	.w2(32'h398f87df),
	.w3(32'h3afeaca2),
	.w4(32'h39d44f72),
	.w5(32'hbb926f81),
	.w6(32'hbb7c874e),
	.w7(32'hbb8758c3),
	.w8(32'hbbe56fc6),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5dc59),
	.w1(32'h3b64f2a5),
	.w2(32'h3b8e8907),
	.w3(32'hbbd2eb6f),
	.w4(32'h3af40bac),
	.w5(32'hbb169301),
	.w6(32'hbb018c83),
	.w7(32'h3b0c2487),
	.w8(32'h3a05a5fe),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2be2e),
	.w1(32'h3911cb7f),
	.w2(32'hbb600e1b),
	.w3(32'hbb359d71),
	.w4(32'hbb673e4b),
	.w5(32'hbb0d3069),
	.w6(32'hbb6a069f),
	.w7(32'hbb40896b),
	.w8(32'hbbd1f839),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1811fb),
	.w1(32'h3a68f36b),
	.w2(32'h3b7654f0),
	.w3(32'hba496f3c),
	.w4(32'h3afcdd9e),
	.w5(32'h3b8e69a2),
	.w6(32'hbb996af6),
	.w7(32'hbb99f259),
	.w8(32'h3b30f8b4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79942c),
	.w1(32'h3bc73802),
	.w2(32'h3b815015),
	.w3(32'h3baf9555),
	.w4(32'h3b73ec70),
	.w5(32'hbb3da6d7),
	.w6(32'h3b06477d),
	.w7(32'h3b28489c),
	.w8(32'hbae223a9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f3846),
	.w1(32'hbb80ab09),
	.w2(32'h3bd89d01),
	.w3(32'hbc45502e),
	.w4(32'h3b9d9487),
	.w5(32'hba263aa7),
	.w6(32'hbb747fb7),
	.w7(32'h3ac4eb81),
	.w8(32'hbbafe6c2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c047d10),
	.w1(32'h3b270fb9),
	.w2(32'hba3d8f05),
	.w3(32'h3adff5da),
	.w4(32'h3a15d84d),
	.w5(32'hbb90cda4),
	.w6(32'h3b9ea29a),
	.w7(32'h3bdd6af5),
	.w8(32'hbace08dd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a5ad),
	.w1(32'h3b07e763),
	.w2(32'hbbc6f6dd),
	.w3(32'h3a32482a),
	.w4(32'hbb712cbe),
	.w5(32'hbbb59194),
	.w6(32'h3b183d63),
	.w7(32'h39b84976),
	.w8(32'hbc0ae9cf),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c4fec),
	.w1(32'h3b4875da),
	.w2(32'h3add00fa),
	.w3(32'h39064142),
	.w4(32'h3a09f054),
	.w5(32'h3a055737),
	.w6(32'hbb84080d),
	.w7(32'hbbb8cbe6),
	.w8(32'h3b217652),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4012d3),
	.w1(32'hb995224a),
	.w2(32'h3b1fc341),
	.w3(32'hb9fed516),
	.w4(32'hbb634d33),
	.w5(32'hba88e9b8),
	.w6(32'h3b423d17),
	.w7(32'h3997a7a4),
	.w8(32'h3b1bfe57),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b713253),
	.w1(32'h3a65a84d),
	.w2(32'h3b2b80b7),
	.w3(32'hbb02af93),
	.w4(32'hb9887ef3),
	.w5(32'hbb01d3f8),
	.w6(32'h3b11b692),
	.w7(32'h3b372361),
	.w8(32'hbafc8ec3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc00ad),
	.w1(32'hbb178462),
	.w2(32'hbb12a6b6),
	.w3(32'hbafb514b),
	.w4(32'hb67e4f59),
	.w5(32'hbadd10bf),
	.w6(32'hbafba16f),
	.w7(32'h3ae63c83),
	.w8(32'h3abda113),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb355729),
	.w1(32'hba09c85d),
	.w2(32'hbbc1c3b0),
	.w3(32'hba8fcd49),
	.w4(32'h3b429c1c),
	.w5(32'hbaf96a53),
	.w6(32'h3c201d70),
	.w7(32'h3c1c3f6c),
	.w8(32'hbb3ae000),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0c5f7),
	.w1(32'h3b30d455),
	.w2(32'h3b6cb0d7),
	.w3(32'h3b83706b),
	.w4(32'h3b981710),
	.w5(32'h3b38970f),
	.w6(32'h3a37a204),
	.w7(32'h3ac17155),
	.w8(32'h3a5a4385),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacea156),
	.w1(32'hbb444c72),
	.w2(32'hbab7ff26),
	.w3(32'h3bec235d),
	.w4(32'h3baa102a),
	.w5(32'hb9005451),
	.w6(32'h3b212979),
	.w7(32'h3b85eeee),
	.w8(32'hba0efcc3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189d2f),
	.w1(32'hba8eda0e),
	.w2(32'h38b5e6c3),
	.w3(32'hbb5dfc0f),
	.w4(32'hba275e42),
	.w5(32'hba8d3c76),
	.w6(32'hb98e0ba0),
	.w7(32'hba0841f5),
	.w8(32'h3b29b2fa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ce84),
	.w1(32'h394f00ee),
	.w2(32'h3b75530e),
	.w3(32'hbc274ecf),
	.w4(32'hbb9cacfe),
	.w5(32'hbb42a888),
	.w6(32'hba8d7264),
	.w7(32'h3a233ea9),
	.w8(32'h3a9a0d8d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18ef28),
	.w1(32'h3baff972),
	.w2(32'h3abe3406),
	.w3(32'hba80f077),
	.w4(32'hbb8724ce),
	.w5(32'hbb2f09cc),
	.w6(32'hb8b31238),
	.w7(32'h38e893a2),
	.w8(32'h395cb0f4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba182034),
	.w1(32'hba6fb551),
	.w2(32'h3a024aff),
	.w3(32'hbb37022a),
	.w4(32'h3a1913de),
	.w5(32'hbba47902),
	.w6(32'h3a56bac6),
	.w7(32'hb993754b),
	.w8(32'hbb87936c),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe4601),
	.w1(32'hbb2ec244),
	.w2(32'hbb90fb0e),
	.w3(32'h3b4cd1d4),
	.w4(32'hbac8008f),
	.w5(32'hba3b99af),
	.w6(32'h3a905547),
	.w7(32'hbab54594),
	.w8(32'h3ba79de0),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb618d2),
	.w1(32'hbb91a512),
	.w2(32'hbb8fc7e4),
	.w3(32'hbac3cc59),
	.w4(32'hbb6fabaf),
	.w5(32'hbbc883a6),
	.w6(32'h3bf6c748),
	.w7(32'h3c0ab2ac),
	.w8(32'h3baaa9ca),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9356d1),
	.w1(32'h3b9f8d47),
	.w2(32'h3b6c9d96),
	.w3(32'hba4c9e9e),
	.w4(32'hbae8c5ef),
	.w5(32'hb940193c),
	.w6(32'h3c089f3e),
	.w7(32'h3b866c7b),
	.w8(32'h3aa97225),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5e381),
	.w1(32'hbb764729),
	.w2(32'h3b19455a),
	.w3(32'hbc1879ec),
	.w4(32'hbbb8bf6a),
	.w5(32'hbb189cb8),
	.w6(32'hbb87df98),
	.w7(32'hbb52a3dc),
	.w8(32'h3c333c34),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be09ec9),
	.w1(32'h3b8707fb),
	.w2(32'h3988255a),
	.w3(32'hb7a0891f),
	.w4(32'hbb67d3fd),
	.w5(32'hbab88fab),
	.w6(32'h3c3cd99d),
	.w7(32'h3c5f9210),
	.w8(32'hbbfda893),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862f6f),
	.w1(32'hbbfeede8),
	.w2(32'hbbab06f4),
	.w3(32'hb960bbe6),
	.w4(32'h3aabcad9),
	.w5(32'h3b5ede75),
	.w6(32'hbc02cdc9),
	.w7(32'hbbac1190),
	.w8(32'hba04f934),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a826ca2),
	.w1(32'h3af3d9f0),
	.w2(32'h3b7eeee5),
	.w3(32'h3bca4568),
	.w4(32'h3b94e388),
	.w5(32'hba9524a9),
	.w6(32'h39f34d5b),
	.w7(32'h3b0943f6),
	.w8(32'hba5b5be3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b124b19),
	.w1(32'h3ab9d434),
	.w2(32'h3ac11832),
	.w3(32'hb9909232),
	.w4(32'hb9ab1557),
	.w5(32'hbb36cdb9),
	.w6(32'h3b4ba73d),
	.w7(32'h39d24f1e),
	.w8(32'h3a8fab37),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad582bc),
	.w1(32'h3af15963),
	.w2(32'h3b2d2249),
	.w3(32'hbb4e19d1),
	.w4(32'hb9528b3c),
	.w5(32'h3b47957e),
	.w6(32'h3b05be15),
	.w7(32'h3a8727d5),
	.w8(32'h3bb06b07),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be852),
	.w1(32'h3b6aed51),
	.w2(32'h3b729872),
	.w3(32'hbafa024d),
	.w4(32'h393e232d),
	.w5(32'hbb52f76b),
	.w6(32'h3bb2ef9b),
	.w7(32'h3bb83af9),
	.w8(32'hbb19797f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68d7ed),
	.w1(32'hbb477d3b),
	.w2(32'hbb909b43),
	.w3(32'hbbcda1b4),
	.w4(32'hbb5c9f59),
	.w5(32'hbb7dbbd2),
	.w6(32'hbb7fb50a),
	.w7(32'hb98c403c),
	.w8(32'hb9b3613f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01f15c),
	.w1(32'h3b4b87ab),
	.w2(32'hba3bb78d),
	.w3(32'hbb920081),
	.w4(32'hbb0b18d6),
	.w5(32'hbb8d77e5),
	.w6(32'hbb85367b),
	.w7(32'hbaa62edc),
	.w8(32'h3b1cf200),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39582d71),
	.w1(32'hbb27b478),
	.w2(32'hba80ab71),
	.w3(32'hbaacb462),
	.w4(32'h39e34fc6),
	.w5(32'hba136f9c),
	.w6(32'h3b26f451),
	.w7(32'h3b4c1c37),
	.w8(32'hbac6ed59),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd0437),
	.w1(32'h3a9faa82),
	.w2(32'h3b52293f),
	.w3(32'hbad5bbef),
	.w4(32'hbb8296d4),
	.w5(32'hbb725b47),
	.w6(32'hbab38c31),
	.w7(32'hbac77f26),
	.w8(32'hbad2a5ed),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad765a5),
	.w1(32'h3bdc4b98),
	.w2(32'h3bb09339),
	.w3(32'h3a0493c2),
	.w4(32'h3a1a94b5),
	.w5(32'hbba8322a),
	.w6(32'h3b6cead4),
	.w7(32'h3bef654f),
	.w8(32'h3c894423),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5dc7ae),
	.w1(32'h3bfd4f83),
	.w2(32'h3bddc607),
	.w3(32'hbc12b16c),
	.w4(32'hbbbca7de),
	.w5(32'hbb2b4505),
	.w6(32'h3c1a03d9),
	.w7(32'h3cb49bc4),
	.w8(32'hbb6764d9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d9ac),
	.w1(32'h3c2497b4),
	.w2(32'h3c3ab857),
	.w3(32'h398ad760),
	.w4(32'h3b8f43f3),
	.w5(32'hbb99e967),
	.w6(32'hbbcfd841),
	.w7(32'hbb935308),
	.w8(32'h387dfed8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07102c),
	.w1(32'h3b677e0e),
	.w2(32'h3b2ea03d),
	.w3(32'h3ae3ca56),
	.w4(32'hbb56f811),
	.w5(32'hbbfecf07),
	.w6(32'h3ac2dc76),
	.w7(32'hbb28bd1b),
	.w8(32'hba1d1b15),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c8983),
	.w1(32'h3b9ea9a4),
	.w2(32'h3b75b54e),
	.w3(32'hbb8a2b06),
	.w4(32'h3a85b119),
	.w5(32'hbb094fbd),
	.w6(32'hb9948d03),
	.w7(32'h3b1b10c1),
	.w8(32'h3b2c2e08),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c591),
	.w1(32'h3b643f41),
	.w2(32'h3b12940b),
	.w3(32'h3bd47501),
	.w4(32'h3aac5fae),
	.w5(32'hb9dc9944),
	.w6(32'h3b4df0c2),
	.w7(32'h3b9ae6da),
	.w8(32'hba9ee0cb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e1556),
	.w1(32'hba9c0db2),
	.w2(32'hbac13c75),
	.w3(32'hbab61867),
	.w4(32'hba338c32),
	.w5(32'hb9e29bdd),
	.w6(32'hbadd4feb),
	.w7(32'h37885d64),
	.w8(32'hbb5d0172),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839046),
	.w1(32'hb90256e6),
	.w2(32'hbacafded),
	.w3(32'h3a877a07),
	.w4(32'h3905fc07),
	.w5(32'hba918ba6),
	.w6(32'h35876c45),
	.w7(32'h3920fcaf),
	.w8(32'h3b29ef83),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25ae8b),
	.w1(32'h3b4e2a72),
	.w2(32'h3b082246),
	.w3(32'hbb8cc11b),
	.w4(32'hbad6fc03),
	.w5(32'hbb70a808),
	.w6(32'h3b562d43),
	.w7(32'h3b857be2),
	.w8(32'h3b3282ef),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae5ecd),
	.w1(32'h3b1836b9),
	.w2(32'h3a658c7d),
	.w3(32'hbb84ea73),
	.w4(32'hbb7c5c1d),
	.w5(32'hbb8169d6),
	.w6(32'hbaba92f0),
	.w7(32'hba1bc860),
	.w8(32'hbab131ee),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e8d62),
	.w1(32'h3b6fa664),
	.w2(32'h3ba7c8fe),
	.w3(32'hbb1b4260),
	.w4(32'hba3a0f70),
	.w5(32'hbb716346),
	.w6(32'hbaf72e3c),
	.w7(32'hba37f8e8),
	.w8(32'hba9a0093),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f04a),
	.w1(32'hbba507e8),
	.w2(32'hbb2fd9de),
	.w3(32'hbc10e02f),
	.w4(32'hbc05e024),
	.w5(32'hba6be7a2),
	.w6(32'hbb86ff0b),
	.w7(32'hbb52c779),
	.w8(32'h3c20b684),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072f6c),
	.w1(32'hbb23679d),
	.w2(32'h39a015c7),
	.w3(32'hbc0595e6),
	.w4(32'hbb860442),
	.w5(32'hbb0b87d2),
	.w6(32'h3b7fecd4),
	.w7(32'h3c1147db),
	.w8(32'h39c3ea70),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cc650),
	.w1(32'h3a25aece),
	.w2(32'hba972d5f),
	.w3(32'h3b37e418),
	.w4(32'h3a27162b),
	.w5(32'hbb672778),
	.w6(32'h3bb62640),
	.w7(32'h3ba0c03d),
	.w8(32'hbb2cf442),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9dfb2),
	.w1(32'hba2072d1),
	.w2(32'h3b487fdd),
	.w3(32'hbb5927ac),
	.w4(32'hbb8a96e1),
	.w5(32'hbb5f1844),
	.w6(32'hbbb5b812),
	.w7(32'hbb657efd),
	.w8(32'hba57619f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0241b),
	.w1(32'h3bf6861f),
	.w2(32'h3bed952c),
	.w3(32'hba28bad7),
	.w4(32'h3b69e08a),
	.w5(32'hbb3ab4de),
	.w6(32'hba8d340c),
	.w7(32'h398b6e2c),
	.w8(32'hbb68aa88),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9c878),
	.w1(32'hbb7236e6),
	.w2(32'hbb54f84d),
	.w3(32'hbaa3cffc),
	.w4(32'hbbbeb816),
	.w5(32'hbb8b735f),
	.w6(32'hbbb55c13),
	.w7(32'hbb8cf302),
	.w8(32'hb897ecfd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe0f6e),
	.w1(32'hba876f36),
	.w2(32'hba94e2f9),
	.w3(32'hbb8a3726),
	.w4(32'hbba7447e),
	.w5(32'hbb4d30f8),
	.w6(32'hbacd7bb8),
	.w7(32'hbab8e845),
	.w8(32'hbbcc49ae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdeec82),
	.w1(32'hbb84e51c),
	.w2(32'h3a3e6509),
	.w3(32'hbb98b69c),
	.w4(32'hb775becc),
	.w5(32'h3a8b3091),
	.w6(32'hbb60e901),
	.w7(32'hbb3bf20f),
	.w8(32'hbb11dc23),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934fa0),
	.w1(32'hbbd7c4cb),
	.w2(32'hbbaf2f0e),
	.w3(32'h3b8285ab),
	.w4(32'h3b1b40b0),
	.w5(32'h3b1a1416),
	.w6(32'hb97a1618),
	.w7(32'hbb8126d2),
	.w8(32'hbb9bfb74),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7419d9),
	.w1(32'hbb7ec099),
	.w2(32'hba97087c),
	.w3(32'hba832f00),
	.w4(32'h3a304e60),
	.w5(32'hbb63a101),
	.w6(32'hbb6ecc13),
	.w7(32'hbbb11ef7),
	.w8(32'h3a855f21),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc81d),
	.w1(32'h3b4a593d),
	.w2(32'h3aac7d65),
	.w3(32'hbb497f01),
	.w4(32'hbb04a0f6),
	.w5(32'hba78d1d0),
	.w6(32'hba372f0e),
	.w7(32'hb9ec9802),
	.w8(32'hba838eb5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0fbcb9),
	.w1(32'hbaebbd49),
	.w2(32'hbb3fb993),
	.w3(32'h3a9abedc),
	.w4(32'h3ba1f4ec),
	.w5(32'h3b4565b9),
	.w6(32'h3a8a5d74),
	.w7(32'h3a52a5bb),
	.w8(32'h3c1292e9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f46a6),
	.w1(32'hb91c2d1d),
	.w2(32'hba907446),
	.w3(32'h39f4afc1),
	.w4(32'h3abd83a0),
	.w5(32'hbb3d7428),
	.w6(32'h3b8dcb12),
	.w7(32'h3c558f1a),
	.w8(32'h39dccd1e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ec1a0),
	.w1(32'h3b34ae60),
	.w2(32'h3b251dc8),
	.w3(32'hb73812c4),
	.w4(32'h3ab94d26),
	.w5(32'h3aa96e9e),
	.w6(32'h3a09565b),
	.w7(32'h3aedb428),
	.w8(32'hbb5ff28b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273d4d),
	.w1(32'h3a8c8e54),
	.w2(32'h3afa516d),
	.w3(32'hbb2ca8f7),
	.w4(32'hbbb9058f),
	.w5(32'h3b086134),
	.w6(32'hb9bd1a81),
	.w7(32'hbb9a28d9),
	.w8(32'h3b953f44),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c041998),
	.w1(32'h39d72e46),
	.w2(32'hbab336ce),
	.w3(32'h3b97bb21),
	.w4(32'hbb0b12a8),
	.w5(32'hbb41a247),
	.w6(32'h3b176d23),
	.w7(32'hbae20e49),
	.w8(32'hbb91d3b4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7837),
	.w1(32'hbaeb2089),
	.w2(32'h3b8cdb39),
	.w3(32'hbb63e2d3),
	.w4(32'h3a984242),
	.w5(32'h3a84f4c8),
	.w6(32'hbb29f5d7),
	.w7(32'hbb0a8e07),
	.w8(32'hbbf5d3ef),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991216),
	.w1(32'hbbf7cf48),
	.w2(32'hbbd3d6dd),
	.w3(32'hba09a81e),
	.w4(32'hba61bade),
	.w5(32'h3bad6013),
	.w6(32'hbbb85cf7),
	.w7(32'hbad83b30),
	.w8(32'h3886b7d0),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a97e3),
	.w1(32'h3b0ecc58),
	.w2(32'h3b17d8b8),
	.w3(32'h3b08b103),
	.w4(32'h3bbfb886),
	.w5(32'h3a006ee6),
	.w6(32'hb9e988c8),
	.w7(32'hbb4a0761),
	.w8(32'hbb0fc5a8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b352839),
	.w1(32'h3b6e4b6d),
	.w2(32'h396831fa),
	.w3(32'hba5fa713),
	.w4(32'hba7e4f4f),
	.w5(32'hba1f97ef),
	.w6(32'hbab790fd),
	.w7(32'hbb379d16),
	.w8(32'hbb2ca1c7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94bdf1),
	.w1(32'hbb166a98),
	.w2(32'hbb6b6147),
	.w3(32'h3a3cf0f1),
	.w4(32'h3a013312),
	.w5(32'hbb2decc6),
	.w6(32'h3b0a91d5),
	.w7(32'h3c0d1707),
	.w8(32'hba9fc70a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af62f5f),
	.w1(32'hba81242a),
	.w2(32'hbacb14f6),
	.w3(32'hbad20b74),
	.w4(32'hbb7059c2),
	.w5(32'h3b170b50),
	.w6(32'hbbcad119),
	.w7(32'hbb9095fc),
	.w8(32'h3b92541a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8d02),
	.w1(32'hbb9c752e),
	.w2(32'hbba474e8),
	.w3(32'h3b0dfc4b),
	.w4(32'hbb7ce6cd),
	.w5(32'hbb682e74),
	.w6(32'h3b5ed6ba),
	.w7(32'h3b22f88f),
	.w8(32'hbb5dbb5c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cec99),
	.w1(32'hba6816fc),
	.w2(32'h3a893ab3),
	.w3(32'hb907f440),
	.w4(32'h3ba9f411),
	.w5(32'hbb23d924),
	.w6(32'hbb3fb43c),
	.w7(32'hbaa024f0),
	.w8(32'hbb83ba27),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc863353),
	.w1(32'hbc022beb),
	.w2(32'hbb1aced8),
	.w3(32'hbc83c878),
	.w4(32'hbb1eec0e),
	.w5(32'hbac7398f),
	.w6(32'hbc201b3d),
	.w7(32'hbb24b465),
	.w8(32'hbb637154),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4c086),
	.w1(32'hbac6c14d),
	.w2(32'hbadddcbc),
	.w3(32'hba878a81),
	.w4(32'h3a9c89c8),
	.w5(32'hbaedda8b),
	.w6(32'hba843c12),
	.w7(32'h3af64d09),
	.w8(32'h39a586d5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f9c17),
	.w1(32'h3b0ba0e7),
	.w2(32'hba555a77),
	.w3(32'h3b696ff6),
	.w4(32'h3a58ec10),
	.w5(32'hba9800cc),
	.w6(32'h3a85fd59),
	.w7(32'hbb3c43da),
	.w8(32'hba6475a8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf64cd),
	.w1(32'hbaa80ad5),
	.w2(32'h3a9bb4d3),
	.w3(32'hbb987104),
	.w4(32'h3b49bcea),
	.w5(32'hbae2241a),
	.w6(32'h39430f24),
	.w7(32'h3b4c530c),
	.w8(32'hbb3c4927),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08088e),
	.w1(32'hbb5eff62),
	.w2(32'hbb85a320),
	.w3(32'hb9a8da8f),
	.w4(32'h3aa79a67),
	.w5(32'hbb21fb2a),
	.w6(32'hbb07f352),
	.w7(32'h3a438f55),
	.w8(32'h3954145f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45aa18),
	.w1(32'hbc6f2dae),
	.w2(32'hbb82f000),
	.w3(32'hbcb5eb1b),
	.w4(32'hbc0bd13a),
	.w5(32'h3b8732de),
	.w6(32'hbbff670f),
	.w7(32'hbb13cb6d),
	.w8(32'hbbf9cab5),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b689eac),
	.w1(32'h3a50bc54),
	.w2(32'h39c8742d),
	.w3(32'h3bc46631),
	.w4(32'h3a680677),
	.w5(32'hbb9c1102),
	.w6(32'h3ba06f6a),
	.w7(32'h3a9bafd2),
	.w8(32'hbbf649ec),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2697c2),
	.w1(32'hbb3b18f1),
	.w2(32'hba92da86),
	.w3(32'hbb6e1622),
	.w4(32'hbb71d2fc),
	.w5(32'h3a32084b),
	.w6(32'hbb8cec97),
	.w7(32'hbaff6b88),
	.w8(32'h3a2d074b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a5b98a),
	.w1(32'h3a9825b5),
	.w2(32'h39e734b5),
	.w3(32'h3af9e45c),
	.w4(32'h3a64db2c),
	.w5(32'hbaebb4df),
	.w6(32'h39839bdd),
	.w7(32'h3a13952f),
	.w8(32'hbb0a955f),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9851b8),
	.w1(32'hbb2aea67),
	.w2(32'hba2f1ae6),
	.w3(32'hbb11ed19),
	.w4(32'hb940f8e6),
	.w5(32'h3a37e4ff),
	.w6(32'hbb40ef5c),
	.w7(32'hbb308750),
	.w8(32'h39eee954),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7628cb),
	.w1(32'h3a341767),
	.w2(32'hba22ceb1),
	.w3(32'h3b1237d9),
	.w4(32'h390a0e5b),
	.w5(32'hbb76f737),
	.w6(32'h3a8c6ae1),
	.w7(32'hb9ab5aa4),
	.w8(32'hbb3db236),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd0c16),
	.w1(32'hba8ab640),
	.w2(32'hbb75c93c),
	.w3(32'h3a1bdd6e),
	.w4(32'h391fabac),
	.w5(32'hbb19de4d),
	.w6(32'h3a147bb2),
	.w7(32'h3a96fc82),
	.w8(32'hbb050776),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab59d8f),
	.w1(32'hba72523f),
	.w2(32'hbb0c36ef),
	.w3(32'hba4f9fee),
	.w4(32'hb9081265),
	.w5(32'h3ab215c0),
	.w6(32'hb93e012d),
	.w7(32'hb9db8cc7),
	.w8(32'h39f05af5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a579991),
	.w1(32'h3b01cf9e),
	.w2(32'h3b310aba),
	.w3(32'h3a12c688),
	.w4(32'h3aa36d1d),
	.w5(32'hb9ddce2a),
	.w6(32'h3a9c6e1b),
	.w7(32'h3b6573b5),
	.w8(32'h3b28c00f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb280784),
	.w1(32'h370640e0),
	.w2(32'h3ae9f4cd),
	.w3(32'hbb951449),
	.w4(32'hbb4f94c0),
	.w5(32'h3b301a57),
	.w6(32'hbaf47def),
	.w7(32'hbae51a90),
	.w8(32'h3a29504d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca72a8),
	.w1(32'hba1a5493),
	.w2(32'hbaca983b),
	.w3(32'h3b040bdd),
	.w4(32'h3ae4709b),
	.w5(32'hbaca4b7c),
	.w6(32'h3b209a79),
	.w7(32'h3942b1f6),
	.w8(32'hbb289107),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bf016),
	.w1(32'hbaadc477),
	.w2(32'hbb29cc5b),
	.w3(32'hba9501fb),
	.w4(32'hba8efccc),
	.w5(32'h3abfd311),
	.w6(32'hb92b81d5),
	.w7(32'hbb1c636a),
	.w8(32'h3a738501),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91b863),
	.w1(32'h3ab73367),
	.w2(32'h3ad8f584),
	.w3(32'h3a365bb1),
	.w4(32'h39aa9be3),
	.w5(32'hb9b0910e),
	.w6(32'hb9a246a7),
	.w7(32'h3a254c61),
	.w8(32'h392f4600),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49bd61),
	.w1(32'hba2e7f2f),
	.w2(32'hb9fbfbdb),
	.w3(32'h38ff61c9),
	.w4(32'hba4c1233),
	.w5(32'hba31eb48),
	.w6(32'h39cc7c61),
	.w7(32'hbae45310),
	.w8(32'hb8b6570e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb44db),
	.w1(32'hbab20bb5),
	.w2(32'h39fe377f),
	.w3(32'hbb24774e),
	.w4(32'hba19da6b),
	.w5(32'hbb6a6251),
	.w6(32'hbb19f1e4),
	.w7(32'hb9f7b827),
	.w8(32'hbb5af881),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae44811),
	.w1(32'hbb82b228),
	.w2(32'hbb9375a7),
	.w3(32'hb977c45e),
	.w4(32'hbb496926),
	.w5(32'h3a4d3203),
	.w6(32'hbad898f1),
	.w7(32'hbba3e63c),
	.w8(32'hba39d95c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2468b7),
	.w1(32'hbb22c5f2),
	.w2(32'hbb595faf),
	.w3(32'hbad87f5c),
	.w4(32'hbaf7b31c),
	.w5(32'hba8a7928),
	.w6(32'hbaa40b89),
	.w7(32'hbafd0c6f),
	.w8(32'hbab4ee87),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b626b),
	.w1(32'hbadcd40e),
	.w2(32'hba74adf3),
	.w3(32'hbb5dba92),
	.w4(32'hb9f457b7),
	.w5(32'h3a5a3d55),
	.w6(32'hbaa1a057),
	.w7(32'hb978924c),
	.w8(32'h3a90211f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacc390),
	.w1(32'h3b974b2f),
	.w2(32'h3a971503),
	.w3(32'h3b8848c1),
	.w4(32'hba6317bc),
	.w5(32'hb9e95a5e),
	.w6(32'h3b309505),
	.w7(32'h38eafedf),
	.w8(32'hb927ea5a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e4b05),
	.w1(32'h3a436dd0),
	.w2(32'hb9a0f64d),
	.w3(32'hb9fda768),
	.w4(32'hb9ec9683),
	.w5(32'h38394dc5),
	.w6(32'h3a914a1c),
	.w7(32'h39d5c528),
	.w8(32'h3a30bf85),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fdb562),
	.w1(32'h3a45e5b7),
	.w2(32'h39638abf),
	.w3(32'hba444641),
	.w4(32'hb9f007f0),
	.w5(32'h36a6383f),
	.w6(32'h3a82a73a),
	.w7(32'h3a400fb1),
	.w8(32'h3a65a2e3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b1608),
	.w1(32'h399efc67),
	.w2(32'h38b01417),
	.w3(32'h39bb6f75),
	.w4(32'hba216d20),
	.w5(32'h3a8d1492),
	.w6(32'h3a3fb250),
	.w7(32'h3946da4d),
	.w8(32'h39e3fb8c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb68d),
	.w1(32'h3a14c04c),
	.w2(32'h3a8c9d02),
	.w3(32'h3a8e7a1a),
	.w4(32'h3a4a1d7f),
	.w5(32'h39dd202b),
	.w6(32'h3a2bdda6),
	.w7(32'hb7e127d8),
	.w8(32'h397691d7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6708a),
	.w1(32'hbb0db24f),
	.w2(32'hbbce8646),
	.w3(32'hb9b6ae0a),
	.w4(32'h39cc4b6f),
	.w5(32'hbbcf043e),
	.w6(32'h3ab15710),
	.w7(32'hbabdc428),
	.w8(32'h3acc81ca),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4b96f),
	.w1(32'h3b0bcaf9),
	.w2(32'h3b8887af),
	.w3(32'hbb3a92ee),
	.w4(32'h3adc68c1),
	.w5(32'h3a4b7e75),
	.w6(32'h383b8985),
	.w7(32'h3aa74c18),
	.w8(32'h3ac116c9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85f1ce9),
	.w1(32'h39330523),
	.w2(32'h3b3d3405),
	.w3(32'hb8c62b42),
	.w4(32'h3a4cbf1b),
	.w5(32'h3a058528),
	.w6(32'h3b00e901),
	.w7(32'h3ae13bbd),
	.w8(32'hb99ae132),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c8c9d),
	.w1(32'hbaebe835),
	.w2(32'hba943bcc),
	.w3(32'hbaac5e6d),
	.w4(32'hbad239ec),
	.w5(32'hbab272d7),
	.w6(32'hba414cdc),
	.w7(32'h395ef605),
	.w8(32'hba0c3158),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986631a),
	.w1(32'hbb0a0519),
	.w2(32'hbafe519b),
	.w3(32'hba84357b),
	.w4(32'hbaaf590f),
	.w5(32'hbb24c1df),
	.w6(32'hbada9bcd),
	.w7(32'hbafe81b6),
	.w8(32'hbb8f95ef),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b716e),
	.w1(32'hbbc76313),
	.w2(32'hbbb31b78),
	.w3(32'hbbb18c77),
	.w4(32'hbb9bc632),
	.w5(32'hba795a6d),
	.w6(32'hbc0aaa44),
	.w7(32'hbbd8d0c5),
	.w8(32'hba3a2faa),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94dbb4b),
	.w1(32'hba9a5b4d),
	.w2(32'hba24b805),
	.w3(32'hbac074be),
	.w4(32'hbb461a9a),
	.w5(32'h3a8eac9e),
	.w6(32'hbb764b20),
	.w7(32'hbb6e4f6e),
	.w8(32'h3a1cf2cc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed1aa),
	.w1(32'hbadf877c),
	.w2(32'h3aa65d88),
	.w3(32'hbbd17d37),
	.w4(32'hbadad841),
	.w5(32'hbb963566),
	.w6(32'hbb504885),
	.w7(32'hba1ae2ad),
	.w8(32'hba825f43),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55585a),
	.w1(32'h39e08189),
	.w2(32'hba752012),
	.w3(32'h3aa79d22),
	.w4(32'h3a01f3ce),
	.w5(32'h3a85ac61),
	.w6(32'hba233dd6),
	.w7(32'hbb39aa9d),
	.w8(32'h3a91f64b),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6de8e),
	.w1(32'h3ababc2d),
	.w2(32'h3b32747a),
	.w3(32'hb8a08b62),
	.w4(32'h3b3524bb),
	.w5(32'hba827f99),
	.w6(32'h3a5bc5e8),
	.w7(32'h3aeba1de),
	.w8(32'hba74d13d),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2df3c),
	.w1(32'hbb044e41),
	.w2(32'hb9a41367),
	.w3(32'hbbbbbcbf),
	.w4(32'hbae88dbe),
	.w5(32'hbb3adced),
	.w6(32'hbb17c85b),
	.w7(32'hbb11d9e4),
	.w8(32'hbac673ba),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98fac60),
	.w1(32'hba3c15a8),
	.w2(32'hb9ae91cb),
	.w3(32'hba9bfc0b),
	.w4(32'hbae14df8),
	.w5(32'h3aa69eab),
	.w6(32'hbb4bf8c2),
	.w7(32'hba6d7014),
	.w8(32'hb9e3d463),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34cb03),
	.w1(32'hb88abe32),
	.w2(32'h3a34e5f4),
	.w3(32'hbb1f327c),
	.w4(32'h3802565a),
	.w5(32'h388e4ba4),
	.w6(32'h38fca8ee),
	.w7(32'h3994addd),
	.w8(32'hb9b86e1d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04c6d2),
	.w1(32'h3a537e36),
	.w2(32'h38d8849b),
	.w3(32'hb997bc88),
	.w4(32'hba31a3ea),
	.w5(32'hbaab0db9),
	.w6(32'h3b0f109d),
	.w7(32'h3a414430),
	.w8(32'hbae930c3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcf4f0),
	.w1(32'hbaf4eadf),
	.w2(32'h3b1231f1),
	.w3(32'h39eac610),
	.w4(32'hba9f2754),
	.w5(32'hba8d55da),
	.w6(32'hb9e5dded),
	.w7(32'hba973c46),
	.w8(32'h3a41905d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb275b6b),
	.w1(32'hbb5feb6d),
	.w2(32'hbb1dd2ac),
	.w3(32'hbb153336),
	.w4(32'hbb2c77db),
	.w5(32'h39da190c),
	.w6(32'hbb107bc5),
	.w7(32'hba9754f3),
	.w8(32'h3a6a5ffc),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fdd764),
	.w1(32'hbacf9fa8),
	.w2(32'h3a34f765),
	.w3(32'hba3e6503),
	.w4(32'hba9a1a25),
	.w5(32'hba154329),
	.w6(32'hb9c62952),
	.w7(32'h3a033a43),
	.w8(32'hba1b55ec),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa4398),
	.w1(32'h3a22298d),
	.w2(32'h3a3901ed),
	.w3(32'h39ceee3a),
	.w4(32'hba1f093b),
	.w5(32'hb84707d3),
	.w6(32'h3a84cd59),
	.w7(32'h3a853992),
	.w8(32'hba3730d8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042413),
	.w1(32'h38e632a9),
	.w2(32'h39faa5ed),
	.w3(32'hb96e5c80),
	.w4(32'hba604c77),
	.w5(32'h39b6966d),
	.w6(32'hb9dba169),
	.w7(32'hb952e584),
	.w8(32'h3ab7d3fc),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae28b2b),
	.w1(32'hba58de1f),
	.w2(32'hba5575cd),
	.w3(32'h36ee700a),
	.w4(32'h3ab5e33e),
	.w5(32'h39b9266c),
	.w6(32'h3acaf237),
	.w7(32'h3a93a8ee),
	.w8(32'hb989ce6a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a705094),
	.w1(32'h39b9b8e5),
	.w2(32'hba1643f6),
	.w3(32'h3a59527f),
	.w4(32'hb9095d7f),
	.w5(32'h3a2d3dd0),
	.w6(32'h3aef45f4),
	.w7(32'h39952a4c),
	.w8(32'h3aea5ff7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab19a74),
	.w1(32'hb8ee70d1),
	.w2(32'h3a4511ab),
	.w3(32'h3a4a0eee),
	.w4(32'h3a1b0f72),
	.w5(32'h3a6ed8d5),
	.w6(32'h3ab17e9c),
	.w7(32'h3ace28ef),
	.w8(32'h3aaa2c4f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b33de),
	.w1(32'h3b481e76),
	.w2(32'h3b3a88a0),
	.w3(32'h3a18ed25),
	.w4(32'h3a8358e2),
	.w5(32'hbaa6754b),
	.w6(32'h39f1100a),
	.w7(32'h3a272d46),
	.w8(32'hbab1c099),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32bcf1),
	.w1(32'hba93cab6),
	.w2(32'hba5bd1a9),
	.w3(32'hb989f1e7),
	.w4(32'hbb193bde),
	.w5(32'hba71efeb),
	.w6(32'h3aa74908),
	.w7(32'hbb23fd2c),
	.w8(32'hba52e60f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4b7b6),
	.w1(32'hbb0a807f),
	.w2(32'hba1f5e41),
	.w3(32'hbb59bc33),
	.w4(32'h37b1a4cc),
	.w5(32'hbabf153c),
	.w6(32'hbad26dc1),
	.w7(32'h38ab2d46),
	.w8(32'hb72ceac7),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87808a),
	.w1(32'h3b869ba6),
	.w2(32'hb9be8dc7),
	.w3(32'h3bcdbbb4),
	.w4(32'h3ba6c853),
	.w5(32'h3a7d7b65),
	.w6(32'h3b587b67),
	.w7(32'h3b03fe46),
	.w8(32'h3b1144f2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac5874),
	.w1(32'h396f7946),
	.w2(32'hbb08ea38),
	.w3(32'h3ae54426),
	.w4(32'hb97e8c39),
	.w5(32'hbab3c3dc),
	.w6(32'h3a943204),
	.w7(32'hbaf48b58),
	.w8(32'hbaa0eda7),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9452e00),
	.w1(32'hba8f66b9),
	.w2(32'hba0d2fb5),
	.w3(32'h3ac97759),
	.w4(32'h3b237140),
	.w5(32'h3b36b5aa),
	.w6(32'h3ae61ef2),
	.w7(32'h3b39d35a),
	.w8(32'h3b2b56db),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47ac13),
	.w1(32'h3a43f5cc),
	.w2(32'h3abb32b3),
	.w3(32'h3a3bd9c7),
	.w4(32'h3abe025b),
	.w5(32'h38811508),
	.w6(32'h3aa07a74),
	.w7(32'h3b4f73be),
	.w8(32'h3ae12e0f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04bde8),
	.w1(32'h39649026),
	.w2(32'hbab6ab4f),
	.w3(32'hb9b367b0),
	.w4(32'hba82f338),
	.w5(32'hbab1ed9b),
	.w6(32'h38883085),
	.w7(32'hbabc5eb8),
	.w8(32'hba5f33a6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bcc71),
	.w1(32'hb94fbd39),
	.w2(32'hba9cec1c),
	.w3(32'hb9903316),
	.w4(32'h39541b1b),
	.w5(32'hba22e594),
	.w6(32'hba042638),
	.w7(32'hb9df3c6e),
	.w8(32'h3919fa82),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fb5e2),
	.w1(32'hbb133501),
	.w2(32'hbaf2be79),
	.w3(32'hbb02b070),
	.w4(32'hbb41a69c),
	.w5(32'h3a77fff1),
	.w6(32'hbb1e6f3e),
	.w7(32'hbb7c28f7),
	.w8(32'h3aa15144),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab41fd),
	.w1(32'hba3b7f96),
	.w2(32'hba5ccfbb),
	.w3(32'h3a9a6c0b),
	.w4(32'hb91a0352),
	.w5(32'hba5b98da),
	.w6(32'h3b0e2649),
	.w7(32'h38027a28),
	.w8(32'hb97cd3f9),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5898e5),
	.w1(32'hbaf4fe3a),
	.w2(32'hba911ab7),
	.w3(32'hba7b223a),
	.w4(32'h3b26a558),
	.w5(32'h39d2221c),
	.w6(32'h3b9b75e3),
	.w7(32'hbb4f8120),
	.w8(32'hb9fd636a),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b85146),
	.w1(32'hb995b75c),
	.w2(32'hb95d3f0f),
	.w3(32'h3a596be8),
	.w4(32'hb9f8b2ab),
	.w5(32'hbaf56ba2),
	.w6(32'h38cb0a6f),
	.w7(32'hb9fa98bf),
	.w8(32'hba78a5d4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d43286),
	.w1(32'h3abdc02e),
	.w2(32'h3a91e4e4),
	.w3(32'h3af154c3),
	.w4(32'h3a9f49a0),
	.w5(32'hbaf5952d),
	.w6(32'hba065673),
	.w7(32'hb9c15301),
	.w8(32'hbaafd489),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9ff42),
	.w1(32'hba3d130b),
	.w2(32'hba6f7833),
	.w3(32'hb9f07add),
	.w4(32'h37f217e1),
	.w5(32'hba9b3def),
	.w6(32'hb8091aa9),
	.w7(32'hbaa009a3),
	.w8(32'h39fcf95c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54f6fc),
	.w1(32'h3a543b3c),
	.w2(32'h39eefd8d),
	.w3(32'h39b66690),
	.w4(32'hba2e01e1),
	.w5(32'hba505d72),
	.w6(32'h3ad44c49),
	.w7(32'hbb47a86b),
	.w8(32'hba247ba2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85b7cbf),
	.w1(32'hba4c31b1),
	.w2(32'hb8d70098),
	.w3(32'hbabcfc85),
	.w4(32'hba048355),
	.w5(32'h3a61f55c),
	.w6(32'hbabf0a55),
	.w7(32'h39e9b692),
	.w8(32'h3a2d2b8a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf235d),
	.w1(32'h3b359149),
	.w2(32'h3b3dba93),
	.w3(32'h3ae8e29b),
	.w4(32'h3a3a17d0),
	.w5(32'hb9d87280),
	.w6(32'h3aa36714),
	.w7(32'h3a0c812d),
	.w8(32'hbacde249),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91e60a),
	.w1(32'hbb481936),
	.w2(32'hba4443a4),
	.w3(32'hbae6a4f1),
	.w4(32'h39453236),
	.w5(32'hbb107e70),
	.w6(32'hbb961a45),
	.w7(32'h3a8a58c5),
	.w8(32'hbb12efa3),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8afe),
	.w1(32'hbb02b9b9),
	.w2(32'hba71b50e),
	.w3(32'hbbadd7a3),
	.w4(32'hb9dd6d19),
	.w5(32'hb81bb3d8),
	.w6(32'hba0fb5b2),
	.w7(32'hb92c2b0e),
	.w8(32'h3b23df20),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fc3f3),
	.w1(32'h3a7f949e),
	.w2(32'h3a58c56e),
	.w3(32'h3b0cf0c5),
	.w4(32'h3a584d56),
	.w5(32'h3a4cf205),
	.w6(32'h3aa8b4a4),
	.w7(32'h3a311ad2),
	.w8(32'h3aa46873),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8715c6),
	.w1(32'h3af6d720),
	.w2(32'h3ae403a8),
	.w3(32'h3b79086f),
	.w4(32'h3af0fc24),
	.w5(32'hbb2d5509),
	.w6(32'h3b8cc97d),
	.w7(32'h3b789331),
	.w8(32'hbb2434dc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb75e3),
	.w1(32'hbb23c03b),
	.w2(32'hba9776d5),
	.w3(32'hbb165228),
	.w4(32'hba7b4dc4),
	.w5(32'hbb1112d0),
	.w6(32'hbaca817b),
	.w7(32'hba61d5be),
	.w8(32'hbac6a314),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3deebc),
	.w1(32'hbaf514ba),
	.w2(32'hbb96dc50),
	.w3(32'hba913283),
	.w4(32'hbb54848c),
	.w5(32'hbb3e6eb6),
	.w6(32'hbae5be5a),
	.w7(32'hbb8ffa07),
	.w8(32'h39756f45),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf13c5),
	.w1(32'h3a910577),
	.w2(32'h3ab73e8b),
	.w3(32'hba05cd54),
	.w4(32'h3b201036),
	.w5(32'h3977f094),
	.w6(32'hb9c0b67d),
	.w7(32'h3ac513b7),
	.w8(32'hb9130ae4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49f403),
	.w1(32'hbadb9d6f),
	.w2(32'h38891435),
	.w3(32'hbb387121),
	.w4(32'hba574c09),
	.w5(32'h3b091b64),
	.w6(32'hbb222f28),
	.w7(32'hba26a325),
	.w8(32'h3b8a0b28),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c7f96),
	.w1(32'h3b2f1b62),
	.w2(32'h3afe7c5e),
	.w3(32'h3b2e3d77),
	.w4(32'h3acfe549),
	.w5(32'h39abc469),
	.w6(32'h3b31ef39),
	.w7(32'h3b4bddc8),
	.w8(32'h3b0e2483),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00a3a4),
	.w1(32'h3b5bc19b),
	.w2(32'h3b6c51da),
	.w3(32'h3a396934),
	.w4(32'h3aa767bc),
	.w5(32'h3b186fe6),
	.w6(32'h3abfd67e),
	.w7(32'h3a9498ea),
	.w8(32'h3b2d3309),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b608),
	.w1(32'h39b825a7),
	.w2(32'h3afcedb4),
	.w3(32'h39902595),
	.w4(32'h3a78192e),
	.w5(32'hbadf0fb9),
	.w6(32'hba75071f),
	.w7(32'h398424e1),
	.w8(32'hbb915072),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5eb77),
	.w1(32'hbb1d7751),
	.w2(32'hbadcf9a9),
	.w3(32'hbb6fc059),
	.w4(32'hba945ba8),
	.w5(32'h3a20fa6b),
	.w6(32'hbb5d907d),
	.w7(32'hba64baad),
	.w8(32'hb9935c9f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b9ea81),
	.w1(32'hba6c0593),
	.w2(32'hbabfc2be),
	.w3(32'hb883b5f7),
	.w4(32'h3aa0f1e7),
	.w5(32'hba2cae44),
	.w6(32'h391d769a),
	.w7(32'hba20d16d),
	.w8(32'hbafe86ea),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc9d3c),
	.w1(32'hb9501c42),
	.w2(32'hb8a10ad4),
	.w3(32'hbafabbf9),
	.w4(32'hbb1385ec),
	.w5(32'hb9ade9a8),
	.w6(32'hbb2de5a9),
	.w7(32'hbb5de737),
	.w8(32'hbafe6b8b),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66a65c),
	.w1(32'hbbc127d5),
	.w2(32'hba5da696),
	.w3(32'hbb9c8b3f),
	.w4(32'hbb00067e),
	.w5(32'h3a4a5694),
	.w6(32'hbb965e95),
	.w7(32'hbaad2673),
	.w8(32'h3a40bac5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398c16bb),
	.w1(32'hb9c45314),
	.w2(32'hbab933a0),
	.w3(32'hb91790fa),
	.w4(32'hba860c35),
	.w5(32'h3706d17b),
	.w6(32'h39aee201),
	.w7(32'hba41e119),
	.w8(32'h3785f19c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a581fe8),
	.w1(32'h3a15521a),
	.w2(32'h38c05b91),
	.w3(32'h3b25d4ed),
	.w4(32'h3ab7587e),
	.w5(32'h39b55c4a),
	.w6(32'h3a208b65),
	.w7(32'hb9d3c8a4),
	.w8(32'hb810d615),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39be913d),
	.w1(32'hbad0cfc1),
	.w2(32'h3af1bb45),
	.w3(32'h3b4adb54),
	.w4(32'h3b47b10a),
	.w5(32'hbafff294),
	.w6(32'h3af9cc2f),
	.w7(32'h3ab3050b),
	.w8(32'hbae23703),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1a097),
	.w1(32'hbb950c48),
	.w2(32'h391fc40a),
	.w3(32'hbc1974de),
	.w4(32'hba6acecd),
	.w5(32'h3b5cb9fc),
	.w6(32'hbbc2bd3c),
	.w7(32'h3950ec92),
	.w8(32'hbb043328),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5b468),
	.w1(32'h37d37681),
	.w2(32'h3ac9f399),
	.w3(32'hb9169196),
	.w4(32'h3aa97205),
	.w5(32'h3a17dd31),
	.w6(32'hba093ed6),
	.w7(32'h3a3f18bf),
	.w8(32'h3a0bf58a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37068a9c),
	.w1(32'h3abfeb55),
	.w2(32'h3a41ab84),
	.w3(32'hb9c22d5e),
	.w4(32'h3b1d1d2b),
	.w5(32'hba9f8615),
	.w6(32'hba8686df),
	.w7(32'h3abdbec8),
	.w8(32'h3aa8d7be),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be43727),
	.w1(32'h3b9bb39a),
	.w2(32'hba63537d),
	.w3(32'h3ba6790c),
	.w4(32'h3b8f2250),
	.w5(32'h395a4298),
	.w6(32'h3aac7bf6),
	.w7(32'h3af2f618),
	.w8(32'h3ac2c604),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ffa40b),
	.w1(32'hba95c8f9),
	.w2(32'hba9b0817),
	.w3(32'hbaab539d),
	.w4(32'hb8f4d934),
	.w5(32'h39b6b510),
	.w6(32'h397b9731),
	.w7(32'hba96513d),
	.w8(32'hbaa65186),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432713),
	.w1(32'hba0668ba),
	.w2(32'hba8fe01c),
	.w3(32'hb9fc6d95),
	.w4(32'hba7da6cf),
	.w5(32'hbaeff06b),
	.w6(32'hbacaa5b9),
	.w7(32'hbb1ec244),
	.w8(32'hbac99447),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5430df),
	.w1(32'hbb2a1f50),
	.w2(32'hba94012e),
	.w3(32'hbadd0140),
	.w4(32'hba4797e9),
	.w5(32'h3a5d3c46),
	.w6(32'hba862398),
	.w7(32'hba9d284d),
	.w8(32'h3a3e7c40),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79bc71e),
	.w1(32'hb9add2ab),
	.w2(32'h3911e2de),
	.w3(32'h3a80acc9),
	.w4(32'h3a2d2742),
	.w5(32'hba003cb9),
	.w6(32'h3a330ec6),
	.w7(32'hb8d45f46),
	.w8(32'hbb0976f4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a1d3d),
	.w1(32'h39938991),
	.w2(32'hbab1bc5d),
	.w3(32'hbb12636c),
	.w4(32'hbadebfa7),
	.w5(32'hbb90b0b5),
	.w6(32'hba8d58ae),
	.w7(32'hbb5b46d9),
	.w8(32'hbb412d35),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf36ef),
	.w1(32'hbafc4b5c),
	.w2(32'hbb22c080),
	.w3(32'hba1e7cf8),
	.w4(32'h39aac06e),
	.w5(32'hbb72205c),
	.w6(32'hb9ecd728),
	.w7(32'hba508e4a),
	.w8(32'hba8d03f8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f111e),
	.w1(32'hbb06eab8),
	.w2(32'hbaf1e4e1),
	.w3(32'hba2e9e3d),
	.w4(32'hbb787f94),
	.w5(32'hb6942c19),
	.w6(32'hbaeef815),
	.w7(32'hbb478a2d),
	.w8(32'hb860ad58),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e82412),
	.w1(32'hbaac51b1),
	.w2(32'hbb63bced),
	.w3(32'h3ac269d1),
	.w4(32'hba2c35e4),
	.w5(32'hbb209df4),
	.w6(32'h3aaff4d2),
	.w7(32'hbb2e5f57),
	.w8(32'hbb8790f4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b133b),
	.w1(32'h39aa3fe9),
	.w2(32'h3afbbd7c),
	.w3(32'hbacfbdbe),
	.w4(32'h3b245849),
	.w5(32'hbb2575d4),
	.w6(32'h3994c77a),
	.w7(32'h3a930c97),
	.w8(32'hba0fb61b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eac574),
	.w1(32'hbb0a8282),
	.w2(32'hbaa8eea2),
	.w3(32'h3a6f72cb),
	.w4(32'h3903a924),
	.w5(32'hba97ee33),
	.w6(32'h3b42d017),
	.w7(32'h39e43a81),
	.w8(32'hba6621a1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b81236),
	.w1(32'hb9efd019),
	.w2(32'h3a9237d5),
	.w3(32'h3a5c1a0d),
	.w4(32'h38bd3da4),
	.w5(32'h3ac0ebf3),
	.w6(32'h39f35419),
	.w7(32'hb96486eb),
	.w8(32'h39c2d3d9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d53db),
	.w1(32'hba93f3c8),
	.w2(32'h3b63cd62),
	.w3(32'hbb2d627e),
	.w4(32'hba81f6da),
	.w5(32'h3a55cc02),
	.w6(32'hb90e69d9),
	.w7(32'hbabbcba8),
	.w8(32'hb8cd0d14),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb916f52d),
	.w1(32'hb8e2666c),
	.w2(32'h3a7ed1ad),
	.w3(32'h39f319ba),
	.w4(32'h3a1d3799),
	.w5(32'hba633bf3),
	.w6(32'hb7c7aca5),
	.w7(32'h39bcb730),
	.w8(32'hba5fc59d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3cc7e8),
	.w1(32'h3a084e3c),
	.w2(32'h3a92030f),
	.w3(32'hbace8542),
	.w4(32'h39d8d4fb),
	.w5(32'hb9fbc0ac),
	.w6(32'h3adb8ef3),
	.w7(32'h3af5358a),
	.w8(32'h393cd4a9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac33aec),
	.w1(32'h3b01eb66),
	.w2(32'hba0b8e5c),
	.w3(32'h3b3d49f6),
	.w4(32'h3a97d429),
	.w5(32'hbad1c33e),
	.w6(32'h3ad9688f),
	.w7(32'h3a4009f8),
	.w8(32'hbb17e46b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba47029e),
	.w1(32'hb99d0a36),
	.w2(32'h3a175031),
	.w3(32'hba223fec),
	.w4(32'hba734b40),
	.w5(32'hbb1000d1),
	.w6(32'h3a4a9b63),
	.w7(32'hb983cc95),
	.w8(32'hbb3e20c3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd3b3a),
	.w1(32'hbabd78fc),
	.w2(32'hbabad6e1),
	.w3(32'hbb5c0d6d),
	.w4(32'hbab76478),
	.w5(32'hbaf8e089),
	.w6(32'hbb21623e),
	.w7(32'hbb28481f),
	.w8(32'hbb1255e6),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50d002),
	.w1(32'hb9286b6f),
	.w2(32'hbac4f424),
	.w3(32'h3aeec725),
	.w4(32'h3a92fd3e),
	.w5(32'hb9c72036),
	.w6(32'hba342538),
	.w7(32'hb9fd957d),
	.w8(32'h38c5b61e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c5874),
	.w1(32'h3ab39980),
	.w2(32'h3b27ec7a),
	.w3(32'hb9d952d3),
	.w4(32'h3a0d9550),
	.w5(32'hb7d5b4a4),
	.w6(32'hb8891e7c),
	.w7(32'hba31b6b3),
	.w8(32'h3acbbca8),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3acae8),
	.w1(32'h3b5509ff),
	.w2(32'h39a6699c),
	.w3(32'h3b53d581),
	.w4(32'h3a895728),
	.w5(32'hba30999a),
	.w6(32'h3b6dcec0),
	.w7(32'h39e3a5ae),
	.w8(32'h3a35869c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba512982),
	.w1(32'hb945337e),
	.w2(32'h3a3be78d),
	.w3(32'h3a37dfb1),
	.w4(32'h3aa205c4),
	.w5(32'hb995c787),
	.w6(32'h3a465992),
	.w7(32'h3a5686fd),
	.w8(32'hba256f28),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65b380),
	.w1(32'hbaf0559f),
	.w2(32'hbb20b906),
	.w3(32'hb9a892bd),
	.w4(32'hbab5fa3c),
	.w5(32'hbab7508f),
	.w6(32'hb745895f),
	.w7(32'hbaced433),
	.w8(32'hb943bd03),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d3520),
	.w1(32'hbb203e5d),
	.w2(32'hbba8362b),
	.w3(32'h3ae4875a),
	.w4(32'hbb07f2ce),
	.w5(32'hbab19e65),
	.w6(32'hbaaede4e),
	.w7(32'hba462fad),
	.w8(32'h3a20c532),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb392367),
	.w1(32'hbb132ede),
	.w2(32'hba33d291),
	.w3(32'hbafd7abe),
	.w4(32'hbadfef70),
	.w5(32'hba735cdf),
	.w6(32'h393bc440),
	.w7(32'hb9abb4a3),
	.w8(32'h3adce406),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35217e),
	.w1(32'h3b4b2725),
	.w2(32'h3a0cdb93),
	.w3(32'h3b844740),
	.w4(32'h3a89b459),
	.w5(32'h3a8c99bb),
	.w6(32'h3b1be6f3),
	.w7(32'hb9b79ed8),
	.w8(32'hb9ce54c1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1345d),
	.w1(32'h3a245eb9),
	.w2(32'h3bca4b65),
	.w3(32'hb962e436),
	.w4(32'h3b8eeb36),
	.w5(32'hbad488ca),
	.w6(32'hbb5cefa7),
	.w7(32'h3a7a876a),
	.w8(32'h382fa91e),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16b2c6),
	.w1(32'h3a442c35),
	.w2(32'hb939e8ab),
	.w3(32'hbab04970),
	.w4(32'hbb3159e3),
	.w5(32'h3a75b57f),
	.w6(32'hba65d712),
	.w7(32'hbaae39d9),
	.w8(32'h3989bae5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c69cd),
	.w1(32'h389dce14),
	.w2(32'h3a8da891),
	.w3(32'hba413ac0),
	.w4(32'hb9de4dff),
	.w5(32'hbadf2fae),
	.w6(32'hb9008063),
	.w7(32'h39c65b01),
	.w8(32'hba55e8fd),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab48fb1),
	.w1(32'hba95039b),
	.w2(32'hbb9801c3),
	.w3(32'hb861e5da),
	.w4(32'hbaa4e979),
	.w5(32'hbb7cde7e),
	.w6(32'h3ac0e0ec),
	.w7(32'hbb9b52b0),
	.w8(32'hbb7bc098),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d7405),
	.w1(32'hbad7b287),
	.w2(32'h39e52f62),
	.w3(32'hbb864b4f),
	.w4(32'hbaa0c937),
	.w5(32'hbac07549),
	.w6(32'hbb2c6e30),
	.w7(32'hb9620dcc),
	.w8(32'h38bd75ee),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3400c),
	.w1(32'hbb12e41c),
	.w2(32'hbae15139),
	.w3(32'hbbb86e63),
	.w4(32'hba6166ff),
	.w5(32'h3a5c8639),
	.w6(32'hba9f82c4),
	.w7(32'hba3cac76),
	.w8(32'h387735ec),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6b4ac),
	.w1(32'hb994a964),
	.w2(32'h39f459ce),
	.w3(32'h394a1cfd),
	.w4(32'hb8e8f660),
	.w5(32'h3aaa7663),
	.w6(32'hb9940554),
	.w7(32'hbaa2e3dc),
	.w8(32'h3a9d4892),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad632d7),
	.w1(32'hba7f3055),
	.w2(32'hbb293b90),
	.w3(32'h3b1a3d2d),
	.w4(32'h3a27273e),
	.w5(32'hbaa9fd24),
	.w6(32'hb8fa1cbd),
	.w7(32'hba01d156),
	.w8(32'hba3559cf),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d17e52),
	.w1(32'hbab9e404),
	.w2(32'hba723432),
	.w3(32'hba8bea11),
	.w4(32'hba80cc39),
	.w5(32'h3aa4146f),
	.w6(32'hba4e4be2),
	.w7(32'hba8f399a),
	.w8(32'h394a4b8d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b4207),
	.w1(32'hb9115be0),
	.w2(32'hba8c62e5),
	.w3(32'hba8bd6e0),
	.w4(32'hb9c9d7cc),
	.w5(32'h3a202f67),
	.w6(32'h3911a0ca),
	.w7(32'h3b0ddc40),
	.w8(32'hba9e0671),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f86bf),
	.w1(32'hb98d0737),
	.w2(32'h3a913aba),
	.w3(32'h38b59b65),
	.w4(32'h3b1b9cb6),
	.w5(32'hbab23ccc),
	.w6(32'hbb2b0a23),
	.w7(32'h3abc8d32),
	.w8(32'hbb20c4b0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1660bb),
	.w1(32'hbad513f8),
	.w2(32'hbb23c57e),
	.w3(32'h3906f27f),
	.w4(32'hba9d7098),
	.w5(32'hb84e267c),
	.w6(32'h3abd90a5),
	.w7(32'hbb2db150),
	.w8(32'hbacf2768),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21283),
	.w1(32'hbbd032cf),
	.w2(32'hbb025f5d),
	.w3(32'hbb42fd9e),
	.w4(32'hbb788545),
	.w5(32'hbb726503),
	.w6(32'hbc35dd6a),
	.w7(32'hbba1a574),
	.w8(32'hbc0e593d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a1096),
	.w1(32'hb9993712),
	.w2(32'h3c34f762),
	.w3(32'hbc039c55),
	.w4(32'hbafd1118),
	.w5(32'hbb577e17),
	.w6(32'hbca10399),
	.w7(32'hba6aa9ee),
	.w8(32'hbb96633b),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c4456),
	.w1(32'hba568840),
	.w2(32'hba37c6fc),
	.w3(32'h39e939ac),
	.w4(32'hbbcfeea4),
	.w5(32'h3ac2c4e6),
	.w6(32'hbc7ad9ec),
	.w7(32'hbc1c9570),
	.w8(32'hbb3d89b4),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46a2cf),
	.w1(32'hbbbdd5dd),
	.w2(32'h39d75bbe),
	.w3(32'hba9192cc),
	.w4(32'hbb84ff4d),
	.w5(32'hbb09cb72),
	.w6(32'hbc0ddf29),
	.w7(32'hbc07b73e),
	.w8(32'hbb858f2f),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49631f),
	.w1(32'hbbbf5a22),
	.w2(32'h3ab985ba),
	.w3(32'hbc7c1f86),
	.w4(32'hbbcc4e3e),
	.w5(32'hbb31a0ee),
	.w6(32'hbc356b6b),
	.w7(32'h3b28544f),
	.w8(32'hbaa5d21a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c77e),
	.w1(32'hb984cb70),
	.w2(32'hbb8e03c9),
	.w3(32'h3ba554cd),
	.w4(32'hba4af125),
	.w5(32'h3b3eba40),
	.w6(32'h3a722fcc),
	.w7(32'hbc04b6ff),
	.w8(32'h3c4ed791),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d02c0),
	.w1(32'h3c4af7a9),
	.w2(32'h3cab027d),
	.w3(32'hbc50a215),
	.w4(32'h3a9e9eae),
	.w5(32'hbacc6763),
	.w6(32'hbc810ebb),
	.w7(32'h378b09f7),
	.w8(32'hbb4f626b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba97333),
	.w1(32'hbb8c1897),
	.w2(32'hbb9ec911),
	.w3(32'hbb6d5e2d),
	.w4(32'hbb6aa2d3),
	.w5(32'h3c4823cd),
	.w6(32'hb9f1d56c),
	.w7(32'hbb794e32),
	.w8(32'h3c03385e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bfbfa),
	.w1(32'hbc4f4826),
	.w2(32'h3a6dc767),
	.w3(32'h3b5b7885),
	.w4(32'h3ab501cd),
	.w5(32'h3b01c3fb),
	.w6(32'hbc7ccfe4),
	.w7(32'hbc2b4081),
	.w8(32'hbab48085),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7b334),
	.w1(32'hba95b5d1),
	.w2(32'h3b2c70cc),
	.w3(32'hbafff89d),
	.w4(32'hbb59dba9),
	.w5(32'hbb6cdb14),
	.w6(32'hbc2f18ed),
	.w7(32'hbb5a9806),
	.w8(32'hbb918342),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cbc6a),
	.w1(32'hbc0cfe90),
	.w2(32'hbac61d15),
	.w3(32'hbb9ceff1),
	.w4(32'hbc0e0887),
	.w5(32'hbb533984),
	.w6(32'hbc6947bf),
	.w7(32'hbbee25e8),
	.w8(32'hbbf917cb),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90231),
	.w1(32'hbc4161b8),
	.w2(32'hbb86be3f),
	.w3(32'hbb9d1288),
	.w4(32'hbb4b80fc),
	.w5(32'h3b8a7380),
	.w6(32'hbc569d47),
	.w7(32'hbc30563b),
	.w8(32'hba0f7718),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d1120),
	.w1(32'hba8e3af2),
	.w2(32'h3bf60b4c),
	.w3(32'hbb811d29),
	.w4(32'h39df390f),
	.w5(32'h3aca500a),
	.w6(32'hbb901172),
	.w7(32'h3b1c6873),
	.w8(32'h3b1c7f0c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dec44),
	.w1(32'h3b68f6fc),
	.w2(32'h3ba2c6af),
	.w3(32'hbba0ceab),
	.w4(32'hbb60c96e),
	.w5(32'h3ab9de0a),
	.w6(32'hbb25bad7),
	.w7(32'h3a9cadba),
	.w8(32'hb9253b93),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0cc62),
	.w1(32'hbb4f91ad),
	.w2(32'hbae43f1b),
	.w3(32'hbb2b36d0),
	.w4(32'h39112c08),
	.w5(32'h3ba9d578),
	.w6(32'hbb276ce6),
	.w7(32'hb8920c29),
	.w8(32'h3b047ad6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae4ccad),
	.w1(32'h3bfa5a86),
	.w2(32'h39ea9bf8),
	.w3(32'h3c089a54),
	.w4(32'h39175581),
	.w5(32'hbb874379),
	.w6(32'h3bf7a4f7),
	.w7(32'hba27ee4e),
	.w8(32'hbb55cc05),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d02f4),
	.w1(32'hbbc8e991),
	.w2(32'hbb8be5eb),
	.w3(32'h3a4065d9),
	.w4(32'h38bbf2a3),
	.w5(32'h3bb43bcc),
	.w6(32'hbc20be19),
	.w7(32'h39ca8910),
	.w8(32'h3b05e07a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9955c4),
	.w1(32'hba0c6a56),
	.w2(32'h3c09ad19),
	.w3(32'hbbbd7b7f),
	.w4(32'hbb119ff1),
	.w5(32'h3bdfa77f),
	.w6(32'hbbb95848),
	.w7(32'h3aa1eb66),
	.w8(32'h3c472a81),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2cde2),
	.w1(32'h3c35d50c),
	.w2(32'h3accb076),
	.w3(32'h3c36cc64),
	.w4(32'h3bc5ddc2),
	.w5(32'hbad90c31),
	.w6(32'h3ca60b62),
	.w7(32'h3bc80805),
	.w8(32'hbacb0f24),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a979ff6),
	.w1(32'hbba718ae),
	.w2(32'hbbfd5b91),
	.w3(32'hbc0ced44),
	.w4(32'h3b35b12b),
	.w5(32'hbb9d1781),
	.w6(32'hbc354bbe),
	.w7(32'hbbabb9c1),
	.w8(32'hbbb99aa2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba875159),
	.w1(32'hbabf5d3c),
	.w2(32'hba8871ec),
	.w3(32'hbbd54cf6),
	.w4(32'h3a2dba1d),
	.w5(32'h3c878bc5),
	.w6(32'hbc278ae3),
	.w7(32'hbbb2f08f),
	.w8(32'h3c5edf6c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21059d),
	.w1(32'h3c3373e8),
	.w2(32'h3bdac465),
	.w3(32'h3c83c1ce),
	.w4(32'h3bbe49d2),
	.w5(32'h3c3c0e6d),
	.w6(32'h3b64c630),
	.w7(32'hb9e08439),
	.w8(32'h3bca933a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a338112),
	.w1(32'h3a20e531),
	.w2(32'h3adf5a26),
	.w3(32'h3bbdf72a),
	.w4(32'h3a8655e3),
	.w5(32'hbaced8d4),
	.w6(32'h3b76645e),
	.w7(32'hba97aca6),
	.w8(32'hbb206d82),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d03b5),
	.w1(32'hbbf1d4b9),
	.w2(32'hbbe08658),
	.w3(32'hbb8a5ae6),
	.w4(32'hbc263881),
	.w5(32'h3ac477e6),
	.w6(32'hbbbbe794),
	.w7(32'hbbac6f03),
	.w8(32'hbb739aa5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2e82b),
	.w1(32'hb93f8ea0),
	.w2(32'h3a93e718),
	.w3(32'h390f68df),
	.w4(32'h3a773d3a),
	.w5(32'hbb9018c0),
	.w6(32'hbc0948b1),
	.w7(32'hbbb9a0ce),
	.w8(32'hbbd688aa),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403025),
	.w1(32'hbb234a9a),
	.w2(32'hbb157242),
	.w3(32'hbb610dd2),
	.w4(32'hbb8868ba),
	.w5(32'h3aae8221),
	.w6(32'hbb18a6eb),
	.w7(32'hbb01b98b),
	.w8(32'hbbe99a62),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392535da),
	.w1(32'hbc0ce6a4),
	.w2(32'hbb78e654),
	.w3(32'h3b4f0eb5),
	.w4(32'h3adaef7f),
	.w5(32'hbb1c8f55),
	.w6(32'hbc0c6068),
	.w7(32'hb9ec2858),
	.w8(32'hb968ca41),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8198f),
	.w1(32'h3b00f79d),
	.w2(32'hbbcb2644),
	.w3(32'h3a719337),
	.w4(32'h3b345ed1),
	.w5(32'h3a84e8d8),
	.w6(32'hbbb6e766),
	.w7(32'hbbb1ed20),
	.w8(32'hba467728),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cd754),
	.w1(32'hbac2ef86),
	.w2(32'h3b5734e6),
	.w3(32'hbb7a036a),
	.w4(32'h3b2278af),
	.w5(32'hba409149),
	.w6(32'hbc79b6df),
	.w7(32'hb9d219fc),
	.w8(32'hba19251c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1baf67),
	.w1(32'h3b1e9132),
	.w2(32'hbacb5d10),
	.w3(32'h3be19619),
	.w4(32'h3baef762),
	.w5(32'hbb5e7573),
	.w6(32'hba6b8903),
	.w7(32'h3b7c8544),
	.w8(32'hbbe229db),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule