module layer_10_featuremap_7(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb180d70),
	.w1(32'h3b3b80bd),
	.w2(32'h3a8d2ef3),
	.w3(32'hbb858562),
	.w4(32'hbb874629),
	.w5(32'h3aa045cf),
	.w6(32'hbaf69de2),
	.w7(32'hbb4556f4),
	.w8(32'hbabf4c3d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb1d90),
	.w1(32'h3b929774),
	.w2(32'h3b584ff9),
	.w3(32'hbba100b5),
	.w4(32'hb9976933),
	.w5(32'hb9f1b1ea),
	.w6(32'hbbfc4775),
	.w7(32'hbb1a8c65),
	.w8(32'hb9feb763),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0de63),
	.w1(32'h3b92e650),
	.w2(32'h389634ee),
	.w3(32'h3ba1431a),
	.w4(32'h3b71b9ae),
	.w5(32'h3a3de78d),
	.w6(32'hbb7d6d8b),
	.w7(32'h3a5e71cc),
	.w8(32'h3b37171d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aab62),
	.w1(32'h3b90ee08),
	.w2(32'h3b522445),
	.w3(32'h3b61436a),
	.w4(32'hb9b1084a),
	.w5(32'h3b3033e2),
	.w6(32'hbb6ef499),
	.w7(32'hb681ab57),
	.w8(32'h3bafd06e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990551),
	.w1(32'h3b368c2f),
	.w2(32'hbb89735e),
	.w3(32'h3b81206a),
	.w4(32'h3bad5db6),
	.w5(32'hbbd89367),
	.w6(32'h3c2df554),
	.w7(32'h3c246923),
	.w8(32'hbbcc94b8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc68d76),
	.w1(32'hbae671cf),
	.w2(32'hbcf84290),
	.w3(32'hbba84f94),
	.w4(32'hbb5716b3),
	.w5(32'hbc888f27),
	.w6(32'hbbc47e6f),
	.w7(32'h38341c07),
	.w8(32'h3be56260),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd42c83c),
	.w1(32'hbd3b084b),
	.w2(32'hbbbc18f4),
	.w3(32'hbcf998e6),
	.w4(32'hbd152d8d),
	.w5(32'hbbf5955b),
	.w6(32'hbaaa59a6),
	.w7(32'h3b5ab2f3),
	.w8(32'h3b63067d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77b550),
	.w1(32'hbbf6bc66),
	.w2(32'h3b209b49),
	.w3(32'hb86790d6),
	.w4(32'hbbb5b441),
	.w5(32'hbcae45ba),
	.w6(32'h3d9a4574),
	.w7(32'h3cbeb511),
	.w8(32'hbc1d7647),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92bfce),
	.w1(32'h3ba5c529),
	.w2(32'hbbc23aba),
	.w3(32'hbb5c08b6),
	.w4(32'hbb3722a7),
	.w5(32'hbbbcda40),
	.w6(32'hbbc67e00),
	.w7(32'hbb79d45a),
	.w8(32'hbb56961a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1949),
	.w1(32'hba8d04d8),
	.w2(32'hbb295dfb),
	.w3(32'hbbc7bdcf),
	.w4(32'hbbcdf3f5),
	.w5(32'hbbd1899f),
	.w6(32'h3c5d2ef5),
	.w7(32'h3b43657f),
	.w8(32'h3aba4e0e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c0745),
	.w1(32'hbc172d39),
	.w2(32'hbaeea48b),
	.w3(32'hbd12c9f9),
	.w4(32'hbcd29885),
	.w5(32'hbb0e1f32),
	.w6(32'hbcc5ce66),
	.w7(32'hbc686f62),
	.w8(32'hbb56995d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf16ae),
	.w1(32'hbbdc114a),
	.w2(32'hbc1bc325),
	.w3(32'h3a06fa52),
	.w4(32'hbbb6ad02),
	.w5(32'hbb0c1ffd),
	.w6(32'h3c068b1e),
	.w7(32'hba2837f2),
	.w8(32'hbaf35f82),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c351d5f),
	.w1(32'h3b5ae2a3),
	.w2(32'hbbd8a95c),
	.w3(32'h3cdd3f68),
	.w4(32'h3c706672),
	.w5(32'hbc886b79),
	.w6(32'h3d065a55),
	.w7(32'h3c8cd48e),
	.w8(32'hbc0de7e3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d3048),
	.w1(32'hbbadf54f),
	.w2(32'h3b71b438),
	.w3(32'hbc2dd6b8),
	.w4(32'hbc3a8a41),
	.w5(32'hbbaa2c25),
	.w6(32'hbbaab41b),
	.w7(32'hba8fbf48),
	.w8(32'hbbae7eeb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d7ba7),
	.w1(32'h3b642fb1),
	.w2(32'h3bd4ec8f),
	.w3(32'hbc290135),
	.w4(32'hbb317ceb),
	.w5(32'h38c7e166),
	.w6(32'hbc4f3a19),
	.w7(32'hbbcf59a4),
	.w8(32'h3b2232d7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46000a),
	.w1(32'hbace3ab7),
	.w2(32'hbd120dfc),
	.w3(32'hbb2abf55),
	.w4(32'hbbda9295),
	.w5(32'hbcf35f52),
	.w6(32'h3b3de7eb),
	.w7(32'hbbbf6703),
	.w8(32'hbcafd4bf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0a34b5),
	.w1(32'hbcc6a79b),
	.w2(32'h3a90d593),
	.w3(32'hbd5df284),
	.w4(32'hbd260b8c),
	.w5(32'h3b2f4fd6),
	.w6(32'hbd067ddb),
	.w7(32'hbcaa5fce),
	.w8(32'h3be19d6a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b76a8),
	.w1(32'hbc83784c),
	.w2(32'hbc5bcbfa),
	.w3(32'h3c041654),
	.w4(32'hbc675504),
	.w5(32'hbc499d05),
	.w6(32'h3d217fcc),
	.w7(32'h3bb29133),
	.w8(32'hbc8ae54d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb758b53),
	.w1(32'hbc1a4780),
	.w2(32'hbbfd40cf),
	.w3(32'hba733544),
	.w4(32'hbbcbd1bc),
	.w5(32'hbc03b2cd),
	.w6(32'h3c7c45ea),
	.w7(32'h3b3947a0),
	.w8(32'hbc051fda),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeae2a9),
	.w1(32'h3b5c5bf9),
	.w2(32'h3b0d5ffd),
	.w3(32'hbb09702a),
	.w4(32'hba85931b),
	.w5(32'h3aef162b),
	.w6(32'hbbb43735),
	.w7(32'hbb9ce2f7),
	.w8(32'hba41e66f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af23be3),
	.w1(32'h3a08367e),
	.w2(32'h3b1cd47a),
	.w3(32'h3a667c8d),
	.w4(32'h3b506880),
	.w5(32'h3adc71cb),
	.w6(32'h3aaa3e56),
	.w7(32'hbae8f596),
	.w8(32'h3a952ba4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b1a58),
	.w1(32'h3b643573),
	.w2(32'h3b7c192f),
	.w3(32'hbbadeef8),
	.w4(32'hbae5669e),
	.w5(32'h3a63b474),
	.w6(32'hbb6e42fa),
	.w7(32'h3a325bd1),
	.w8(32'h3a33c4d2),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfee2b),
	.w1(32'hbbe7e628),
	.w2(32'hbcbc0c72),
	.w3(32'h3bf1764a),
	.w4(32'hbc14999f),
	.w5(32'hbc0d3523),
	.w6(32'h3c614717),
	.w7(32'h3c830122),
	.w8(32'h3c2cf843),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9016da),
	.w1(32'h3c93f9df),
	.w2(32'hbab336d3),
	.w3(32'h3c17d7dc),
	.w4(32'h3c42d0f1),
	.w5(32'h3b40c6fd),
	.w6(32'h3adc234b),
	.w7(32'h3c148348),
	.w8(32'h3ba08b97),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabf979),
	.w1(32'h3c163743),
	.w2(32'h3c4a9439),
	.w3(32'hbc422f52),
	.w4(32'h3c65149d),
	.w5(32'h3c6d322e),
	.w6(32'hbc8ed19a),
	.w7(32'h3aece8bc),
	.w8(32'h3c84dd4b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a375f),
	.w1(32'h3b7329c3),
	.w2(32'h3b9dea1a),
	.w3(32'h39d28919),
	.w4(32'hbacb8ff4),
	.w5(32'h39d9bced),
	.w6(32'h3b4b1a9e),
	.w7(32'h3b652774),
	.w8(32'h3b824ce2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba176a33),
	.w1(32'h39dee533),
	.w2(32'hb9519a46),
	.w3(32'hba8f6e2b),
	.w4(32'h3a51eb1c),
	.w5(32'hba62ae1d),
	.w6(32'hbb1b6e4d),
	.w7(32'hbab4eeab),
	.w8(32'h3a305b87),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb281a43),
	.w1(32'h3c9272a8),
	.w2(32'h3b5c0675),
	.w3(32'hbc05aeae),
	.w4(32'h3c7a6aa0),
	.w5(32'h3c7fc8a0),
	.w6(32'hbc9d4cdf),
	.w7(32'hba3d2ff4),
	.w8(32'hbb8ca722),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f777),
	.w1(32'hbc3a1587),
	.w2(32'h3b8d7c57),
	.w3(32'hbc24af47),
	.w4(32'hbc80cb08),
	.w5(32'h3b0a19c3),
	.w6(32'hbbebabd5),
	.w7(32'hbc5dbdca),
	.w8(32'hbbddd0bf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba454c3),
	.w1(32'h3cc45128),
	.w2(32'h3c6f4e77),
	.w3(32'hbc6e3896),
	.w4(32'h3c987c63),
	.w5(32'h3c4f207b),
	.w6(32'hbca69661),
	.w7(32'h3b9d8166),
	.w8(32'h3b781008),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94f129),
	.w1(32'h3ba54305),
	.w2(32'hbabf497b),
	.w3(32'hbbc12b9c),
	.w4(32'h3b9e339f),
	.w5(32'hbc2b57e6),
	.w6(32'hbba0a072),
	.w7(32'h3bcca876),
	.w8(32'hbc5d1903),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb981d7),
	.w1(32'h3c8c9117),
	.w2(32'hbbd06f96),
	.w3(32'h3b1688bb),
	.w4(32'h3ca66b2b),
	.w5(32'hbbcfa4a9),
	.w6(32'h3b1b99e3),
	.w7(32'h3c84208b),
	.w8(32'hbb7b31b1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba650fe4),
	.w1(32'hbb9e6674),
	.w2(32'h3afe3681),
	.w3(32'hbb6d2266),
	.w4(32'h3b931941),
	.w5(32'h3c0a1866),
	.w6(32'h3c4f25bf),
	.w7(32'h3bc0d971),
	.w8(32'h3c2ea7f2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba770571),
	.w1(32'hbb1abe4e),
	.w2(32'hb901934e),
	.w3(32'hb8ad80cb),
	.w4(32'h3939d981),
	.w5(32'hbb23d5ba),
	.w6(32'hb9e0c461),
	.w7(32'hbab5b5d9),
	.w8(32'hbba49d48),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3876),
	.w1(32'h3aeb8eae),
	.w2(32'h3bdb3ee9),
	.w3(32'h3b98eec8),
	.w4(32'h3bf9a689),
	.w5(32'h3c95d004),
	.w6(32'h3bca1474),
	.w7(32'h3b6dc834),
	.w8(32'h3c80b0e0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab333b9),
	.w1(32'hbc8b0a92),
	.w2(32'hbbcbd062),
	.w3(32'h3c4790be),
	.w4(32'hbc61ea86),
	.w5(32'hbb5f5bec),
	.w6(32'h3c862a3e),
	.w7(32'hbb5f5106),
	.w8(32'h3beaa61a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7915f6),
	.w1(32'h3c28ccf6),
	.w2(32'hbd145da2),
	.w3(32'hbc34bc3b),
	.w4(32'h3bb84007),
	.w5(32'hbd27ae36),
	.w6(32'h3c4b3513),
	.w7(32'h3c45e957),
	.w8(32'hbc9f4ffe),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab92d0),
	.w1(32'h3caedb00),
	.w2(32'h3d000bf8),
	.w3(32'hbc918332),
	.w4(32'h3cbb5195),
	.w5(32'h3d02d008),
	.w6(32'hbd03c3c3),
	.w7(32'h3b85f7bb),
	.w8(32'h3c8ad325),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc707402),
	.w1(32'h3c28ef02),
	.w2(32'h3cad0d7b),
	.w3(32'hbc2240c5),
	.w4(32'h3c229dde),
	.w5(32'h3cefed76),
	.w6(32'hbca247e5),
	.w7(32'h3ac0eedb),
	.w8(32'h3cb5ba9d),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc233a48),
	.w1(32'hbbac4bdc),
	.w2(32'h3c323a48),
	.w3(32'hbc6b44ef),
	.w4(32'hbc0fcb37),
	.w5(32'h3cae304a),
	.w6(32'hbc69d6a7),
	.w7(32'hbc1ab745),
	.w8(32'h3c87158a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba431777),
	.w1(32'hbbd71c9c),
	.w2(32'h3b03d6c9),
	.w3(32'h3c0923e6),
	.w4(32'hbc005935),
	.w5(32'h3ac3dabb),
	.w6(32'h3af40557),
	.w7(32'hbb91aa91),
	.w8(32'h3b5af8eb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966931),
	.w1(32'hba25ce3b),
	.w2(32'h3b99825e),
	.w3(32'h3b68619a),
	.w4(32'hbb53f882),
	.w5(32'hbb61b258),
	.w6(32'h3b5ea0de),
	.w7(32'h3b40b8ba),
	.w8(32'hbc618afb),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2caf8),
	.w1(32'h3c044356),
	.w2(32'h3bf0dff0),
	.w3(32'h3b0ed8bb),
	.w4(32'h3c64baf3),
	.w5(32'h3c348525),
	.w6(32'h3b818c2a),
	.w7(32'h3be4671c),
	.w8(32'h3c17716c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b2f81),
	.w1(32'hbc006742),
	.w2(32'hbbc583f5),
	.w3(32'h3c267094),
	.w4(32'h3ae031fe),
	.w5(32'h3c8cd87d),
	.w6(32'h3cca0bed),
	.w7(32'h3c605012),
	.w8(32'h3b6dc497),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a97e74e),
	.w1(32'h3c0b759c),
	.w2(32'h3c5341ee),
	.w3(32'hbb5ad77b),
	.w4(32'h3c5696c5),
	.w5(32'h3c24726b),
	.w6(32'hbba39241),
	.w7(32'h3c50265f),
	.w8(32'h3b9e55d5),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa92212),
	.w1(32'h3b22cb50),
	.w2(32'hbb924b9d),
	.w3(32'hb9fd098c),
	.w4(32'h3bb75846),
	.w5(32'hbbdffd9e),
	.w6(32'h3bfb4910),
	.w7(32'h3c969f03),
	.w8(32'h3bc182c4),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dac4cc),
	.w1(32'h3c74253f),
	.w2(32'hbb903551),
	.w3(32'hbbdfd9bc),
	.w4(32'h3c44785e),
	.w5(32'h3c0913af),
	.w6(32'hbb15cae9),
	.w7(32'h3c07270b),
	.w8(32'h3c159ab7),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87ab58),
	.w1(32'hbb80d491),
	.w2(32'hbca42e2e),
	.w3(32'h3ca8fc9a),
	.w4(32'hbc0029e1),
	.w5(32'hbcd0a61f),
	.w6(32'h3d472fca),
	.w7(32'h3bd93cce),
	.w8(32'hbc898e61),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7034f),
	.w1(32'hbaf5f98a),
	.w2(32'hba89c957),
	.w3(32'hbb38afa8),
	.w4(32'h388730d0),
	.w5(32'hbc0fbe07),
	.w6(32'hbb479a84),
	.w7(32'hbac11e98),
	.w8(32'hbbef1326),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf8e52),
	.w1(32'hb8051dfb),
	.w2(32'h3c266dd4),
	.w3(32'hba8e83f8),
	.w4(32'h3a69323f),
	.w5(32'h3b11ac1c),
	.w6(32'hbbd839cd),
	.w7(32'hbb3abba3),
	.w8(32'hbb156dc7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2113a1),
	.w1(32'h3c22c1d8),
	.w2(32'hbb35f548),
	.w3(32'h3bcd7ecc),
	.w4(32'h3c19eee2),
	.w5(32'hbc6575af),
	.w6(32'h3b9ab919),
	.w7(32'h3c0326cd),
	.w8(32'hbc5678de),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dc3c0),
	.w1(32'h3bc9cec2),
	.w2(32'h3bb2e29f),
	.w3(32'hbc55c802),
	.w4(32'h3b33d123),
	.w5(32'h3c28ab47),
	.w6(32'hbc2e874b),
	.w7(32'h3c5e41ad),
	.w8(32'h3c60d08d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15d802),
	.w1(32'h3aa0b668),
	.w2(32'h3bd38302),
	.w3(32'h3c1cafaa),
	.w4(32'h3c57958a),
	.w5(32'hbafd41fb),
	.w6(32'h3c1fa6aa),
	.w7(32'h3bdfabfd),
	.w8(32'hbb6ab385),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4fdfbd),
	.w1(32'h3af84df1),
	.w2(32'hbc8c3032),
	.w3(32'h3bc768d8),
	.w4(32'hbc062399),
	.w5(32'hbcbbe26d),
	.w6(32'h3d0cbea3),
	.w7(32'h3c157155),
	.w8(32'hbc98a963),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78707c),
	.w1(32'hbb921a9c),
	.w2(32'hbb5b573d),
	.w3(32'hbbcfe221),
	.w4(32'hb8cd5b1f),
	.w5(32'h3b6050de),
	.w6(32'hbb7ed0bb),
	.w7(32'hba40465d),
	.w8(32'h3bada86c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee3564),
	.w1(32'hbb3bf36f),
	.w2(32'hbac9eb2e),
	.w3(32'hbb232a02),
	.w4(32'hbb68406d),
	.w5(32'hbb079850),
	.w6(32'h3af2ac1e),
	.w7(32'hbb4e95e8),
	.w8(32'hbad17806),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb747705),
	.w1(32'h3b212434),
	.w2(32'h3c19f27c),
	.w3(32'hbc50c5e6),
	.w4(32'hb63e4264),
	.w5(32'h3be97fec),
	.w6(32'hbb280649),
	.w7(32'hba8cc77d),
	.w8(32'h3a8056a1),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a5c20),
	.w1(32'h3abf9f78),
	.w2(32'h3b6f1c98),
	.w3(32'hbb16036c),
	.w4(32'h3aac8731),
	.w5(32'h3c0111ba),
	.w6(32'hbbd14c33),
	.w7(32'h3b1545be),
	.w8(32'h3c5a7d00),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac89000),
	.w1(32'hbc701161),
	.w2(32'h3bcdf1f1),
	.w3(32'h39c45ac9),
	.w4(32'hbc6cf38f),
	.w5(32'h3b0d6002),
	.w6(32'h3b49c426),
	.w7(32'hbc19c328),
	.w8(32'hbb961d46),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f0924),
	.w1(32'h3ae2d153),
	.w2(32'h3a1f79eb),
	.w3(32'h3779e1f7),
	.w4(32'hba374831),
	.w5(32'h3b4b5fb6),
	.w6(32'hbb8d0ed6),
	.w7(32'h39bf1356),
	.w8(32'h38f0a02e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad12f9c),
	.w1(32'hbc18a19e),
	.w2(32'hbc56a83f),
	.w3(32'hbbbe4948),
	.w4(32'hbc00e590),
	.w5(32'hbce8ae59),
	.w6(32'h3bda99be),
	.w7(32'hb78e3684),
	.w8(32'hbcb4a4ce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06f0b6),
	.w1(32'h3bde1545),
	.w2(32'hbad95be5),
	.w3(32'hbc361118),
	.w4(32'h3c4010e5),
	.w5(32'h3c99e5e2),
	.w6(32'hbbf295e8),
	.w7(32'h3c4d2d2c),
	.w8(32'h3c098e6a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b2e6e),
	.w1(32'hbbe995e9),
	.w2(32'hbbae2a4b),
	.w3(32'hba92de94),
	.w4(32'hbc1067b4),
	.w5(32'hbc5633a7),
	.w6(32'h3bc82533),
	.w7(32'hbb74feb2),
	.w8(32'hbc0204fa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab964d7),
	.w1(32'h3bab9e12),
	.w2(32'h3840c821),
	.w3(32'hbb7feddb),
	.w4(32'h3b71421a),
	.w5(32'h3c361baf),
	.w6(32'hbbf64e7c),
	.w7(32'h3a3b16c8),
	.w8(32'h3c4425f2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5512ea),
	.w1(32'hbbb8e970),
	.w2(32'hbb8d2312),
	.w3(32'hb9de2e2f),
	.w4(32'hbc001895),
	.w5(32'hbb8f5b51),
	.w6(32'h3c525da0),
	.w7(32'hbba4cf91),
	.w8(32'hbb311f1f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2431c),
	.w1(32'hb9dd48e6),
	.w2(32'hbb9d4efd),
	.w3(32'hbb22e21b),
	.w4(32'hba6a4a73),
	.w5(32'hbba9d673),
	.w6(32'hba3a951a),
	.w7(32'hb885f6b4),
	.w8(32'hbb215600),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a8c51),
	.w1(32'hbc117966),
	.w2(32'hbcffab05),
	.w3(32'hbce93729),
	.w4(32'hbcad0a9a),
	.w5(32'hbc19837a),
	.w6(32'h3cae051f),
	.w7(32'hbc81f321),
	.w8(32'hbd237d84),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a1af1),
	.w1(32'hbc86b9b6),
	.w2(32'hbbd74ab5),
	.w3(32'h3b8b957c),
	.w4(32'hbc4b9db3),
	.w5(32'h3b837272),
	.w6(32'h3cc0524a),
	.w7(32'h3cd5f008),
	.w8(32'h3ca95ed5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb990ac4),
	.w1(32'hbcc04dfc),
	.w2(32'hbc97fc24),
	.w3(32'h3b4b24de),
	.w4(32'hbc818fd6),
	.w5(32'hbc772f08),
	.w6(32'h3b3a60e5),
	.w7(32'hbb034beb),
	.w8(32'hbc438f08),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c146fa),
	.w1(32'h3caf03bb),
	.w2(32'h3c414e5b),
	.w3(32'hbc31d051),
	.w4(32'h3cacb0e1),
	.w5(32'h3c74927f),
	.w6(32'hbcc4415f),
	.w7(32'h3c47faf8),
	.w8(32'h3c832958),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b04b2),
	.w1(32'hbb2d53eb),
	.w2(32'h3b157a74),
	.w3(32'hbbaa2fc5),
	.w4(32'hbb83460d),
	.w5(32'h39c1ef26),
	.w6(32'hbb4aad6b),
	.w7(32'hbb804831),
	.w8(32'hba9bf398),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac19d3),
	.w1(32'h3bbfa323),
	.w2(32'h3bc706dc),
	.w3(32'h3b999f01),
	.w4(32'h3ba6d405),
	.w5(32'h3be64c27),
	.w6(32'h3b4fc678),
	.w7(32'h3bd4d75d),
	.w8(32'h3b47c7cd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03b592),
	.w1(32'hbb7ac506),
	.w2(32'hbc98724a),
	.w3(32'h3b36d1d8),
	.w4(32'hbab7dd8b),
	.w5(32'hbcdaab6f),
	.w6(32'hba44d739),
	.w7(32'hbb04ee45),
	.w8(32'hbc95cfb6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93a1fb),
	.w1(32'h3c22e471),
	.w2(32'hbbd137f4),
	.w3(32'hbcae6e8b),
	.w4(32'h3c6c0fc6),
	.w5(32'hbc0ff7aa),
	.w6(32'hbbd54c08),
	.w7(32'h3c981972),
	.w8(32'hbbfcaf25),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab74c7e),
	.w1(32'hbb5f6150),
	.w2(32'h3ce11121),
	.w3(32'hbb816c7f),
	.w4(32'hba641013),
	.w5(32'h3d4a6aa7),
	.w6(32'hba842454),
	.w7(32'hbae4887e),
	.w8(32'h3d331b54),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1c5a9),
	.w1(32'hbcd62492),
	.w2(32'hbc5819b1),
	.w3(32'h3cd63ccc),
	.w4(32'hbcca0aa3),
	.w5(32'hbc52dce2),
	.w6(32'h3d28ceb6),
	.w7(32'hbc49780a),
	.w8(32'hbc15a0d4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3367c9),
	.w1(32'h3b5439db),
	.w2(32'hbc5b0911),
	.w3(32'h3bbe3a1f),
	.w4(32'hbb44f7dc),
	.w5(32'hbcbed319),
	.w6(32'h3d12b921),
	.w7(32'h3c40136a),
	.w8(32'hbc675d8a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc03e0),
	.w1(32'h3cb7d999),
	.w2(32'h3c4a66a0),
	.w3(32'h3b0b8903),
	.w4(32'h3caf3f57),
	.w5(32'h3b2dfbe7),
	.w6(32'hbb72f543),
	.w7(32'h3c238ea1),
	.w8(32'hbae1c1ca),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f0177),
	.w1(32'h3c2eb7bc),
	.w2(32'hbb99e6ff),
	.w3(32'h3c82302c),
	.w4(32'h3c5e49b8),
	.w5(32'hbbc92d2c),
	.w6(32'h3c8bdb7d),
	.w7(32'h3c885b2a),
	.w8(32'hbbaf95d7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c048138),
	.w1(32'h3bb7d23e),
	.w2(32'hbc194f94),
	.w3(32'hbbb667b4),
	.w4(32'hbb7ce9ac),
	.w5(32'hbbed041a),
	.w6(32'h3c8a19d9),
	.w7(32'h3a9a2d07),
	.w8(32'hbc55e316),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dba6a),
	.w1(32'h3b4af746),
	.w2(32'h39cd7c3d),
	.w3(32'hbc08ec6e),
	.w4(32'h3b5dbfa1),
	.w5(32'h3bf351ab),
	.w6(32'hbc033023),
	.w7(32'h3b1e5c81),
	.w8(32'h3b8cbdea),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2e994),
	.w1(32'hbb729c88),
	.w2(32'hbbb9f19e),
	.w3(32'h3b1ee96d),
	.w4(32'hbb91ee0f),
	.w5(32'hbbd2a56c),
	.w6(32'h3c548c3f),
	.w7(32'h3bb3ad30),
	.w8(32'hbb95cb49),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1c827),
	.w1(32'h3a83ce22),
	.w2(32'hbbdcacca),
	.w3(32'hbb63f029),
	.w4(32'hbaa7f78c),
	.w5(32'hbbb65b9a),
	.w6(32'hbb63b711),
	.w7(32'hbbead3a6),
	.w8(32'hbb259100),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25dfd9),
	.w1(32'h3c327a92),
	.w2(32'hbb5285eb),
	.w3(32'hbae1c53e),
	.w4(32'h3c0a5347),
	.w5(32'hb93ee253),
	.w6(32'h3a098906),
	.w7(32'h3b8d8597),
	.w8(32'hbbee4f6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bf9ce),
	.w1(32'h3ba9a55f),
	.w2(32'h3b99c7af),
	.w3(32'h3c01b337),
	.w4(32'h3abe860a),
	.w5(32'hbb744477),
	.w6(32'h3b1a0d71),
	.w7(32'hba187cbb),
	.w8(32'hbbeebaf9),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e7c5),
	.w1(32'hba259f50),
	.w2(32'h3b165705),
	.w3(32'hbc806022),
	.w4(32'hbb815c1a),
	.w5(32'h3a941930),
	.w6(32'hbc6cca26),
	.w7(32'hbb5b5923),
	.w8(32'h3ac8c4c6),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf5b878),
	.w1(32'hb906e2b1),
	.w2(32'h3ba24603),
	.w3(32'hbbed9ddc),
	.w4(32'h3b1cf335),
	.w5(32'h3bb65e46),
	.w6(32'hbc4a021a),
	.w7(32'hbb575440),
	.w8(32'h3bd1d68d),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba745724),
	.w1(32'hbb4bd45f),
	.w2(32'h3a8a4690),
	.w3(32'h3b15baed),
	.w4(32'hbb1a141a),
	.w5(32'h3922d057),
	.w6(32'h39bfe44f),
	.w7(32'hbac54d43),
	.w8(32'hbbbbc051),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b5735),
	.w1(32'h3b9c5cf6),
	.w2(32'h3a4d6b69),
	.w3(32'h3b8f7b51),
	.w4(32'h3c8c266b),
	.w5(32'hbad2e470),
	.w6(32'hbb16f9b8),
	.w7(32'h3c8c1480),
	.w8(32'hbafe4322),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5a64),
	.w1(32'hbc35bc77),
	.w2(32'hbae86ef9),
	.w3(32'hbb3dd1ae),
	.w4(32'hbc8dffec),
	.w5(32'h3b40ac2d),
	.w6(32'h3cb298c0),
	.w7(32'h3ba80e10),
	.w8(32'hba83975f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7c8a1),
	.w1(32'hbbdc4696),
	.w2(32'h3ba2d19d),
	.w3(32'hbc023d15),
	.w4(32'hbb895cd6),
	.w5(32'h3c35f5c5),
	.w6(32'hbc510eae),
	.w7(32'hbc05e1e9),
	.w8(32'h3c38c1a8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb631955),
	.w1(32'hbbcda39c),
	.w2(32'hbcddbf64),
	.w3(32'hba8ed24c),
	.w4(32'hbc353f73),
	.w5(32'hbc6c6f7c),
	.w6(32'h3c187c22),
	.w7(32'hbc0c6968),
	.w8(32'hbc16bdee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6623d),
	.w1(32'h3bf45064),
	.w2(32'h3c65ff07),
	.w3(32'h3a1f14db),
	.w4(32'h3c2dd795),
	.w5(32'h3c8ada31),
	.w6(32'hba8ae8de),
	.w7(32'h3c3cde62),
	.w8(32'h3c9f8e42),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b881b03),
	.w1(32'hbbf2fc6c),
	.w2(32'hbbdb6e88),
	.w3(32'hbc02a163),
	.w4(32'hbc2abf8b),
	.w5(32'h3c04e987),
	.w6(32'h3c0ffa4e),
	.w7(32'hbb3b1e71),
	.w8(32'hbc0c3071),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa03823),
	.w1(32'hbadf5fea),
	.w2(32'hbbc55d61),
	.w3(32'h3811b0eb),
	.w4(32'hbbcab715),
	.w5(32'h3b168445),
	.w6(32'h3ad64897),
	.w7(32'hbc1c0528),
	.w8(32'hbb877cb2),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca93d7),
	.w1(32'h3c351c98),
	.w2(32'h3cab207e),
	.w3(32'hbc08112c),
	.w4(32'h3c05c5ec),
	.w5(32'h3d1b053b),
	.w6(32'hbc0e4c4e),
	.w7(32'hba5bec55),
	.w8(32'h3cd0a15c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e19c9),
	.w1(32'hbc82735b),
	.w2(32'hb851902a),
	.w3(32'h3c1038b5),
	.w4(32'hbc8fc097),
	.w5(32'h3b8b5577),
	.w6(32'h3be6962e),
	.w7(32'hbbcf49b0),
	.w8(32'h3c333d8b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baade34),
	.w1(32'h3b8eb598),
	.w2(32'hbcae4123),
	.w3(32'h3bfa2fcc),
	.w4(32'h3bd93db2),
	.w5(32'hbcafc10b),
	.w6(32'h3cbcf20d),
	.w7(32'h3c923713),
	.w8(32'hbc6e4eea),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3e510),
	.w1(32'h3b8e1bb8),
	.w2(32'hbb25b1fa),
	.w3(32'hbb8edbda),
	.w4(32'h3c93c9a6),
	.w5(32'h3c8a8036),
	.w6(32'h3c26eaf2),
	.w7(32'h3c583808),
	.w8(32'h3c595ac3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ba80f),
	.w1(32'hbb8d9912),
	.w2(32'hbcf3d47e),
	.w3(32'h3cb6a778),
	.w4(32'h39c073b7),
	.w5(32'hbcde51cb),
	.w6(32'h3ca1cea4),
	.w7(32'h3c7092e1),
	.w8(32'h3c83a498),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc70a5),
	.w1(32'h3bae9894),
	.w2(32'h3bf5a2fe),
	.w3(32'hbaf1e38f),
	.w4(32'h3c1396c4),
	.w5(32'h3ca2c55c),
	.w6(32'hbc48c7c4),
	.w7(32'h3bf7995f),
	.w8(32'h3c880c7f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57edc3),
	.w1(32'h3c215f3b),
	.w2(32'h3bc2e5e8),
	.w3(32'hba103afd),
	.w4(32'h3c7ca173),
	.w5(32'h3b892f9e),
	.w6(32'hba8f5f96),
	.w7(32'h3c41283c),
	.w8(32'h3aa46d27),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e3a81),
	.w1(32'h3a7a0886),
	.w2(32'hbc33cdc2),
	.w3(32'hbc032c22),
	.w4(32'hbc000252),
	.w5(32'hbc4f2d57),
	.w6(32'h3a872acd),
	.w7(32'hbb2b68ec),
	.w8(32'hbbe02cd1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8ab30),
	.w1(32'h3c087558),
	.w2(32'hbbc6847a),
	.w3(32'h3b6816ba),
	.w4(32'h3bd11bab),
	.w5(32'hbbe63a49),
	.w6(32'hb9ed003c),
	.w7(32'h3bab3aa2),
	.w8(32'hbbc78818),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc171f29),
	.w1(32'h3cbd4174),
	.w2(32'hbc5c0f44),
	.w3(32'hbbf9cc38),
	.w4(32'h3c072481),
	.w5(32'hbd033420),
	.w6(32'h3bf45cae),
	.w7(32'h3c9c6f29),
	.w8(32'hbb1f9ed0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68dc38),
	.w1(32'h3c410567),
	.w2(32'hbb06b317),
	.w3(32'h3c037250),
	.w4(32'h3c564f23),
	.w5(32'hbbc41a1c),
	.w6(32'h3bdcafaf),
	.w7(32'h3c4615cc),
	.w8(32'h3b3027b4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ad82),
	.w1(32'h3b3dea35),
	.w2(32'hb8bd7b87),
	.w3(32'hbba184e0),
	.w4(32'h39e31362),
	.w5(32'hbbafc53a),
	.w6(32'hbb904c03),
	.w7(32'hba603b90),
	.w8(32'h3b44b9cd),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f3f6e),
	.w1(32'h3c164192),
	.w2(32'hbc40f11e),
	.w3(32'hbb8912cf),
	.w4(32'h3bbba3b4),
	.w5(32'hb9ea6d79),
	.w6(32'hbc0d1a51),
	.w7(32'h3ba524b8),
	.w8(32'hba98a0c9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf5b7),
	.w1(32'h3ba5d9eb),
	.w2(32'h3a47deac),
	.w3(32'h3ace7775),
	.w4(32'h3b078115),
	.w5(32'hbc4be947),
	.w6(32'h3c8738e0),
	.w7(32'h3c5b7188),
	.w8(32'hbc12363e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c358a),
	.w1(32'h3cc669e8),
	.w2(32'h3c7211d7),
	.w3(32'h3ae351f9),
	.w4(32'h3cd2a98b),
	.w5(32'h3bf810fd),
	.w6(32'h3aaefd58),
	.w7(32'h3ca33834),
	.w8(32'h3c1c8f7a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0460b4),
	.w1(32'h3bb3adc8),
	.w2(32'hbbb9d477),
	.w3(32'hbbbe4d23),
	.w4(32'h3c56dd19),
	.w5(32'hbc4242fb),
	.w6(32'hbc259958),
	.w7(32'h3c02ecf8),
	.w8(32'hbc5bbeb3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd05c1),
	.w1(32'h3c58f7bf),
	.w2(32'h3bc07155),
	.w3(32'hbc57115c),
	.w4(32'h3ca88375),
	.w5(32'h3bf28ef0),
	.w6(32'hbc0b3264),
	.w7(32'h3cba3d3b),
	.w8(32'h3b714f14),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4bb218),
	.w1(32'hbbf3c49e),
	.w2(32'hbc27dd0b),
	.w3(32'h3b85a0c5),
	.w4(32'hb7a7016b),
	.w5(32'hbce76e65),
	.w6(32'h3b351066),
	.w7(32'h3b987126),
	.w8(32'hbc9b417a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca34ef9),
	.w1(32'h3c5f37b7),
	.w2(32'hbca045ab),
	.w3(32'hbbaed1f1),
	.w4(32'h3c440c68),
	.w5(32'hbc080277),
	.w6(32'hb913a8f4),
	.w7(32'h3bda0528),
	.w8(32'hbbcedf0d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e029),
	.w1(32'hb94ecd98),
	.w2(32'h3b52c456),
	.w3(32'hbba89ef7),
	.w4(32'hbb74aee6),
	.w5(32'h3bc86e87),
	.w6(32'h398baf49),
	.w7(32'h3b934717),
	.w8(32'h3c0f7a85),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b354884),
	.w1(32'h3b12400e),
	.w2(32'h3895c279),
	.w3(32'h3af4db28),
	.w4(32'hba3dffa2),
	.w5(32'h3975c570),
	.w6(32'h3b992c98),
	.w7(32'h3b432b1d),
	.w8(32'hba2044c6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c2294),
	.w1(32'h3a8586fd),
	.w2(32'hb9e9e55f),
	.w3(32'hbbcc2e3a),
	.w4(32'hbaad623b),
	.w5(32'h3a4dffc3),
	.w6(32'hbc12a135),
	.w7(32'hbbdd265f),
	.w8(32'hbb9009b4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b597ebf),
	.w1(32'h3b9107a9),
	.w2(32'hbb12d9ee),
	.w3(32'h3b5fe9ea),
	.w4(32'h3b524d5f),
	.w5(32'hbbb9ae0e),
	.w6(32'h3b291701),
	.w7(32'h3b86fe2b),
	.w8(32'hbc065ccb),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09d7cb),
	.w1(32'h3c7cf561),
	.w2(32'hbbb480d4),
	.w3(32'h3ba5535f),
	.w4(32'h3cb0d7f7),
	.w5(32'hbbbb883d),
	.w6(32'hbb7858b4),
	.w7(32'h3c107f9f),
	.w8(32'hbaf285bb),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00a1b2),
	.w1(32'hba9c4486),
	.w2(32'h3beac88a),
	.w3(32'h3ad98e54),
	.w4(32'hbbbd83a6),
	.w5(32'h3c96fa8b),
	.w6(32'hba5917ca),
	.w7(32'h3b38469b),
	.w8(32'h3c8aa493),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7195),
	.w1(32'hbc26f763),
	.w2(32'hbb7c7b86),
	.w3(32'h3b890e6b),
	.w4(32'hbc2cc336),
	.w5(32'hbbdaa90e),
	.w6(32'h3c047136),
	.w7(32'hbadd30de),
	.w8(32'hbbe21dba),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad97d0b),
	.w1(32'hbaf0dde0),
	.w2(32'hbb1673d3),
	.w3(32'hbac4e8a9),
	.w4(32'hbbbafee8),
	.w5(32'h3b4028e4),
	.w6(32'h3c01283c),
	.w7(32'h3a871679),
	.w8(32'h3b8095a3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a8a99),
	.w1(32'h3bbc813c),
	.w2(32'h3c75b389),
	.w3(32'h3b9146d5),
	.w4(32'h3c2291d0),
	.w5(32'h3ca2c7d9),
	.w6(32'hbb9d4742),
	.w7(32'h3b3f17e7),
	.w8(32'h3c52f4b8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d8d6d),
	.w1(32'h3b7bb107),
	.w2(32'hbb064ded),
	.w3(32'h3bf7c0ec),
	.w4(32'h3bd04f84),
	.w5(32'hbb807a3a),
	.w6(32'hb9a35025),
	.w7(32'h3ba8f48c),
	.w8(32'hbbc4c118),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1dd11),
	.w1(32'h3a985bbc),
	.w2(32'hbc1d23db),
	.w3(32'hbaf528ed),
	.w4(32'hbacf88cd),
	.w5(32'hbc5e2488),
	.w6(32'hbb6021a8),
	.w7(32'hbb2a443e),
	.w8(32'hbc5e06f5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b3ac9),
	.w1(32'h3c2ad9cd),
	.w2(32'hbb464440),
	.w3(32'hbb4307d2),
	.w4(32'h3cb28212),
	.w5(32'hbba15fe2),
	.w6(32'h39a48e27),
	.w7(32'h3ca698cb),
	.w8(32'hbbea56f3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be90bda),
	.w1(32'h3be219e2),
	.w2(32'hbbcec812),
	.w3(32'h38e9223e),
	.w4(32'h3c20091d),
	.w5(32'hbae48c14),
	.w6(32'hbb91faca),
	.w7(32'h3ba7b17f),
	.w8(32'hbada43d5),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a5be8),
	.w1(32'hbca7b317),
	.w2(32'hbca155e0),
	.w3(32'h3c2faeba),
	.w4(32'hbc5c242f),
	.w5(32'hbc25a6b1),
	.w6(32'h3c2071ed),
	.w7(32'h3c2a2a25),
	.w8(32'h3c5d2104),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b036d8f),
	.w1(32'hbbd649fa),
	.w2(32'hbb807819),
	.w3(32'h3b25ad0c),
	.w4(32'hbc110827),
	.w5(32'hbba1e13b),
	.w6(32'h3ca0b909),
	.w7(32'h3bc07649),
	.w8(32'hbb93ccd2),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58f49),
	.w1(32'hbc477523),
	.w2(32'hbc33f137),
	.w3(32'hbc62623f),
	.w4(32'hbc1a80fd),
	.w5(32'hbbcefe40),
	.w6(32'hbb85ed4f),
	.w7(32'hbbf78b44),
	.w8(32'hbb7a646d),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dcc2b),
	.w1(32'hbb91f55d),
	.w2(32'h3a62be5e),
	.w3(32'h3bae2f34),
	.w4(32'h3ad64596),
	.w5(32'hbb66cc49),
	.w6(32'h3c5f4dcb),
	.w7(32'h3bdfd01a),
	.w8(32'h3ac1ae7b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac0e7),
	.w1(32'hbb4dcf26),
	.w2(32'h39e1444a),
	.w3(32'hbb47b5b9),
	.w4(32'hbae88f93),
	.w5(32'hbb8d6e33),
	.w6(32'h3bf5bf00),
	.w7(32'h3b912dde),
	.w8(32'hba29139f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4930d0),
	.w1(32'h3b56cb2a),
	.w2(32'h3c02584a),
	.w3(32'hbb9db75e),
	.w4(32'hbbc37cde),
	.w5(32'h3c62b90f),
	.w6(32'h3bac5585),
	.w7(32'hba1b27d5),
	.w8(32'hbb1b3821),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca50a),
	.w1(32'h3b4f8456),
	.w2(32'h3b22bcfd),
	.w3(32'hbc1e5cd1),
	.w4(32'hbaa87454),
	.w5(32'h3c111fc3),
	.w6(32'hbc2d8402),
	.w7(32'hbaf6d3d4),
	.w8(32'hbb03cc36),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28ab47),
	.w1(32'hbc5b8358),
	.w2(32'hbcb21e86),
	.w3(32'hbb1fd32b),
	.w4(32'hbc9d33b3),
	.w5(32'hbc801186),
	.w6(32'h3cacf40c),
	.w7(32'hbaaccb0c),
	.w8(32'hbc67664c),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cb12b),
	.w1(32'h3c4e1d97),
	.w2(32'h3b040e72),
	.w3(32'hbab60c63),
	.w4(32'h3c3d1ff8),
	.w5(32'hbb38d922),
	.w6(32'hbb8de501),
	.w7(32'h3bc811a2),
	.w8(32'hbbbb7a78),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ce468),
	.w1(32'h38c3119d),
	.w2(32'h3c8f1fa8),
	.w3(32'hb82428b2),
	.w4(32'hbb7a15a4),
	.w5(32'h3d509378),
	.w6(32'hbb86ab2a),
	.w7(32'hba08c050),
	.w8(32'h3d339907),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f272c),
	.w1(32'hbce98d71),
	.w2(32'hbc2c9693),
	.w3(32'h3cd8c0b3),
	.w4(32'hbd06f578),
	.w5(32'hbba128b7),
	.w6(32'h3d1070b7),
	.w7(32'hbc92335f),
	.w8(32'hb9dc9a76),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50fdd9),
	.w1(32'hbade3d51),
	.w2(32'hbc1ef201),
	.w3(32'h3b07b727),
	.w4(32'h3a84618c),
	.w5(32'hbb9225b3),
	.w6(32'h3abd2603),
	.w7(32'h3b8ae2a2),
	.w8(32'h3b368000),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac57f2),
	.w1(32'hbb3d3856),
	.w2(32'hbc1450e2),
	.w3(32'hbbc0a264),
	.w4(32'hbbd257cb),
	.w5(32'hbbcc557a),
	.w6(32'h3c95c859),
	.w7(32'h3b8cc776),
	.w8(32'hbb8abf04),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba943ac),
	.w1(32'hbb7f1e91),
	.w2(32'h3b4a2acd),
	.w3(32'hbb5e13f4),
	.w4(32'hbb22e147),
	.w5(32'h3b7ad225),
	.w6(32'hbab48268),
	.w7(32'hbad72902),
	.w8(32'h3bcd11f6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11de94),
	.w1(32'h3d005d8d),
	.w2(32'h3d063467),
	.w3(32'hba4f6334),
	.w4(32'h3cfd0b2e),
	.w5(32'h3d08698b),
	.w6(32'hbc2e44b2),
	.w7(32'h3cad8628),
	.w8(32'h3c44b9b2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e0199),
	.w1(32'h3c09c5b5),
	.w2(32'h3b5b1a2d),
	.w3(32'h3c45bf6d),
	.w4(32'h3c39fb8c),
	.w5(32'h3b95d759),
	.w6(32'h3c2e8de5),
	.w7(32'h3c198219),
	.w8(32'h3ad22bd9),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe4e0b),
	.w1(32'h3b280395),
	.w2(32'hbaa81d1a),
	.w3(32'h3b44a3da),
	.w4(32'h3b5316e3),
	.w5(32'hbaca7f70),
	.w6(32'hbad751bc),
	.w7(32'h39372ca0),
	.w8(32'hbae4c18b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3791d3),
	.w1(32'hba225e6e),
	.w2(32'hbbbb9167),
	.w3(32'hbb45b994),
	.w4(32'h39967fb0),
	.w5(32'hbc164d8a),
	.w6(32'hbb055c25),
	.w7(32'h3a186d23),
	.w8(32'hbc1929dd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace8b7),
	.w1(32'h3bbb1070),
	.w2(32'hbb8a8680),
	.w3(32'hbaca3df9),
	.w4(32'h3b4b602b),
	.w5(32'hbbde3d7b),
	.w6(32'h3ab683e8),
	.w7(32'h3c0e808f),
	.w8(32'hba4b876d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8601),
	.w1(32'h3c053489),
	.w2(32'h3b67e30a),
	.w3(32'hbbe75f98),
	.w4(32'h3bc57549),
	.w5(32'h3a2c617b),
	.w6(32'hbb6e95a0),
	.w7(32'h3b501ef4),
	.w8(32'hba44906f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5000df),
	.w1(32'h3b854492),
	.w2(32'hba87bbef),
	.w3(32'h3c1bfbff),
	.w4(32'h3c5d67fd),
	.w5(32'hbaf9c853),
	.w6(32'h3cb7f013),
	.w7(32'h3c880d27),
	.w8(32'hbb05a97e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae740c1),
	.w1(32'h3b62a5d6),
	.w2(32'hb9a8aea5),
	.w3(32'hba8fb638),
	.w4(32'h3b74e46f),
	.w5(32'hb9af5ff7),
	.w6(32'hba54522b),
	.w7(32'h3ad3adcc),
	.w8(32'h3b08eff7),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bff23),
	.w1(32'h3bcc76f1),
	.w2(32'hbc75a94b),
	.w3(32'hba927a1e),
	.w4(32'h3c11b80e),
	.w5(32'hbc1442a2),
	.w6(32'h3c5b6ef5),
	.w7(32'h3c5e044e),
	.w8(32'hbc2970d9),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06e887),
	.w1(32'h3b0d5069),
	.w2(32'h3bf3b24d),
	.w3(32'hbc278b48),
	.w4(32'h3beb2308),
	.w5(32'h3c171cf6),
	.w6(32'hbb66a289),
	.w7(32'h3b1d056f),
	.w8(32'h3bcb1426),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93bf2),
	.w1(32'hbc0a1499),
	.w2(32'hbc817857),
	.w3(32'h3b6bd2cf),
	.w4(32'hbc26c1f6),
	.w5(32'hbc97111e),
	.w6(32'h3c06e102),
	.w7(32'hbc1b872a),
	.w8(32'hbc36e5b3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba41ca4),
	.w1(32'h3ca52a35),
	.w2(32'h3bf74a3d),
	.w3(32'hbc355682),
	.w4(32'h3c9402ea),
	.w5(32'h3c81cefc),
	.w6(32'hbc6f624a),
	.w7(32'h3bb9f878),
	.w8(32'h3b0d3aab),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983f95b),
	.w1(32'hbb9c45f6),
	.w2(32'hbbe9ac26),
	.w3(32'h3b64c173),
	.w4(32'h3b00c77d),
	.w5(32'h3baf89dc),
	.w6(32'hb9546a3d),
	.w7(32'h3aa68afc),
	.w8(32'hbb2afd44),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda5fdd),
	.w1(32'h3c14c5fe),
	.w2(32'h3a4a755f),
	.w3(32'h3b81e8ff),
	.w4(32'h3c5b807c),
	.w5(32'hbb92b5f5),
	.w6(32'hba1447fe),
	.w7(32'h3be56b26),
	.w8(32'hbb2f92d7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48b8f2),
	.w1(32'h3ae99889),
	.w2(32'h3bb784ff),
	.w3(32'hbce05bd5),
	.w4(32'hbb9dd20c),
	.w5(32'h3c11830e),
	.w6(32'hbcb5dff8),
	.w7(32'hbb5c2403),
	.w8(32'h3bc75f07),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e952),
	.w1(32'hbbbd2290),
	.w2(32'hbabd1b3b),
	.w3(32'hbb3131b5),
	.w4(32'hbc2f73d9),
	.w5(32'hba27b46d),
	.w6(32'hbc2f3793),
	.w7(32'hbc5daa3d),
	.w8(32'h3ae68f71),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0209d1),
	.w1(32'h3b87e55a),
	.w2(32'h3c3a981b),
	.w3(32'hb98e9856),
	.w4(32'h3c1947a5),
	.w5(32'h3bf58272),
	.w6(32'hbc47360f),
	.w7(32'hbb652c00),
	.w8(32'h3bd724e9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6b01),
	.w1(32'h3aea3e04),
	.w2(32'hbbba8651),
	.w3(32'hbbf5b954),
	.w4(32'hbbe663c6),
	.w5(32'hbbc21fc8),
	.w6(32'hbb901e89),
	.w7(32'hbb9bea47),
	.w8(32'hbc172398),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc155de),
	.w1(32'hbb82c621),
	.w2(32'h3b451184),
	.w3(32'hbb7f58a9),
	.w4(32'hbade23b3),
	.w5(32'hba70279b),
	.w6(32'hbc1949c6),
	.w7(32'hbbf1fa5a),
	.w8(32'h3b383a62),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cbf38),
	.w1(32'h3ae43d8e),
	.w2(32'hbb7381e0),
	.w3(32'hba32ec00),
	.w4(32'hbb12cb6c),
	.w5(32'hbbb80bac),
	.w6(32'h3c00a859),
	.w7(32'h3ae86881),
	.w8(32'h3ac29f91),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5454),
	.w1(32'hba34a162),
	.w2(32'hbb4774c6),
	.w3(32'hbbb58c73),
	.w4(32'hbbb2ae8b),
	.w5(32'hbc18ff6b),
	.w6(32'hba746747),
	.w7(32'hbacc0758),
	.w8(32'hbc2fcb6c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafbe71),
	.w1(32'hb9e0e0ee),
	.w2(32'h3bfb1b43),
	.w3(32'hbc014f6f),
	.w4(32'h3978d6b9),
	.w5(32'h3c7fe031),
	.w6(32'hbc1006bf),
	.w7(32'h3bccdf02),
	.w8(32'h3c73001f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c92a8),
	.w1(32'h3babb14f),
	.w2(32'hbba54d5b),
	.w3(32'h3cae6387),
	.w4(32'h3c60bce2),
	.w5(32'hbba11a11),
	.w6(32'h3ca007a8),
	.w7(32'h3c6fcd88),
	.w8(32'h3b5a6526),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36d9c4),
	.w1(32'h39b49fd9),
	.w2(32'hb99f2966),
	.w3(32'hbb1bafdf),
	.w4(32'hbb97bbd4),
	.w5(32'h3b578541),
	.w6(32'h3bf38145),
	.w7(32'h3bbfef83),
	.w8(32'h3c305e52),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85c8ff),
	.w1(32'h3a1e62a8),
	.w2(32'hbadb140a),
	.w3(32'h3ae0de5e),
	.w4(32'h3b9e4f29),
	.w5(32'hbb8a754e),
	.w6(32'h3bc5ce2e),
	.w7(32'h3c000fee),
	.w8(32'hba83379f),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bd3b2),
	.w1(32'hba10e810),
	.w2(32'h3b68b9af),
	.w3(32'hbb6ede77),
	.w4(32'hbbb55e78),
	.w5(32'hb8c5c4fc),
	.w6(32'hbbdef408),
	.w7(32'hbac3b110),
	.w8(32'hbb9da116),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8b493),
	.w1(32'hbba6bf9b),
	.w2(32'h3a675878),
	.w3(32'hbc0536fe),
	.w4(32'hbbd44343),
	.w5(32'hbaa0e755),
	.w6(32'hbc8fb328),
	.w7(32'hbc3f361d),
	.w8(32'hba8e0f1e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b1f6b),
	.w1(32'hbc0ae8b0),
	.w2(32'hbb48774b),
	.w3(32'h3bd3dcf2),
	.w4(32'hbb9db260),
	.w5(32'hbbf66409),
	.w6(32'h3c9d6d1f),
	.w7(32'h3c91401c),
	.w8(32'h3c41cd70),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b772235),
	.w1(32'h3bab2ec4),
	.w2(32'h3b9c8240),
	.w3(32'h3af54174),
	.w4(32'h3abafce8),
	.w5(32'h38d074c1),
	.w6(32'h3b9068fb),
	.w7(32'h3ad16d76),
	.w8(32'hbadb8804),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940fb3c),
	.w1(32'h3c066102),
	.w2(32'h3bd0d85a),
	.w3(32'hbb7d58d1),
	.w4(32'h3bfe2b15),
	.w5(32'h3b0e6cdf),
	.w6(32'hbc43427e),
	.w7(32'h3a26063c),
	.w8(32'h3b4d16a6),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8fb57),
	.w1(32'hbb752f0a),
	.w2(32'h3b8cc9c5),
	.w3(32'hbcb829e0),
	.w4(32'hbc572f1e),
	.w5(32'h3c088786),
	.w6(32'hbc887440),
	.w7(32'hbc2f8a77),
	.w8(32'h3b9ed34b),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2292e2),
	.w1(32'hbb45a7b1),
	.w2(32'hbba12355),
	.w3(32'h3bd00b3e),
	.w4(32'h3b021782),
	.w5(32'h3a5b74af),
	.w6(32'h3bc5f164),
	.w7(32'h3be2b50b),
	.w8(32'h39d5828e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135e0d),
	.w1(32'hbb448d14),
	.w2(32'hbbba606f),
	.w3(32'h3b0f2881),
	.w4(32'h3b7cd82f),
	.w5(32'hbbb13789),
	.w6(32'h3c1dda63),
	.w7(32'h3bbb6118),
	.w8(32'hbb4379be),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb7dc1),
	.w1(32'hbc03a0df),
	.w2(32'hbc03a923),
	.w3(32'hbbb6fb7c),
	.w4(32'hbb2063bf),
	.w5(32'hbc58f4dc),
	.w6(32'h3c1b1308),
	.w7(32'h3b01817d),
	.w8(32'hbc28275a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc111167),
	.w1(32'hbaad5411),
	.w2(32'h39281c71),
	.w3(32'hbc48423c),
	.w4(32'h39e01396),
	.w5(32'h3c364d70),
	.w6(32'hbbaae56e),
	.w7(32'hbaefad33),
	.w8(32'h3c0dac4c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebdfcf),
	.w1(32'h3aa63a2c),
	.w2(32'hba6c926d),
	.w3(32'h3c977c2d),
	.w4(32'h3c6051d0),
	.w5(32'h3aed906d),
	.w6(32'h3cba4c23),
	.w7(32'h3c31fbf8),
	.w8(32'hbb955999),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6777c3),
	.w1(32'hbbc3b92c),
	.w2(32'h3ad70f23),
	.w3(32'hbb5760dc),
	.w4(32'hbbbda257),
	.w5(32'h3b07b333),
	.w6(32'h3bb787a2),
	.w7(32'h3a4985c6),
	.w8(32'h3b9c7a07),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ff1f),
	.w1(32'h3a9a56c7),
	.w2(32'hb86a87e7),
	.w3(32'h3b6689b5),
	.w4(32'hbb908dc1),
	.w5(32'h3ae98d24),
	.w6(32'h3bbb430e),
	.w7(32'h3b6eb053),
	.w8(32'h3b1bcfe6),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ca1e0),
	.w1(32'h3ae022da),
	.w2(32'hbb2309e8),
	.w3(32'h3ba68812),
	.w4(32'h3bc1d509),
	.w5(32'h3b11a953),
	.w6(32'h3b0013eb),
	.w7(32'hbb683046),
	.w8(32'hb913a15e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be167cd),
	.w1(32'hbbf8d15b),
	.w2(32'hbb5e193e),
	.w3(32'hbb5ad667),
	.w4(32'hbb886d60),
	.w5(32'h3b7fb961),
	.w6(32'hbb1fec43),
	.w7(32'hbbf8bb02),
	.w8(32'hbba2b3be),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981e220),
	.w1(32'h3a82d1ec),
	.w2(32'h3b9c2ee9),
	.w3(32'h3a87dc89),
	.w4(32'h3b92957e),
	.w5(32'h3becfc4a),
	.w6(32'h3b8636a3),
	.w7(32'h3b2b42fa),
	.w8(32'h3b695084),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e800dd),
	.w1(32'hbb140b48),
	.w2(32'h3a9e4b41),
	.w3(32'h3c1ac3d0),
	.w4(32'h3b71507e),
	.w5(32'h3a98bade),
	.w6(32'h388735fd),
	.w7(32'hb90ed2cb),
	.w8(32'hb9f5e5d0),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a75c3),
	.w1(32'hbb2891ef),
	.w2(32'hbb50aaea),
	.w3(32'hbb5e3cc3),
	.w4(32'h396b3958),
	.w5(32'hbb5f6413),
	.w6(32'hbb6c631a),
	.w7(32'hba880405),
	.w8(32'hbb03a1b4),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a8403),
	.w1(32'hbb9893ba),
	.w2(32'hbc3abee7),
	.w3(32'hbc79e72b),
	.w4(32'hbc3948a0),
	.w5(32'h3abbfd83),
	.w6(32'hbc278bf2),
	.w7(32'hbc4e2711),
	.w8(32'h3b266137),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4d28b),
	.w1(32'h3b97fd9d),
	.w2(32'hbc0f45d9),
	.w3(32'h3b02b78f),
	.w4(32'h3a833a18),
	.w5(32'hbc1692b9),
	.w6(32'h3c3fa39b),
	.w7(32'h3bed5350),
	.w8(32'hbb74b07c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba833ae4),
	.w1(32'hbba29530),
	.w2(32'h3b4bb62d),
	.w3(32'hbbde1c37),
	.w4(32'hbc358ef8),
	.w5(32'h3ba9f54a),
	.w6(32'hbc555678),
	.w7(32'hbc92f2cd),
	.w8(32'h3b8cf339),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc13f94),
	.w1(32'hbca80fbe),
	.w2(32'hbcb5e5a5),
	.w3(32'h3c0b567b),
	.w4(32'hbcc7571b),
	.w5(32'hbcfa0163),
	.w6(32'h3c7ffddd),
	.w7(32'hbc2b27d7),
	.w8(32'hbcec16f1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc897480),
	.w1(32'hbc04a4d5),
	.w2(32'hbb4f5867),
	.w3(32'hbc9ffb94),
	.w4(32'h3af40d68),
	.w5(32'h3c02c33a),
	.w6(32'hbca12234),
	.w7(32'hbc7a375c),
	.w8(32'hbb19a1d0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4107a9),
	.w1(32'hbafce0ff),
	.w2(32'hbb981095),
	.w3(32'hbb9403ac),
	.w4(32'hbb2e9e88),
	.w5(32'hbbed7afe),
	.w6(32'h3b5b4b41),
	.w7(32'h3a1a0627),
	.w8(32'hbbe6f790),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83fa94),
	.w1(32'hbb0ed0d2),
	.w2(32'h3b229b69),
	.w3(32'hbbc9fdda),
	.w4(32'hbbbe0dfb),
	.w5(32'hbb152a77),
	.w6(32'hbbf9b2f7),
	.w7(32'hbb448e4a),
	.w8(32'h3aeb4eb4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2058a),
	.w1(32'h3b2de6d5),
	.w2(32'hbaa2b1aa),
	.w3(32'hba8c151d),
	.w4(32'hbb886565),
	.w5(32'hbb5367ff),
	.w6(32'h3a84fc11),
	.w7(32'h392d9ce0),
	.w8(32'h3a9dc4a7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f1477),
	.w1(32'hbadf5a53),
	.w2(32'hbafc4bfb),
	.w3(32'hbb95ba24),
	.w4(32'hbb7d42ea),
	.w5(32'hba4a925c),
	.w6(32'hba4f38b7),
	.w7(32'hbaa71608),
	.w8(32'h3acc233a),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4d976),
	.w1(32'hbc2bdd04),
	.w2(32'hbcb58fcf),
	.w3(32'h399f057a),
	.w4(32'hbc19021c),
	.w5(32'hbd0e0f7c),
	.w6(32'h3bc7f2f0),
	.w7(32'h38923106),
	.w8(32'hbcc0d334),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1af68e),
	.w1(32'hbceba1dd),
	.w2(32'hbae4d2e7),
	.w3(32'hbd8af4df),
	.w4(32'hbd53c8e9),
	.w5(32'hba9ab198),
	.w6(32'hbd59f0a3),
	.w7(32'hbd10d3b8),
	.w8(32'h3c0905fa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb873a7e),
	.w1(32'h3bcc05dd),
	.w2(32'hbaccdfcb),
	.w3(32'hbba5b012),
	.w4(32'h3c0a9372),
	.w5(32'h39dcd0cd),
	.w6(32'hbafd8d04),
	.w7(32'h3baea473),
	.w8(32'hbb6ce482),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc05ed4),
	.w1(32'hbb2f5965),
	.w2(32'h3a863fd4),
	.w3(32'hba8bb69c),
	.w4(32'h3a39f148),
	.w5(32'h3b117ab0),
	.w6(32'hbb976b01),
	.w7(32'hbb11ba1c),
	.w8(32'hba5edd0e),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0099db),
	.w1(32'hbb8fd18c),
	.w2(32'hbb7ae9b5),
	.w3(32'h3b37ee29),
	.w4(32'hbb9d74f0),
	.w5(32'hbb4742b3),
	.w6(32'h3c143781),
	.w7(32'h3baed859),
	.w8(32'h3b7b6622),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953d7d3),
	.w1(32'h3bb14798),
	.w2(32'hbafc5d56),
	.w3(32'h3b3b131a),
	.w4(32'h3c185ff0),
	.w5(32'hbab925d9),
	.w6(32'h3b924d3e),
	.w7(32'h3bcaf349),
	.w8(32'h3ad32eec),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b119968),
	.w1(32'h3abc2562),
	.w2(32'h3a9d0570),
	.w3(32'h3a8c2201),
	.w4(32'hb99c342f),
	.w5(32'hbada8eb1),
	.w6(32'h3acae29d),
	.w7(32'hb9b73cdb),
	.w8(32'h3ae1105b),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dcd4f),
	.w1(32'hbba6e488),
	.w2(32'hbad5a062),
	.w3(32'hbbf16f30),
	.w4(32'hbb8ad734),
	.w5(32'h3a891c27),
	.w6(32'h3afaed2b),
	.w7(32'h3b771b67),
	.w8(32'hbad85d8e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c0303c),
	.w1(32'hba8343b3),
	.w2(32'hbc839dc9),
	.w3(32'h3aa87137),
	.w4(32'hbbab7480),
	.w5(32'hbbc7982b),
	.w6(32'hbbf9135a),
	.w7(32'hbbc5fe5b),
	.w8(32'hbc22bee3),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb383115),
	.w1(32'hbc41e26c),
	.w2(32'hbb9fce09),
	.w3(32'h3c350e5c),
	.w4(32'h3a969e67),
	.w5(32'hbb7114fa),
	.w6(32'h3c50545d),
	.w7(32'h3bb8b3d2),
	.w8(32'h3aed0150),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306d22),
	.w1(32'hbba6e832),
	.w2(32'hbb700c86),
	.w3(32'hbc546a87),
	.w4(32'hbbf0437e),
	.w5(32'hbbc02f98),
	.w6(32'hbc85dc16),
	.w7(32'hbc13a719),
	.w8(32'hbbc984fc),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f579),
	.w1(32'hbb84c2f2),
	.w2(32'h3b5e465e),
	.w3(32'hbb8c7cc0),
	.w4(32'hbb45dfc8),
	.w5(32'h3b8c3d21),
	.w6(32'hbc36a3f8),
	.w7(32'hba12a514),
	.w8(32'hbb131838),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f78001),
	.w1(32'hb9de24c4),
	.w2(32'h3ac1565d),
	.w3(32'hbb933c16),
	.w4(32'hbaaec057),
	.w5(32'hb9ee921e),
	.w6(32'hbb77cfe6),
	.w7(32'hbb4b6f26),
	.w8(32'hbb164f34),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fdca9),
	.w1(32'h3bb3e067),
	.w2(32'h3bd7059c),
	.w3(32'hbc2daecf),
	.w4(32'h3bd3ffac),
	.w5(32'h3bdb765d),
	.w6(32'hbc2d447c),
	.w7(32'hba6e8419),
	.w8(32'hbaee5593),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2ecab),
	.w1(32'h38dda0de),
	.w2(32'hbba90e14),
	.w3(32'hbc764375),
	.w4(32'hbbcb70dc),
	.w5(32'hbbde7235),
	.w6(32'hbb8880fb),
	.w7(32'hbb90331c),
	.w8(32'hbc1d0dd9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3710f),
	.w1(32'h3b36b91f),
	.w2(32'hbc87c845),
	.w3(32'h3bb45d71),
	.w4(32'h3b5ed661),
	.w5(32'hbd1aedb3),
	.w6(32'h3c2006fc),
	.w7(32'h3c043439),
	.w8(32'hbd03140f),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd344468),
	.w1(32'hbcf44040),
	.w2(32'hbbac0df4),
	.w3(32'hbda26b1c),
	.w4(32'hbd6f6c55),
	.w5(32'hbb045a20),
	.w6(32'hbd93e1b3),
	.w7(32'hbd50f864),
	.w8(32'hbb186fd1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac174a1),
	.w1(32'hba02e84c),
	.w2(32'h39b6913a),
	.w3(32'hba71aaf0),
	.w4(32'h3be12a3b),
	.w5(32'hba2efe58),
	.w6(32'h3b43722b),
	.w7(32'h3b51b960),
	.w8(32'h3aebeeee),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28aa65),
	.w1(32'hbbe153fc),
	.w2(32'hbbf94f36),
	.w3(32'h3987cbe1),
	.w4(32'h3b9e1985),
	.w5(32'hbc34270d),
	.w6(32'h3c144d28),
	.w7(32'h3cac0c71),
	.w8(32'h3a0dd5fa),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1214a6),
	.w1(32'hbc2e25e7),
	.w2(32'hbc19efaf),
	.w3(32'hba836a5c),
	.w4(32'hbbd98090),
	.w5(32'hbc1ba664),
	.w6(32'h3c1d5c30),
	.w7(32'h3c0ab36c),
	.w8(32'hbaf77e52),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc040a71),
	.w1(32'hbc10eaf5),
	.w2(32'h3a03c261),
	.w3(32'hbca72604),
	.w4(32'hbc21929e),
	.w5(32'h3b47a96d),
	.w6(32'hbc17b440),
	.w7(32'h3a984600),
	.w8(32'h3ba39fe2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebfa1e),
	.w1(32'hbbd37430),
	.w2(32'hbca9dde8),
	.w3(32'hbcb8c898),
	.w4(32'hbca099d7),
	.w5(32'hbc83cbf5),
	.w6(32'h3b99b96f),
	.w7(32'hbc799302),
	.w8(32'hbcb00953),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8d07),
	.w1(32'h3a41a3f5),
	.w2(32'h3ba41c77),
	.w3(32'hbb7c9791),
	.w4(32'hbb17082a),
	.w5(32'h3b72e1ce),
	.w6(32'hbb901c58),
	.w7(32'hba21610f),
	.w8(32'hba98dcfa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a2b9),
	.w1(32'h3ae5851a),
	.w2(32'h3bb452d3),
	.w3(32'h3b2fee58),
	.w4(32'hbaa85fc3),
	.w5(32'hba4f66aa),
	.w6(32'h3ba32e63),
	.w7(32'h3afc1b3d),
	.w8(32'h3a5c1c91),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafac22f),
	.w1(32'hbc06bf1e),
	.w2(32'hbcbaa0dd),
	.w3(32'h3c4709c6),
	.w4(32'h3ac33a87),
	.w5(32'hbc895be4),
	.w6(32'h3c7d7968),
	.w7(32'h3cc4cadf),
	.w8(32'h3c89ce95),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0fb5),
	.w1(32'hbcc31928),
	.w2(32'hbcbda14e),
	.w3(32'hbc0bfa96),
	.w4(32'hbca993bb),
	.w5(32'hbcdb573c),
	.w6(32'h3cbef1ec),
	.w7(32'h3bcdd649),
	.w8(32'hbcb906dd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca17a49),
	.w1(32'hbca799b1),
	.w2(32'hbc92351b),
	.w3(32'hbb71d71e),
	.w4(32'hbca8cdbf),
	.w5(32'hbc82b020),
	.w6(32'hbb09fcfa),
	.w7(32'hbc749806),
	.w8(32'hbacb5865),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27c02),
	.w1(32'h3ad6d488),
	.w2(32'h3c696766),
	.w3(32'hbbcd0b64),
	.w4(32'h3b878320),
	.w5(32'h3c54c6ec),
	.w6(32'hbc2531ff),
	.w7(32'h3906af13),
	.w8(32'h3c23ccaf),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb834417),
	.w1(32'h3beab395),
	.w2(32'h3b1eb056),
	.w3(32'hbcd72cee),
	.w4(32'hbb882621),
	.w5(32'h3bfdfa85),
	.w6(32'hbcf56ce1),
	.w7(32'hbc3c6536),
	.w8(32'hba7d8720),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb81518c),
	.w1(32'hbbe57fd9),
	.w2(32'h3a6a389e),
	.w3(32'hbbf62573),
	.w4(32'hbadd2253),
	.w5(32'hbc462f59),
	.w6(32'hbb13ecdf),
	.w7(32'hbb929239),
	.w8(32'hbb4f8cab),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe37d54),
	.w1(32'hbc16cf38),
	.w2(32'h3b13cd92),
	.w3(32'hbc8b175d),
	.w4(32'hbc5b1f8c),
	.w5(32'h39f3915a),
	.w6(32'hb907ada5),
	.w7(32'hb8d00f1a),
	.w8(32'h3b41e28e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195089),
	.w1(32'hbbeea765),
	.w2(32'hbb0f054b),
	.w3(32'hbbfedf96),
	.w4(32'hbc29188d),
	.w5(32'h388040c1),
	.w6(32'h3b61ab62),
	.w7(32'hbad7bd62),
	.w8(32'h3aa4c580),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22bf1),
	.w1(32'hbb20ce3c),
	.w2(32'h3a472f0e),
	.w3(32'h3a2938d9),
	.w4(32'h378694b2),
	.w5(32'h3b589acd),
	.w6(32'hbb8d9ce6),
	.w7(32'hbb94e646),
	.w8(32'h3b95a449),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54a1b1),
	.w1(32'hbacd9da6),
	.w2(32'hbb810fd3),
	.w3(32'h3b39fc63),
	.w4(32'hbb4727c3),
	.w5(32'hbc02f3a2),
	.w6(32'h3ad1d1f2),
	.w7(32'h3a439ab2),
	.w8(32'hbc080fd3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31db06),
	.w1(32'hbc20952b),
	.w2(32'hbc310e10),
	.w3(32'hbb6bb1a1),
	.w4(32'hbb21a351),
	.w5(32'hbc62def0),
	.w6(32'h39fd5574),
	.w7(32'h3be85335),
	.w8(32'h3ac3d7aa),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb712338),
	.w1(32'hbb32ea2d),
	.w2(32'hba8ce34e),
	.w3(32'hbbd0f4c5),
	.w4(32'hbb8268ff),
	.w5(32'hbb2cd6c4),
	.w6(32'hbb241a93),
	.w7(32'h3b2474b3),
	.w8(32'h3b235f1a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02365b),
	.w1(32'hbba822a6),
	.w2(32'h3b8447b2),
	.w3(32'hbbcbdf19),
	.w4(32'hbb58d00e),
	.w5(32'h3a84f19d),
	.w6(32'hbbbf9419),
	.w7(32'hbbd6afd6),
	.w8(32'hbac8aa96),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc370c82),
	.w1(32'hbbb93039),
	.w2(32'hbc9b2eaf),
	.w3(32'h3a4eab52),
	.w4(32'hbc3ca334),
	.w5(32'hbcc3381f),
	.w6(32'h3c9b0f77),
	.w7(32'h3bf74525),
	.w8(32'hbb5d809c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bd4e3),
	.w1(32'hbb76938b),
	.w2(32'hbc13e910),
	.w3(32'hb955f668),
	.w4(32'hbb12d144),
	.w5(32'hbc298bf4),
	.w6(32'h3c18c513),
	.w7(32'h3c3ba77f),
	.w8(32'hbbed4f18),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb14b97),
	.w1(32'hbbec89d6),
	.w2(32'h3a906a01),
	.w3(32'hbb33c0a7),
	.w4(32'hbbb84dad),
	.w5(32'h3b6cb8c7),
	.w6(32'hbc03585b),
	.w7(32'hbb7dabb6),
	.w8(32'h3a8595aa),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c526a),
	.w1(32'hbab6fb03),
	.w2(32'hbba04a2b),
	.w3(32'h3c270318),
	.w4(32'hbb6a23a5),
	.w5(32'h3b00c7d2),
	.w6(32'h3c52bcd0),
	.w7(32'h3ba4a25c),
	.w8(32'h3bb2373d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0aa44e),
	.w1(32'hbb46e8e8),
	.w2(32'hbb631405),
	.w3(32'h3b1c1caf),
	.w4(32'hbb7a6314),
	.w5(32'hbb111ae1),
	.w6(32'h3b5a0eae),
	.w7(32'hbb047f30),
	.w8(32'hbb817656),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0afe68),
	.w1(32'h3bd5406a),
	.w2(32'h3b1f6311),
	.w3(32'hbb70d950),
	.w4(32'h3bb522a8),
	.w5(32'h38908f2e),
	.w6(32'hbb2837b3),
	.w7(32'h3956ea05),
	.w8(32'h3a7f6dfb),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3eb2cd),
	.w1(32'hb95b5382),
	.w2(32'h3b858c9d),
	.w3(32'hba92d140),
	.w4(32'h3b691cb8),
	.w5(32'hba5f8d81),
	.w6(32'hba62c3e7),
	.w7(32'h39eeca57),
	.w8(32'h3b9dd247),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6441c0),
	.w1(32'hba056600),
	.w2(32'h39bcb47e),
	.w3(32'hbb0a808c),
	.w4(32'h3ab0cf23),
	.w5(32'h3aa9a1e7),
	.w6(32'h3b378db8),
	.w7(32'h3b574b66),
	.w8(32'hbafbea98),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acf568),
	.w1(32'h3b443ccc),
	.w2(32'h39bf9e65),
	.w3(32'hbb69fc78),
	.w4(32'h3b394c96),
	.w5(32'hbab5ea41),
	.w6(32'hbbb931e4),
	.w7(32'h3b177990),
	.w8(32'h3b61f3ef),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba081a8),
	.w1(32'hbc0eaff6),
	.w2(32'hbc656678),
	.w3(32'hbc7bde03),
	.w4(32'hbba73ee9),
	.w5(32'h39943b14),
	.w6(32'h3b17006a),
	.w7(32'hbbf6e830),
	.w8(32'hbc2260fd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacebd78),
	.w1(32'hbbb694e1),
	.w2(32'hba826a99),
	.w3(32'hbb86cd78),
	.w4(32'hbb66e489),
	.w5(32'hbad50669),
	.w6(32'h3bcbc2d1),
	.w7(32'h3bb587f9),
	.w8(32'hbbb69c90),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d275d),
	.w1(32'h3a8aa339),
	.w2(32'hbbc9724d),
	.w3(32'hbb3c5d75),
	.w4(32'hbba03f2a),
	.w5(32'h3b5d62cc),
	.w6(32'h3c14c0bc),
	.w7(32'h3a754da2),
	.w8(32'hbb5d9225),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89ca79),
	.w1(32'h3c00387e),
	.w2(32'h3b1af1f7),
	.w3(32'h3bad6ac6),
	.w4(32'hba1c45b6),
	.w5(32'h3a4a9c0d),
	.w6(32'h3b164d2d),
	.w7(32'hbb2449f7),
	.w8(32'hbb124f44),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba106f9),
	.w1(32'h3baa18b4),
	.w2(32'h3c39ea8d),
	.w3(32'h3b2943b3),
	.w4(32'h3b6e814f),
	.w5(32'h3c578a0f),
	.w6(32'h39b117cb),
	.w7(32'hb920a203),
	.w8(32'h3c1e3a44),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ca061),
	.w1(32'h3b3801de),
	.w2(32'h3b5898d3),
	.w3(32'h3c2b5fb6),
	.w4(32'h3c102cb0),
	.w5(32'h3aebe969),
	.w6(32'h3bc1cadd),
	.w7(32'h3bb0562f),
	.w8(32'hbb6eca13),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9883),
	.w1(32'h3b1b1def),
	.w2(32'h3b435883),
	.w3(32'h39602a96),
	.w4(32'hba6a8522),
	.w5(32'hbafcf906),
	.w6(32'hbbae1b06),
	.w7(32'hbbc23e1f),
	.w8(32'hbb33c745),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e7163),
	.w1(32'hbbbb3326),
	.w2(32'hbb9bb929),
	.w3(32'hbc3ee617),
	.w4(32'hbc7435de),
	.w5(32'hbbe1bc18),
	.w6(32'hbb65d5c4),
	.w7(32'hbb99b6ff),
	.w8(32'hbc0eaf3f),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac434a1),
	.w1(32'h3a57d013),
	.w2(32'hba9cc530),
	.w3(32'hbab07ba0),
	.w4(32'hbba4b489),
	.w5(32'hbb37a9a4),
	.w6(32'hb9e7eb8b),
	.w7(32'hbbbcb7a0),
	.w8(32'hbb12dc93),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a3bac),
	.w1(32'hbad19444),
	.w2(32'hbb29ec72),
	.w3(32'hbb08e37d),
	.w4(32'hbbe1cc6e),
	.w5(32'h3b41f4f2),
	.w6(32'hbb58a34b),
	.w7(32'hbbb036fc),
	.w8(32'h3b59df2e),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bae5b),
	.w1(32'h3b4c4a3b),
	.w2(32'h3a9d0e70),
	.w3(32'h3c318773),
	.w4(32'h3c5d96a7),
	.w5(32'h39c3cde3),
	.w6(32'h3c4ad52d),
	.w7(32'h3c2c6b83),
	.w8(32'h3b4886e2),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52d97c),
	.w1(32'h3ba159fb),
	.w2(32'h393822e0),
	.w3(32'h3bbbd8bd),
	.w4(32'h3bafb120),
	.w5(32'h3bae99df),
	.w6(32'h3bcc5364),
	.w7(32'h3bbbd2d7),
	.w8(32'h3b7098b5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66cec2),
	.w1(32'hbae14cce),
	.w2(32'h3b0843f9),
	.w3(32'h3bac33e6),
	.w4(32'hbb8ecefc),
	.w5(32'h3b3b031a),
	.w6(32'h3b6402f3),
	.w7(32'hbad54166),
	.w8(32'h3a7b1a3d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b774697),
	.w1(32'hbb80b8ad),
	.w2(32'h3c106891),
	.w3(32'h3b33cf72),
	.w4(32'hbb46140e),
	.w5(32'h3b8dadd3),
	.w6(32'hb9b9e863),
	.w7(32'hbba03c2d),
	.w8(32'h3a256eef),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24cd9e),
	.w1(32'hbc16ba7e),
	.w2(32'hbce5b494),
	.w3(32'hbc2c8c8e),
	.w4(32'hbbbfac75),
	.w5(32'hbc2b8403),
	.w6(32'hbbe27bcc),
	.w7(32'hbc0f7a73),
	.w8(32'hbcee7045),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4714c),
	.w1(32'hb7c6bc5a),
	.w2(32'hbb5892ef),
	.w3(32'hbbddb4cf),
	.w4(32'hbb151166),
	.w5(32'hbbc8c607),
	.w6(32'hbba1d1ff),
	.w7(32'h3a34363b),
	.w8(32'hbb97d4c4),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc576270),
	.w1(32'hbc1fb4a6),
	.w2(32'hbb29ce35),
	.w3(32'hbbd5228e),
	.w4(32'h39a796b2),
	.w5(32'hbb3beece),
	.w6(32'h3a9d16bb),
	.w7(32'h3bef7183),
	.w8(32'h3b9b9be1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule