module layer_10_featuremap_97(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ee591),
	.w1(32'h3b29cbd1),
	.w2(32'h3a4f2206),
	.w3(32'hb99c7ea2),
	.w4(32'h3c01aa36),
	.w5(32'h3c1ea368),
	.w6(32'hbbadaf66),
	.w7(32'hbc174986),
	.w8(32'hbc40ae38),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba54c77),
	.w1(32'hbb18f2f5),
	.w2(32'hbad5386f),
	.w3(32'h3953ff1f),
	.w4(32'hbb06b3e8),
	.w5(32'hb9d81891),
	.w6(32'hba8a598a),
	.w7(32'hba8cb59a),
	.w8(32'h389017e9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dda0df),
	.w1(32'h3b311be1),
	.w2(32'h3b1cd443),
	.w3(32'h3a832e69),
	.w4(32'h3b6996ca),
	.w5(32'h3b94a45f),
	.w6(32'h3b807b46),
	.w7(32'h3b92cc1d),
	.w8(32'h3ba8eaff),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b750264),
	.w1(32'h3b641fb6),
	.w2(32'h3b76b766),
	.w3(32'h3b880de9),
	.w4(32'hbbdf20a2),
	.w5(32'hbbac7abe),
	.w6(32'h3bca35b2),
	.w7(32'h3c2ade5b),
	.w8(32'h3c060178),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad9367),
	.w1(32'hbbc93144),
	.w2(32'h3a0b4cc7),
	.w3(32'hba12a754),
	.w4(32'hbb14c1b4),
	.w5(32'h397db196),
	.w6(32'hbb512a8a),
	.w7(32'h3b001ad8),
	.w8(32'h3c02590b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17e0e0),
	.w1(32'h3c0f4f39),
	.w2(32'h3cb4486b),
	.w3(32'h3bb002fc),
	.w4(32'h39afe1e6),
	.w5(32'h3c60ed1b),
	.w6(32'hb8c323fb),
	.w7(32'h3c467403),
	.w8(32'h3b8e0b00),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61cdfa),
	.w1(32'hbbbbf0c3),
	.w2(32'hbb25fa0c),
	.w3(32'h3bfec849),
	.w4(32'hbb05ba19),
	.w5(32'h3a662506),
	.w6(32'hbb5bf967),
	.w7(32'hbb1e38a4),
	.w8(32'h3b27a87d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b775937),
	.w1(32'h39defeed),
	.w2(32'h3b6b2567),
	.w3(32'h3bbe6c18),
	.w4(32'hbb457c04),
	.w5(32'hb80f491e),
	.w6(32'hbb7eeac4),
	.w7(32'h391a592f),
	.w8(32'hbaff5aab),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa67799),
	.w1(32'h3b614671),
	.w2(32'h3ad7ccdb),
	.w3(32'hba8ddcd4),
	.w4(32'h3ac411ec),
	.w5(32'hb93cdb1e),
	.w6(32'h3a52a89b),
	.w7(32'h39398b98),
	.w8(32'hb996a142),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaebeab),
	.w1(32'hbc0aba4d),
	.w2(32'hbb99dc7f),
	.w3(32'hb9f399e1),
	.w4(32'hbbe5094b),
	.w5(32'hbaf0a7dc),
	.w6(32'hbbdf5f23),
	.w7(32'hbb97220e),
	.w8(32'hbab576ac),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4be3c0),
	.w1(32'hb9b942f1),
	.w2(32'hbafd7a7e),
	.w3(32'h3a74e253),
	.w4(32'hbb0201c3),
	.w5(32'hbb2660ae),
	.w6(32'h3ab44c4b),
	.w7(32'h3ac7692e),
	.w8(32'h3aa485cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178901),
	.w1(32'hbb050eea),
	.w2(32'hbb199bc9),
	.w3(32'hbb9b1a01),
	.w4(32'hbb927e2d),
	.w5(32'hbb80ef73),
	.w6(32'h3a8d4c6e),
	.w7(32'h3b4d5832),
	.w8(32'h3aa53926),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ce2cb),
	.w1(32'h3b0eb41e),
	.w2(32'h3b4a25cf),
	.w3(32'hbaa4534f),
	.w4(32'h3b128417),
	.w5(32'h3b565924),
	.w6(32'h3abc1ae8),
	.w7(32'h3b507281),
	.w8(32'h3a7027bc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a934f),
	.w1(32'hbc9bf6a2),
	.w2(32'hbc51811b),
	.w3(32'h3a5e8f6c),
	.w4(32'hbcb5db6f),
	.w5(32'hbc8cf482),
	.w6(32'hbcd245fd),
	.w7(32'hbca63ef0),
	.w8(32'hbcc31756),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9320e1),
	.w1(32'hbb06b612),
	.w2(32'hbb4930e5),
	.w3(32'hbcb14c8b),
	.w4(32'hbbd9942a),
	.w5(32'hbb9c8886),
	.w6(32'h3b91f0c0),
	.w7(32'h3be0648d),
	.w8(32'h3b930dc1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3902dae5),
	.w1(32'h37d55393),
	.w2(32'h3b265960),
	.w3(32'hbbdbadfb),
	.w4(32'hbb7f2feb),
	.w5(32'hba925bb7),
	.w6(32'hbb8eba18),
	.w7(32'hb9e8a22e),
	.w8(32'hbb46dd74),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba507e9f),
	.w1(32'hbb9a3d7c),
	.w2(32'hbaaa0d32),
	.w3(32'hbb104733),
	.w4(32'hbb7a4ac6),
	.w5(32'hba9b3d2f),
	.w6(32'hbbcf2a19),
	.w7(32'hbba1ee4e),
	.w8(32'hbb8db1b4),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a2e3b),
	.w1(32'hbc096db8),
	.w2(32'hbbc28d72),
	.w3(32'hbb02554a),
	.w4(32'hbbbfe048),
	.w5(32'hbb3eb555),
	.w6(32'hbbb0a474),
	.w7(32'hbb916145),
	.w8(32'hbac44ec9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a8974),
	.w1(32'h3b1646c9),
	.w2(32'h3b50d5ce),
	.w3(32'h395775a4),
	.w4(32'h3b3f43a8),
	.w5(32'h3b8e1aa3),
	.w6(32'h3b6dcce9),
	.w7(32'h3b728a5b),
	.w8(32'h3ba72795),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae6264),
	.w1(32'h3b807fb3),
	.w2(32'hba5e94dd),
	.w3(32'h3bb94afa),
	.w4(32'h3acee5f5),
	.w5(32'hbad1e5af),
	.w6(32'h3aa9c208),
	.w7(32'hbabdb391),
	.w8(32'hbb25c9f0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae994d7),
	.w1(32'h3983de95),
	.w2(32'h3a522fe6),
	.w3(32'hbb2ae7f7),
	.w4(32'hbb09cade),
	.w5(32'hbb46d8d1),
	.w6(32'hbb353d7e),
	.w7(32'h389210e2),
	.w8(32'hbb1cff65),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15057d),
	.w1(32'h3a6b12b7),
	.w2(32'hbb0e7d97),
	.w3(32'hbb19aa81),
	.w4(32'h3c68eead),
	.w5(32'h3c03c671),
	.w6(32'hbb0727ea),
	.w7(32'hbb3eda5a),
	.w8(32'hbb82134f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8decaf),
	.w1(32'h39d0dfbd),
	.w2(32'hbb80c4cb),
	.w3(32'h3b4eb137),
	.w4(32'hb8582900),
	.w5(32'hbb4b4f23),
	.w6(32'h3a9cb362),
	.w7(32'hbaf83517),
	.w8(32'hba73f2cc),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b7b47),
	.w1(32'h3a47e265),
	.w2(32'h3ae5e0a1),
	.w3(32'hbacbcaf5),
	.w4(32'hbb252eb5),
	.w5(32'hbaa54d61),
	.w6(32'hbb572447),
	.w7(32'hba8d6029),
	.w8(32'hbb34bb72),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7e01c),
	.w1(32'h3c09041f),
	.w2(32'h3c196398),
	.w3(32'hba9cc833),
	.w4(32'hbabc739c),
	.w5(32'hbab36a8e),
	.w6(32'h3b82adf2),
	.w7(32'h3c0078c9),
	.w8(32'h3b297984),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b609e4a),
	.w1(32'h3a574138),
	.w2(32'hbae37cff),
	.w3(32'hbb5588f4),
	.w4(32'h3adf0b22),
	.w5(32'h3a2a703d),
	.w6(32'h3c0addea),
	.w7(32'h3c0c9e25),
	.w8(32'h3bbc2020),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd8725),
	.w1(32'h3b42eb3f),
	.w2(32'h39dcb4ab),
	.w3(32'hbb29a94b),
	.w4(32'h39639eb0),
	.w5(32'hbad5fee9),
	.w6(32'h3a6214ab),
	.w7(32'h39b2c2c3),
	.w8(32'hb8d5b288),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5080f2),
	.w1(32'hbc1d3e3b),
	.w2(32'hbc2d0fb3),
	.w3(32'hbaed6a62),
	.w4(32'hbc5feee3),
	.w5(32'hbc4d36b0),
	.w6(32'hbc27bf14),
	.w7(32'hbc107083),
	.w8(32'hbc2e3c0c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc474404),
	.w1(32'hbbef5aa9),
	.w2(32'hbc56e259),
	.w3(32'hbc6b49c4),
	.w4(32'hbb98c152),
	.w5(32'hbc33d895),
	.w6(32'hbbb3e3d8),
	.w7(32'hbc3db629),
	.w8(32'hbb746ba3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1a81e),
	.w1(32'h3ab906e0),
	.w2(32'h3b24be71),
	.w3(32'hbb65542d),
	.w4(32'h3a9eeb38),
	.w5(32'h3afa14c3),
	.w6(32'h3a50b02a),
	.w7(32'h3addd9f1),
	.w8(32'h3a528fb3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aad754),
	.w1(32'h3b232ea4),
	.w2(32'h3b4f66dc),
	.w3(32'h394a4c5f),
	.w4(32'hb99f8ccb),
	.w5(32'hb99af55d),
	.w6(32'h39b6d4d0),
	.w7(32'h3b05ee78),
	.w8(32'hbabde4d2),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ad761),
	.w1(32'h39dd9eb4),
	.w2(32'h39cce670),
	.w3(32'hbafb3a74),
	.w4(32'hba0fe01e),
	.w5(32'hb9cace7d),
	.w6(32'hba2ca5e4),
	.w7(32'h39e4f7e6),
	.w8(32'h3869aacb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b6b08),
	.w1(32'h3bc42d0d),
	.w2(32'hbbad050a),
	.w3(32'hb98bab16),
	.w4(32'h3bdd69f9),
	.w5(32'hbb2f5ee4),
	.w6(32'h3baa0144),
	.w7(32'hba97f496),
	.w8(32'hba9ef864),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ecb8),
	.w1(32'hbaf2df0a),
	.w2(32'hbb955a54),
	.w3(32'hbb8c2aab),
	.w4(32'hb83c7c7c),
	.w5(32'hba25c58c),
	.w6(32'hbabae378),
	.w7(32'h39c139f7),
	.w8(32'h3b1c3fe3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b3f7c),
	.w1(32'hbb6988f9),
	.w2(32'hbb64ef0f),
	.w3(32'h39a51ca8),
	.w4(32'hbb39f598),
	.w5(32'hbaa36402),
	.w6(32'hbb0da8cf),
	.w7(32'hbac8ac61),
	.w8(32'h3a9a539f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943c7ef),
	.w1(32'h3b2426ed),
	.w2(32'h3a9c32a7),
	.w3(32'h3b0d1666),
	.w4(32'hba735bd4),
	.w5(32'hba8e02ae),
	.w6(32'h3b1005b3),
	.w7(32'h3b8a7436),
	.w8(32'h3ad10fd6),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b347c),
	.w1(32'hbb1be039),
	.w2(32'h3b56fd12),
	.w3(32'hbab7ebcb),
	.w4(32'hbb938bbe),
	.w5(32'h3a87a637),
	.w6(32'h3aa4e9c5),
	.w7(32'h3bcfef3e),
	.w8(32'h3c05b90d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf5534),
	.w1(32'hbb5443e7),
	.w2(32'hba370a2c),
	.w3(32'h3b5b09ca),
	.w4(32'hb9cdb3ab),
	.w5(32'h3af77b7b),
	.w6(32'hbae6c9ee),
	.w7(32'hbaf01a08),
	.w8(32'h3ac6b109),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa02c3),
	.w1(32'h3b695cc7),
	.w2(32'h3b8039ad),
	.w3(32'h3b8f56ff),
	.w4(32'hb908fab9),
	.w5(32'h3a773b22),
	.w6(32'h3981b452),
	.w7(32'h3a40fb42),
	.w8(32'h3a0023a0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35385b),
	.w1(32'h39239973),
	.w2(32'hba8647e2),
	.w3(32'h37d19754),
	.w4(32'h3a2743cd),
	.w5(32'hb96a9011),
	.w6(32'h3afe23d2),
	.w7(32'h3aab1eac),
	.w8(32'h3b8452a8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2650),
	.w1(32'hbb0c111c),
	.w2(32'hbb8fbf0f),
	.w3(32'h3af3bbb8),
	.w4(32'hb8b54612),
	.w5(32'hbb2af876),
	.w6(32'h38d84326),
	.w7(32'hbac6186c),
	.w8(32'hbaf2e9f9),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba42cf4),
	.w1(32'hbb922fb2),
	.w2(32'hbbf183c3),
	.w3(32'hbb543504),
	.w4(32'hbbf71cc3),
	.w5(32'hbc081a6d),
	.w6(32'hb9e4d87b),
	.w7(32'h38b7668d),
	.w8(32'hbb43ff03),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba15e6b),
	.w1(32'h3a23ad74),
	.w2(32'hb931cd33),
	.w3(32'hbbe16864),
	.w4(32'h3a83efc7),
	.w5(32'h3a4a7f04),
	.w6(32'hb9083780),
	.w7(32'hb8d304e0),
	.w8(32'h3ac012dd),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af35603),
	.w1(32'hbc3d3bf2),
	.w2(32'hba688afa),
	.w3(32'h3970526c),
	.w4(32'hbc0b8c14),
	.w5(32'h3b12c37d),
	.w6(32'hbc56ce5f),
	.w7(32'hbbd88b6b),
	.w8(32'hbae54e21),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cfd0f),
	.w1(32'hbcac36a6),
	.w2(32'hbcbfdfff),
	.w3(32'h3bc2c2e5),
	.w4(32'hbc8c77cd),
	.w5(32'hbcac466a),
	.w6(32'hbcaec421),
	.w7(32'hbcb8f6b4),
	.w8(32'hbca19607),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9fe118),
	.w1(32'hbc2ab76f),
	.w2(32'hbc486ddc),
	.w3(32'hbc98d2fc),
	.w4(32'hbc199968),
	.w5(32'hbc31b5a3),
	.w6(32'hbc087baf),
	.w7(32'hbc0fafc4),
	.w8(32'hbc24106d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40b004),
	.w1(32'h3b2f02ee),
	.w2(32'h3b68f2fe),
	.w3(32'hbc2b594d),
	.w4(32'hbb72c52a),
	.w5(32'hbb42c443),
	.w6(32'h3c0ae49a),
	.w7(32'h3c310168),
	.w8(32'h3c6a0c4c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b3fea),
	.w1(32'hba8b1943),
	.w2(32'hbba27427),
	.w3(32'h3be6df02),
	.w4(32'h3a232f22),
	.w5(32'hbb36e165),
	.w6(32'h3ace9b49),
	.w7(32'hbb0ced64),
	.w8(32'h3ada068a),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ece09),
	.w1(32'hb884e0e0),
	.w2(32'hbac11433),
	.w3(32'hba058a81),
	.w4(32'hb92a63e0),
	.w5(32'hba6a6b45),
	.w6(32'hba8a3d93),
	.w7(32'hbac2c15d),
	.w8(32'hba816717),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a81559),
	.w1(32'hbb3b5647),
	.w2(32'h3a370dad),
	.w3(32'hba38b20a),
	.w4(32'hbba92838),
	.w5(32'hbb0c236b),
	.w6(32'hbbc5dd97),
	.w7(32'hbb1fb845),
	.w8(32'hbbadddb1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032aac),
	.w1(32'hbc63dd03),
	.w2(32'hbc39c6ad),
	.w3(32'hbb916eda),
	.w4(32'hbc4e83c4),
	.w5(32'hbc22d18c),
	.w6(32'hbc3e637b),
	.w7(32'hbc3e9049),
	.w8(32'hbc3b98d1),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46edf3),
	.w1(32'h3c565001),
	.w2(32'h39bb9c0d),
	.w3(32'hbc410ab9),
	.w4(32'h3b505109),
	.w5(32'hbbc1c95d),
	.w6(32'h3bbdbf92),
	.w7(32'h3b9e1008),
	.w8(32'h3ae090fb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1755ab),
	.w1(32'h3c96fbbf),
	.w2(32'h3d053261),
	.w3(32'hba343609),
	.w4(32'h3ba72044),
	.w5(32'h3c9ae4aa),
	.w6(32'h3bbfcce2),
	.w7(32'h3ca14441),
	.w8(32'h3ba9d0d3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c852102),
	.w1(32'hbbffb14a),
	.w2(32'h3a66116d),
	.w3(32'h3c052731),
	.w4(32'hbbfdbf9c),
	.w5(32'hbb865189),
	.w6(32'hbbbd8c3b),
	.w7(32'h3ac7809b),
	.w8(32'h3bdc84bd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15ad74),
	.w1(32'h3c0ddccc),
	.w2(32'h3bdaaa59),
	.w3(32'h3aa9e7b4),
	.w4(32'h3bf4a209),
	.w5(32'h3bd93c03),
	.w6(32'h3c08ed68),
	.w7(32'h3bde3830),
	.w8(32'h3bfe4763),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd08816),
	.w1(32'hba518ce4),
	.w2(32'hbc2ed4f1),
	.w3(32'h3bdbeb4a),
	.w4(32'h3b0c268e),
	.w5(32'hbbf4133a),
	.w6(32'h3b6d2292),
	.w7(32'hbb95fc11),
	.w8(32'h37a2551a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a989),
	.w1(32'hbc912064),
	.w2(32'hbc6a5353),
	.w3(32'hbb0f1061),
	.w4(32'hbc9829a7),
	.w5(32'hbc819024),
	.w6(32'hbc8e9d55),
	.w7(32'hbc758583),
	.w8(32'hbc7d8504),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72b7f8),
	.w1(32'hbbbe5670),
	.w2(32'h3b639005),
	.w3(32'hbc8c0da2),
	.w4(32'hbb203901),
	.w5(32'h3b99c082),
	.w6(32'hbb4f35fd),
	.w7(32'h3b2e080f),
	.w8(32'h3b0228ac),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0763c3),
	.w1(32'hba5a755a),
	.w2(32'hbb8683d9),
	.w3(32'h3ac6f31f),
	.w4(32'hba328000),
	.w5(32'hbae8fa71),
	.w6(32'hba1a354a),
	.w7(32'hbb50e4e4),
	.w8(32'h3a37e380),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba592692),
	.w1(32'h3af6e057),
	.w2(32'h3a8cae49),
	.w3(32'h3a72e605),
	.w4(32'hbaa740a7),
	.w5(32'hbabccab3),
	.w6(32'hbb186fa7),
	.w7(32'hbae2ee49),
	.w8(32'hbb1f5deb),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e851),
	.w1(32'h3b9031e8),
	.w2(32'h3b63d0cf),
	.w3(32'hbad478f0),
	.w4(32'h3ba055ee),
	.w5(32'h3bad08d6),
	.w6(32'h3be02557),
	.w7(32'h3bc33732),
	.w8(32'h3bf2b23d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb09fc2),
	.w1(32'h3a33b8c0),
	.w2(32'hb9f4e43f),
	.w3(32'h3bd17eec),
	.w4(32'hbaaa481d),
	.w5(32'hbb126be3),
	.w6(32'hbb37ac6b),
	.w7(32'hbb489ab0),
	.w8(32'hbb69d182),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaade4d7),
	.w1(32'h3c460a62),
	.w2(32'hbbb8e113),
	.w3(32'hbb70b79e),
	.w4(32'h3caa3721),
	.w5(32'h39c5a6bd),
	.w6(32'h3c2d7c4d),
	.w7(32'hbb16eacc),
	.w8(32'h3980dccc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c2af5),
	.w1(32'hbbef11c7),
	.w2(32'hba894118),
	.w3(32'hba464b70),
	.w4(32'hbbb71195),
	.w5(32'h3a844798),
	.w6(32'hbbfe2985),
	.w7(32'hbb8fd1cd),
	.w8(32'hba13f98e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c0f00),
	.w1(32'hbb33bce0),
	.w2(32'hbb66108a),
	.w3(32'h3b850325),
	.w4(32'hbb1e8b9f),
	.w5(32'hba8aca8c),
	.w6(32'hbacd996e),
	.w7(32'hb990fba5),
	.w8(32'h3ad5ef55),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a294de),
	.w1(32'h3ae0814d),
	.w2(32'h3c766756),
	.w3(32'hba624875),
	.w4(32'h3b24cf5c),
	.w5(32'h3c83e29e),
	.w6(32'h3ab89a36),
	.w7(32'h3c5bcd37),
	.w8(32'h3b2b2fc3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4753ed),
	.w1(32'h3a234bde),
	.w2(32'hbaa5b463),
	.w3(32'h3b5f56fb),
	.w4(32'hb901c0f7),
	.w5(32'hbb2894dd),
	.w6(32'h3b870935),
	.w7(32'h3af7b648),
	.w8(32'hbb7315fb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2d12d),
	.w1(32'hbb159921),
	.w2(32'hba92b4ff),
	.w3(32'hbbfe09e2),
	.w4(32'hbadc51f0),
	.w5(32'hb9ede2c0),
	.w6(32'h3a716f4b),
	.w7(32'h3b2605d5),
	.w8(32'h389e1212),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e05b9),
	.w1(32'h3ac4aaff),
	.w2(32'h3b822288),
	.w3(32'hba9eb4ce),
	.w4(32'hbba4dbbb),
	.w5(32'hbb4a977b),
	.w6(32'hbb467a38),
	.w7(32'h3b0413a3),
	.w8(32'hbae062b7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381bfba7),
	.w1(32'hbd0d9598),
	.w2(32'hbcfc244f),
	.w3(32'hbb688e86),
	.w4(32'hbd08f4e4),
	.w5(32'hbcf7ed0f),
	.w6(32'hbcf770c1),
	.w7(32'hbce24afe),
	.w8(32'hbd011e51),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1154c2),
	.w1(32'hbb4097ba),
	.w2(32'hbbad1fec),
	.w3(32'hbd120426),
	.w4(32'hbaff5bcd),
	.w5(32'hbb1282be),
	.w6(32'hbb0d6e19),
	.w7(32'hbb933c29),
	.w8(32'hbafaa570),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb112b8f),
	.w1(32'hb9f01c73),
	.w2(32'h39b0c587),
	.w3(32'h39947f45),
	.w4(32'hbb50a0c8),
	.w5(32'hbaca2bf1),
	.w6(32'hbb6ed3eb),
	.w7(32'hba96c7e8),
	.w8(32'hbb29db58),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f4eca),
	.w1(32'h3b36b8d9),
	.w2(32'h3b1a5f69),
	.w3(32'hbadb40c5),
	.w4(32'hba3b1668),
	.w5(32'hb9539256),
	.w6(32'hba1bc27e),
	.w7(32'h385bbb7d),
	.w8(32'hba1c69b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b120588),
	.w1(32'h3adce15b),
	.w2(32'h3ae47ee8),
	.w3(32'hb8fdd1dc),
	.w4(32'hb9446222),
	.w5(32'hb92dcc28),
	.w6(32'h3836d7fa),
	.w7(32'h3b3c7c51),
	.w8(32'h3a868ad1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cfe02),
	.w1(32'hbb41ae24),
	.w2(32'hbb505c93),
	.w3(32'h3a56d798),
	.w4(32'hbbb80d87),
	.w5(32'hbb803d9c),
	.w6(32'hbacf025a),
	.w7(32'h3967bbf5),
	.w8(32'h3a606bff),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b1143),
	.w1(32'hbae15104),
	.w2(32'hbba10680),
	.w3(32'hbb1f1fc7),
	.w4(32'h39eb3c3c),
	.w5(32'h3ac77eae),
	.w6(32'h3c105e04),
	.w7(32'h3b99b58f),
	.w8(32'h3ad1668f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7328b0),
	.w1(32'hbb4ce297),
	.w2(32'h3b9fb8ff),
	.w3(32'h3b4e5edf),
	.w4(32'hbbba6ca8),
	.w5(32'h3ab4f02b),
	.w6(32'hbc1d7811),
	.w7(32'hbb1b2bb5),
	.w8(32'hbbbf1210),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a782bb8),
	.w1(32'h3b995c3d),
	.w2(32'hbb58ec08),
	.w3(32'hbb10f504),
	.w4(32'h3b91c265),
	.w5(32'hbb567cec),
	.w6(32'h3b8fd115),
	.w7(32'hbadb28f4),
	.w8(32'h3b0d3e94),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed8876),
	.w1(32'hba9e1277),
	.w2(32'hbb09676b),
	.w3(32'h3ae01749),
	.w4(32'hb968cc32),
	.w5(32'h3a5042e9),
	.w6(32'hba201c2f),
	.w7(32'h3a58bd99),
	.w8(32'h3b3cd553),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bd10e),
	.w1(32'h3b83c069),
	.w2(32'h3bd145a9),
	.w3(32'h3a8062ac),
	.w4(32'h39f4931e),
	.w5(32'h3acff3cd),
	.w6(32'h3a5337cd),
	.w7(32'h3b7488c8),
	.w8(32'hbb14cd0a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebc0c4),
	.w1(32'hbaf0c932),
	.w2(32'hbb0a0b11),
	.w3(32'hbb348154),
	.w4(32'hbadebe12),
	.w5(32'hbb400954),
	.w6(32'h3b72ea1f),
	.w7(32'h3b5897ee),
	.w8(32'hbb2da818),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde10ba),
	.w1(32'hbc13803d),
	.w2(32'hbc018071),
	.w3(32'hbbd9efb4),
	.w4(32'hbc472c27),
	.w5(32'hbc3e87d9),
	.w6(32'hbc3b4bd7),
	.w7(32'hbc2e1864),
	.w8(32'hbc2d438f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc195acb),
	.w1(32'h3c58d288),
	.w2(32'h3c18fac1),
	.w3(32'hbc36582f),
	.w4(32'h3ba692f2),
	.w5(32'h3a612694),
	.w6(32'h3c496a49),
	.w7(32'h3c2dccad),
	.w8(32'h3b7c736d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06fd96),
	.w1(32'hba986ad2),
	.w2(32'hbb73a2bb),
	.w3(32'hbb6b43c8),
	.w4(32'h3a3a6a64),
	.w5(32'hb9f3d877),
	.w6(32'hbb052395),
	.w7(32'hbba64d0c),
	.w8(32'hbb844df1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb358360),
	.w1(32'h3b1de9d7),
	.w2(32'h3bb71491),
	.w3(32'h3780cf62),
	.w4(32'h3a421863),
	.w5(32'h3b6b5ed0),
	.w6(32'h3b9da84a),
	.w7(32'h3bb951bd),
	.w8(32'h3af318c7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fddea),
	.w1(32'hbc237c43),
	.w2(32'hbc14bb00),
	.w3(32'hbb88e62e),
	.w4(32'hbc19cae9),
	.w5(32'hbc0f0a97),
	.w6(32'hbc215924),
	.w7(32'hbc201b9a),
	.w8(32'hbc2ef46e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c7bdb),
	.w1(32'hbc13d30a),
	.w2(32'hbc2c1e06),
	.w3(32'hbc179f4b),
	.w4(32'hbc09e048),
	.w5(32'hbc188d33),
	.w6(32'hbbeeab6b),
	.w7(32'hbc28a555),
	.w8(32'hbc2b0c36),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e6c76),
	.w1(32'h3b1d51ce),
	.w2(32'h3b08880e),
	.w3(32'hbc2134c4),
	.w4(32'hb96cebe4),
	.w5(32'hbaa3540c),
	.w6(32'h393bb903),
	.w7(32'h3a987cea),
	.w8(32'hb996ec24),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e7289),
	.w1(32'h3bea77ca),
	.w2(32'h3bcdf22f),
	.w3(32'hba484925),
	.w4(32'h3bad6da5),
	.w5(32'h3ba15f7e),
	.w6(32'h3bbe3f97),
	.w7(32'h3b98465d),
	.w8(32'h3b89df22),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81057c),
	.w1(32'h3a8164e9),
	.w2(32'h3ad216d3),
	.w3(32'h3b6a0884),
	.w4(32'hba8dd198),
	.w5(32'hba98ad04),
	.w6(32'hba381d7a),
	.w7(32'h3a923a0d),
	.w8(32'hb9cba356),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bacc6),
	.w1(32'h3b3931e9),
	.w2(32'h3b50fe94),
	.w3(32'hba7bfac2),
	.w4(32'h3a88dbdd),
	.w5(32'h39f709d2),
	.w6(32'h378ab568),
	.w7(32'h3af0dd0d),
	.w8(32'h3a2e4d9d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0461af),
	.w1(32'hbc4cad23),
	.w2(32'hbbf7176f),
	.w3(32'h3902cbd9),
	.w4(32'hbc231acc),
	.w5(32'hbbaf1ba6),
	.w6(32'hbc257f2d),
	.w7(32'hbc0eb8ee),
	.w8(32'hbbbfab6b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb93f98),
	.w1(32'h3ba9f0ee),
	.w2(32'h3b9fb6fa),
	.w3(32'hbb7d2a92),
	.w4(32'h3b489487),
	.w5(32'h3ba41343),
	.w6(32'h3a241d9f),
	.w7(32'h3742f67b),
	.w8(32'h381623d6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36dfb0),
	.w1(32'hbbd9d8ac),
	.w2(32'hbc739029),
	.w3(32'h3b9e189d),
	.w4(32'hbb6f1f00),
	.w5(32'hbc4e9fa4),
	.w6(32'h3a45aa3f),
	.w7(32'hbbf6e8fd),
	.w8(32'hbae36520),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd323ff),
	.w1(32'h3b9e3fd6),
	.w2(32'h3b32f1f1),
	.w3(32'hbb5a26d4),
	.w4(32'h3bd00db1),
	.w5(32'h3bb8a14d),
	.w6(32'h3c0c9af4),
	.w7(32'h3beac65c),
	.w8(32'h3bd13b13),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49b04c),
	.w1(32'hbb446ca4),
	.w2(32'h3bf01ac2),
	.w3(32'h3b8e0bdb),
	.w4(32'hbb124c9f),
	.w5(32'h3c2c103c),
	.w6(32'hbc1728f9),
	.w7(32'hbb0ed7e7),
	.w8(32'hbc30e0c0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d24c5),
	.w1(32'h3b388d65),
	.w2(32'h3adc6a89),
	.w3(32'h3aad0b0a),
	.w4(32'h3b552715),
	.w5(32'h3b35814c),
	.w6(32'h3b85c05d),
	.w7(32'h3aec75b5),
	.w8(32'hbab96ee8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb989d099),
	.w1(32'h3c09dfb1),
	.w2(32'hbb8a4d47),
	.w3(32'h3a8bf0af),
	.w4(32'h3c02af42),
	.w5(32'h382e29be),
	.w6(32'h3bd27671),
	.w7(32'h381985b0),
	.w8(32'hbb76de8c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc3c3),
	.w1(32'h3b29ae73),
	.w2(32'h3a600490),
	.w3(32'hbb9e9b9c),
	.w4(32'h3b10766e),
	.w5(32'h39c63416),
	.w6(32'h3b82ed83),
	.w7(32'h3b234ac8),
	.w8(32'h3b683bca),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b456309),
	.w1(32'h3c7a11d7),
	.w2(32'h3cda11d1),
	.w3(32'h398e24f1),
	.w4(32'h3b946146),
	.w5(32'h3c794912),
	.w6(32'h3bc62573),
	.w7(32'h3c92c0ba),
	.w8(32'h3baac597),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c226efa),
	.w1(32'hbb950af0),
	.w2(32'hbaf06ae1),
	.w3(32'h3bba754c),
	.w4(32'hbb3c6c0e),
	.w5(32'h3b11129f),
	.w6(32'h392a90c1),
	.w7(32'h3bc7edb9),
	.w8(32'h3c41ee8d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd22b94),
	.w1(32'hbbadb21c),
	.w2(32'hbbcfdab3),
	.w3(32'h3b0ab07c),
	.w4(32'hbaaa84c3),
	.w5(32'hbb7b2270),
	.w6(32'hbba86dca),
	.w7(32'hbb828a71),
	.w8(32'hb9738910),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37bdd7),
	.w1(32'hbb891ebe),
	.w2(32'h3bfaa2ee),
	.w3(32'h3907e737),
	.w4(32'hbc13be80),
	.w5(32'h3b0eca99),
	.w6(32'hbc7c48f4),
	.w7(32'hbb88b099),
	.w8(32'hbc1aa59d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d564f),
	.w1(32'hb8ced5a5),
	.w2(32'h3b39ec22),
	.w3(32'hbb83d281),
	.w4(32'hbb821f66),
	.w5(32'hba24f3c9),
	.w6(32'hbb3a8a56),
	.w7(32'h3acde219),
	.w8(32'hba9e8bcc),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab238ac),
	.w1(32'hbb0292bb),
	.w2(32'h3b543844),
	.w3(32'hbb06e12e),
	.w4(32'hbb979d6b),
	.w5(32'h3a043a3a),
	.w6(32'hbbf41b6a),
	.w7(32'hbb0c417a),
	.w8(32'hbb8f0de0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c131a),
	.w1(32'h3b9053d3),
	.w2(32'h380b7b78),
	.w3(32'hbae25738),
	.w4(32'h3af595f8),
	.w5(32'hba803485),
	.w6(32'h3ae456a5),
	.w7(32'h37fb8cba),
	.w8(32'hb96a4edd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3945979f),
	.w1(32'h3bcdb025),
	.w2(32'h3b6b355d),
	.w3(32'hbaa322ad),
	.w4(32'h3beb7b9e),
	.w5(32'h3bd03b3a),
	.w6(32'h3bc89615),
	.w7(32'h3bb9a84c),
	.w8(32'h3bc88a68),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ef5fc),
	.w1(32'h3b4ef866),
	.w2(32'h3b37f4f7),
	.w3(32'h3b597b06),
	.w4(32'hb94e51a9),
	.w5(32'hbacac06a),
	.w6(32'hb9cb8af3),
	.w7(32'h3abd8631),
	.w8(32'hba965391),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5a6c),
	.w1(32'hbb0cb6a2),
	.w2(32'h3b92a369),
	.w3(32'hbafb27e8),
	.w4(32'hbb837aa9),
	.w5(32'h3b00d0db),
	.w6(32'hbbf4b4b5),
	.w7(32'hba878ddc),
	.w8(32'hbb7f9bad),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c4270),
	.w1(32'hbc2034ea),
	.w2(32'hbc245734),
	.w3(32'hbaa55f17),
	.w4(32'hbc0a5dd6),
	.w5(32'hbc194551),
	.w6(32'hbbd22dce),
	.w7(32'hbbedae26),
	.w8(32'hbc0366ca),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d8994),
	.w1(32'h3b6d6170),
	.w2(32'h3b72fc06),
	.w3(32'hbc157c1f),
	.w4(32'hbad98d73),
	.w5(32'hbb01728f),
	.w6(32'hba8dfc10),
	.w7(32'h3afcf348),
	.w8(32'hbab18075),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f24f10),
	.w1(32'h3b9340b1),
	.w2(32'hbc1b027b),
	.w3(32'hbb1b9447),
	.w4(32'h3c2752c4),
	.w5(32'hbb2400e0),
	.w6(32'h3b97bfa5),
	.w7(32'hbbba7af4),
	.w8(32'hbbb52c53),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f0677),
	.w1(32'h3b87d519),
	.w2(32'h3c19889a),
	.w3(32'hbb082516),
	.w4(32'hbb83b3ee),
	.w5(32'h3a1eec42),
	.w6(32'hba692b78),
	.w7(32'h3b9d49a0),
	.w8(32'hb951de25),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79b224),
	.w1(32'h39f91d89),
	.w2(32'hbb22b42f),
	.w3(32'hbab0c4eb),
	.w4(32'hb8af92fd),
	.w5(32'hbaf80cc0),
	.w6(32'h3ba47f08),
	.w7(32'h3b27c6bc),
	.w8(32'h3ad4b8c7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd09ea),
	.w1(32'hbc17291d),
	.w2(32'hbbecf364),
	.w3(32'hba6c248c),
	.w4(32'hbc1cd366),
	.w5(32'hbc11801c),
	.w6(32'hbc2a2b41),
	.w7(32'hbc10d10d),
	.w8(32'hbc20fa71),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0755c9),
	.w1(32'hbb561c04),
	.w2(32'h3bbb3f91),
	.w3(32'hbc2d9a79),
	.w4(32'hbbd4c85a),
	.w5(32'h3ad206d6),
	.w6(32'hbc38267f),
	.w7(32'hbb3e6e31),
	.w8(32'hbbd74d02),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64df1a),
	.w1(32'h39e5b790),
	.w2(32'h3b7ae03a),
	.w3(32'hbb315588),
	.w4(32'hbb454c48),
	.w5(32'h39b7bcd0),
	.w6(32'hbb8a16b0),
	.w7(32'hb8b0c14e),
	.w8(32'hbb2df544),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7e98f),
	.w1(32'h3a2e399f),
	.w2(32'h3bb117ca),
	.w3(32'hbac55a8d),
	.w4(32'hbb7024f9),
	.w5(32'h3aac98bc),
	.w6(32'hbbb40a3c),
	.w7(32'h391b0ddc),
	.w8(32'hbb2a024a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17e10b),
	.w1(32'hbae2b84c),
	.w2(32'hbb6a8ac2),
	.w3(32'hba45eca5),
	.w4(32'h3a9022e6),
	.w5(32'hbaa99b26),
	.w6(32'hbba1ab16),
	.w7(32'hbbb4a2c6),
	.w8(32'hbbd4cc86),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b4084),
	.w1(32'h3b08a3b9),
	.w2(32'h3ba92400),
	.w3(32'hbbb7f034),
	.w4(32'h3b2a7f8b),
	.w5(32'h3bb88b88),
	.w6(32'h3b9ef541),
	.w7(32'h3bcfd4ac),
	.w8(32'h3b9df190),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d3ff9),
	.w1(32'hbbec6be6),
	.w2(32'hb94ddb9b),
	.w3(32'h3b815299),
	.w4(32'hbc4e682e),
	.w5(32'hbbe7ba1a),
	.w6(32'hbc30ad38),
	.w7(32'hbaf039ab),
	.w8(32'hbc0acfcd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cc307),
	.w1(32'hb86d4262),
	.w2(32'h39d40105),
	.w3(32'hbc28a005),
	.w4(32'hbbe55be1),
	.w5(32'hbb60ec90),
	.w6(32'hbc138152),
	.w7(32'hbbce583c),
	.w8(32'hbc639cc6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ada34),
	.w1(32'h3a63ae84),
	.w2(32'h3ae7851e),
	.w3(32'hbc225e92),
	.w4(32'hbb0fc33f),
	.w5(32'hba883750),
	.w6(32'hbb73ff4c),
	.w7(32'hbaeec5cc),
	.w8(32'hbb5a8161),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c64207),
	.w1(32'hbba9e7a6),
	.w2(32'hbbff2dbe),
	.w3(32'hbaf902c8),
	.w4(32'h3a64fa7d),
	.w5(32'hbb25401a),
	.w6(32'hbc1a7bf9),
	.w7(32'hbc496b8d),
	.w8(32'hbc0b4aeb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1560b),
	.w1(32'h3c979547),
	.w2(32'h3d2c2b93),
	.w3(32'hbb3bfd0a),
	.w4(32'h3bb0490b),
	.w5(32'h3ce67f9b),
	.w6(32'h3b45dbf2),
	.w7(32'h3cc0e6b3),
	.w8(32'h3b85469a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab829b),
	.w1(32'h3c0ebea0),
	.w2(32'h3bf58536),
	.w3(32'h3c48526d),
	.w4(32'h3b6e6332),
	.w5(32'h3ae50c96),
	.w6(32'h3b4e5bfa),
	.w7(32'h3baa8b27),
	.w8(32'h3aa59c2d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844806),
	.w1(32'hbb08d88d),
	.w2(32'h3bc4a095),
	.w3(32'h3a3413d0),
	.w4(32'hbad7cf73),
	.w5(32'h3ba74a8a),
	.w6(32'hbb348744),
	.w7(32'h3b708932),
	.w8(32'h39b2c1ec),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bb2b2),
	.w1(32'hba8dafe5),
	.w2(32'h3b2824ec),
	.w3(32'hb9efcc3b),
	.w4(32'hbafee0f9),
	.w5(32'h3ac0ddc0),
	.w6(32'hba88791a),
	.w7(32'h3ac9cc4e),
	.w8(32'h3b652090),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e960c),
	.w1(32'hba95319e),
	.w2(32'h3b790f63),
	.w3(32'h3b364439),
	.w4(32'h39e2e383),
	.w5(32'h3a82b507),
	.w6(32'hbb07e71b),
	.w7(32'h3a862083),
	.w8(32'hbb337c24),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac2429),
	.w1(32'hb92940fc),
	.w2(32'hbaf5d745),
	.w3(32'h3b4cb260),
	.w4(32'hb922fcf0),
	.w5(32'hbaeee81e),
	.w6(32'hb9e5d446),
	.w7(32'hbaa273c8),
	.w8(32'h39dfe23f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac02e64),
	.w1(32'hbae82c8b),
	.w2(32'hbb01e87d),
	.w3(32'h3926c8f1),
	.w4(32'hbb5d081f),
	.w5(32'hbb3bc18d),
	.w6(32'hbb5de46c),
	.w7(32'hbb261081),
	.w8(32'h3979ffab),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab697bf),
	.w1(32'h3b26e7ac),
	.w2(32'h3bbb00c0),
	.w3(32'h3a5ed86f),
	.w4(32'hbba58e01),
	.w5(32'hbacf7ecc),
	.w6(32'hba9a3e58),
	.w7(32'hb9d61005),
	.w8(32'hb942339d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9b223),
	.w1(32'h3a92d406),
	.w2(32'h3b56dc03),
	.w3(32'hbb61875a),
	.w4(32'h3b13c5e2),
	.w5(32'h3b897302),
	.w6(32'h3b03bfaf),
	.w7(32'h3b494b2c),
	.w8(32'h3b82a7e2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75aef5),
	.w1(32'hba85a425),
	.w2(32'h3b5adce9),
	.w3(32'h3b13a797),
	.w4(32'hbabfa957),
	.w5(32'h3ac6c8b0),
	.w6(32'hba8988b0),
	.w7(32'h3a30ffc1),
	.w8(32'h3bf00caf),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083943),
	.w1(32'h3a0d5203),
	.w2(32'hbb5a03fb),
	.w3(32'h3bc0c5ae),
	.w4(32'hba65814b),
	.w5(32'hbad0c1fd),
	.w6(32'hbaa2f2d8),
	.w7(32'hba64dcd0),
	.w8(32'h39258eba),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a129e48),
	.w1(32'hb98ac922),
	.w2(32'h3a8da457),
	.w3(32'h3a0110a9),
	.w4(32'hba9e98a6),
	.w5(32'h3aac3e4b),
	.w6(32'hb9bf1889),
	.w7(32'h3a380c4e),
	.w8(32'h3ae30072),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addd970),
	.w1(32'hb98ce70f),
	.w2(32'h3b150d24),
	.w3(32'h3b0293a9),
	.w4(32'h39d10cae),
	.w5(32'h3b2f2355),
	.w6(32'hba90a4f7),
	.w7(32'h3ad324dc),
	.w8(32'h3a80b656),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac51c86),
	.w1(32'hba533f5f),
	.w2(32'hbab2f3c0),
	.w3(32'h3ac9d8f8),
	.w4(32'hbac0b081),
	.w5(32'hbb2894a4),
	.w6(32'hbb270a09),
	.w7(32'hbac850a8),
	.w8(32'h3b8b9674),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3be332),
	.w1(32'hbba0c199),
	.w2(32'hbb890d56),
	.w3(32'h3a88bcc0),
	.w4(32'hbbda45f1),
	.w5(32'hbb486472),
	.w6(32'hbb01fadf),
	.w7(32'hb9c4c8d6),
	.w8(32'h3a265e21),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72e1fe),
	.w1(32'h3980bc02),
	.w2(32'h3b0913c4),
	.w3(32'hbb30e1d6),
	.w4(32'hbb62ba71),
	.w5(32'hba361943),
	.w6(32'hba29d9ad),
	.w7(32'h3a78f376),
	.w8(32'h3b938a33),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77ae8b),
	.w1(32'hbb366baf),
	.w2(32'hbb0f957c),
	.w3(32'h3b503d7c),
	.w4(32'hbb11a6fc),
	.w5(32'hba9a8cd1),
	.w6(32'hbb2da039),
	.w7(32'hbb0d8606),
	.w8(32'hbac9275d),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f6cd3),
	.w1(32'h3af2a571),
	.w2(32'h395565db),
	.w3(32'hb91ad39c),
	.w4(32'hbac54842),
	.w5(32'hba65a130),
	.w6(32'h3a5cbfba),
	.w7(32'hba0835d0),
	.w8(32'hb92131f3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186731),
	.w1(32'h3b851df8),
	.w2(32'h3b69e798),
	.w3(32'hb897242b),
	.w4(32'h3bd2a97b),
	.w5(32'h3b78fa4e),
	.w6(32'h3b8edf04),
	.w7(32'h3b044f4f),
	.w8(32'h3b696d54),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87a561),
	.w1(32'hb9842cfd),
	.w2(32'h3b172e8f),
	.w3(32'h3ad8edfb),
	.w4(32'h397c3296),
	.w5(32'h3ae0b6fb),
	.w6(32'hba4638fe),
	.w7(32'h3aab3946),
	.w8(32'h3b379c83),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c025),
	.w1(32'hbb8c9809),
	.w2(32'h3af4a8f6),
	.w3(32'h3b34604c),
	.w4(32'hba879286),
	.w5(32'h3afc4f6b),
	.w6(32'hbbc0737f),
	.w7(32'hbaca171c),
	.w8(32'hbbbacaaa),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad7842),
	.w1(32'h3a81bcae),
	.w2(32'hba100dbf),
	.w3(32'hbbb11f15),
	.w4(32'hba93de51),
	.w5(32'hbac89096),
	.w6(32'hbae4e783),
	.w7(32'hba307bf2),
	.w8(32'h382b4866),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a230c19),
	.w1(32'h3a85b06c),
	.w2(32'h3afa4ac0),
	.w3(32'hbabbed86),
	.w4(32'h3a274902),
	.w5(32'h3b22ba64),
	.w6(32'h3a736a72),
	.w7(32'h3b3874e3),
	.w8(32'h3b1df23f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241d7c),
	.w1(32'h3a93538a),
	.w2(32'h3af56de8),
	.w3(32'h3af1d969),
	.w4(32'h3a4bb555),
	.w5(32'h3b093e49),
	.w6(32'hb8a1f261),
	.w7(32'h3ad851be),
	.w8(32'h3acf5ae9),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4dbd29),
	.w1(32'hbafd4845),
	.w2(32'h3aafa99a),
	.w3(32'h3a99532d),
	.w4(32'hbbe4e1c5),
	.w5(32'hbb5aa0b6),
	.w6(32'hbb870c46),
	.w7(32'hba5f53cd),
	.w8(32'hbb50c4c2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8eb71),
	.w1(32'h3aa3f4b9),
	.w2(32'hb9cc1e0b),
	.w3(32'hbb2e9482),
	.w4(32'h3b0e5a2f),
	.w5(32'hba557b8b),
	.w6(32'hbb09da55),
	.w7(32'hbaa03da3),
	.w8(32'h394f6b3b),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa38850),
	.w1(32'h3c14f7ce),
	.w2(32'h3be13dd0),
	.w3(32'h3b21bac1),
	.w4(32'h3a672d23),
	.w5(32'hb9d598f3),
	.w6(32'hb8658bb0),
	.w7(32'hbaac5118),
	.w8(32'hbbe44437),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade8545),
	.w1(32'hb815c393),
	.w2(32'h3a788e83),
	.w3(32'hbb9c804a),
	.w4(32'hba1b5876),
	.w5(32'h3a78507e),
	.w6(32'hb91f1279),
	.w7(32'h3a203042),
	.w8(32'h3a7fd586),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa436db),
	.w1(32'hbb4a598c),
	.w2(32'hbb063713),
	.w3(32'h3ad211e6),
	.w4(32'hbb96de6a),
	.w5(32'hbb9305b2),
	.w6(32'hbb55898f),
	.w7(32'hbb022cc3),
	.w8(32'hba2ee510),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb934c590),
	.w1(32'hbc2aee2b),
	.w2(32'hbbd11746),
	.w3(32'hbaaaf218),
	.w4(32'hbba3d732),
	.w5(32'hbbb96ebd),
	.w6(32'hbc9c2450),
	.w7(32'hbbfdfe3f),
	.w8(32'h3aa9d741),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1eae2),
	.w1(32'h3a6a867e),
	.w2(32'hba47efce),
	.w3(32'hbba4d633),
	.w4(32'h3a441579),
	.w5(32'hb9ca6bb7),
	.w6(32'h39ab32b7),
	.w7(32'hb9b67af6),
	.w8(32'h3a1768b4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11857c),
	.w1(32'hb9add450),
	.w2(32'hbb47ef45),
	.w3(32'hb98b1e30),
	.w4(32'hba874e1e),
	.w5(32'hbba41595),
	.w6(32'hbab81fa7),
	.w7(32'hbb1a025b),
	.w8(32'hba632c47),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0db889),
	.w1(32'h3c493f2b),
	.w2(32'h3c9a99a5),
	.w3(32'hbabcc00b),
	.w4(32'h3bd1e484),
	.w5(32'h3c63beec),
	.w6(32'h3c13509f),
	.w7(32'h3c53b989),
	.w8(32'hb9dcc516),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6de1f),
	.w1(32'h3c18e9d0),
	.w2(32'h3b8d4c9a),
	.w3(32'h3b3f5167),
	.w4(32'h3c110d08),
	.w5(32'h3b5d5d88),
	.w6(32'h3bb04116),
	.w7(32'h3ae4a64b),
	.w8(32'hbb0c9d07),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e192),
	.w1(32'hba632d2a),
	.w2(32'h3a82f6e2),
	.w3(32'hbb35dc26),
	.w4(32'hbaf8c146),
	.w5(32'hba086598),
	.w6(32'hba86bdbf),
	.w7(32'h3a1af492),
	.w8(32'hbaa68940),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07303f),
	.w1(32'hbaa9e30d),
	.w2(32'h398263ba),
	.w3(32'hba679ccb),
	.w4(32'hbb2eb875),
	.w5(32'hba6fc821),
	.w6(32'hbae8b88e),
	.w7(32'hba4ffa49),
	.w8(32'hba5cf095),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8baaeaf),
	.w1(32'h3a633404),
	.w2(32'hbc127b48),
	.w3(32'hba4c9589),
	.w4(32'hbae5afad),
	.w5(32'hbc080acf),
	.w6(32'hba920ed2),
	.w7(32'hbc353df6),
	.w8(32'hbba1e5d7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb195e),
	.w1(32'h3c684cf5),
	.w2(32'hba9a7c66),
	.w3(32'hbbbed531),
	.w4(32'h3c91b1c3),
	.w5(32'h3c41b874),
	.w6(32'h3c1ae0f1),
	.w7(32'h3bba8987),
	.w8(32'hbc54e9fe),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b343),
	.w1(32'hbb1597ee),
	.w2(32'hbb7b1914),
	.w3(32'hbc339cf1),
	.w4(32'hbb38bd54),
	.w5(32'hbb8754ec),
	.w6(32'hbb7b74d6),
	.w7(32'hbb2493cc),
	.w8(32'h38f12974),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a29ca),
	.w1(32'hba85666b),
	.w2(32'hb7f7a49a),
	.w3(32'hbb348653),
	.w4(32'hbb41314d),
	.w5(32'hbb1659c4),
	.w6(32'hba9a5dfe),
	.w7(32'hb9d4c9f3),
	.w8(32'hbb05e211),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a9fbe),
	.w1(32'hb9c248c2),
	.w2(32'hbb2dcf28),
	.w3(32'hba2c65c6),
	.w4(32'h38828051),
	.w5(32'hbaca610c),
	.w6(32'hba972acd),
	.w7(32'hba5e5506),
	.w8(32'h3ad2d652),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab57d05),
	.w1(32'h3b2abdda),
	.w2(32'hbb1d5b14),
	.w3(32'hbae78659),
	.w4(32'h3af9e43a),
	.w5(32'hbae53e09),
	.w6(32'h3aad4924),
	.w7(32'hba8fb707),
	.w8(32'hba025750),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a57b26),
	.w1(32'hb9000d2d),
	.w2(32'h3aae4f6e),
	.w3(32'hba257453),
	.w4(32'hba0bb224),
	.w5(32'h3a0e61b9),
	.w6(32'h3882407b),
	.w7(32'h3a80f411),
	.w8(32'h3aca2f74),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b077c4d),
	.w1(32'h39e01c7d),
	.w2(32'hba2cb1e6),
	.w3(32'h3acc531f),
	.w4(32'h397214d5),
	.w5(32'h399c19c4),
	.w6(32'hb9078d31),
	.w7(32'h3ae17905),
	.w8(32'h3b223db7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b247a0d),
	.w1(32'h3ca9584e),
	.w2(32'h3c08cd71),
	.w3(32'h3a7ccbc4),
	.w4(32'h3cc69685),
	.w5(32'h3c12ab69),
	.w6(32'h3c90c14d),
	.w7(32'h3b9af5b7),
	.w8(32'hbb8f36ad),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cb55b),
	.w1(32'hbb2a0d7b),
	.w2(32'hba30b9bb),
	.w3(32'h3b420d26),
	.w4(32'hbb72899b),
	.w5(32'hba936a44),
	.w6(32'hbac5abdb),
	.w7(32'hb8efeb7a),
	.w8(32'h3b0e055e),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a87b887),
	.w1(32'hbb48d4e8),
	.w2(32'hbb8ba66d),
	.w3(32'h385a14f8),
	.w4(32'hbb1b677a),
	.w5(32'hbb3f2095),
	.w6(32'hbb730dd3),
	.w7(32'hbb8b169b),
	.w8(32'hbafcd415),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae47c9d),
	.w1(32'hb962b1d8),
	.w2(32'hba2a44ae),
	.w3(32'hbab70d85),
	.w4(32'hb9bdca75),
	.w5(32'h395edc83),
	.w6(32'hba9d9cad),
	.w7(32'h3a4b27f8),
	.w8(32'h3b63de63),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a228756),
	.w1(32'h3934e4aa),
	.w2(32'h3b824696),
	.w3(32'hb9210674),
	.w4(32'hbab241ea),
	.w5(32'h3b2af60c),
	.w6(32'hba2f799f),
	.w7(32'h3a808c8c),
	.w8(32'hbaa37448),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a3755),
	.w1(32'hba70aa5d),
	.w2(32'hba887b1e),
	.w3(32'h3b0039eb),
	.w4(32'hbb0d13d2),
	.w5(32'hb9644bf9),
	.w6(32'hbaa466a9),
	.w7(32'hb9ab4c57),
	.w8(32'hb981a0bb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdc122),
	.w1(32'h3c07bb89),
	.w2(32'h3bb5f48c),
	.w3(32'h3b131b2b),
	.w4(32'h3ba2b6bb),
	.w5(32'h3ba87b8f),
	.w6(32'h3bc3ac8a),
	.w7(32'h3b8bc600),
	.w8(32'h3b9be80f),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6e1ca2),
	.w1(32'h3c242d34),
	.w2(32'h3cca7db1),
	.w3(32'hba5a112c),
	.w4(32'h3bc393e1),
	.w5(32'h3cc2a2dc),
	.w6(32'h3bc1c3d6),
	.w7(32'h3ccc8b7d),
	.w8(32'hbb70c1b9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963e11a),
	.w1(32'hbacf7161),
	.w2(32'hbb872c39),
	.w3(32'hbb8bc625),
	.w4(32'hbad4029a),
	.w5(32'hbb341721),
	.w6(32'hbb4be9fc),
	.w7(32'hbb93512b),
	.w8(32'hbaade0e4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41480),
	.w1(32'h3ab4bf24),
	.w2(32'h3addd414),
	.w3(32'hba738ae8),
	.w4(32'h39e094b4),
	.w5(32'h3aab82d7),
	.w6(32'h3acee6dc),
	.w7(32'h3aace7ad),
	.w8(32'h3ae40f9c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1fe7e),
	.w1(32'h3b4964f7),
	.w2(32'h3b36357d),
	.w3(32'h3af6089d),
	.w4(32'h3b35386d),
	.w5(32'h3b77ce1d),
	.w6(32'h39015b43),
	.w7(32'h3b469425),
	.w8(32'h3b3b91f0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2a15),
	.w1(32'h3b3030de),
	.w2(32'h3b82dacd),
	.w3(32'h3b20fe72),
	.w4(32'h3a9de78e),
	.w5(32'hbb38f507),
	.w6(32'hb8ea7cd4),
	.w7(32'h3a269d47),
	.w8(32'h3af753cc),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a546e03),
	.w1(32'hb7e89428),
	.w2(32'hb90adcc5),
	.w3(32'hbb433989),
	.w4(32'hb9f7dd24),
	.w5(32'hba5df2c1),
	.w6(32'hba782db5),
	.w7(32'hbaeab719),
	.w8(32'h3b43a6b5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ecb1),
	.w1(32'hbb864be5),
	.w2(32'h3b19bc4a),
	.w3(32'h3b09f888),
	.w4(32'hbb06734c),
	.w5(32'h3b05a2e3),
	.w6(32'hbb23d088),
	.w7(32'h3aa274e7),
	.w8(32'h3b736023),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4c31),
	.w1(32'hbba0868e),
	.w2(32'hbb2cad36),
	.w3(32'h3b4c267c),
	.w4(32'hbad5795a),
	.w5(32'hbaa1975d),
	.w6(32'hbb908486),
	.w7(32'hbb6dc272),
	.w8(32'hba19bfd5),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0c1b),
	.w1(32'h3a083407),
	.w2(32'hbc34e369),
	.w3(32'h3b0e168f),
	.w4(32'h3bcf3eea),
	.w5(32'hbbff7646),
	.w6(32'h3ab0122f),
	.w7(32'hbc6b762e),
	.w8(32'hbc0180aa),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb623bbd),
	.w1(32'h3b0a442e),
	.w2(32'hbb7ad4ce),
	.w3(32'h390797b5),
	.w4(32'h3b1cb5af),
	.w5(32'hbb93ecd8),
	.w6(32'h39bceaf2),
	.w7(32'hbb5edb8e),
	.w8(32'hbbc49604),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2084b6),
	.w1(32'hb987b6c9),
	.w2(32'h3a366b08),
	.w3(32'hbbd44731),
	.w4(32'h39a1c827),
	.w5(32'h3b6e84ec),
	.w6(32'hba1740c7),
	.w7(32'h3a26f2eb),
	.w8(32'h3b1ac7f8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad74580),
	.w1(32'h368eb27a),
	.w2(32'hb98da1a1),
	.w3(32'h3b3bc4b1),
	.w4(32'hb6e16e78),
	.w5(32'h39115a3e),
	.w6(32'hb926ed67),
	.w7(32'hb95d3889),
	.w8(32'h3a0918dc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeba8e8),
	.w1(32'h39aca231),
	.w2(32'h3a77b1d2),
	.w3(32'h3abd5f3d),
	.w4(32'hb9e1e505),
	.w5(32'hb9094a29),
	.w6(32'h3a85bdb0),
	.w7(32'h3b07b018),
	.w8(32'h3abd57d5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d8227),
	.w1(32'hbadf46ee),
	.w2(32'h3ab06cfe),
	.w3(32'h3a0f49e7),
	.w4(32'hba824da2),
	.w5(32'h3a9472c4),
	.w6(32'hbad4041b),
	.w7(32'h3b1bd1ec),
	.w8(32'h3ba65d29),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f17db),
	.w1(32'h3aef72f7),
	.w2(32'h3ad48d07),
	.w3(32'h3b6d673e),
	.w4(32'h3b4eca71),
	.w5(32'h3ab13962),
	.w6(32'h3a58eabf),
	.w7(32'h39dbff4a),
	.w8(32'h3a132cc2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91caf51),
	.w1(32'h3aefd59e),
	.w2(32'hbb8ce0c5),
	.w3(32'h3a5be089),
	.w4(32'h3b397ca3),
	.w5(32'hbb1ccf9b),
	.w6(32'h3a1b71ca),
	.w7(32'hbbb1966b),
	.w8(32'h3b2975ca),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e824),
	.w1(32'hbaa27671),
	.w2(32'hba2fc381),
	.w3(32'hb6e592a9),
	.w4(32'hba8396e0),
	.w5(32'hb8ec35a2),
	.w6(32'hbad60e64),
	.w7(32'h3a038a4c),
	.w8(32'h3b435919),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e8c3b),
	.w1(32'hb9d92598),
	.w2(32'hba76296e),
	.w3(32'h38d53d50),
	.w4(32'hba711fac),
	.w5(32'hba3cfa37),
	.w6(32'hba9f3c6e),
	.w7(32'hbb3d2567),
	.w8(32'h3a932f1b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01acb1),
	.w1(32'h391547f0),
	.w2(32'hbb1ec19a),
	.w3(32'h3b2e4763),
	.w4(32'h3a3187d3),
	.w5(32'h3ba82ef9),
	.w6(32'h37612608),
	.w7(32'h3a1d1748),
	.w8(32'hba67a41f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4340),
	.w1(32'h3cd03bee),
	.w2(32'h39e011a2),
	.w3(32'hba49420f),
	.w4(32'h3cdddfd5),
	.w5(32'h3a1fbb90),
	.w6(32'h3cb4bb9f),
	.w7(32'hbaa9f982),
	.w8(32'hb94af0bc),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb142f98),
	.w1(32'h3ccd8bae),
	.w2(32'h3ccf52c1),
	.w3(32'h3a86b371),
	.w4(32'h3caed73e),
	.w5(32'h3cc46967),
	.w6(32'h3c879f07),
	.w7(32'h3cad4792),
	.w8(32'hbb49b428),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37222a09),
	.w1(32'h3a6e5cf6),
	.w2(32'h3abdb1c8),
	.w3(32'h3b2d7897),
	.w4(32'h3833bf8a),
	.w5(32'h39416010),
	.w6(32'h39d8bcd3),
	.w7(32'h39aab471),
	.w8(32'h3b2fac48),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dfc51),
	.w1(32'h3b5d3143),
	.w2(32'h3b3798b7),
	.w3(32'h3b38f398),
	.w4(32'h3aea7d38),
	.w5(32'h3bafc527),
	.w6(32'h3a960fc5),
	.w7(32'h3b21d49b),
	.w8(32'h3b0aa53b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10b06e),
	.w1(32'hba446203),
	.w2(32'hbb084559),
	.w3(32'h3b84c029),
	.w4(32'hbb09ffff),
	.w5(32'hbb127d63),
	.w6(32'hbae39303),
	.w7(32'hbac1293e),
	.w8(32'hbae369ab),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab711e8),
	.w1(32'h39933fb6),
	.w2(32'h3b2a100a),
	.w3(32'hbb5050a9),
	.w4(32'hba70657a),
	.w5(32'h3af9ab77),
	.w6(32'h39c3f458),
	.w7(32'h3a2b668f),
	.w8(32'h3a01acf3),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8934fd),
	.w1(32'hb7a93e18),
	.w2(32'h3a968cc5),
	.w3(32'h3aa011df),
	.w4(32'hba4aa0ea),
	.w5(32'h38cdf579),
	.w6(32'h38586f36),
	.w7(32'h3a4da626),
	.w8(32'h3a797205),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2165a),
	.w1(32'hbac66858),
	.w2(32'hb9926390),
	.w3(32'h3a7be0c6),
	.w4(32'hbb8d367e),
	.w5(32'hbb26111c),
	.w6(32'hbaf28346),
	.w7(32'hba283305),
	.w8(32'hbb29e69f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b7946),
	.w1(32'h3a0fcaa1),
	.w2(32'h3b4cc72a),
	.w3(32'hbb0544ea),
	.w4(32'h3a43b29a),
	.w5(32'h3a68fee0),
	.w6(32'h3a800ca9),
	.w7(32'h3aea31a6),
	.w8(32'h3ab823d5),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27ffcb),
	.w1(32'hbb826d98),
	.w2(32'hbafe89ed),
	.w3(32'h3a267518),
	.w4(32'hbb34faae),
	.w5(32'h399dca97),
	.w6(32'hbbd65b60),
	.w7(32'hbbaaa15e),
	.w8(32'h3906a772),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f391ca),
	.w1(32'h3a17914c),
	.w2(32'h3981ddee),
	.w3(32'hba89eb9a),
	.w4(32'hba4665b2),
	.w5(32'hb7d03b55),
	.w6(32'h3a400d07),
	.w7(32'hba09401b),
	.w8(32'h3a2b2678),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6502b),
	.w1(32'hba022ce1),
	.w2(32'h3baa4253),
	.w3(32'h3a31b9df),
	.w4(32'hba1860ba),
	.w5(32'h3b5f9eb2),
	.w6(32'h39e1af54),
	.w7(32'h3b2c4e1a),
	.w8(32'h3bb14831),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3a56c),
	.w1(32'hbc6d0dd4),
	.w2(32'hbbbd5c48),
	.w3(32'h3b63176b),
	.w4(32'hbc1d9ea2),
	.w5(32'hbbd39146),
	.w6(32'hbc84e451),
	.w7(32'hbbd4d66c),
	.w8(32'hbb8e5791),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8653ab),
	.w1(32'hb9b9b56f),
	.w2(32'h3b5d7c61),
	.w3(32'hbb783226),
	.w4(32'hbb25d097),
	.w5(32'h3a6e2cff),
	.w6(32'hb9bcda9e),
	.w7(32'h3b565f92),
	.w8(32'hba954ecd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec3eb8),
	.w1(32'h3cd86a1a),
	.w2(32'h3c85ff6c),
	.w3(32'hba635315),
	.w4(32'h3cf58765),
	.w5(32'h3cae9388),
	.w6(32'h3ccf22f1),
	.w7(32'h3c888f76),
	.w8(32'hbc0bfab4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4aacf),
	.w1(32'h3acfa87e),
	.w2(32'h3b75b3fe),
	.w3(32'h3b6ce61d),
	.w4(32'h39a43fe2),
	.w5(32'h3b1cf19c),
	.w6(32'h3a1cbab3),
	.w7(32'h3b2d55d7),
	.w8(32'h3b2dd92b),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4481ba),
	.w1(32'hbb5f5624),
	.w2(32'hbaae61e2),
	.w3(32'h3b259645),
	.w4(32'hbb8d5458),
	.w5(32'hbb7bf3e5),
	.w6(32'hbb652922),
	.w7(32'hbb1735b9),
	.w8(32'hbae4af38),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba590a5f),
	.w1(32'h3af34b56),
	.w2(32'h3b3f8f94),
	.w3(32'hbb42d80c),
	.w4(32'h3a5d3665),
	.w5(32'h3ab19fcd),
	.w6(32'h3adc36d1),
	.w7(32'h3af25e3c),
	.w8(32'h3aa831ea),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ced13),
	.w1(32'h3bc12de6),
	.w2(32'h3cc75d8a),
	.w3(32'h3b3c14e8),
	.w4(32'h3b204f05),
	.w5(32'h3cf2c0a6),
	.w6(32'h3bbdd4d9),
	.w7(32'h3cde1770),
	.w8(32'hbc8edd63),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6766),
	.w1(32'h3bd08854),
	.w2(32'h3ae71a6f),
	.w3(32'hbc07d708),
	.w4(32'h3b9abab0),
	.w5(32'h3a213309),
	.w6(32'h3ba2b59a),
	.w7(32'h3b04b487),
	.w8(32'h3b78480e),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ee65a),
	.w1(32'hbb5e5d07),
	.w2(32'hba546682),
	.w3(32'h3b47b008),
	.w4(32'hbbb2e26d),
	.w5(32'hba194adb),
	.w6(32'hbb8e3fca),
	.w7(32'hbaff59e0),
	.w8(32'hbb10d0a6),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3703ec),
	.w1(32'hba82cf6d),
	.w2(32'h3a4dc8f0),
	.w3(32'hbb2ebf4d),
	.w4(32'hbb157682),
	.w5(32'hba3c84d5),
	.w6(32'hba5a67d5),
	.w7(32'h3a2fb346),
	.w8(32'hbaacebea),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f2bdd),
	.w1(32'hbb04d5de),
	.w2(32'hbacc499f),
	.w3(32'hba341819),
	.w4(32'h38cfb0ba),
	.w5(32'hba244150),
	.w6(32'hbace6290),
	.w7(32'hbb04cece),
	.w8(32'h39b9ee04),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f31231),
	.w1(32'hbaf477eb),
	.w2(32'h3a6c3291),
	.w3(32'h3ad0ef2c),
	.w4(32'hbb5560c1),
	.w5(32'hbad5dd72),
	.w6(32'hbb101bef),
	.w7(32'hb98babcb),
	.w8(32'hbaa1d381),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8612bf9),
	.w1(32'hba7be6fb),
	.w2(32'h39d157c3),
	.w3(32'hba66a2a0),
	.w4(32'hbb923327),
	.w5(32'hbb44627f),
	.w6(32'hbab1e499),
	.w7(32'h3959e936),
	.w8(32'hba26c9bd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a9bda),
	.w1(32'h3b328526),
	.w2(32'hbaecbff8),
	.w3(32'hbb17904e),
	.w4(32'h3ae6bc63),
	.w5(32'hb9c3a4bf),
	.w6(32'h3a77c566),
	.w7(32'hbaaa4ea0),
	.w8(32'h39019e27),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf9766),
	.w1(32'hbb12f119),
	.w2(32'hbb2348ca),
	.w3(32'h38b9e8dd),
	.w4(32'hbb5669a7),
	.w5(32'hbb85836f),
	.w6(32'hba4114e1),
	.w7(32'hbb29a005),
	.w8(32'hbae77f42),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba932b9f),
	.w1(32'h3ca5cd95),
	.w2(32'h3b80f053),
	.w3(32'hbb109863),
	.w4(32'h3cbd81ec),
	.w5(32'h3befd188),
	.w6(32'h3cb26757),
	.w7(32'h3b1720e7),
	.w8(32'hbbd46d1d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8489a1),
	.w1(32'hbac812a2),
	.w2(32'hbae0b023),
	.w3(32'h3bb5ec30),
	.w4(32'hbb325ad9),
	.w5(32'hbb0a65d1),
	.w6(32'hbb82192b),
	.w7(32'hbb0c1952),
	.w8(32'h3aa04935),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b438c0a),
	.w1(32'hba93ed3c),
	.w2(32'h3b88f573),
	.w3(32'h3aa0bdfb),
	.w4(32'h3a16e49a),
	.w5(32'h3b86a833),
	.w6(32'hbb25fad5),
	.w7(32'hbabf756c),
	.w8(32'h3b0b0bc4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5d210),
	.w1(32'h3c6f002f),
	.w2(32'h3c945397),
	.w3(32'h3bad0cdd),
	.w4(32'h3c00d81a),
	.w5(32'h3c518fdc),
	.w6(32'h3b583ede),
	.w7(32'h3c162c9c),
	.w8(32'hbb79602f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50aac4),
	.w1(32'h3a492ef5),
	.w2(32'hbc13e467),
	.w3(32'hbb25f220),
	.w4(32'hba1439c1),
	.w5(32'hbc0d92a1),
	.w6(32'hbaaeb37e),
	.w7(32'hbbfe88a1),
	.w8(32'hbb5d9cfc),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc96659),
	.w1(32'hb90c5e79),
	.w2(32'h3b07a39f),
	.w3(32'hbb9b6972),
	.w4(32'hba876827),
	.w5(32'h3aba02a9),
	.w6(32'hb9fb7ac8),
	.w7(32'h3b1013fc),
	.w8(32'h3b937b95),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a9fd5),
	.w1(32'h3a0adebe),
	.w2(32'hba8b5d5f),
	.w3(32'h3b857833),
	.w4(32'hba7f5259),
	.w5(32'hbb222233),
	.w6(32'hb9e026e6),
	.w7(32'hba70f296),
	.w8(32'hbb376049),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a539f),
	.w1(32'h3a1f979e),
	.w2(32'hbc2ddaeb),
	.w3(32'hbb975aee),
	.w4(32'hba958856),
	.w5(32'hbbd81c8b),
	.w6(32'hbb33f9a3),
	.w7(32'hbc0d7280),
	.w8(32'hbaee3cae),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03aaeb),
	.w1(32'hba5a4c4c),
	.w2(32'hba21f149),
	.w3(32'hbb3aaab2),
	.w4(32'hb89ad9e4),
	.w5(32'hb9ba2e73),
	.w6(32'h3a533f3b),
	.w7(32'hba9a6460),
	.w8(32'h3afd7c90),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc159d),
	.w1(32'h3a8715f5),
	.w2(32'h39cadc3e),
	.w3(32'h3b1d2397),
	.w4(32'hba8a3bb5),
	.w5(32'h394c1ebc),
	.w6(32'h3a7c72f5),
	.w7(32'hba878f97),
	.w8(32'h3a634ca0),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a1cdd),
	.w1(32'h3872cb12),
	.w2(32'h3b05657c),
	.w3(32'h3a216a74),
	.w4(32'hba34acdf),
	.w5(32'h3a55d76a),
	.w6(32'h3a313a35),
	.w7(32'h381bf557),
	.w8(32'h3b1a4fb0),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ee540),
	.w1(32'h396cf30d),
	.w2(32'h3a0c489c),
	.w3(32'h3af72082),
	.w4(32'hba55794d),
	.w5(32'hb7325497),
	.w6(32'h39b18262),
	.w7(32'hb9a23bc6),
	.w8(32'h3a10c24b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be225c),
	.w1(32'h3a517449),
	.w2(32'hba8cee82),
	.w3(32'h399ca823),
	.w4(32'h39c56890),
	.w5(32'hba54916d),
	.w6(32'hba072cc9),
	.w7(32'hba6b8de9),
	.w8(32'hba278b4d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fc3c6),
	.w1(32'hbb0592ef),
	.w2(32'hb9529816),
	.w3(32'h374c29f0),
	.w4(32'hbb2c7f59),
	.w5(32'hb90a212c),
	.w6(32'hbb76d73f),
	.w7(32'hbae24f17),
	.w8(32'h3a653271),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4ac4),
	.w1(32'hba56817c),
	.w2(32'hb7a1fe0c),
	.w3(32'h3ad0f99f),
	.w4(32'hbbdbeb87),
	.w5(32'hbba45dbc),
	.w6(32'hbb256431),
	.w7(32'hba89c93a),
	.w8(32'hbb3ac328),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85caf5),
	.w1(32'h3a1b2e18),
	.w2(32'h383568e3),
	.w3(32'hbb86ebc7),
	.w4(32'hba072e41),
	.w5(32'h385cecfc),
	.w6(32'h3a3988d4),
	.w7(32'hba1e0be7),
	.w8(32'h3a0244f5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9df3366),
	.w1(32'h3b3dea6c),
	.w2(32'h3bd31c15),
	.w3(32'h3a027b84),
	.w4(32'h3a8db76a),
	.w5(32'h3b7e9232),
	.w6(32'h3b14ebf4),
	.w7(32'h3b47c594),
	.w8(32'h3af68b86),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4bfa2c),
	.w1(32'h3ac665ae),
	.w2(32'h3a71a5cf),
	.w3(32'h3b7ac875),
	.w4(32'hba1a2436),
	.w5(32'hba93b8ad),
	.w6(32'h396285ed),
	.w7(32'h39e26d2f),
	.w8(32'h3b036e86),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c90f0),
	.w1(32'hbb3b7990),
	.w2(32'h3b26e4d0),
	.w3(32'h3af88668),
	.w4(32'hbab7a08a),
	.w5(32'hba84bd2b),
	.w6(32'hbb2d82b4),
	.w7(32'h3af2c702),
	.w8(32'h3b51684f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a477fe4),
	.w1(32'hb8a40308),
	.w2(32'h3b280723),
	.w3(32'h3b0912dc),
	.w4(32'hba132b1e),
	.w5(32'h3a672ae9),
	.w6(32'h39989037),
	.w7(32'h3b32e640),
	.w8(32'h3b4cb210),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b740da4),
	.w1(32'hbb967c13),
	.w2(32'hbb3a8723),
	.w3(32'h3b0d6642),
	.w4(32'hbb699ad2),
	.w5(32'hbaa308e7),
	.w6(32'hbb8339b1),
	.w7(32'hbae8c9f4),
	.w8(32'h3a7b8e1d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8d811),
	.w1(32'hbb7735e8),
	.w2(32'hbc10ed4e),
	.w3(32'h3ac5bbac),
	.w4(32'hbb2e8e2c),
	.w5(32'hbbbbe52d),
	.w6(32'hbb9a00f1),
	.w7(32'hbbf98692),
	.w8(32'hbbccbfea),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08f69c),
	.w1(32'h3a34e31a),
	.w2(32'h39f176c5),
	.w3(32'hbbc88f7d),
	.w4(32'hba636682),
	.w5(32'h38c7a4f9),
	.w6(32'h3a6063ba),
	.w7(32'hba3e2d1c),
	.w8(32'h3a4bff59),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1b52a),
	.w1(32'hba58936e),
	.w2(32'h3a3739f4),
	.w3(32'h3a37fcfd),
	.w4(32'hbab3b5cb),
	.w5(32'h39667139),
	.w6(32'hb9c6d74d),
	.w7(32'h393d6cb5),
	.w8(32'h3ae39fcb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9e4d5),
	.w1(32'hbaa2905e),
	.w2(32'h3ae29fbb),
	.w3(32'h3aa42d37),
	.w4(32'hbaf4fe93),
	.w5(32'h3a17b29d),
	.w6(32'hba473a0f),
	.w7(32'h3a4d8c16),
	.w8(32'h3afec88a),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae76748),
	.w1(32'hba881787),
	.w2(32'h3ad26204),
	.w3(32'h3a9429dc),
	.w4(32'h3adc4c91),
	.w5(32'h39db5431),
	.w6(32'hbb5c3ea6),
	.w7(32'hb9d5b7fc),
	.w8(32'h399b79fa),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25c050),
	.w1(32'h3bb6d7a2),
	.w2(32'h3b89fcde),
	.w3(32'h3b35ce9e),
	.w4(32'h3baaa494),
	.w5(32'h3bdba5c9),
	.w6(32'h3b529257),
	.w7(32'h3bc9b5ca),
	.w8(32'hbac858c7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6f5a),
	.w1(32'hb9f3e8da),
	.w2(32'h3b153ac5),
	.w3(32'hba14cf22),
	.w4(32'hbb170df4),
	.w5(32'h38af3965),
	.w6(32'hbac9ba05),
	.w7(32'h39ba2a39),
	.w8(32'h3a38d6ef),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad786cd),
	.w1(32'hba1f5225),
	.w2(32'h3b04aa03),
	.w3(32'hba851f74),
	.w4(32'hba4982a8),
	.w5(32'h3a66c4dc),
	.w6(32'hbad61363),
	.w7(32'h3aec9a97),
	.w8(32'h3aebb797),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae288d0),
	.w1(32'hb90aa482),
	.w2(32'h3a8da81f),
	.w3(32'hb9ddb33f),
	.w4(32'hba15aac6),
	.w5(32'h3a431c1e),
	.w6(32'hb95b6699),
	.w7(32'h39dc0e7a),
	.w8(32'h3a9aeff0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc525f),
	.w1(32'h3a83bb89),
	.w2(32'h3bb562ad),
	.w3(32'h3abb6647),
	.w4(32'h3b1473a0),
	.w5(32'h3b8491cd),
	.w6(32'hba2161a4),
	.w7(32'h3a50a992),
	.w8(32'h3aab64eb),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d6ec5),
	.w1(32'h3a7d01bb),
	.w2(32'h3b614230),
	.w3(32'h3bf466fc),
	.w4(32'h39d20cfe),
	.w5(32'h3af87daa),
	.w6(32'h390e8fdf),
	.w7(32'h3a8dba51),
	.w8(32'h3b6569d2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88a0d7),
	.w1(32'hbaeeff28),
	.w2(32'h3b6e1c03),
	.w3(32'h3b142a2f),
	.w4(32'hbb8c9aab),
	.w5(32'h3a96e8b0),
	.w6(32'hba8d3454),
	.w7(32'h3b942b17),
	.w8(32'hba8a7da3),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9629c56),
	.w1(32'hbb374c46),
	.w2(32'hbc822564),
	.w3(32'hbaa21037),
	.w4(32'hbc44544b),
	.w5(32'hbc62a4e2),
	.w6(32'hbc3f6c9c),
	.w7(32'hbc9bd408),
	.w8(32'hbb773817),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5b1f7),
	.w1(32'h3bbd6aa7),
	.w2(32'h3ac85350),
	.w3(32'hb930b4fc),
	.w4(32'hbc31b127),
	.w5(32'hba2d174d),
	.w6(32'h3a1a8cce),
	.w7(32'hbb3b6de1),
	.w8(32'hb9c5030a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule