module layer_10_featuremap_45(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad0dc4),
	.w1(32'h3b94599f),
	.w2(32'hbc8e9cb0),
	.w3(32'hbb6b82f5),
	.w4(32'hbb143619),
	.w5(32'h3b0c59a8),
	.w6(32'hbc204702),
	.w7(32'hbc392263),
	.w8(32'h3c4f0c03),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31433f),
	.w1(32'h3a690118),
	.w2(32'h3bdb3e67),
	.w3(32'hbc52465d),
	.w4(32'hbc06407c),
	.w5(32'h3c3c7568),
	.w6(32'h3c8f2092),
	.w7(32'h3b84c127),
	.w8(32'h3bf1de55),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27a172),
	.w1(32'h3c0705ec),
	.w2(32'hbbd5db0d),
	.w3(32'h3c081267),
	.w4(32'hbab5b6b7),
	.w5(32'hbb61dd8d),
	.w6(32'hbb8b3722),
	.w7(32'hbb0affcf),
	.w8(32'hbb492bdc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4be1d7),
	.w1(32'h3bc976bc),
	.w2(32'h39c6a4be),
	.w3(32'hba505034),
	.w4(32'hbbba32b5),
	.w5(32'h3c99de61),
	.w6(32'h3a9035d6),
	.w7(32'hba8f8a7d),
	.w8(32'h390dd6f8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb502f99),
	.w1(32'hbb8bc270),
	.w2(32'hbb8b24b6),
	.w3(32'h3cef9ee4),
	.w4(32'h3c83deed),
	.w5(32'h3b4ce311),
	.w6(32'h3c90b4e5),
	.w7(32'hb8f63a89),
	.w8(32'hbb10fdba),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4cfe5),
	.w1(32'h3b96deba),
	.w2(32'hbb831310),
	.w3(32'h3a35d1d3),
	.w4(32'h3ae8671d),
	.w5(32'hbaba3ffc),
	.w6(32'h3bd5c287),
	.w7(32'h3be36bdf),
	.w8(32'hbbd3f1c3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2282b),
	.w1(32'h3aa68cd7),
	.w2(32'hbc2ec4a5),
	.w3(32'hbaf17359),
	.w4(32'h3bb3de2b),
	.w5(32'hba4d55ea),
	.w6(32'hbbd09c1c),
	.w7(32'hba5dc340),
	.w8(32'hbbfaa8f8),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2c696),
	.w1(32'hbc3251c8),
	.w2(32'h3a28912b),
	.w3(32'h3c41d484),
	.w4(32'h3c029add),
	.w5(32'h3ac4b4fb),
	.w6(32'h3a9d9e3a),
	.w7(32'h3be8d944),
	.w8(32'hbc69fe8b),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c40dbaf),
	.w1(32'h3bcdb680),
	.w2(32'h3c036c22),
	.w3(32'h3bfa06ad),
	.w4(32'hbac515ca),
	.w5(32'h3c448aa9),
	.w6(32'hbc5415f2),
	.w7(32'hbc434720),
	.w8(32'h3bfc5030),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c200cff),
	.w1(32'h3c3d0667),
	.w2(32'h3bd50711),
	.w3(32'h3b6fe5c8),
	.w4(32'h3b50070c),
	.w5(32'h3b63d36d),
	.w6(32'hbb52bfb1),
	.w7(32'hbbd4b0d1),
	.w8(32'h3b92f09e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77438),
	.w1(32'h3c2c7a21),
	.w2(32'hba1b096d),
	.w3(32'hbb8155d0),
	.w4(32'hbaf66545),
	.w5(32'hbb82af45),
	.w6(32'hbb38adee),
	.w7(32'hba99d0f8),
	.w8(32'h3a67e7d5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f8c2d),
	.w1(32'h3c09f6d0),
	.w2(32'h3a3a5322),
	.w3(32'hbae572a1),
	.w4(32'hb9d0a6fe),
	.w5(32'h3b308bc0),
	.w6(32'h39998aaa),
	.w7(32'hbafd2e75),
	.w8(32'h3aa1b935),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893ab70),
	.w1(32'h3aecfb87),
	.w2(32'h3c3d53fa),
	.w3(32'hbad90901),
	.w4(32'h3af66fe0),
	.w5(32'h3c35b177),
	.w6(32'hbb3b150e),
	.w7(32'h3a565464),
	.w8(32'h3bf03994),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a9e25),
	.w1(32'h3c263de1),
	.w2(32'hbc160a91),
	.w3(32'h3c4f6a30),
	.w4(32'h3c62d3eb),
	.w5(32'hbba6e73f),
	.w6(32'h3c2963a0),
	.w7(32'h3b8278ce),
	.w8(32'hbba98a4f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2dace),
	.w1(32'h3ba26d50),
	.w2(32'hbc585196),
	.w3(32'h3bd7aabf),
	.w4(32'h3b87bc85),
	.w5(32'hbbfb60c0),
	.w6(32'hbb9e7697),
	.w7(32'hbc30249b),
	.w8(32'h3bab2b08),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a5e1f),
	.w1(32'hbc46897e),
	.w2(32'h3be93231),
	.w3(32'hbc4fedff),
	.w4(32'hbc81134a),
	.w5(32'h3af9d2d7),
	.w6(32'h3c918601),
	.w7(32'h3c7abfef),
	.w8(32'h3b8bbcf8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc566ec),
	.w1(32'h3bcf243c),
	.w2(32'h3c14b1d2),
	.w3(32'hbb8c9323),
	.w4(32'hbb3b0dc2),
	.w5(32'hbba67184),
	.w6(32'hbb131cc3),
	.w7(32'h3b1c3657),
	.w8(32'hbce5805a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1df760),
	.w1(32'h3c8d95a0),
	.w2(32'h3c2ae301),
	.w3(32'h3bc230b5),
	.w4(32'h3cc01b0e),
	.w5(32'h3beab07d),
	.w6(32'hbd06966f),
	.w7(32'hbcbcd563),
	.w8(32'h3b23958a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0215c4),
	.w1(32'h3c2b0b3c),
	.w2(32'hbb437249),
	.w3(32'h3c66e551),
	.w4(32'h3c1e8f6a),
	.w5(32'h3b1ace23),
	.w6(32'h3adb7088),
	.w7(32'h3b5d498b),
	.w8(32'h3bc6b334),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fa71a),
	.w1(32'hbabc99dd),
	.w2(32'h3b5ec0ab),
	.w3(32'h3c010198),
	.w4(32'h3a126a08),
	.w5(32'h3b4f1258),
	.w6(32'h3bc07f30),
	.w7(32'hbb6279a7),
	.w8(32'h39921276),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82b287),
	.w1(32'h3b56ea5d),
	.w2(32'hbb211edb),
	.w3(32'h3c03044a),
	.w4(32'hbb0fc27f),
	.w5(32'h3b7b04c6),
	.w6(32'h39a91d75),
	.w7(32'hbc069b03),
	.w8(32'h39cd7086),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0b352),
	.w1(32'h3b79538c),
	.w2(32'hbbfd63f8),
	.w3(32'h3c2c5f18),
	.w4(32'hbaf49e45),
	.w5(32'h3bef324f),
	.w6(32'h3bc652c4),
	.w7(32'hbbe59ef6),
	.w8(32'hbb9b1b52),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2857eb),
	.w1(32'h3b97f34f),
	.w2(32'h3afa2548),
	.w3(32'hb95eb496),
	.w4(32'h3ba61c52),
	.w5(32'h3b88c7fa),
	.w6(32'h3b42bff6),
	.w7(32'hba9d0ed6),
	.w8(32'h3b581f41),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39359069),
	.w1(32'h3b32e47b),
	.w2(32'h3b05218c),
	.w3(32'hb9d8a780),
	.w4(32'h3b0bbc83),
	.w5(32'h3b10925d),
	.w6(32'h398b095e),
	.w7(32'h3b20ebf5),
	.w8(32'h39bba8f8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b35eb),
	.w1(32'hbbb4a248),
	.w2(32'hbc4c267e),
	.w3(32'h3c39bf20),
	.w4(32'h3a87fb59),
	.w5(32'h3bbd5c9f),
	.w6(32'h3c644a7d),
	.w7(32'h3bbeeedf),
	.w8(32'hbb9c2b3d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87c135),
	.w1(32'hbc35692c),
	.w2(32'h3b30d7fd),
	.w3(32'h3cd1493a),
	.w4(32'h3bb68840),
	.w5(32'hbc117af9),
	.w6(32'hbc09b04d),
	.w7(32'hbc478b6d),
	.w8(32'hbc0e6807),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50b6ef),
	.w1(32'hbb4a63b9),
	.w2(32'h3ad6280d),
	.w3(32'hbabb5aec),
	.w4(32'h3ada2cd9),
	.w5(32'hb93509e2),
	.w6(32'hbbed9950),
	.w7(32'h3a9f3952),
	.w8(32'h3a9936fc),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e27782),
	.w1(32'h3a69ac9a),
	.w2(32'h3b670589),
	.w3(32'hbb50d111),
	.w4(32'hba659e36),
	.w5(32'hbc1b2353),
	.w6(32'h3b7341ea),
	.w7(32'h3bb00d63),
	.w8(32'h3a1a3b52),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d407),
	.w1(32'hbb3dc524),
	.w2(32'h3bb953cd),
	.w3(32'hbc1b0d66),
	.w4(32'hbbb451e3),
	.w5(32'hbbf71cd4),
	.w6(32'h3bfba17d),
	.w7(32'h3a7ef4d7),
	.w8(32'h3b965c49),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8956),
	.w1(32'hbc25fa39),
	.w2(32'hbb1b11eb),
	.w3(32'hbc7377db),
	.w4(32'hbc817317),
	.w5(32'hb99e4670),
	.w6(32'h3bc6730a),
	.w7(32'h3c5077c3),
	.w8(32'hbc36c6cb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b3398),
	.w1(32'h3bb5bb00),
	.w2(32'h3bf5ac50),
	.w3(32'h3b770ba1),
	.w4(32'h3b6e9b75),
	.w5(32'hbbdb93cf),
	.w6(32'hbc6bf326),
	.w7(32'hbbf1224a),
	.w8(32'hbc337e68),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe39bc),
	.w1(32'hbaf98655),
	.w2(32'hbbd83d6c),
	.w3(32'hbca1c8ca),
	.w4(32'hbcdb4d82),
	.w5(32'hbc932a62),
	.w6(32'hbc9a92d9),
	.w7(32'hbc80cd5e),
	.w8(32'hbc50f97b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bd298),
	.w1(32'h3a560039),
	.w2(32'hbac6d5ea),
	.w3(32'hbc8cca27),
	.w4(32'hbc87cdc8),
	.w5(32'hbaf4f576),
	.w6(32'hbcb95614),
	.w7(32'hbc2f920d),
	.w8(32'h3ad6515e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c2577),
	.w1(32'hbbadaadf),
	.w2(32'h3bac1701),
	.w3(32'h3a968d26),
	.w4(32'h3aeab480),
	.w5(32'h3ca63c8b),
	.w6(32'h3c05c035),
	.w7(32'h3bcfb639),
	.w8(32'h3b65abae),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccac1fc),
	.w1(32'h3cfd3024),
	.w2(32'hbb103470),
	.w3(32'h3cddcb2f),
	.w4(32'h3b7a5f9f),
	.w5(32'hbb9d2c43),
	.w6(32'h3bfcbee3),
	.w7(32'h3c9020a8),
	.w8(32'h3b1b66d1),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc085a0b),
	.w1(32'hbba308e4),
	.w2(32'h3a886b7e),
	.w3(32'hbbe58214),
	.w4(32'hb98a7b3d),
	.w5(32'hbb487456),
	.w6(32'h3b78bc88),
	.w7(32'h3a9c4d3f),
	.w8(32'hbc2d05cd),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1754ff),
	.w1(32'h3ac2b807),
	.w2(32'hbb15acb9),
	.w3(32'hbc20a68c),
	.w4(32'hbc1326ca),
	.w5(32'hba52a61f),
	.w6(32'hbc28863e),
	.w7(32'h3b4b4c33),
	.w8(32'h3c1982d5),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2b58c3),
	.w1(32'hbc08a112),
	.w2(32'hbc5b4be9),
	.w3(32'h3b35e326),
	.w4(32'h3adda627),
	.w5(32'hbb9bfe3b),
	.w6(32'h3ca5c8f2),
	.w7(32'h3c2d65e0),
	.w8(32'h3c803818),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c39db),
	.w1(32'hbcb068f8),
	.w2(32'h3bac0254),
	.w3(32'hbc82f486),
	.w4(32'h3c163df4),
	.w5(32'hbc8c4bce),
	.w6(32'h3d21d45f),
	.w7(32'h3d06b5e4),
	.w8(32'hbc8c6cc1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074a85),
	.w1(32'h3c4d8496),
	.w2(32'hbb8fe720),
	.w3(32'h3b77b057),
	.w4(32'h3b081ccd),
	.w5(32'hbb696dd6),
	.w6(32'hbc24481f),
	.w7(32'hbbe9c7d0),
	.w8(32'h3ac59fca),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c60a7),
	.w1(32'h39202287),
	.w2(32'h3b0a775c),
	.w3(32'hb9723c4c),
	.w4(32'h3b6b3965),
	.w5(32'hbca59fdd),
	.w6(32'h3b4b8819),
	.w7(32'h3bfba2a5),
	.w8(32'hbb739010),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093f85),
	.w1(32'h3be0b028),
	.w2(32'hbc28e76b),
	.w3(32'hbcef262d),
	.w4(32'hbc6693c9),
	.w5(32'hbc51ea63),
	.w6(32'hbc0e4117),
	.w7(32'hbb0e9eaf),
	.w8(32'hbad1cc0e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca6481),
	.w1(32'h3991d2a9),
	.w2(32'hbb114bba),
	.w3(32'hbc96d750),
	.w4(32'hbc9596d8),
	.w5(32'hbbbbc6db),
	.w6(32'hbb8a7d14),
	.w7(32'h3b37b8b0),
	.w8(32'h3c13f118),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9049c),
	.w1(32'h39f7600b),
	.w2(32'hba2ace8f),
	.w3(32'hbb806028),
	.w4(32'h3b61848f),
	.w5(32'h3b42a5c8),
	.w6(32'h3c9a6275),
	.w7(32'h3c5fd175),
	.w8(32'h39176161),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3094ee),
	.w1(32'hb8ca9e2d),
	.w2(32'hbbdab477),
	.w3(32'h3b8e3664),
	.w4(32'hbbfda68f),
	.w5(32'hbc57d2ed),
	.w6(32'hbc020e5f),
	.w7(32'hbbfa949b),
	.w8(32'hbac90c57),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232476),
	.w1(32'hbb4d2e95),
	.w2(32'h3b85a97a),
	.w3(32'hbbd2e839),
	.w4(32'hb8755379),
	.w5(32'hbb95f522),
	.w6(32'h3b93525e),
	.w7(32'hbb21cbbd),
	.w8(32'hba56001b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b245b74),
	.w1(32'hbb393329),
	.w2(32'h3b9a832a),
	.w3(32'h39dc2a11),
	.w4(32'hbc7ec2a0),
	.w5(32'h3a46d8f3),
	.w6(32'hbb8732fd),
	.w7(32'hbb18fda7),
	.w8(32'h3a0757d6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4cb71),
	.w1(32'h3c66acd1),
	.w2(32'h392ccf7d),
	.w3(32'h3c0a4265),
	.w4(32'h3bb48217),
	.w5(32'h3a174fe3),
	.w6(32'hbc0c4526),
	.w7(32'hbbda13c2),
	.w8(32'h3c226280),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6c8b7),
	.w1(32'hbbcb1b57),
	.w2(32'hbae0c3ea),
	.w3(32'hbb889bb0),
	.w4(32'hbbab8d03),
	.w5(32'hbc5c14bc),
	.w6(32'h3c0caf40),
	.w7(32'h3b8a3a8e),
	.w8(32'h3b5582f5),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c4e78),
	.w1(32'h3be3b9e6),
	.w2(32'h3c0fc551),
	.w3(32'hbd013ded),
	.w4(32'hbc8bb7e2),
	.w5(32'h3b7201f7),
	.w6(32'h3b8b54d2),
	.w7(32'h3c19ac94),
	.w8(32'hba96e635),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085fd7),
	.w1(32'h3a64886d),
	.w2(32'hbb25db3a),
	.w3(32'hbb59e69f),
	.w4(32'h3b3a0d9e),
	.w5(32'h3b92e364),
	.w6(32'hbb887492),
	.w7(32'h3a3274ed),
	.w8(32'hbc6c5a99),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf856a4),
	.w1(32'hbc3187ed),
	.w2(32'h3a2ee071),
	.w3(32'hbbc92c03),
	.w4(32'hba01bd13),
	.w5(32'hba8d457b),
	.w6(32'hbc3e922d),
	.w7(32'hbabef01e),
	.w8(32'h3b6c204f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b092dab),
	.w1(32'h3b81a546),
	.w2(32'hbbd1d802),
	.w3(32'hbbb47f31),
	.w4(32'h3ba31759),
	.w5(32'h3b25bb14),
	.w6(32'h3a2f6d24),
	.w7(32'h3b953852),
	.w8(32'hb9dffa6b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1265bf),
	.w1(32'h3b9a3a7a),
	.w2(32'hbc042ba2),
	.w3(32'h3c3dcae8),
	.w4(32'h3c4811d3),
	.w5(32'hbbc8f87d),
	.w6(32'h3b8a500b),
	.w7(32'h3c08eab9),
	.w8(32'h3bf9d442),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b2aa2),
	.w1(32'hbc0c5db1),
	.w2(32'h3b4e8da8),
	.w3(32'hbbd502bd),
	.w4(32'h3a97a9e6),
	.w5(32'h3c78aa22),
	.w6(32'h3c15593d),
	.w7(32'h3b49eef0),
	.w8(32'h37a6d6e7),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5928a7),
	.w1(32'h3c80cb8f),
	.w2(32'hbb2b61df),
	.w3(32'h3cae1ded),
	.w4(32'h3c130978),
	.w5(32'hbbcf4d4b),
	.w6(32'hbc3fa973),
	.w7(32'hbbc0a191),
	.w8(32'hbab7fbd1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfd98a),
	.w1(32'hbb3d5205),
	.w2(32'h3b3e7552),
	.w3(32'hbc34f429),
	.w4(32'h39d6a989),
	.w5(32'hbb905d0c),
	.w6(32'hbc1247fa),
	.w7(32'hbbeadff2),
	.w8(32'hbc0ed865),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c361df1),
	.w1(32'h3c3a1d84),
	.w2(32'hba622776),
	.w3(32'hbc101a2b),
	.w4(32'hbc043b3d),
	.w5(32'hbb3e6773),
	.w6(32'hbc55f3fb),
	.w7(32'h3ab843a2),
	.w8(32'h3c022ac9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96df0ba),
	.w1(32'hbb8a3ed7),
	.w2(32'h3bcdfe73),
	.w3(32'hbb3fc26f),
	.w4(32'hbb850e4b),
	.w5(32'hbc91f06b),
	.w6(32'h3c52ec5e),
	.w7(32'h3c219a59),
	.w8(32'hbc7ab4a4),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86ef48),
	.w1(32'h3c47db76),
	.w2(32'h3c927866),
	.w3(32'hbd1a6fab),
	.w4(32'hbcc866d2),
	.w5(32'h3c1d42e8),
	.w6(32'hbc81a4e2),
	.w7(32'hbb3ba27b),
	.w8(32'hbc2caad5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfd790a),
	.w1(32'h3ca78611),
	.w2(32'h3af3ef36),
	.w3(32'h3c709e7a),
	.w4(32'h3c0cc3f3),
	.w5(32'hbb8b7e10),
	.w6(32'hbcb5ec7f),
	.w7(32'hbc70abf4),
	.w8(32'h3b9295f8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9466a97),
	.w1(32'h3b3a65e6),
	.w2(32'hbb804a45),
	.w3(32'hbb86b6fb),
	.w4(32'h38157e1c),
	.w5(32'h3b99d82a),
	.w6(32'h3c0b9282),
	.w7(32'h3c617aed),
	.w8(32'hba9986c1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2add3b),
	.w1(32'hbad93e85),
	.w2(32'h3b05821a),
	.w3(32'h3a9a711f),
	.w4(32'hb8f8b226),
	.w5(32'hbc4f5fc4),
	.w6(32'h3b4b6ab3),
	.w7(32'hbb4f9b6b),
	.w8(32'hbaaf6b5e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ceac2),
	.w1(32'h3b9636a5),
	.w2(32'h3c15a1c1),
	.w3(32'hbc831b6d),
	.w4(32'hbb7eac6c),
	.w5(32'h3b836cb5),
	.w6(32'hbb445511),
	.w7(32'h3bdf2bb5),
	.w8(32'hbc0d94f7),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31dd34),
	.w1(32'h3c61067f),
	.w2(32'h3b998730),
	.w3(32'hbb71e52b),
	.w4(32'hbc3c8c5b),
	.w5(32'h3c56965f),
	.w6(32'hbc67efc1),
	.w7(32'hbc44032a),
	.w8(32'h3b9695f5),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6cb1f),
	.w1(32'h3b8674c7),
	.w2(32'h3a26d7ce),
	.w3(32'h3c7c588c),
	.w4(32'h3c54ab05),
	.w5(32'hbba6a6ff),
	.w6(32'h3bdaf54d),
	.w7(32'h3ad01e47),
	.w8(32'h3b7d66b2),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a556d7e),
	.w1(32'h3b6b5a0c),
	.w2(32'hbb509945),
	.w3(32'h3a09550f),
	.w4(32'h3ab31093),
	.w5(32'h3abd4420),
	.w6(32'h3c68a988),
	.w7(32'h3c365fdf),
	.w8(32'h3c075522),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be954f9),
	.w1(32'h3b8f5a97),
	.w2(32'h3a82de39),
	.w3(32'hbb7737a0),
	.w4(32'h3ba72e9d),
	.w5(32'h3b23e1eb),
	.w6(32'hbc682f37),
	.w7(32'hbb32c5fb),
	.w8(32'h3ae98210),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb59e55),
	.w1(32'h3add97d0),
	.w2(32'h3ba0a816),
	.w3(32'h39590e48),
	.w4(32'h3c0fc7ff),
	.w5(32'h3aeebf9b),
	.w6(32'h3b39ec2a),
	.w7(32'h39e29dc1),
	.w8(32'hbb297d4d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc81f24),
	.w1(32'hb89bae08),
	.w2(32'hbbd2f860),
	.w3(32'h3b5ee0ef),
	.w4(32'hbb5c527a),
	.w5(32'hbc15ab9b),
	.w6(32'hba201bfb),
	.w7(32'hbb1e110d),
	.w8(32'hbbc17bae),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f697),
	.w1(32'h3c0e484c),
	.w2(32'h3b7c33b2),
	.w3(32'h3b94b9e1),
	.w4(32'h3b94afd9),
	.w5(32'h3c386dea),
	.w6(32'h39632131),
	.w7(32'hbb9f48bd),
	.w8(32'hbb5c6431),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96cbab),
	.w1(32'hbc164553),
	.w2(32'hbb32a112),
	.w3(32'h3c758c01),
	.w4(32'h3bd952da),
	.w5(32'h3b1b0d47),
	.w6(32'h3b50153a),
	.w7(32'h3b625959),
	.w8(32'h3b031546),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28091a),
	.w1(32'h3aa5c172),
	.w2(32'h3b943b17),
	.w3(32'h3b80181e),
	.w4(32'hbb2ed500),
	.w5(32'hbaf30141),
	.w6(32'hbb12135b),
	.w7(32'hbb4c4cf3),
	.w8(32'h3ae75957),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14410a),
	.w1(32'h3c062ad9),
	.w2(32'h3bcd34c5),
	.w3(32'hbc270ea2),
	.w4(32'h3987b460),
	.w5(32'h3bb6b59c),
	.w6(32'h3bbea724),
	.w7(32'h3bf3964c),
	.w8(32'h3bc4319d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a376b),
	.w1(32'h3b95e0d8),
	.w2(32'hbba89b1d),
	.w3(32'hbbd95512),
	.w4(32'h3b490eb5),
	.w5(32'hbc42cedf),
	.w6(32'hbb53a847),
	.w7(32'h3b15890f),
	.w8(32'hbb729c30),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70ab78),
	.w1(32'hb8840f42),
	.w2(32'hbae2a660),
	.w3(32'hbc60ed8d),
	.w4(32'hbc30c5f5),
	.w5(32'h3b822674),
	.w6(32'h3b25edeb),
	.w7(32'h3b7ab6de),
	.w8(32'hbbe422b2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a07d034),
	.w1(32'hbac0f624),
	.w2(32'hbaa6a87d),
	.w3(32'hbc6e984f),
	.w4(32'hbc63e3e2),
	.w5(32'hbc62ee65),
	.w6(32'hbc8d4d0e),
	.w7(32'hbba42092),
	.w8(32'hbbe7cfa0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b2b6d),
	.w1(32'hbc6ec99a),
	.w2(32'hbbd2b598),
	.w3(32'hbcdd517b),
	.w4(32'hbcc6ffe9),
	.w5(32'h3bb941f3),
	.w6(32'hbbe83c05),
	.w7(32'hbc28707d),
	.w8(32'h3bff1d21),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15f089),
	.w1(32'hbb3e8e50),
	.w2(32'h3b2d9729),
	.w3(32'hbb8fa647),
	.w4(32'hbbce3df8),
	.w5(32'hb7b29736),
	.w6(32'hbb9ebcb5),
	.w7(32'hbb26b048),
	.w8(32'h3b2ddba7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b200),
	.w1(32'h3af493f4),
	.w2(32'h3a8bd668),
	.w3(32'hbbcc911b),
	.w4(32'hb90813a1),
	.w5(32'h3b8eec05),
	.w6(32'hbb885193),
	.w7(32'h3b7ff60a),
	.w8(32'h3b8bc091),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49d711),
	.w1(32'h3af437ee),
	.w2(32'h3b2db800),
	.w3(32'h3afddf66),
	.w4(32'h3b14c6ed),
	.w5(32'hbb668c31),
	.w6(32'hb9d52e19),
	.w7(32'h3b84365d),
	.w8(32'hbc1b23bf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39405b),
	.w1(32'h3bb5a5ba),
	.w2(32'hbadf1dfa),
	.w3(32'hba9c018e),
	.w4(32'h3a565bff),
	.w5(32'h3b4bd9c2),
	.w6(32'hbc2952d8),
	.w7(32'hbba80d4c),
	.w8(32'h3a9fbc14),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55fae3),
	.w1(32'hbc2fb598),
	.w2(32'h3b145ad6),
	.w3(32'hbaecf223),
	.w4(32'h3c024460),
	.w5(32'h3c4e0d3b),
	.w6(32'h3b24944f),
	.w7(32'h3c21a891),
	.w8(32'h3a1adc21),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54366a),
	.w1(32'h3bb45673),
	.w2(32'h3bebc1e5),
	.w3(32'h3c3ee4cd),
	.w4(32'h3ab24c6a),
	.w5(32'h3adcb55b),
	.w6(32'h3cbc5139),
	.w7(32'h3be3a7c4),
	.w8(32'hb8edd197),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73682c),
	.w1(32'h3b71cbf6),
	.w2(32'h3c35f140),
	.w3(32'hbb553cd0),
	.w4(32'h3bb74e1c),
	.w5(32'hbc2d55b2),
	.w6(32'hbb19705b),
	.w7(32'h3b361879),
	.w8(32'h3baa755c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2aec5),
	.w1(32'h3c3e8142),
	.w2(32'h393ffec0),
	.w3(32'h3b456762),
	.w4(32'h3bf324f6),
	.w5(32'h3b1ff248),
	.w6(32'h3c9b1452),
	.w7(32'h3c3a6961),
	.w8(32'h3b34aebf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accb8a4),
	.w1(32'h3ba16af1),
	.w2(32'hbb9e5526),
	.w3(32'h3be90173),
	.w4(32'h3c0608e3),
	.w5(32'hbb72e4cc),
	.w6(32'h3c4318a3),
	.w7(32'h3bc66663),
	.w8(32'hbb4b780f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b074e57),
	.w1(32'h3b4fcfed),
	.w2(32'h3bf7e933),
	.w3(32'hbad29212),
	.w4(32'h39d5d0c7),
	.w5(32'h3aa3261c),
	.w6(32'hbb0ba467),
	.w7(32'h3b1cf8e8),
	.w8(32'hbc55a2c8),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc6b07),
	.w1(32'hbbbddf9a),
	.w2(32'h3b8e272d),
	.w3(32'hbc638e88),
	.w4(32'hbc2b19eb),
	.w5(32'h3c80ec8e),
	.w6(32'hbc64af90),
	.w7(32'h3a28fa3a),
	.w8(32'h3c2fa62e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cdf93),
	.w1(32'h3c772929),
	.w2(32'h3b35649f),
	.w3(32'h3d16407e),
	.w4(32'h3c8ccbea),
	.w5(32'h3c5c6b32),
	.w6(32'h3cc8f83c),
	.w7(32'h3c88c698),
	.w8(32'hbb5189cb),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2ba28b),
	.w1(32'h3a8cf478),
	.w2(32'h3bb2b627),
	.w3(32'h3cd994d1),
	.w4(32'h3ca139e3),
	.w5(32'h3b64dcb1),
	.w6(32'h3b4d7cf1),
	.w7(32'hbc70ea46),
	.w8(32'hbc45d3bc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca8bd6),
	.w1(32'h3b5450ab),
	.w2(32'h3b55c2c7),
	.w3(32'h3b31c21a),
	.w4(32'hbb1c4027),
	.w5(32'hba05ae03),
	.w6(32'hbca6bbcd),
	.w7(32'hbcb57824),
	.w8(32'h3ab9c94c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94d131),
	.w1(32'h3bdc2ad7),
	.w2(32'h3b993afc),
	.w3(32'hbb21af91),
	.w4(32'h3b438a30),
	.w5(32'hbade4665),
	.w6(32'h3a5696a9),
	.w7(32'h3c082d86),
	.w8(32'hbc595833),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c815325),
	.w1(32'h3c77a2a1),
	.w2(32'h3c13d9e9),
	.w3(32'h3aba5552),
	.w4(32'h3b073d12),
	.w5(32'h3ba2b63c),
	.w6(32'hbc862b6d),
	.w7(32'hbc0b363f),
	.w8(32'h3b158e90),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b645754),
	.w1(32'hbb2528e9),
	.w2(32'h399cdaba),
	.w3(32'h3b484f27),
	.w4(32'h3b570156),
	.w5(32'h3c01cd34),
	.w6(32'h3b9612fc),
	.w7(32'hbb31d01b),
	.w8(32'h3b8b46f4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cd9e9),
	.w1(32'hbb1c990d),
	.w2(32'hbbc5c80a),
	.w3(32'h3bb98e76),
	.w4(32'hba215feb),
	.w5(32'hbc609f30),
	.w6(32'h3a707dc2),
	.w7(32'h3c092d96),
	.w8(32'h3c62315d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc038b6e),
	.w1(32'hbbc30881),
	.w2(32'hbb3bafd4),
	.w3(32'hbc8dc529),
	.w4(32'h39b67bd5),
	.w5(32'hbb40cc25),
	.w6(32'h3cd2a76f),
	.w7(32'h3c9457c4),
	.w8(32'hbb532bd4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0aec0),
	.w1(32'h3b613328),
	.w2(32'h3c2def1f),
	.w3(32'hbb6b7eaa),
	.w4(32'h3a15cf25),
	.w5(32'hbbd9662e),
	.w6(32'hbbb0cefa),
	.w7(32'hb9082f46),
	.w8(32'hbb024894),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d0336),
	.w1(32'hbbecf310),
	.w2(32'h3ac3c196),
	.w3(32'hbc703d7f),
	.w4(32'hbcc68e3f),
	.w5(32'hb9c151e0),
	.w6(32'hbb977ee6),
	.w7(32'h3bc08291),
	.w8(32'h3bed5ccb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6015d8),
	.w1(32'h3b4f2332),
	.w2(32'h3b3230f3),
	.w3(32'hb89cd35c),
	.w4(32'h3bda1265),
	.w5(32'hbc5840d3),
	.w6(32'h3c11b3cf),
	.w7(32'hb9b3f229),
	.w8(32'hb9fc4784),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5299),
	.w1(32'hbb108a32),
	.w2(32'h3c188e52),
	.w3(32'hbd056d5f),
	.w4(32'hbc97f65a),
	.w5(32'hbc768de3),
	.w6(32'hbb87ca69),
	.w7(32'h3ae8391c),
	.w8(32'hbc2c8425),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30eb15),
	.w1(32'h3c1eed18),
	.w2(32'h3b99ccf9),
	.w3(32'hbcc1e5ae),
	.w4(32'hbcfa20ad),
	.w5(32'hbc57a2dc),
	.w6(32'h3ae81cd6),
	.w7(32'h3a7b2ea4),
	.w8(32'hbb002162),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c195c67),
	.w1(32'h3b6ca88d),
	.w2(32'h3abb3901),
	.w3(32'hbccee123),
	.w4(32'hbc84e07d),
	.w5(32'h3c6e1a05),
	.w6(32'h3a0c3456),
	.w7(32'h3bf7d5c8),
	.w8(32'h3b0fb656),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75948f),
	.w1(32'h3ad6305d),
	.w2(32'h3bcd684b),
	.w3(32'h3c515eb9),
	.w4(32'h3c67a003),
	.w5(32'h3a8b0adf),
	.w6(32'h3c093f61),
	.w7(32'h39ef8cb6),
	.w8(32'hbb8c00af),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b223e6c),
	.w1(32'hba2ecdd9),
	.w2(32'h3a6b87d3),
	.w3(32'hbb1fde2a),
	.w4(32'h3aa5bc20),
	.w5(32'hbbe7501d),
	.w6(32'hbb7ed53a),
	.w7(32'hbb96caee),
	.w8(32'hbbac627d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4fe33f),
	.w1(32'hbb890e99),
	.w2(32'h3b601678),
	.w3(32'hbc6f75aa),
	.w4(32'hbc05d21c),
	.w5(32'h3baf80c0),
	.w6(32'h39d8f295),
	.w7(32'hba79fd48),
	.w8(32'h3bb890fc),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f2af9),
	.w1(32'h3a70f86e),
	.w2(32'h3aaeaab9),
	.w3(32'h39d14d6e),
	.w4(32'h3b52b2be),
	.w5(32'hbbfed304),
	.w6(32'h3b85ac4f),
	.w7(32'h3b9d4a60),
	.w8(32'hbb80acc7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2b91d),
	.w1(32'h3ba4c2a3),
	.w2(32'hba8d2a9a),
	.w3(32'hbcd2099b),
	.w4(32'hbc8840e0),
	.w5(32'hbb1ab408),
	.w6(32'h3b4d203b),
	.w7(32'h3be52d2d),
	.w8(32'hb73f68d5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814db5),
	.w1(32'h38aed8ff),
	.w2(32'hbb9b9c42),
	.w3(32'hbb542c93),
	.w4(32'hbb3e3dec),
	.w5(32'hbc821283),
	.w6(32'hbb7083b9),
	.w7(32'hbb54aad2),
	.w8(32'hbc2a8006),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e9508),
	.w1(32'hbbe881f8),
	.w2(32'hbc0fe4a6),
	.w3(32'hbcb85f10),
	.w4(32'hbcb5c5ea),
	.w5(32'hba298aad),
	.w6(32'hbbc7ad59),
	.w7(32'h3a3258f2),
	.w8(32'hbb34b32b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd678),
	.w1(32'h3bc9914d),
	.w2(32'h3a2fe4cb),
	.w3(32'hba97e339),
	.w4(32'hbad359c8),
	.w5(32'hbb041348),
	.w6(32'h39e9d8b0),
	.w7(32'h3b8e8072),
	.w8(32'h3bf88b7e),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fce28),
	.w1(32'h3af8ef1f),
	.w2(32'h3b57eb5b),
	.w3(32'hb9da25b3),
	.w4(32'h3b87034e),
	.w5(32'hbbc85f26),
	.w6(32'h3b79c6c6),
	.w7(32'hba315aa8),
	.w8(32'hbc182e79),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345e86),
	.w1(32'h3bdf9546),
	.w2(32'h3c1d6b43),
	.w3(32'hbbda1800),
	.w4(32'h3b7ac413),
	.w5(32'hbc13a1c0),
	.w6(32'hbc7f5ddf),
	.w7(32'hbc57c60c),
	.w8(32'hbb98fc24),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca85d1e),
	.w1(32'h3c241b45),
	.w2(32'h3c8867d0),
	.w3(32'hbc8d0c8f),
	.w4(32'hbc9c90b3),
	.w5(32'h3c9d3716),
	.w6(32'hba7fe41d),
	.w7(32'h39e5737e),
	.w8(32'hbb872944),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ceb9bfb),
	.w1(32'h3c923844),
	.w2(32'hbba24aa9),
	.w3(32'h3c390976),
	.w4(32'hbca5125a),
	.w5(32'hbc4e8fe7),
	.w6(32'hbcf93f0c),
	.w7(32'hbcc7a47d),
	.w8(32'h3aa31f65),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15c766),
	.w1(32'hbb9756af),
	.w2(32'hbbba2a02),
	.w3(32'hbca4d739),
	.w4(32'hbc10cbcc),
	.w5(32'h3cbab4e2),
	.w6(32'h3a3e1087),
	.w7(32'h3c21dd20),
	.w8(32'h3af818b0),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab4c38),
	.w1(32'h3b2c5ebf),
	.w2(32'h3c0ef496),
	.w3(32'h3d21ea51),
	.w4(32'h3cfeddd5),
	.w5(32'hbc5c93ad),
	.w6(32'h3b782e35),
	.w7(32'h3b32bcc5),
	.w8(32'hbb8ccc05),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24b795),
	.w1(32'h3c23881c),
	.w2(32'hbb5fd71e),
	.w3(32'hbca9db60),
	.w4(32'hbc910cd5),
	.w5(32'hbcae5b0f),
	.w6(32'hb7c672b3),
	.w7(32'h3bb98b9b),
	.w8(32'hbaf7cb15),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f34f3),
	.w1(32'hbac475e6),
	.w2(32'h3aed43b0),
	.w3(32'hbd1256ab),
	.w4(32'hbcc2bb63),
	.w5(32'hbbbef32f),
	.w6(32'h3aae027e),
	.w7(32'h3c8b95f5),
	.w8(32'h3b1052dc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880aa1f),
	.w1(32'h3ba76b07),
	.w2(32'hbae2f405),
	.w3(32'hbcb1abba),
	.w4(32'hbc468975),
	.w5(32'h3a62e07f),
	.w6(32'hbc097fc5),
	.w7(32'hbb8ae6c9),
	.w8(32'hbb3f1f81),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b628777),
	.w1(32'hbb317722),
	.w2(32'h3a90158b),
	.w3(32'h3b62c64d),
	.w4(32'h3be48557),
	.w5(32'hba79e6e9),
	.w6(32'hbb7738fc),
	.w7(32'h392c5c85),
	.w8(32'hbad0ad86),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa127d),
	.w1(32'h3b2646f4),
	.w2(32'hbb62231b),
	.w3(32'hb9420c3d),
	.w4(32'hba4bafc8),
	.w5(32'hbb128016),
	.w6(32'hbb5b7c6e),
	.w7(32'hbb25e8d2),
	.w8(32'hbbe9e0e3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d55a8a),
	.w1(32'hba32863b),
	.w2(32'hbad67ff8),
	.w3(32'hbac394cd),
	.w4(32'hbb83925c),
	.w5(32'hbb4a3d35),
	.w6(32'hbc178ed0),
	.w7(32'hbb658a74),
	.w8(32'h3b3959ce),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd10eb2),
	.w1(32'hbc313fdc),
	.w2(32'h3a0fd326),
	.w3(32'hbc9d7114),
	.w4(32'hbcc3326a),
	.w5(32'hbc293947),
	.w6(32'h3be2b5f6),
	.w7(32'h3c0a6402),
	.w8(32'hbae6563a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cf9ee),
	.w1(32'h3bb54944),
	.w2(32'hbb173a24),
	.w3(32'hbc1ad327),
	.w4(32'hbbacd258),
	.w5(32'hbc2bf764),
	.w6(32'h39e73b12),
	.w7(32'h39cc171b),
	.w8(32'hbc22845c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacbb70),
	.w1(32'hbc13852a),
	.w2(32'h3badec20),
	.w3(32'hbcabdcaf),
	.w4(32'hbc538e7f),
	.w5(32'hbb30f141),
	.w6(32'hbc7bf71d),
	.w7(32'hbc2e0a4f),
	.w8(32'hbc0eb530),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28c317),
	.w1(32'hbb197ff4),
	.w2(32'h3b132d45),
	.w3(32'hbb3caffc),
	.w4(32'h3b817c9c),
	.w5(32'h3b2b5c7e),
	.w6(32'hbc346d51),
	.w7(32'hba5f4ed2),
	.w8(32'h3c1ccf62),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16b96a),
	.w1(32'h3bac86b9),
	.w2(32'h3cc8f2bd),
	.w3(32'h3b394fbf),
	.w4(32'hbab571bf),
	.w5(32'h3c69cf1f),
	.w6(32'hbb173db8),
	.w7(32'h3abf5e0c),
	.w8(32'hbbf35927),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c899371),
	.w1(32'h3c261440),
	.w2(32'h3b30a77c),
	.w3(32'h3c3b09a2),
	.w4(32'h3b05de16),
	.w5(32'hbc6d999e),
	.w6(32'hbc4d77b2),
	.w7(32'h3b2f53a3),
	.w8(32'hbc507f7b),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880a48a),
	.w1(32'hbb0a21cd),
	.w2(32'h3b79c272),
	.w3(32'hbc13f3f2),
	.w4(32'hbbd5a438),
	.w5(32'h3c37ef44),
	.w6(32'hbc52e21c),
	.w7(32'h3bb1e124),
	.w8(32'hbb0ae0a4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15b517),
	.w1(32'h3c44c936),
	.w2(32'hbc010e92),
	.w3(32'h3c85f739),
	.w4(32'h3ca6493a),
	.w5(32'hbba1a172),
	.w6(32'hbb84ce0b),
	.w7(32'h3b2f96b9),
	.w8(32'h3bf0e740),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e56eb),
	.w1(32'h3b62438b),
	.w2(32'h3ac2f8ae),
	.w3(32'hbc36fde3),
	.w4(32'hbb54cf74),
	.w5(32'hbbe7fc16),
	.w6(32'hbbea9a0c),
	.w7(32'hbb83c815),
	.w8(32'h3d003438),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb300afb),
	.w1(32'hbc574386),
	.w2(32'h3bc04a69),
	.w3(32'h3c1422a8),
	.w4(32'h3cdf9bab),
	.w5(32'h3b4ec9a4),
	.w6(32'h3d606cb8),
	.w7(32'h3d1efb61),
	.w8(32'h3b407dc3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1ff4),
	.w1(32'h3c13aab3),
	.w2(32'h3bc96c89),
	.w3(32'h3ba7c6e3),
	.w4(32'h3c220acf),
	.w5(32'hbaecea1b),
	.w6(32'h3b21cc6e),
	.w7(32'h3bf81033),
	.w8(32'h3a5c053c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa914c),
	.w1(32'h3c19381a),
	.w2(32'h3c1de772),
	.w3(32'hbc304976),
	.w4(32'h3b9a75e4),
	.w5(32'hbc004ad2),
	.w6(32'hbc0f8f30),
	.w7(32'h3b15f0ab),
	.w8(32'h3c4e0fa1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c209231),
	.w1(32'hbacc5fce),
	.w2(32'h3b20a7a0),
	.w3(32'hbcc44760),
	.w4(32'hbc7dec2a),
	.w5(32'h3ca7a598),
	.w6(32'h3ca9650a),
	.w7(32'h3cd77642),
	.w8(32'h3bb24641),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb76498),
	.w1(32'h3a618d1c),
	.w2(32'hbb52ad53),
	.w3(32'h3cc0bf3d),
	.w4(32'h3c89eccf),
	.w5(32'h3b653e54),
	.w6(32'h3c86a575),
	.w7(32'h3b806b82),
	.w8(32'hbb675e54),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd74790),
	.w1(32'hba848fe0),
	.w2(32'h39099521),
	.w3(32'h3c004749),
	.w4(32'h3c57f475),
	.w5(32'hb97a86d0),
	.w6(32'hba597180),
	.w7(32'hbacd2b89),
	.w8(32'hbc108148),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ee389),
	.w1(32'h3b2958e3),
	.w2(32'h3b634873),
	.w3(32'h3af0e51d),
	.w4(32'h3a3ec84e),
	.w5(32'hbb2cee98),
	.w6(32'hbc607088),
	.w7(32'hbc32aa02),
	.w8(32'hbbd4c4b7),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae01fd),
	.w1(32'h3c2af71a),
	.w2(32'h3bccf0d7),
	.w3(32'hba022c8f),
	.w4(32'h3c0912cc),
	.w5(32'h3b2ff0cb),
	.w6(32'hbc17170e),
	.w7(32'hbb26c388),
	.w8(32'hbad9de58),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02fd55),
	.w1(32'h3bd858c6),
	.w2(32'hbab8e60c),
	.w3(32'hba59fbac),
	.w4(32'h39e80160),
	.w5(32'hbb3018b4),
	.w6(32'hbbe871d9),
	.w7(32'h38fdc3b3),
	.w8(32'hbbccd6ab),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe49827),
	.w1(32'hb9c14562),
	.w2(32'h3a73bc5e),
	.w3(32'hbaab6e48),
	.w4(32'hbb2af82d),
	.w5(32'hbc4b0e4a),
	.w6(32'hba70eb77),
	.w7(32'hbbfa7dab),
	.w8(32'hbc009554),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb986992),
	.w1(32'h3b651b04),
	.w2(32'h3b8de893),
	.w3(32'hbc538929),
	.w4(32'h3b83c958),
	.w5(32'hbc60fcf3),
	.w6(32'hbb7d5cda),
	.w7(32'hbbcc5b34),
	.w8(32'hbc2cb844),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b566),
	.w1(32'h3bd39de8),
	.w2(32'h3b64a46e),
	.w3(32'hbcb95ef9),
	.w4(32'hbc6f0847),
	.w5(32'hb9695c16),
	.w6(32'hbc2ff244),
	.w7(32'hbb86397c),
	.w8(32'hbc478299),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ce86d),
	.w1(32'h3bcd0ff5),
	.w2(32'h3bbdd831),
	.w3(32'h3b056441),
	.w4(32'h393fb541),
	.w5(32'h3c0ed235),
	.w6(32'hbc70f0b1),
	.w7(32'hbc308fe6),
	.w8(32'h3b854a2b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3af39c),
	.w1(32'hba6c7103),
	.w2(32'h3a866e15),
	.w3(32'h3c1abb5e),
	.w4(32'h3c1ea175),
	.w5(32'h3b921fff),
	.w6(32'h3c11cdea),
	.w7(32'h3ba35595),
	.w8(32'hb98e1159),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77d225),
	.w1(32'hbbe6e5d1),
	.w2(32'hbbdff297),
	.w3(32'hbb22842f),
	.w4(32'h3a6bc804),
	.w5(32'hbc3aad2c),
	.w6(32'h39aead2a),
	.w7(32'hbab91581),
	.w8(32'hbbe42b34),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c4823),
	.w1(32'hba8c7ba2),
	.w2(32'hbb4e34ce),
	.w3(32'hbc038bf1),
	.w4(32'h3b98e5ee),
	.w5(32'h3c01ccfe),
	.w6(32'hbc293442),
	.w7(32'hbbfd0d01),
	.w8(32'h3ba8d26b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d0ffd),
	.w1(32'h3a541f7f),
	.w2(32'hbbd0c8bd),
	.w3(32'h3c3dd84b),
	.w4(32'h3c457863),
	.w5(32'h3bad6d91),
	.w6(32'h3bd8ddb5),
	.w7(32'h3b810459),
	.w8(32'h3abf87d0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5982e7),
	.w1(32'h3bd24c84),
	.w2(32'h3c2fc75d),
	.w3(32'h3bbd6c44),
	.w4(32'h3bb3c4cb),
	.w5(32'hbbc333ae),
	.w6(32'h396957a5),
	.w7(32'hbba4e661),
	.w8(32'h3bc08db1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c947b18),
	.w1(32'h3c01e588),
	.w2(32'hbaf9f85c),
	.w3(32'hbbfbd4c7),
	.w4(32'hba1e4e12),
	.w5(32'h3a0abc51),
	.w6(32'h3c4e32be),
	.w7(32'h3c7be24a),
	.w8(32'hbbb370f2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b281bed),
	.w1(32'h3b8a69c3),
	.w2(32'h3b5019aa),
	.w3(32'hba0bf17d),
	.w4(32'h3b0ac05a),
	.w5(32'h3abcd9e2),
	.w6(32'hbc20cc1a),
	.w7(32'h3a065e30),
	.w8(32'hb9fd5a86),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe99aa9),
	.w1(32'hbb813027),
	.w2(32'hbbe2c6d8),
	.w3(32'hbb9918da),
	.w4(32'h3a2f95b4),
	.w5(32'hbb8490a6),
	.w6(32'h3ae50424),
	.w7(32'h3a54fd80),
	.w8(32'hb8a843ee),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4fd9c),
	.w1(32'hbbbd43da),
	.w2(32'hbbe6854f),
	.w3(32'hbb692a4e),
	.w4(32'h3b76661b),
	.w5(32'hbafe94e5),
	.w6(32'h3c43fac8),
	.w7(32'h3c86414a),
	.w8(32'hbc586d7b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b27f23),
	.w1(32'hbc1bfa03),
	.w2(32'hbad397e9),
	.w3(32'hbcc2e17c),
	.w4(32'hbca5d0a4),
	.w5(32'hb90d1166),
	.w6(32'h3b9a02e6),
	.w7(32'hbb41e265),
	.w8(32'hbb09da1f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb712c54),
	.w1(32'hbb85e406),
	.w2(32'h3be54e8a),
	.w3(32'h39d1199e),
	.w4(32'hbb19c738),
	.w5(32'h3c93438c),
	.w6(32'hbb271996),
	.w7(32'hbae00c7c),
	.w8(32'h3cb28bc3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96b559),
	.w1(32'h3b9ea76a),
	.w2(32'h3b8028c0),
	.w3(32'h3cce5f30),
	.w4(32'h3bd1307c),
	.w5(32'h3b60a703),
	.w6(32'h3cd0c3ae),
	.w7(32'h3bb8d61b),
	.w8(32'h3b9b8057),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e8ad8),
	.w1(32'hbbb41028),
	.w2(32'hbd742740),
	.w3(32'h3b962be0),
	.w4(32'hb9ec4a12),
	.w5(32'hbdcfc214),
	.w6(32'hbb050790),
	.w7(32'h3be02695),
	.w8(32'hbd95c694),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83b566),
	.w1(32'h3d705099),
	.w2(32'h3c21dd7a),
	.w3(32'h3c06cc0b),
	.w4(32'h3dfdd24a),
	.w5(32'hbb813e5a),
	.w6(32'hbbf5f68b),
	.w7(32'h3d8b8e89),
	.w8(32'h394fddcd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f414a),
	.w1(32'hba16fd72),
	.w2(32'h3bb77967),
	.w3(32'hbac0a846),
	.w4(32'hbb1ce326),
	.w5(32'h3b72cc8b),
	.w6(32'h388da68a),
	.w7(32'h3b506dee),
	.w8(32'h3b14e0cc),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66f2a5),
	.w1(32'h3b02a28f),
	.w2(32'hbd8327e4),
	.w3(32'hbbae1d68),
	.w4(32'hbbcf3efa),
	.w5(32'hbde3c4d1),
	.w6(32'hbb1bd295),
	.w7(32'hbb5e19b3),
	.w8(32'hbd9ad7c1),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c0b41),
	.w1(32'h3d423472),
	.w2(32'h3c0594d4),
	.w3(32'hbb8cbf7b),
	.w4(32'h3deb1cda),
	.w5(32'h3ba890f4),
	.w6(32'hbc9cbb60),
	.w7(32'h3d612d56),
	.w8(32'h396846c5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f23ceb),
	.w1(32'h3a715af0),
	.w2(32'h3cf4b853),
	.w3(32'h3bc301b5),
	.w4(32'h3ba9c131),
	.w5(32'h3d573d4f),
	.w6(32'hbb97d670),
	.w7(32'hbb30ecad),
	.w8(32'h3d24f8b2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb872e1f5),
	.w1(32'hbcd3f270),
	.w2(32'h3aa230e8),
	.w3(32'hbb22d1dc),
	.w4(32'hbd832f8b),
	.w5(32'h3bf4273d),
	.w6(32'h3ba490c3),
	.w7(32'hbd16feac),
	.w8(32'h3c3fd3e7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd09e18),
	.w1(32'hba82df36),
	.w2(32'hbd10e722),
	.w3(32'hbb558382),
	.w4(32'h3bbd2470),
	.w5(32'hbd9d582a),
	.w6(32'hbaeab2f7),
	.w7(32'h3b0da8d8),
	.w8(32'hbd3cdd6a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e2c6f),
	.w1(32'h3d26a328),
	.w2(32'hbbbc25e6),
	.w3(32'hbb70c9f1),
	.w4(32'h3dc92676),
	.w5(32'hbbf5cb7a),
	.w6(32'hbc75e44d),
	.w7(32'h3d354861),
	.w8(32'hbaf833d8),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6af1f3),
	.w1(32'hbbfd7a75),
	.w2(32'h3aa4edde),
	.w3(32'hbaa2fa3f),
	.w4(32'hbae510c0),
	.w5(32'h3b75c525),
	.w6(32'h3ac16bac),
	.w7(32'h3b532bd9),
	.w8(32'hbb925945),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ccd59),
	.w1(32'hbab9cf80),
	.w2(32'h3a9560f8),
	.w3(32'hbbaaafda),
	.w4(32'h3a86e664),
	.w5(32'hbb5186a8),
	.w6(32'hbc10d220),
	.w7(32'hbb88b80b),
	.w8(32'hbac96c03),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaead99b),
	.w1(32'h3c0745f8),
	.w2(32'h3b2eb3e0),
	.w3(32'hbadb53ee),
	.w4(32'h3c23f29e),
	.w5(32'h3aa0789e),
	.w6(32'hbb6aa6f8),
	.w7(32'h3b2ee5e0),
	.w8(32'h3b4f248f),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb840624),
	.w1(32'hbb26d421),
	.w2(32'h3b9306a7),
	.w3(32'hbc0bcc86),
	.w4(32'hbb714fe8),
	.w5(32'h3b54c466),
	.w6(32'hbc09c4be),
	.w7(32'h3b8556ad),
	.w8(32'hbb8da750),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933af8),
	.w1(32'hbb12b18e),
	.w2(32'h3d8e5bcd),
	.w3(32'h3a67ff47),
	.w4(32'hbbd65ed5),
	.w5(32'h3de89e3d),
	.w6(32'hbba55705),
	.w7(32'hbb80b0f7),
	.w8(32'h3da2f50f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb960d13),
	.w1(32'hbd8c77b4),
	.w2(32'h3bb0f828),
	.w3(32'hbc38c2dd),
	.w4(32'hbe03d5a6),
	.w5(32'h3b68b369),
	.w6(32'h3c1e727e),
	.w7(32'hbd890461),
	.w8(32'h39e2636f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5060e8),
	.w1(32'h3b787608),
	.w2(32'hbab33e68),
	.w3(32'hbada21ea),
	.w4(32'h3b6ea980),
	.w5(32'h3bab4d6d),
	.w6(32'h3b8cc9cb),
	.w7(32'h3c1a072d),
	.w8(32'h3bdb8e83),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca0c2),
	.w1(32'hba6e1e4a),
	.w2(32'h3c0bc87d),
	.w3(32'h3ba529a9),
	.w4(32'hb9e118cb),
	.w5(32'h3bbc2054),
	.w6(32'h3bbe50e8),
	.w7(32'h3c14b771),
	.w8(32'h3be3932c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ceb0d),
	.w1(32'hbb020df4),
	.w2(32'h3bd6be8f),
	.w3(32'h3bc82a90),
	.w4(32'hbb7d882c),
	.w5(32'h3b81fe05),
	.w6(32'hb9f28e83),
	.w7(32'hbbf7bdb4),
	.w8(32'hbb1111e7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b0fb6),
	.w1(32'hbba02bf2),
	.w2(32'h3d8ec492),
	.w3(32'hbc437b74),
	.w4(32'hbbe806b0),
	.w5(32'h3dedf963),
	.w6(32'hbc82eae9),
	.w7(32'hbc1b2175),
	.w8(32'h3da7dbe5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d047ca),
	.w1(32'hbd81db42),
	.w2(32'hbbf04a1f),
	.w3(32'hbb80ee8f),
	.w4(32'hbe05fd04),
	.w5(32'hbbd605a4),
	.w6(32'h3c28d34c),
	.w7(32'hbd9627a1),
	.w8(32'h3a88fa11),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda56b9),
	.w1(32'hbbcdad56),
	.w2(32'h3ac8e12c),
	.w3(32'hbc18d80b),
	.w4(32'h3b5d8c6a),
	.w5(32'h3a6a9b3e),
	.w6(32'h3b94b814),
	.w7(32'h3baa0979),
	.w8(32'h395be2c7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b851165),
	.w1(32'h3a8242b8),
	.w2(32'h3b7fd303),
	.w3(32'h3c192790),
	.w4(32'hbadd2d22),
	.w5(32'hbb4ff8e4),
	.w6(32'hbb5946df),
	.w7(32'hba7969b2),
	.w8(32'h3b15347f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacce24),
	.w1(32'h3c3fed84),
	.w2(32'h3a23b97b),
	.w3(32'hbba3381a),
	.w4(32'h3b9d8291),
	.w5(32'h3b9cd3da),
	.w6(32'hbbd0a6fe),
	.w7(32'hba2a1877),
	.w8(32'hbb252edf),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0595ad),
	.w1(32'hbba0974a),
	.w2(32'h3b85e7f9),
	.w3(32'hba871576),
	.w4(32'h3ab53c73),
	.w5(32'h3b348fe9),
	.w6(32'hbba575fc),
	.w7(32'hbb436f21),
	.w8(32'hbb1d0238),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8cad6),
	.w1(32'hbb529f22),
	.w2(32'hbb6e608e),
	.w3(32'h38a6991a),
	.w4(32'h3a62b93d),
	.w5(32'hbb76f059),
	.w6(32'hb9dd860a),
	.w7(32'hbb1e2192),
	.w8(32'h3a101097),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15ef6b),
	.w1(32'hbb299db7),
	.w2(32'hb8d5eac3),
	.w3(32'h3c244233),
	.w4(32'h3a711d58),
	.w5(32'hbbdcd56b),
	.w6(32'h3b76b77d),
	.w7(32'h3b49e4ef),
	.w8(32'hbbc9183a),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d06b),
	.w1(32'h3bada5e3),
	.w2(32'hbb0c79d4),
	.w3(32'h3a5d2267),
	.w4(32'hb9c0d225),
	.w5(32'h3c0cd3ee),
	.w6(32'hbb927bc5),
	.w7(32'hba530b6c),
	.w8(32'hbb3f7808),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17156f),
	.w1(32'h3c005e79),
	.w2(32'h3a41e5b9),
	.w3(32'hb997500e),
	.w4(32'h3a0d2a62),
	.w5(32'h3b40392a),
	.w6(32'h3bf4aa87),
	.w7(32'h3a56597d),
	.w8(32'h3b8a7e09),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5121),
	.w1(32'hbba9a573),
	.w2(32'hba85bf06),
	.w3(32'h3a68c070),
	.w4(32'h3a7d3ade),
	.w5(32'hbb855464),
	.w6(32'hbb9bb8aa),
	.w7(32'hbbb09ae6),
	.w8(32'hba9af26c),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76ab84),
	.w1(32'h3c865f60),
	.w2(32'h3c018eee),
	.w3(32'hbc23c088),
	.w4(32'h3c943ad0),
	.w5(32'hbae00f79),
	.w6(32'hbc354f13),
	.w7(32'h3c2f850b),
	.w8(32'hbae16370),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be6ba),
	.w1(32'h3c126a0c),
	.w2(32'h3c59498b),
	.w3(32'hba74b45f),
	.w4(32'h3bd772c1),
	.w5(32'h3c7b419b),
	.w6(32'hbc0b12fc),
	.w7(32'hbace355a),
	.w8(32'h3c16b9cc),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b75e398),
	.w1(32'h3987148d),
	.w2(32'h3c029a36),
	.w3(32'h3bd8da50),
	.w4(32'h3be5c350),
	.w5(32'hba97d4ec),
	.w6(32'h3c3e9cc1),
	.w7(32'h3c1ddcf1),
	.w8(32'hbb9e4164),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10145a),
	.w1(32'hbadc44f1),
	.w2(32'h3bd28b4b),
	.w3(32'hbb818580),
	.w4(32'hbc014705),
	.w5(32'h3b29cad8),
	.w6(32'hbc0f1b9c),
	.w7(32'hbbb9975a),
	.w8(32'hba05a440),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb626),
	.w1(32'h3c08b354),
	.w2(32'hbb7725c3),
	.w3(32'h3bb807c5),
	.w4(32'h3b03adcb),
	.w5(32'hbbd9bee4),
	.w6(32'h3b254bf4),
	.w7(32'hba78e865),
	.w8(32'hbc06a1e6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82462b),
	.w1(32'hbbb2ddde),
	.w2(32'h3ba45898),
	.w3(32'hbc2beb75),
	.w4(32'hbc0921e1),
	.w5(32'h3c08836d),
	.w6(32'hbbc901d5),
	.w7(32'hbb576fe1),
	.w8(32'h3c0c54fd),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c980),
	.w1(32'h3badd9e7),
	.w2(32'h3b711831),
	.w3(32'h3b582d29),
	.w4(32'h3987b4d8),
	.w5(32'h3b93d793),
	.w6(32'h3b44aa68),
	.w7(32'hba7c3645),
	.w8(32'h3b89c578),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0167fc),
	.w1(32'h3b9e6198),
	.w2(32'h3bd47c91),
	.w3(32'h3c0cbd6a),
	.w4(32'h3bf2b3c4),
	.w5(32'h3b45c782),
	.w6(32'h3bbb6701),
	.w7(32'h3bb8c0ab),
	.w8(32'h39404cb0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecc0be),
	.w1(32'hbbf5579a),
	.w2(32'h3b5a0253),
	.w3(32'hbc148966),
	.w4(32'hbbc79e20),
	.w5(32'h3bbe548b),
	.w6(32'hbc18f5a8),
	.w7(32'hbba7c047),
	.w8(32'hb986d127),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43fe9e),
	.w1(32'hbb9ca282),
	.w2(32'hbaa3887b),
	.w3(32'hbbeb308e),
	.w4(32'hbae6f5f9),
	.w5(32'hbb99e4b6),
	.w6(32'hbbe25781),
	.w7(32'hbc00b274),
	.w8(32'h3afe3118),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba802de),
	.w1(32'h3b17e1c4),
	.w2(32'hbb53da0e),
	.w3(32'hbb42f1ff),
	.w4(32'hbba0975c),
	.w5(32'hbbb6708d),
	.w6(32'h3bb75d26),
	.w7(32'h3900780c),
	.w8(32'h3a0d5256),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f480c),
	.w1(32'hbad88b6d),
	.w2(32'hbae94bf1),
	.w3(32'h3a807621),
	.w4(32'hbb1ebb66),
	.w5(32'hbc3e889a),
	.w6(32'h3b9b32d4),
	.w7(32'h3a846476),
	.w8(32'hbbbdc86a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e64a4),
	.w1(32'h3c097d0b),
	.w2(32'hbb9d9e65),
	.w3(32'hbc6ec380),
	.w4(32'h3b8b0f78),
	.w5(32'hb998b5d7),
	.w6(32'hbbd43d22),
	.w7(32'hbab7863f),
	.w8(32'h3a0fe8b3),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2e7f),
	.w1(32'hb95e0137),
	.w2(32'h3b998cc8),
	.w3(32'hbc042fdf),
	.w4(32'hbb3fa53e),
	.w5(32'h3bc9233a),
	.w6(32'hbc010d2f),
	.w7(32'hbb8ee051),
	.w8(32'h3b7d61b2),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22f2dc),
	.w1(32'hbaf61455),
	.w2(32'h3bce2d20),
	.w3(32'hbbb6f6d8),
	.w4(32'hbb1907f8),
	.w5(32'h3c7a1869),
	.w6(32'h3a57b414),
	.w7(32'hbb80621f),
	.w8(32'h3c33b95d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35005c),
	.w1(32'h3b9acf18),
	.w2(32'h3d3c1647),
	.w3(32'h3c0df36e),
	.w4(32'h3c066cc3),
	.w5(32'h3da61d92),
	.w6(32'h3bd46288),
	.w7(32'h3c02ed9a),
	.w8(32'h3d747f68),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb562c83),
	.w1(32'hbd507ff1),
	.w2(32'h3bc88e95),
	.w3(32'hbb15cc88),
	.w4(32'hbdbaceac),
	.w5(32'h3b88a3ea),
	.w6(32'h3c2f97a7),
	.w7(32'hbd50565a),
	.w8(32'h3c1dd31d),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dfd26),
	.w1(32'hb9963e79),
	.w2(32'h3b8343ba),
	.w3(32'h3b24156d),
	.w4(32'hba3df8cd),
	.w5(32'h397ab9b2),
	.w6(32'h3bc2fdd4),
	.w7(32'h3b7221f6),
	.w8(32'hbb6a9b46),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d3051),
	.w1(32'h3bdc457f),
	.w2(32'hb98f1cf8),
	.w3(32'h3b5df06e),
	.w4(32'hbad3f8c2),
	.w5(32'h3baa1966),
	.w6(32'h3a2899ef),
	.w7(32'hbb942299),
	.w8(32'h3a402624),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21dc8),
	.w1(32'h3b1d7ec1),
	.w2(32'h3b809a54),
	.w3(32'hbb87df43),
	.w4(32'hbb7cddc4),
	.w5(32'h3c3de094),
	.w6(32'hbbbc66fa),
	.w7(32'hbc0d9770),
	.w8(32'h3c328ede),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb70890),
	.w1(32'hbc0a7794),
	.w2(32'hbb8fc6a1),
	.w3(32'h3b992ef8),
	.w4(32'hbbdcfe98),
	.w5(32'hbc46a541),
	.w6(32'hbaaed472),
	.w7(32'h3afcc608),
	.w8(32'hbb83ed71),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b8a0),
	.w1(32'hba4bdf9a),
	.w2(32'h3aef68d6),
	.w3(32'h3b916b14),
	.w4(32'hbb7b5975),
	.w5(32'h3a05588c),
	.w6(32'h3c0ad962),
	.w7(32'hbab939d5),
	.w8(32'hb92c15fd),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb18c2a),
	.w1(32'h3b9c05c2),
	.w2(32'hbc87e72c),
	.w3(32'hbc7686ac),
	.w4(32'h3a4c1472),
	.w5(32'hbd145931),
	.w6(32'hbc299ef0),
	.w7(32'h3a7f2183),
	.w8(32'hbcac4193),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63acdb),
	.w1(32'h3cbe662e),
	.w2(32'hbb99835d),
	.w3(32'h3bd3b424),
	.w4(32'h3d7e5e69),
	.w5(32'hba988c93),
	.w6(32'hbb1092c2),
	.w7(32'h3d017248),
	.w8(32'hbb48382a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc145961),
	.w1(32'hbb61fedb),
	.w2(32'h3c0e6c51),
	.w3(32'hbc16a107),
	.w4(32'hbb27fba7),
	.w5(32'h3c193a31),
	.w6(32'hbb191497),
	.w7(32'hbc312cc5),
	.w8(32'h3ac92729),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f10d9),
	.w1(32'h3a53a6f5),
	.w2(32'h3b82f7b6),
	.w3(32'hba038ba1),
	.w4(32'h3aa9533f),
	.w5(32'h3bfbed6f),
	.w6(32'hbb7bdf41),
	.w7(32'hbbeb9d56),
	.w8(32'h3a86e1e9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9741a9),
	.w1(32'hba7631ba),
	.w2(32'hbbc47104),
	.w3(32'h3c0c1005),
	.w4(32'h3aaf1b7f),
	.w5(32'hbbb19f0f),
	.w6(32'hba0117e0),
	.w7(32'hbbf976b1),
	.w8(32'hbbd89725),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10c360),
	.w1(32'hbbac8576),
	.w2(32'h3b4e50ea),
	.w3(32'hbc5ae5a1),
	.w4(32'hbc4206ab),
	.w5(32'h3bb68e02),
	.w6(32'hbc8c35ae),
	.w7(32'hbbbd8d25),
	.w8(32'h3bd19e7a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb5510),
	.w1(32'h3bec3069),
	.w2(32'hbad33093),
	.w3(32'hbc39eae0),
	.w4(32'h3bd88588),
	.w5(32'h3ab707cf),
	.w6(32'hbbbaf7f7),
	.w7(32'h3bb964b3),
	.w8(32'h3bd69d95),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69c3f8),
	.w1(32'hbb2957d1),
	.w2(32'h39d093af),
	.w3(32'h3b0dcd29),
	.w4(32'hbbbde146),
	.w5(32'h3baa91ba),
	.w6(32'hba5e3686),
	.w7(32'hbbf6d3f2),
	.w8(32'hb83c950e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad21a7c),
	.w1(32'h3b251c11),
	.w2(32'h3acb4e13),
	.w3(32'h3b45fa30),
	.w4(32'h3b585899),
	.w5(32'hbb2c79eb),
	.w6(32'hbb9f1591),
	.w7(32'hbb828603),
	.w8(32'hbae40329),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c28bf),
	.w1(32'hbb9b908b),
	.w2(32'h3c8d9298),
	.w3(32'hbc20f692),
	.w4(32'h3c067a21),
	.w5(32'h3c257c8b),
	.w6(32'hbc02268c),
	.w7(32'hbbdb6c3f),
	.w8(32'hbc339638),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b8df1),
	.w1(32'hbbd5b115),
	.w2(32'h3c6c334b),
	.w3(32'hbba0d47e),
	.w4(32'hbc288285),
	.w5(32'h3c78ddd7),
	.w6(32'hbc23ad62),
	.w7(32'hbabfab75),
	.w8(32'h3c3a7d9c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8857e1),
	.w1(32'h3b98caca),
	.w2(32'hbaa805a5),
	.w3(32'hbb36ede6),
	.w4(32'hbbb47b1a),
	.w5(32'hbc03642d),
	.w6(32'hbb862202),
	.w7(32'hbb9ae166),
	.w8(32'hbb8b7791),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf738fd),
	.w1(32'h3b61104c),
	.w2(32'h3b275d88),
	.w3(32'hbb2f9b36),
	.w4(32'h3b2ab70f),
	.w5(32'h3c85d042),
	.w6(32'h3a89e556),
	.w7(32'h3b5f9928),
	.w8(32'h3c213c30),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf81792),
	.w1(32'hbc8c299e),
	.w2(32'hbc0723e0),
	.w3(32'hbb6f7ac7),
	.w4(32'hbcd52b5f),
	.w5(32'hbb8dcdb3),
	.w6(32'h3b2944d5),
	.w7(32'hbc425f54),
	.w8(32'hbafde822),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3b17a),
	.w1(32'hbacb76d3),
	.w2(32'h3bdfe631),
	.w3(32'hb985bb6c),
	.w4(32'h3ac5071a),
	.w5(32'h3c0e5ae3),
	.w6(32'hbb150aae),
	.w7(32'hbb351cbd),
	.w8(32'h3c09c683),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8242b1),
	.w1(32'h3baf6aef),
	.w2(32'hbbeb4d01),
	.w3(32'hbbad7e21),
	.w4(32'hbad20c6a),
	.w5(32'h3b43ee34),
	.w6(32'h3c0bfedf),
	.w7(32'h3c352ca0),
	.w8(32'h3b5417a7),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba72b87),
	.w1(32'h3b1059a8),
	.w2(32'hbae265f2),
	.w3(32'hbbd059c5),
	.w4(32'h3b6ed6bc),
	.w5(32'h3b4d2b3e),
	.w6(32'hbb0ef1f9),
	.w7(32'h3b7a35ef),
	.w8(32'hbb39d7d0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e50ab),
	.w1(32'hbb5a7593),
	.w2(32'h3bbd28f3),
	.w3(32'hbb0dfc93),
	.w4(32'h3b643d74),
	.w5(32'h3b17e99e),
	.w6(32'hbb07f304),
	.w7(32'hbb974d38),
	.w8(32'h3b26e939),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c034ce1),
	.w1(32'h3b675f0f),
	.w2(32'h3840f69a),
	.w3(32'h3c36bb1b),
	.w4(32'hbb605791),
	.w5(32'hbc1560e8),
	.w6(32'hbb558a2f),
	.w7(32'hbc0cdad3),
	.w8(32'hbb7755a9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd29534f),
	.w1(32'hbc76568b),
	.w2(32'h3b4005ff),
	.w3(32'hbd5985c7),
	.w4(32'hbc9e6247),
	.w5(32'h3aee235f),
	.w6(32'hbd22bafe),
	.w7(32'hbc4857f6),
	.w8(32'h3c1044ce),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf64d58),
	.w1(32'hbb73b8ce),
	.w2(32'h3c433755),
	.w3(32'hbabe9dad),
	.w4(32'hbb73a63f),
	.w5(32'hbb115ab7),
	.w6(32'hbb929b20),
	.w7(32'h3aa266d9),
	.w8(32'h3b4529b2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafba61),
	.w1(32'h3b8bf29b),
	.w2(32'h3b3b9cd9),
	.w3(32'hbb18a964),
	.w4(32'hbb285dd4),
	.w5(32'h3c08c8d0),
	.w6(32'hbb808651),
	.w7(32'hba98e299),
	.w8(32'h3ac0e828),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26d3e5),
	.w1(32'h3b9ff6f9),
	.w2(32'hbb0dd687),
	.w3(32'hbc3f0d2b),
	.w4(32'hbb31cadc),
	.w5(32'hbc278ebc),
	.w6(32'hbc6b4692),
	.w7(32'hbbe8a9ec),
	.w8(32'hbc955b39),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bb444),
	.w1(32'hbb90d66c),
	.w2(32'h3bcd518c),
	.w3(32'hbcf3c9dc),
	.w4(32'hbc61796e),
	.w5(32'hbae7b224),
	.w6(32'hbca10c82),
	.w7(32'hbbcf2485),
	.w8(32'hbb52cbd3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c8fff),
	.w1(32'hbae34fd9),
	.w2(32'hbb557ddb),
	.w3(32'h3b91e10f),
	.w4(32'hbc4c65d9),
	.w5(32'h3a0c0741),
	.w6(32'hbbcfa51c),
	.w7(32'hbc4ecf5d),
	.w8(32'hbb77ad30),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb904c),
	.w1(32'hbb3e6ae3),
	.w2(32'h3b527e73),
	.w3(32'hbc6c6d64),
	.w4(32'hb96b94a9),
	.w5(32'h3b49f473),
	.w6(32'hbc1cb5c8),
	.w7(32'hbbec76a2),
	.w8(32'h39f225f1),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b404bd1),
	.w1(32'h3b413795),
	.w2(32'hbbc545fe),
	.w3(32'hbb6df58e),
	.w4(32'h3b57dfad),
	.w5(32'hbbc25176),
	.w6(32'h39f95b5c),
	.w7(32'h3a5fedcf),
	.w8(32'h3c30ac4e),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdab690),
	.w1(32'hbb880129),
	.w2(32'h3a825ac4),
	.w3(32'hbcaaf892),
	.w4(32'hbba8b21d),
	.w5(32'h3ae739a5),
	.w6(32'hbbb9fbaf),
	.w7(32'hbbe0c8b3),
	.w8(32'h3baa4a48),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcd310),
	.w1(32'hbb44e627),
	.w2(32'hba71ca5b),
	.w3(32'h3a05563e),
	.w4(32'hba83fbcd),
	.w5(32'hba2d5b83),
	.w6(32'hbb659463),
	.w7(32'hbb52d3bf),
	.w8(32'h3a8669e4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb715cd3),
	.w1(32'hbc10362d),
	.w2(32'h3b75b096),
	.w3(32'hbab02491),
	.w4(32'h3a10c222),
	.w5(32'h3b83be9c),
	.w6(32'hbbd448da),
	.w7(32'h3b7b9fb6),
	.w8(32'hba130b32),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a831b26),
	.w1(32'h3a3fc56a),
	.w2(32'h3b27719c),
	.w3(32'h3ba39b9d),
	.w4(32'h3b6552ee),
	.w5(32'h3c355918),
	.w6(32'hbba5d912),
	.w7(32'hbbbf47ce),
	.w8(32'h3b78d4d1),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde256d),
	.w1(32'h3ad04d5b),
	.w2(32'h3b65ba6b),
	.w3(32'h3bdf8b3b),
	.w4(32'h3c4426ab),
	.w5(32'h39a58c59),
	.w6(32'h3a908d84),
	.w7(32'h3b412339),
	.w8(32'hbbb5fe2a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf62b1e),
	.w1(32'h3b7a3092),
	.w2(32'h3c251bc2),
	.w3(32'hbb9c2f5c),
	.w4(32'h3b96101b),
	.w5(32'h3bb32ee3),
	.w6(32'hbb2e2912),
	.w7(32'hbb5a1438),
	.w8(32'h3bd702b1),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb35c1e),
	.w1(32'h3b458fd0),
	.w2(32'h3b9a51ee),
	.w3(32'hbbbc62cf),
	.w4(32'hbb5ca973),
	.w5(32'h3bd138e7),
	.w6(32'hbb7fed63),
	.w7(32'hbbc5f32e),
	.w8(32'h3b80c729),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f4ac),
	.w1(32'h3b01e7ef),
	.w2(32'hbbe00878),
	.w3(32'h3bdd84c5),
	.w4(32'h3ab1e976),
	.w5(32'hbbaa5260),
	.w6(32'hbb2adf28),
	.w7(32'hbb58330c),
	.w8(32'h3b944f79),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf60aa),
	.w1(32'hbb360291),
	.w2(32'h3b8d3a5a),
	.w3(32'hbb95bf0e),
	.w4(32'h3b2ed0b0),
	.w5(32'h3aadc3b7),
	.w6(32'h3b070e1d),
	.w7(32'h39132105),
	.w8(32'h3c51505f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3adcf),
	.w1(32'h3b81f210),
	.w2(32'h3a49522c),
	.w3(32'h3b3344ee),
	.w4(32'h3c17e0a2),
	.w5(32'h3a8d8751),
	.w6(32'h3c0970eb),
	.w7(32'h3c39e05d),
	.w8(32'h3c12b9e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6acca8),
	.w1(32'hbb1e348f),
	.w2(32'h3af097dc),
	.w3(32'h3a9a682e),
	.w4(32'hbb312c0a),
	.w5(32'h3b77a54d),
	.w6(32'h3bbdd60c),
	.w7(32'hbb36cc9d),
	.w8(32'h3c066d89),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09ba44),
	.w1(32'h3a9203a2),
	.w2(32'h3c002be1),
	.w3(32'hbb931b3e),
	.w4(32'h3ba8d3e7),
	.w5(32'h3bac349d),
	.w6(32'hbc02abed),
	.w7(32'hbba17707),
	.w8(32'h3ba30fce),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301635),
	.w1(32'h3bda0cab),
	.w2(32'h3bf01431),
	.w3(32'hbb6d80d8),
	.w4(32'hbbc6f5b6),
	.w5(32'h3b357bd6),
	.w6(32'h3a57decb),
	.w7(32'hbaa05707),
	.w8(32'hba8dad0d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b092736),
	.w1(32'h3b0e7976),
	.w2(32'hbc3c51ca),
	.w3(32'h3c04fac1),
	.w4(32'h3c17d940),
	.w5(32'hbcb4f1ee),
	.w6(32'h3c21b433),
	.w7(32'h3c028798),
	.w8(32'hbc424823),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1cfd4),
	.w1(32'h3cb7eb87),
	.w2(32'hbca31372),
	.w3(32'h3c3b09b3),
	.w4(32'h3d0fc3ec),
	.w5(32'hbd1fa342),
	.w6(32'h3c06de3f),
	.w7(32'h3cdc2f61),
	.w8(32'hbcb3876f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc32f5a),
	.w1(32'h3cfe2bb3),
	.w2(32'h3c2eabca),
	.w3(32'h3c45d7ee),
	.w4(32'h3d7bfb3d),
	.w5(32'h3c77f313),
	.w6(32'h3b837ee5),
	.w7(32'h3d17be1c),
	.w8(32'h3c22aa8c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf95b2d),
	.w1(32'hbc7c21ab),
	.w2(32'h3b326882),
	.w3(32'hbc813e3a),
	.w4(32'hbc4a9943),
	.w5(32'h3b2eee9b),
	.w6(32'hbc3152ce),
	.w7(32'hbcb3ea5c),
	.w8(32'h3bf8c210),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd975d9),
	.w1(32'h3be3579d),
	.w2(32'h3c34764d),
	.w3(32'h3bc85b4b),
	.w4(32'h3bbf7ea3),
	.w5(32'h3c3d4a34),
	.w6(32'h3bdb6e15),
	.w7(32'h3b1b9980),
	.w8(32'h3b72d998),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c054cde),
	.w1(32'h3bf2547a),
	.w2(32'h3bd67dfb),
	.w3(32'h3c13a6ca),
	.w4(32'h3b93e087),
	.w5(32'h3bb1a187),
	.w6(32'hbb56e1a1),
	.w7(32'h3a706bda),
	.w8(32'h3c030c58),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accd044),
	.w1(32'hbac22be5),
	.w2(32'h3c1524e5),
	.w3(32'h3b40956a),
	.w4(32'h3a6c6157),
	.w5(32'h3c07d56c),
	.w6(32'h3b0fd702),
	.w7(32'hbb153d79),
	.w8(32'h3c1f611e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb908311),
	.w1(32'hbbf89263),
	.w2(32'hbb90ac08),
	.w3(32'hbbda2a7b),
	.w4(32'h3a779b48),
	.w5(32'hbb833ad8),
	.w6(32'hbc145896),
	.w7(32'hbb9204ac),
	.w8(32'hbbd470a8),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule