module layer_10_featuremap_154(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37084ab1),
	.w1(32'h3a41688e),
	.w2(32'hba15c478),
	.w3(32'h39a4ed24),
	.w4(32'h3a6b5765),
	.w5(32'h38f32a74),
	.w6(32'h3aa61d46),
	.w7(32'h3a71115d),
	.w8(32'h3a74b2ad),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a215ccd),
	.w1(32'h3986d542),
	.w2(32'h3aa55e05),
	.w3(32'h3a5c93ea),
	.w4(32'h3930aedb),
	.w5(32'h3a9f2b32),
	.w6(32'hba0d0eed),
	.w7(32'h3a56f07a),
	.w8(32'h3a00fed0),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a8718d),
	.w1(32'h38c65da4),
	.w2(32'h39745085),
	.w3(32'h39192dba),
	.w4(32'hba93b4a6),
	.w5(32'hba010e3e),
	.w6(32'hba8e2bee),
	.w7(32'hb995bdbe),
	.w8(32'hb8a935fe),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cbc938),
	.w1(32'hbacbc81b),
	.w2(32'hbb679875),
	.w3(32'hba016c9c),
	.w4(32'hba8f3eaf),
	.w5(32'hbb336c57),
	.w6(32'h3941c7cc),
	.w7(32'hb9a3bdd9),
	.w8(32'hba2c7b97),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc9bd9),
	.w1(32'h3a89d32c),
	.w2(32'hb906502a),
	.w3(32'hbac8d778),
	.w4(32'h3b16a26d),
	.w5(32'h3a0297cd),
	.w6(32'h3a9b18dc),
	.w7(32'hb998860e),
	.w8(32'h3a73826a),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa27ef3),
	.w1(32'h379bd893),
	.w2(32'h396232c6),
	.w3(32'h3a53268c),
	.w4(32'h3a2ed2f9),
	.w5(32'h3a85bdea),
	.w6(32'h39509465),
	.w7(32'hb9d58a7d),
	.w8(32'hba308c0d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8120c41),
	.w1(32'hba04ea82),
	.w2(32'hb9549ddf),
	.w3(32'h39adedf9),
	.w4(32'hb8ba9fc5),
	.w5(32'hb9e34b8d),
	.w6(32'hba5dd651),
	.w7(32'hb995a437),
	.w8(32'hb981b131),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9becb25),
	.w1(32'hba355535),
	.w2(32'hbaaa7041),
	.w3(32'h38c978b6),
	.w4(32'h393c4281),
	.w5(32'h36f4f867),
	.w6(32'h3a9cc2d2),
	.w7(32'hb9d42154),
	.w8(32'hba8d61c6),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a927d3),
	.w1(32'hb98cef78),
	.w2(32'hba5415a0),
	.w3(32'h397deb8f),
	.w4(32'h39c26971),
	.w5(32'hb9662d40),
	.w6(32'h39a8f6e7),
	.w7(32'hb9c5f6c2),
	.w8(32'hb98291a1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90547e1),
	.w1(32'hb9a48679),
	.w2(32'h3a60cd6d),
	.w3(32'h39771329),
	.w4(32'h38e27cbd),
	.w5(32'h3ad43042),
	.w6(32'hba96bef0),
	.w7(32'h3886672b),
	.w8(32'hba6b0b59),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9718c8c),
	.w1(32'h3af9d67d),
	.w2(32'h3ad98853),
	.w3(32'h389eec32),
	.w4(32'hb8e29edc),
	.w5(32'h39df671c),
	.w6(32'h3a1294ec),
	.w7(32'h3a3db269),
	.w8(32'h39ed675d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a968e),
	.w1(32'h3923d9bc),
	.w2(32'h390ccb99),
	.w3(32'h3a7ef663),
	.w4(32'h398302d3),
	.w5(32'h38ba724f),
	.w6(32'h3a4d2bb7),
	.w7(32'hb9858424),
	.w8(32'hba38e43c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b6d9b),
	.w1(32'hb9892c20),
	.w2(32'hb9fdcb61),
	.w3(32'h3a6ad32e),
	.w4(32'h38aa751c),
	.w5(32'h386eb2b4),
	.w6(32'h39aaaa63),
	.w7(32'hb9c66271),
	.w8(32'h37d182a2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a85305),
	.w1(32'h39c31474),
	.w2(32'hb9b6e5c9),
	.w3(32'hb99427a9),
	.w4(32'h3aa4d603),
	.w5(32'h3a817c2b),
	.w6(32'h3a6486f2),
	.w7(32'hb9cdc3d3),
	.w8(32'hb95763c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5baa9db),
	.w1(32'h3a84faa4),
	.w2(32'h3aa4ae7f),
	.w3(32'h39983d6b),
	.w4(32'h3af9378a),
	.w5(32'h3a1b5ff5),
	.w6(32'h3adb0454),
	.w7(32'h3aa6173a),
	.w8(32'h3b502837),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ff465),
	.w1(32'hb957137e),
	.w2(32'hb992f5bf),
	.w3(32'h3acc3e65),
	.w4(32'h39abe225),
	.w5(32'h39579e29),
	.w6(32'h3a17c7c5),
	.w7(32'h387855dc),
	.w8(32'h39aa5493),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c8683),
	.w1(32'h39d5bfd0),
	.w2(32'h3b35d0fb),
	.w3(32'h39acf599),
	.w4(32'hbad410fb),
	.w5(32'h3ae21435),
	.w6(32'hbb30a6ea),
	.w7(32'h3a8a5f00),
	.w8(32'hbb3511da),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93451e),
	.w1(32'hbae28b26),
	.w2(32'hb9bc7173),
	.w3(32'hbb6cd9e4),
	.w4(32'hbb237c5c),
	.w5(32'hbab402aa),
	.w6(32'hba85103c),
	.w7(32'hba25a0a4),
	.w8(32'hbb0e7b8f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9b70),
	.w1(32'hba500e7e),
	.w2(32'hb993acce),
	.w3(32'hbaa02551),
	.w4(32'hba8352b9),
	.w5(32'hba4aa6ef),
	.w6(32'hb9cb09d6),
	.w7(32'hb8660af8),
	.w8(32'hb9ec2534),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a36d7),
	.w1(32'hb9b2f4ea),
	.w2(32'hba67a8de),
	.w3(32'h390e1218),
	.w4(32'h39520bd4),
	.w5(32'hb99dee88),
	.w6(32'h38be6ccd),
	.w7(32'hba224e5c),
	.w8(32'hba232662),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba01a122),
	.w1(32'h39fac2a7),
	.w2(32'hbab17f0b),
	.w3(32'hb817f218),
	.w4(32'h3a82c4f8),
	.w5(32'hb99af21b),
	.w6(32'h3b3216c4),
	.w7(32'h3a2994ca),
	.w8(32'hb881b0fa),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53ce47),
	.w1(32'hb9165f9a),
	.w2(32'h398255f8),
	.w3(32'hba687f2c),
	.w4(32'hba15bab6),
	.w5(32'hb96270ea),
	.w6(32'hba80dc1a),
	.w7(32'hba21ccae),
	.w8(32'hb997177f),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6940e),
	.w1(32'h3c07376e),
	.w2(32'h3be7633d),
	.w3(32'hbb43f444),
	.w4(32'h3b252152),
	.w5(32'h3b468c33),
	.w6(32'h3c0c7a29),
	.w7(32'h3bd144ac),
	.w8(32'hba391651),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d9d5e),
	.w1(32'hba15c613),
	.w2(32'hbaaaa6bb),
	.w3(32'hbafa7be7),
	.w4(32'h3a3a82e5),
	.w5(32'h3957686c),
	.w6(32'h3a510032),
	.w7(32'hba1e8d49),
	.w8(32'h39f71c45),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7cb81),
	.w1(32'h3a85a1e2),
	.w2(32'h3a3272a7),
	.w3(32'h39f5c10c),
	.w4(32'h3ad01426),
	.w5(32'h3af5a1b4),
	.w6(32'h3b08c332),
	.w7(32'h3ae86fb0),
	.w8(32'h3a0d478e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65d56b),
	.w1(32'hba44f470),
	.w2(32'h39aacaaf),
	.w3(32'hb93cdb31),
	.w4(32'hbabe8467),
	.w5(32'hba0bbbd0),
	.w6(32'hbb843dda),
	.w7(32'hbb670b8f),
	.w8(32'hbb58eba8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ddb96),
	.w1(32'hba037228),
	.w2(32'hbad1480c),
	.w3(32'hbafc1ccc),
	.w4(32'h38b658a5),
	.w5(32'hba6c8eeb),
	.w6(32'h39afca18),
	.w7(32'hba7c328c),
	.w8(32'hba3190f9),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4430a0),
	.w1(32'hb9f63afb),
	.w2(32'hba9afdca),
	.w3(32'hba3477b3),
	.w4(32'h37f6b678),
	.w5(32'hb9dd4598),
	.w6(32'hba1cf50e),
	.w7(32'hba04b309),
	.w8(32'hb93c2ca9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83ce7f),
	.w1(32'h3b832fde),
	.w2(32'h3b833ad7),
	.w3(32'h392929a3),
	.w4(32'h3b434c46),
	.w5(32'h3b855dcc),
	.w6(32'h3bbeaccb),
	.w7(32'h3be7c423),
	.w8(32'h3b912978),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b458bdb),
	.w1(32'h3af6df27),
	.w2(32'h3bb6f394),
	.w3(32'h3a49a068),
	.w4(32'hb9ba1246),
	.w5(32'h3b98e867),
	.w6(32'h3a96102a),
	.w7(32'h3bd3eb17),
	.w8(32'h3a72115c),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77780c),
	.w1(32'h37ecccff),
	.w2(32'hba875ee3),
	.w3(32'hb9348249),
	.w4(32'h3a15f7eb),
	.w5(32'hb996f578),
	.w6(32'h3aad6c6d),
	.w7(32'hb82eed67),
	.w8(32'hb976dcfb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66fc64),
	.w1(32'hb9588f9f),
	.w2(32'hba2fb101),
	.w3(32'hba0f0716),
	.w4(32'h39bb3302),
	.w5(32'hb91ffe73),
	.w6(32'h3a66fed3),
	.w7(32'h390a7561),
	.w8(32'h3890ecc0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b0c59),
	.w1(32'hba9fa637),
	.w2(32'h3899da6e),
	.w3(32'hb9906280),
	.w4(32'hba005d60),
	.w5(32'h3a47248a),
	.w6(32'hbae31482),
	.w7(32'hba2f5857),
	.w8(32'hba626c0c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8838797),
	.w1(32'hbb858c24),
	.w2(32'hbaac51b0),
	.w3(32'h3a4ba6b3),
	.w4(32'hbb044ca1),
	.w5(32'hbaa5d715),
	.w6(32'hbb0efcf9),
	.w7(32'h3a55d7e9),
	.w8(32'h39b08f77),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd3e02),
	.w1(32'hba9a12e3),
	.w2(32'hb97da616),
	.w3(32'hba148dec),
	.w4(32'hbaa91acd),
	.w5(32'hb9c8e75b),
	.w6(32'hbaddd8d6),
	.w7(32'hba2bd667),
	.w8(32'hbac104a5),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba876501),
	.w1(32'hb9ceb99d),
	.w2(32'hba97e364),
	.w3(32'hba30570e),
	.w4(32'h39d4be3a),
	.w5(32'hba2ae19d),
	.w6(32'h3ad28d6b),
	.w7(32'hb907d9e5),
	.w8(32'h384986ce),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fef45f),
	.w1(32'hba49a87d),
	.w2(32'h3a6569cf),
	.w3(32'hb9f60b73),
	.w4(32'hb9448508),
	.w5(32'h39c9163a),
	.w6(32'hba64bc27),
	.w7(32'hb9cea3e7),
	.w8(32'hba0a5901),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd7c7a),
	.w1(32'h39b4e964),
	.w2(32'h3a9ea4c3),
	.w3(32'h3aaf0c2b),
	.w4(32'h3a00529b),
	.w5(32'h3a9a184c),
	.w6(32'hb9f7c2d8),
	.w7(32'h3ac1c4da),
	.w8(32'h3aa8a356),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8ce5d),
	.w1(32'h399f714e),
	.w2(32'hba212a42),
	.w3(32'hb9cdfa40),
	.w4(32'h3a8ea620),
	.w5(32'h3992d729),
	.w6(32'h3a1aa1d8),
	.w7(32'h36f14d72),
	.w8(32'h3a9088f6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38507dad),
	.w1(32'h39c2079d),
	.w2(32'h3a01f4b0),
	.w3(32'h39ac0908),
	.w4(32'h3a3ea942),
	.w5(32'h3a152f6b),
	.w6(32'h38bad907),
	.w7(32'h3a1e49b0),
	.w8(32'h3a2f43ee),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7644b),
	.w1(32'hb917e978),
	.w2(32'h3b9b873b),
	.w3(32'h3a03e3e0),
	.w4(32'hbb3fc6b8),
	.w5(32'h3b745d57),
	.w6(32'h3b775900),
	.w7(32'h3c24ef9b),
	.w8(32'h3b5815d3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6bc043),
	.w1(32'h3a157408),
	.w2(32'h3a19d906),
	.w3(32'hbaa746a0),
	.w4(32'hb976602c),
	.w5(32'hb8b9840c),
	.w6(32'hb9192515),
	.w7(32'h39c2a528),
	.w8(32'hb9abd08a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ff2200),
	.w1(32'h39dcecac),
	.w2(32'hb925f1f2),
	.w3(32'h386e996a),
	.w4(32'h3a3d9f43),
	.w5(32'h38d94c4e),
	.w6(32'h3a97dd86),
	.w7(32'h3995ad9a),
	.w8(32'hb93e6e48),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98dce4d),
	.w1(32'hb90f0893),
	.w2(32'h3ac2e05a),
	.w3(32'hba129afe),
	.w4(32'h398fdad8),
	.w5(32'h3b2cc2c5),
	.w6(32'hbab66017),
	.w7(32'h3a050fc0),
	.w8(32'hbafe35bb),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba372598),
	.w1(32'hb8b7ae96),
	.w2(32'hb9f36bd7),
	.w3(32'h39981d99),
	.w4(32'h3a50e8ca),
	.w5(32'h3a90c250),
	.w6(32'hba08a953),
	.w7(32'hb9514c05),
	.w8(32'h39a35bb4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba575456),
	.w1(32'hba221e8d),
	.w2(32'hba40135d),
	.w3(32'hb9cbbce5),
	.w4(32'h39daf468),
	.w5(32'hb90173eb),
	.w6(32'hba820d5b),
	.w7(32'hba544241),
	.w8(32'h3949d3e3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2257ff),
	.w1(32'h39ab9da6),
	.w2(32'h3a89a7f5),
	.w3(32'hb9a31a14),
	.w4(32'h3ae8e4e7),
	.w5(32'h3ac3308c),
	.w6(32'h3b24ba72),
	.w7(32'h3af6ea62),
	.w8(32'h3ad2d94b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68620b),
	.w1(32'h3b355ecf),
	.w2(32'h3b4cfe99),
	.w3(32'hb92c4f65),
	.w4(32'h3a80259e),
	.w5(32'h3b013736),
	.w6(32'h3b544141),
	.w7(32'h3ba65627),
	.w8(32'h3a93271e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b625027),
	.w1(32'hb9716f2e),
	.w2(32'hba822f29),
	.w3(32'h3b0cea4f),
	.w4(32'h3916707b),
	.w5(32'hba3bfc8f),
	.w6(32'h39fe50c4),
	.w7(32'hba10f0e4),
	.w8(32'hba1eeb80),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba432ebf),
	.w1(32'h39b91f52),
	.w2(32'hb97a8e2b),
	.w3(32'hba863c68),
	.w4(32'h3a68d12a),
	.w5(32'h39e3ad9c),
	.w6(32'h3a740c84),
	.w7(32'h36dbfa6b),
	.w8(32'h39ffc140),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39867fff),
	.w1(32'hb86ec7c9),
	.w2(32'h38fd9575),
	.w3(32'h3a05a6ab),
	.w4(32'hb91b67c8),
	.w5(32'hb99c32e6),
	.w6(32'hb80d34cb),
	.w7(32'h3a4201cd),
	.w8(32'h3a46ac96),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2de4e),
	.w1(32'hb926b203),
	.w2(32'hb9284202),
	.w3(32'hb9e26a98),
	.w4(32'hba29ebbb),
	.w5(32'hba0178e8),
	.w6(32'h39bf4cbc),
	.w7(32'hba4eb85c),
	.w8(32'hba294803),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba559bc8),
	.w1(32'h397f65e2),
	.w2(32'h3a54beb2),
	.w3(32'h3af7d808),
	.w4(32'h39943bc0),
	.w5(32'h3a9ffff1),
	.w6(32'h3a8384f1),
	.w7(32'h3a5721fb),
	.w8(32'hba447c5f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab177ee),
	.w1(32'h39f99598),
	.w2(32'hb82a44b6),
	.w3(32'hba52baac),
	.w4(32'h3a85c470),
	.w5(32'hb96388b2),
	.w6(32'h3a4a48e1),
	.w7(32'hba42da03),
	.w8(32'hb9ebd7dd),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fa7a0),
	.w1(32'hbb10f04d),
	.w2(32'hb992dbfe),
	.w3(32'h3a5bfe34),
	.w4(32'hbb435b4e),
	.w5(32'hba539c1f),
	.w6(32'hbb0fb10c),
	.w7(32'h38b6e843),
	.w8(32'hbb1947bc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152f01),
	.w1(32'h3a891dcd),
	.w2(32'hb95ac584),
	.w3(32'hbb4cf7ca),
	.w4(32'hbaf0e0a4),
	.w5(32'hbabe065c),
	.w6(32'h3bf59e1a),
	.w7(32'h3bd12af2),
	.w8(32'h3b2c3b74),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ef2e4),
	.w1(32'hba5845a6),
	.w2(32'h3acedbc9),
	.w3(32'hbb984781),
	.w4(32'hbb2bec54),
	.w5(32'h38ad7762),
	.w6(32'hba070e93),
	.w7(32'h3b060a6c),
	.w8(32'h38d243eb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75d3a98),
	.w1(32'hb89d702f),
	.w2(32'hbb05954a),
	.w3(32'hbababb42),
	.w4(32'h3a24f2fc),
	.w5(32'hbac4d48e),
	.w6(32'hba926cc5),
	.w7(32'hbaecd581),
	.w8(32'h391e28c9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb975d34f),
	.w1(32'h39c64bf6),
	.w2(32'h39e7ea64),
	.w3(32'hb80ff797),
	.w4(32'h3a270b05),
	.w5(32'h3a026008),
	.w6(32'h39f2709e),
	.w7(32'h3a446d0a),
	.w8(32'h364d7e79),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05ca57),
	.w1(32'hb9c94753),
	.w2(32'hba8cbbe1),
	.w3(32'hb95389a4),
	.w4(32'h39c20468),
	.w5(32'hb98c5d40),
	.w6(32'h3a0c8f01),
	.w7(32'hb9f4b525),
	.w8(32'h392e8ac4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba101ab5),
	.w1(32'h38855017),
	.w2(32'h39d706c0),
	.w3(32'hb98a185c),
	.w4(32'h389f3ba7),
	.w5(32'h39ae11e5),
	.w6(32'h391a2284),
	.w7(32'h3a1af63a),
	.w8(32'hb8d45fed),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8463282),
	.w1(32'hba0c4aa1),
	.w2(32'hba833b9f),
	.w3(32'hb9ff423b),
	.w4(32'hb9ffeeec),
	.w5(32'hb96e928d),
	.w6(32'h39a8d4ca),
	.w7(32'hba0efca2),
	.w8(32'hb94cd902),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c5a45),
	.w1(32'hbae77000),
	.w2(32'hb995e11c),
	.w3(32'hb8b23d5b),
	.w4(32'hba8e9695),
	.w5(32'h38ad5c1a),
	.w6(32'hbb213332),
	.w7(32'hb8c01603),
	.w8(32'h399fd61a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5e3f1),
	.w1(32'hb6c77898),
	.w2(32'h3a7cb029),
	.w3(32'h3ad50e05),
	.w4(32'h399e12e9),
	.w5(32'h3ae39976),
	.w6(32'hba82c5d2),
	.w7(32'h39c170ff),
	.w8(32'hba9b143b),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0df44e),
	.w1(32'hba8abd6b),
	.w2(32'hba0f9372),
	.w3(32'h399eaee5),
	.w4(32'hb9f50a25),
	.w5(32'hb96c46eb),
	.w6(32'hba92b9aa),
	.w7(32'hb9fb091b),
	.w8(32'hb94ce028),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2d0f),
	.w1(32'hba39e899),
	.w2(32'hbaab5fe2),
	.w3(32'hb9e704a5),
	.w4(32'h38d26b1e),
	.w5(32'hbac68164),
	.w6(32'hbaea2c8b),
	.w7(32'hbaa64f25),
	.w8(32'hba60d6b7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b4f9),
	.w1(32'hba9b14eb),
	.w2(32'h3b83ad61),
	.w3(32'hba8bd622),
	.w4(32'hbb8d1568),
	.w5(32'h39b98711),
	.w6(32'hbb060c83),
	.w7(32'h3b226d24),
	.w8(32'hba870a01),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e38567),
	.w1(32'h3b2f8013),
	.w2(32'h3ba7035f),
	.w3(32'hbb1e1eba),
	.w4(32'h3a390e29),
	.w5(32'h3bb903ba),
	.w6(32'h3bb2f5d1),
	.w7(32'h3c33d398),
	.w8(32'h3bb7928d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb255ef),
	.w1(32'hba178719),
	.w2(32'hb99514ed),
	.w3(32'h3ad1af59),
	.w4(32'hb99cf8d7),
	.w5(32'h39a986bd),
	.w6(32'h3ab43918),
	.w7(32'h39f9216b),
	.w8(32'hb9ab9cd2),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f47351),
	.w1(32'h3a80bc98),
	.w2(32'h398650ec),
	.w3(32'h3a01b9b1),
	.w4(32'h3b4c9348),
	.w5(32'h3ade76a2),
	.w6(32'h39b407f9),
	.w7(32'h39c2115b),
	.w8(32'h3aed48dc),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b70ca),
	.w1(32'hb990613c),
	.w2(32'h39b1deb3),
	.w3(32'h39b24dcc),
	.w4(32'hb9e0e61b),
	.w5(32'h389992e4),
	.w6(32'hba2e0d1e),
	.w7(32'h3a056061),
	.w8(32'hb9bd4a8e),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d5266),
	.w1(32'hb9005f1f),
	.w2(32'hba29f47c),
	.w3(32'hb9f64cc9),
	.w4(32'h393836f0),
	.w5(32'hb9ac4c86),
	.w6(32'h39e7a95a),
	.w7(32'hb9b84903),
	.w8(32'hb9f06117),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba393640),
	.w1(32'hb94823cb),
	.w2(32'hba49b7bc),
	.w3(32'hba2d067a),
	.w4(32'h39b61fc2),
	.w5(32'hb9764e26),
	.w6(32'h3a303cd8),
	.w7(32'hb965ca61),
	.w8(32'h39a5ec8f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef5e62),
	.w1(32'hb9039832),
	.w2(32'hba7dd059),
	.w3(32'hb8e55256),
	.w4(32'h39b29ccd),
	.w5(32'hb9e3190c),
	.w6(32'h3ad6061f),
	.w7(32'h38cf1f67),
	.w8(32'h38eaae6a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95ba1f5),
	.w1(32'h3a4e0c95),
	.w2(32'h3a710b1c),
	.w3(32'hb9a73754),
	.w4(32'h3a5df1a5),
	.w5(32'h3a3b9acf),
	.w6(32'h3a58fa2b),
	.w7(32'h3a9eeb9e),
	.w8(32'h3a2e46a8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980114c),
	.w1(32'hbabd2465),
	.w2(32'h3a8663d2),
	.w3(32'h3a0f4c0d),
	.w4(32'hbb334db9),
	.w5(32'hbaa2ee3a),
	.w6(32'hbabea315),
	.w7(32'hb9a119d7),
	.w8(32'hbacc781e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2e51),
	.w1(32'hba4af3f8),
	.w2(32'hba1f3be4),
	.w3(32'hb9cc44ac),
	.w4(32'hb92fda80),
	.w5(32'h392c3156),
	.w6(32'h3a38402f),
	.w7(32'hba803c38),
	.w8(32'hbab8654b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00477f),
	.w1(32'hba4c9b3b),
	.w2(32'h395eeee8),
	.w3(32'hb70a8a16),
	.w4(32'hba601ae5),
	.w5(32'h397149f0),
	.w6(32'hba8ea726),
	.w7(32'h3a37b72b),
	.w8(32'h39e2ab6b),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e3cc07),
	.w1(32'hbb10b8c7),
	.w2(32'hb9f7c4e7),
	.w3(32'hb9008e40),
	.w4(32'hbb0ab82e),
	.w5(32'hb9cecb66),
	.w6(32'hbb7c5bf1),
	.w7(32'hbad0ac32),
	.w8(32'hbb6e9728),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bc54e),
	.w1(32'h397a5ae7),
	.w2(32'hbae3de9d),
	.w3(32'hbb836f3f),
	.w4(32'h3aa0f982),
	.w5(32'hba4ab96f),
	.w6(32'h3b13a8b8),
	.w7(32'hb993ecb8),
	.w8(32'hba16daeb),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94b1ef),
	.w1(32'h3b2e654b),
	.w2(32'h3bab4383),
	.w3(32'hba988821),
	.w4(32'hba3051c1),
	.w5(32'h3b5443b0),
	.w6(32'h3bf1fb57),
	.w7(32'h3c3d7c98),
	.w8(32'h3bce17d4),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b724f6f),
	.w1(32'hba1eb95a),
	.w2(32'h397bcacc),
	.w3(32'hba6f82ab),
	.w4(32'hbab219b4),
	.w5(32'hba82e612),
	.w6(32'hb8ccd86e),
	.w7(32'hb983709e),
	.w8(32'hbaa4b31c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cf7fa6),
	.w1(32'h3b00e18c),
	.w2(32'h3b00fb21),
	.w3(32'hb9bfc77d),
	.w4(32'h399ec144),
	.w5(32'h3a7573c6),
	.w6(32'h3b0d69ae),
	.w7(32'h3b480f27),
	.w8(32'h3a8a6cf7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b5fe32),
	.w1(32'h388649c5),
	.w2(32'h3a0574a3),
	.w3(32'hba0eaf12),
	.w4(32'h390671bf),
	.w5(32'h39aa76ad),
	.w6(32'h3911f8b1),
	.w7(32'h3a1c528a),
	.w8(32'hb8539a3a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca397a),
	.w1(32'h3b83e86f),
	.w2(32'h3bb79b05),
	.w3(32'hb9bcf584),
	.w4(32'h3ad3e3b2),
	.w5(32'h3b99cde0),
	.w6(32'hbb56424e),
	.w7(32'h3b014241),
	.w8(32'hba3f202e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd9102),
	.w1(32'hb9dbbf1d),
	.w2(32'h3ada4428),
	.w3(32'h3b8a7d8c),
	.w4(32'hbab4133d),
	.w5(32'h39c2ded6),
	.w6(32'hb9e2300a),
	.w7(32'h3ab8a41b),
	.w8(32'h39180466),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a551d2b),
	.w1(32'h39a541d7),
	.w2(32'h399f7e40),
	.w3(32'hba0f6bb2),
	.w4(32'h3a165db1),
	.w5(32'h39059095),
	.w6(32'h39a7d2dd),
	.w7(32'h3a877888),
	.w8(32'h3a1939ae),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a2205),
	.w1(32'h36935d47),
	.w2(32'hba3d9c24),
	.w3(32'h3680499a),
	.w4(32'h39db2ba2),
	.w5(32'hb88fc07d),
	.w6(32'h3acd1fd1),
	.w7(32'h3a0dd008),
	.w8(32'h39833b3a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb992143f),
	.w1(32'hbaff5381),
	.w2(32'hb96faef3),
	.w3(32'hb9a929c9),
	.w4(32'hbb2b2426),
	.w5(32'hb9fb8921),
	.w6(32'hbad5a9ef),
	.w7(32'h38814b95),
	.w8(32'hbb0069c9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245ff3),
	.w1(32'hb956da68),
	.w2(32'hbad544fb),
	.w3(32'hbb2d08c9),
	.w4(32'h38c94d0b),
	.w5(32'hba5b06c3),
	.w6(32'h3b392c79),
	.w7(32'h393b951b),
	.w8(32'hba8dca97),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba866917),
	.w1(32'h39524739),
	.w2(32'hb9003a5a),
	.w3(32'hba289b5d),
	.w4(32'h396b5703),
	.w5(32'h398ce10b),
	.w6(32'h3ab58db6),
	.w7(32'h3a608c51),
	.w8(32'h3a80413c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc8d90),
	.w1(32'hb9badc1b),
	.w2(32'h3ac19010),
	.w3(32'h39c69fa3),
	.w4(32'hba73b393),
	.w5(32'h3a0c672b),
	.w6(32'hbaab5884),
	.w7(32'h385a933f),
	.w8(32'hba9abe86),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e914ba),
	.w1(32'h38eba4ad),
	.w2(32'h3adbbae4),
	.w3(32'hba99eca1),
	.w4(32'hba5925b5),
	.w5(32'h3aab48c6),
	.w6(32'hb9f1bad6),
	.w7(32'h3a9a595e),
	.w8(32'hb9f60cab),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c8f814),
	.w1(32'h3ba60922),
	.w2(32'h3baed9ff),
	.w3(32'hb996ae96),
	.w4(32'h3a87000b),
	.w5(32'h3b5719cb),
	.w6(32'h3c31abef),
	.w7(32'h3c33fea2),
	.w8(32'h3bc0acc7),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64efbe),
	.w1(32'h3a4a0073),
	.w2(32'h3a30c7ac),
	.w3(32'hbac9ec5b),
	.w4(32'hb9eb8d54),
	.w5(32'h36e736ee),
	.w6(32'hba150252),
	.w7(32'hb96ec55c),
	.w8(32'h3812a78c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8174d5),
	.w1(32'hb78b53be),
	.w2(32'h39b7bbb6),
	.w3(32'h377f6805),
	.w4(32'h3a457e31),
	.w5(32'h3a3eb7fa),
	.w6(32'h39dbfad2),
	.w7(32'hb9e5b6fe),
	.w8(32'h3a1c22ab),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9463e1b),
	.w1(32'h3b5b8c30),
	.w2(32'h3b8e61cc),
	.w3(32'hb89af14b),
	.w4(32'h3b5dcf4b),
	.w5(32'h3baa4f39),
	.w6(32'h3b907d32),
	.w7(32'h3bfee0f6),
	.w8(32'h3a78d7ca),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a0dd6),
	.w1(32'hbb2a1d79),
	.w2(32'hbb401816),
	.w3(32'hbaa1e3bb),
	.w4(32'hbb35162d),
	.w5(32'hbb15896a),
	.w6(32'hbb0d5abe),
	.w7(32'hbaf49595),
	.w8(32'hba3dc623),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad53838),
	.w1(32'hba1576a7),
	.w2(32'h39dbb538),
	.w3(32'hb858861f),
	.w4(32'hb9b04bb3),
	.w5(32'h39d4c2fb),
	.w6(32'hb9e7b2d3),
	.w7(32'h39bfaff1),
	.w8(32'hb97344b7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec552),
	.w1(32'h38fa6740),
	.w2(32'h3a17e7e0),
	.w3(32'hb9bed74e),
	.w4(32'hba798136),
	.w5(32'h36951436),
	.w6(32'h3a98d3fb),
	.w7(32'h3a426df7),
	.w8(32'hbb0e5ab9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07c865),
	.w1(32'hbaeb6a7f),
	.w2(32'hba9122ef),
	.w3(32'hba1ee94b),
	.w4(32'hba0c2812),
	.w5(32'hba8b4c42),
	.w6(32'hbb406a43),
	.w7(32'hb9aed1bc),
	.w8(32'h3a20a4bf),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9379e26),
	.w1(32'hba2bce36),
	.w2(32'hba6f7344),
	.w3(32'hb75841b8),
	.w4(32'hb99c7d4e),
	.w5(32'hb98248bd),
	.w6(32'hba0dbf91),
	.w7(32'hba824845),
	.w8(32'hba0170bc),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5e9fb),
	.w1(32'hba69dae4),
	.w2(32'hbad074fc),
	.w3(32'hba8df5d9),
	.w4(32'h3a034724),
	.w5(32'hb7168e76),
	.w6(32'h3a6b1e16),
	.w7(32'hbade9db0),
	.w8(32'hbac75d31),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90656f),
	.w1(32'hb786f846),
	.w2(32'hba1a6489),
	.w3(32'hb96510ea),
	.w4(32'h3a0768bc),
	.w5(32'hb8e7eb9d),
	.w6(32'h3a72ac26),
	.w7(32'hb9bfed92),
	.w8(32'hb9867673),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99347c6),
	.w1(32'hb980c188),
	.w2(32'h3979c007),
	.w3(32'hbaa43dc8),
	.w4(32'hbae65d14),
	.w5(32'hba1ce4fe),
	.w6(32'h39830a06),
	.w7(32'hb96543c8),
	.w8(32'h3992d2df),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ddce25),
	.w1(32'hb926e9e7),
	.w2(32'hba8b25a8),
	.w3(32'h396ca734),
	.w4(32'h3a01bdcb),
	.w5(32'hb9b6f626),
	.w6(32'h3a0298c6),
	.w7(32'hb9973a13),
	.w8(32'hb8bd219c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e90428),
	.w1(32'h397875b6),
	.w2(32'h3a005f60),
	.w3(32'hb7aae708),
	.w4(32'hba618fae),
	.w5(32'hb9cbad24),
	.w6(32'hba0e8445),
	.w7(32'hb94eda05),
	.w8(32'hb9ac7ec2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24f1ec),
	.w1(32'h3a286491),
	.w2(32'hb9c5ec00),
	.w3(32'hb7b64a5d),
	.w4(32'h39dcd458),
	.w5(32'hb7d2fcb3),
	.w6(32'h3b0eb231),
	.w7(32'h3a831b78),
	.w8(32'h3a43e1c5),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3966705b),
	.w1(32'hb93de06f),
	.w2(32'hba4761de),
	.w3(32'hb9b6a8f8),
	.w4(32'h3a40873b),
	.w5(32'h3a16c409),
	.w6(32'h39b6268f),
	.w7(32'hba2b7946),
	.w8(32'hb9d54c48),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99adef0),
	.w1(32'hbac1fb68),
	.w2(32'hbaa38a7c),
	.w3(32'hb85a28b3),
	.w4(32'hba6825cc),
	.w5(32'hba662e85),
	.w6(32'hbacf2aab),
	.w7(32'hba82335d),
	.w8(32'hb98ccbf3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6f32),
	.w1(32'hb9fa7912),
	.w2(32'hba52d389),
	.w3(32'hbac168ae),
	.w4(32'h380ca01f),
	.w5(32'hb90a6f5f),
	.w6(32'h3a2ebc21),
	.w7(32'hb90cd382),
	.w8(32'h3a21735f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392df34f),
	.w1(32'hba77132b),
	.w2(32'hba420561),
	.w3(32'h3a0e5464),
	.w4(32'hb9ea0d95),
	.w5(32'hb808d31e),
	.w6(32'hb9f297a0),
	.w7(32'hba0082da),
	.w8(32'h3a80e83b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b6096),
	.w1(32'hb9e3da6c),
	.w2(32'hba914aba),
	.w3(32'h3a28487f),
	.w4(32'h39985289),
	.w5(32'hb9ab34b4),
	.w6(32'h3ab376bd),
	.w7(32'hb90f1b42),
	.w8(32'h39688819),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399786ee),
	.w1(32'h39d4f7be),
	.w2(32'h3976653c),
	.w3(32'h3a604047),
	.w4(32'hb9550da2),
	.w5(32'hba023737),
	.w6(32'h397e6b10),
	.w7(32'h393431de),
	.w8(32'hb91fbe4e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9365418),
	.w1(32'hbab7b514),
	.w2(32'hbadb5508),
	.w3(32'hb9b4fffb),
	.w4(32'hbab75381),
	.w5(32'hbab9359d),
	.w6(32'hb98d64ae),
	.w7(32'hba8b74bb),
	.w8(32'hba9581d8),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5c991),
	.w1(32'hb8de2d86),
	.w2(32'hba68aad5),
	.w3(32'hbaddee59),
	.w4(32'h3a90af92),
	.w5(32'h3a550c2e),
	.w6(32'h3a1b1e66),
	.w7(32'hba42c70f),
	.w8(32'hba3f86dc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f6257),
	.w1(32'h378b9949),
	.w2(32'hb9bb4b98),
	.w3(32'hb90c2f25),
	.w4(32'h3a05ee8f),
	.w5(32'h3990867a),
	.w6(32'h398ae0c1),
	.w7(32'hb9aec47a),
	.w8(32'hb9776135),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e3666),
	.w1(32'hb5a64738),
	.w2(32'hba0d6617),
	.w3(32'h3918a92b),
	.w4(32'h3a366540),
	.w5(32'h39be6078),
	.w6(32'h39c74e53),
	.w7(32'hb9e34e7f),
	.w8(32'hb90ca773),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9169258),
	.w1(32'hb9519b1b),
	.w2(32'hb9f3cff6),
	.w3(32'h39f2a4c1),
	.w4(32'h39df42c9),
	.w5(32'h3a5d9d18),
	.w6(32'hb92a4b6e),
	.w7(32'hb80edd63),
	.w8(32'h39f23a69),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0803a9),
	.w1(32'hba77d2bf),
	.w2(32'hba9b0985),
	.w3(32'h39cc95be),
	.w4(32'hb95ae35c),
	.w5(32'hba23b5c2),
	.w6(32'hba39f671),
	.w7(32'h39c7335e),
	.w8(32'h3a110399),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8720),
	.w1(32'h3a8eaa49),
	.w2(32'hba54e5c0),
	.w3(32'hb9c8f9eb),
	.w4(32'h3ace7c6b),
	.w5(32'hb95e4497),
	.w6(32'h3aa69c32),
	.w7(32'hba9aa698),
	.w8(32'hba14c6ab),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0197d1),
	.w1(32'hba2b2bd8),
	.w2(32'hba7875ca),
	.w3(32'hb9396e5c),
	.w4(32'h38a00348),
	.w5(32'hb9ff8be1),
	.w6(32'h3a04193e),
	.w7(32'hba0c74c0),
	.w8(32'hba838a5c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dd5b98),
	.w1(32'h371c255e),
	.w2(32'hba441391),
	.w3(32'h3a107069),
	.w4(32'h3a59f55e),
	.w5(32'h39e603db),
	.w6(32'h39d8be22),
	.w7(32'hb9c306f3),
	.w8(32'h3a75361d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb929df5d),
	.w1(32'hb9ec71a2),
	.w2(32'hba39c68e),
	.w3(32'h393bb18b),
	.w4(32'h39809c5d),
	.w5(32'hb8642568),
	.w6(32'h3800887d),
	.w7(32'h3979643e),
	.w8(32'hb9d262b8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace9c81),
	.w1(32'h3817f158),
	.w2(32'h3a270660),
	.w3(32'hba24a77c),
	.w4(32'h39e7014c),
	.w5(32'h3abe46b5),
	.w6(32'h39e582a7),
	.w7(32'h380e42df),
	.w8(32'hbaafa080),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03f041),
	.w1(32'h3a4735f2),
	.w2(32'hbadf22de),
	.w3(32'hb9933f80),
	.w4(32'h3b037367),
	.w5(32'hb958e249),
	.w6(32'h3b5309f0),
	.w7(32'h3a25bec1),
	.w8(32'h3a02953f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba436a78),
	.w1(32'hba222b3a),
	.w2(32'hba8dc3a3),
	.w3(32'hb985d6f6),
	.w4(32'hba7e7fdd),
	.w5(32'hba5f40d7),
	.w6(32'hba78f4ed),
	.w7(32'hbaba75f6),
	.w8(32'hb9b6a819),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c04eed),
	.w1(32'h39ee8648),
	.w2(32'h3a1404ee),
	.w3(32'hba234df5),
	.w4(32'h3794e901),
	.w5(32'h39f78c2d),
	.w6(32'h3a4f1005),
	.w7(32'h39bc6e83),
	.w8(32'hb8e6a7c2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57643d),
	.w1(32'h3ae537bf),
	.w2(32'hbb238a08),
	.w3(32'h3a50cf57),
	.w4(32'h38a460f1),
	.w5(32'hba585a15),
	.w6(32'h399a6d0a),
	.w7(32'hbb1c4475),
	.w8(32'hb9b7e6f8),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bff2a6),
	.w1(32'hba6bda47),
	.w2(32'hba4fddb9),
	.w3(32'hbadf858c),
	.w4(32'hb9d83d25),
	.w5(32'hba4e66c9),
	.w6(32'hbaa19a0f),
	.w7(32'hba9cfc7b),
	.w8(32'hbae1630a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb52fa),
	.w1(32'hba1b71ce),
	.w2(32'hb77571fd),
	.w3(32'hba87b292),
	.w4(32'h399b9352),
	.w5(32'hb9c220b8),
	.w6(32'h35f06294),
	.w7(32'hba1cdfa7),
	.w8(32'hbad9f043),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba408121),
	.w1(32'h3a499ef7),
	.w2(32'h3ab83dbd),
	.w3(32'h3805f0f1),
	.w4(32'h3b1d4c4a),
	.w5(32'h3b57b8c5),
	.w6(32'h3aafddfb),
	.w7(32'h3adce23f),
	.w8(32'h3afe7a9f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36e851),
	.w1(32'h3b24b3a8),
	.w2(32'hba155e25),
	.w3(32'h3b6078af),
	.w4(32'h3ad7592e),
	.w5(32'hba10cf9f),
	.w6(32'h3b58658e),
	.w7(32'h3a47e4fb),
	.w8(32'h39b76544),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af93dd8),
	.w1(32'h3ad32778),
	.w2(32'h3aa38ccc),
	.w3(32'h3b17219b),
	.w4(32'h3aeec374),
	.w5(32'h3ac83b66),
	.w6(32'h3a9de124),
	.w7(32'h3a36c446),
	.w8(32'h3a7b5a8e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7148c0f),
	.w1(32'hbaa587d9),
	.w2(32'hbabd983e),
	.w3(32'h39d07404),
	.w4(32'hbb15877b),
	.w5(32'hbb1088c2),
	.w6(32'hbac23cff),
	.w7(32'hbb095ca4),
	.w8(32'hbb56b53f),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11f6a4),
	.w1(32'hb93ab110),
	.w2(32'h39a907a7),
	.w3(32'hbae60186),
	.w4(32'hba0165fd),
	.w5(32'h3971fb85),
	.w6(32'h3894082d),
	.w7(32'hb968c263),
	.w8(32'hb8fe5217),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8df0ff8),
	.w1(32'h3a5d7453),
	.w2(32'h3a57758b),
	.w3(32'hb9594a13),
	.w4(32'h38504202),
	.w5(32'h39a3d6ed),
	.w6(32'h3a1bf213),
	.w7(32'hb9864cd1),
	.w8(32'hb9995978),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0153d),
	.w1(32'hbb42d1c9),
	.w2(32'hbb22047b),
	.w3(32'hba4186ef),
	.w4(32'hbb44dd46),
	.w5(32'hbb1eb447),
	.w6(32'hbb37431b),
	.w7(32'hbac1b53e),
	.w8(32'hbacb42c0),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820d75),
	.w1(32'h3ad4e93b),
	.w2(32'h3a8c4b1c),
	.w3(32'hbaa9fd46),
	.w4(32'h3abd1222),
	.w5(32'h39cf5205),
	.w6(32'h3b0c13b2),
	.w7(32'h39e1bad1),
	.w8(32'hba66cc4b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba459683),
	.w1(32'h3ac0d548),
	.w2(32'h3a24be7e),
	.w3(32'hba7b4d83),
	.w4(32'hb9d9c2e4),
	.w5(32'hbaa5a23f),
	.w6(32'h3a89e026),
	.w7(32'h3aa22936),
	.w8(32'h3aae682e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7fe1ad),
	.w1(32'hb90df171),
	.w2(32'hb7f4ed63),
	.w3(32'h38eb84d8),
	.w4(32'hb98e4a9d),
	.w5(32'h370071e2),
	.w6(32'hb9a49092),
	.w7(32'hba05dff6),
	.w8(32'hb81755a3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab289),
	.w1(32'hba2d59be),
	.w2(32'h359e43f9),
	.w3(32'h38807935),
	.w4(32'hbaabdf51),
	.w5(32'hba7b8e86),
	.w6(32'hba358990),
	.w7(32'hba886337),
	.w8(32'hba3e4573),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3c86c),
	.w1(32'h3b30e2a1),
	.w2(32'hb8ae2b12),
	.w3(32'hbab64863),
	.w4(32'h3afaeb0f),
	.w5(32'hb9a6fec2),
	.w6(32'h3b087537),
	.w7(32'h3ac6cfc0),
	.w8(32'hb9cb830f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae51f57),
	.w1(32'h3a52540e),
	.w2(32'h3aaa91cf),
	.w3(32'h3a9208ff),
	.w4(32'h39c99f6d),
	.w5(32'h39fe6d33),
	.w6(32'h39f78f6a),
	.w7(32'h3a108e5b),
	.w8(32'hb69f14ff),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9552b1d),
	.w1(32'hba0b13e5),
	.w2(32'h3aa48178),
	.w3(32'h39a7cd76),
	.w4(32'h3a87f0b1),
	.w5(32'h3a2a4c15),
	.w6(32'h39df1da4),
	.w7(32'h3a4d0862),
	.w8(32'h3a83bf53),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29f3dc),
	.w1(32'hbae15482),
	.w2(32'hbacfb2ff),
	.w3(32'h39e5cc79),
	.w4(32'hbadca34f),
	.w5(32'hba7789b7),
	.w6(32'hbb103c44),
	.w7(32'hba9bf7b3),
	.w8(32'hbab8e15b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7d51),
	.w1(32'hb8bf9cea),
	.w2(32'hb9c7cdd8),
	.w3(32'hba7901aa),
	.w4(32'hb937e197),
	.w5(32'h39970ecc),
	.w6(32'hb9a3e0b2),
	.w7(32'h38f2ed24),
	.w8(32'h390257b7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c83f8),
	.w1(32'h3a83c581),
	.w2(32'h3a6ef0f8),
	.w3(32'h39bdcbc4),
	.w4(32'h390a1f8d),
	.w5(32'h39e50799),
	.w6(32'h39b384da),
	.w7(32'h3a10a12f),
	.w8(32'h398e8ade),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9202d),
	.w1(32'hba7e0b76),
	.w2(32'hb9e59546),
	.w3(32'h397f372b),
	.w4(32'hba90c08b),
	.w5(32'hba5e798e),
	.w6(32'hbabcccbb),
	.w7(32'hbac8566d),
	.w8(32'hbaba2efd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cb674),
	.w1(32'h3af77894),
	.w2(32'h3b2676ac),
	.w3(32'hba8b5ee2),
	.w4(32'h3a55e145),
	.w5(32'hb717a808),
	.w6(32'h3aa149f1),
	.w7(32'h393fb8b4),
	.w8(32'h39aff9f5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b743e3),
	.w1(32'hba3427a3),
	.w2(32'hb9c405d6),
	.w3(32'hbaf7580f),
	.w4(32'h3ae3aa92),
	.w5(32'h3abd823b),
	.w6(32'h38d0e708),
	.w7(32'hba515b13),
	.w8(32'h3a1ffeb4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0049b),
	.w1(32'hba4615d1),
	.w2(32'hb94934c2),
	.w3(32'h3abef5da),
	.w4(32'hbacf7c49),
	.w5(32'hbaa89f05),
	.w6(32'hb8bdefc2),
	.w7(32'hba90edb8),
	.w8(32'hbadb4906),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38194fa3),
	.w1(32'h3ad962ff),
	.w2(32'h3a2785ce),
	.w3(32'hb9790ff8),
	.w4(32'h3a5c842e),
	.w5(32'h390a8468),
	.w6(32'h3a6af09f),
	.w7(32'h3a8a05b7),
	.w8(32'h39a94787),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899abf5),
	.w1(32'h3a824ddc),
	.w2(32'h39921508),
	.w3(32'h39808ef8),
	.w4(32'h3af52ba9),
	.w5(32'h3ad249f1),
	.w6(32'h3a1f03d7),
	.w7(32'h39de54ed),
	.w8(32'h3ab349b3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a765e11),
	.w1(32'h3a544dff),
	.w2(32'h3a8118ef),
	.w3(32'h3a91afff),
	.w4(32'h38849aca),
	.w5(32'h3992c94f),
	.w6(32'h39d578c7),
	.w7(32'h39b608ed),
	.w8(32'hb8ae0d17),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4d0cd),
	.w1(32'h3adb91be),
	.w2(32'hba00a624),
	.w3(32'h37f6bd4d),
	.w4(32'h3a19d3ea),
	.w5(32'h38bdda98),
	.w6(32'h3ab7b8e6),
	.w7(32'h3aeffe31),
	.w8(32'h3987f991),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45b901),
	.w1(32'h3a873786),
	.w2(32'h3b0f7390),
	.w3(32'h3ae3c707),
	.w4(32'h388356dd),
	.w5(32'h3aa7de57),
	.w6(32'hb6aab51f),
	.w7(32'h3a821f08),
	.w8(32'hb99a8490),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb999f81c),
	.w1(32'hba579248),
	.w2(32'hba99c640),
	.w3(32'hb8459e86),
	.w4(32'h38aa9cdd),
	.w5(32'hba7a6f8c),
	.w6(32'hb949686e),
	.w7(32'hbacd304f),
	.w8(32'hba852150),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e4bb1),
	.w1(32'hb928b021),
	.w2(32'h3962ec64),
	.w3(32'hba09db98),
	.w4(32'hba0b9ff8),
	.w5(32'hba33fb9e),
	.w6(32'hb993e6a5),
	.w7(32'hba6af285),
	.w8(32'hba4ccffe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca2490),
	.w1(32'hba01d3ea),
	.w2(32'h3914fb05),
	.w3(32'hba24e195),
	.w4(32'hba6fcee8),
	.w5(32'hb9eb800b),
	.w6(32'hba2308de),
	.w7(32'hba2d0076),
	.w8(32'hba0a5640),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9e83d),
	.w1(32'h3af68b59),
	.w2(32'h3a3d1efe),
	.w3(32'hba6f0bf2),
	.w4(32'h39bebbda),
	.w5(32'h39f220e5),
	.w6(32'h3acd27e0),
	.w7(32'h3a67c572),
	.w8(32'h3b105e83),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10aec9),
	.w1(32'h3ab43310),
	.w2(32'h39abd393),
	.w3(32'h3aaac8a6),
	.w4(32'h39d71afa),
	.w5(32'h3adc1bb5),
	.w6(32'h39ef7e04),
	.w7(32'h39b15507),
	.w8(32'h3a965394),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1a092),
	.w1(32'hba8db3a2),
	.w2(32'hbafa9257),
	.w3(32'h3a9db0a2),
	.w4(32'hba0ae3c8),
	.w5(32'hba1858c7),
	.w6(32'hba81fd13),
	.w7(32'hba46df34),
	.w8(32'hba633333),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94f2a9),
	.w1(32'h3a18f2fc),
	.w2(32'h3a60129e),
	.w3(32'hba19748c),
	.w4(32'hb98e3813),
	.w5(32'hb9e5f229),
	.w6(32'h39b4b346),
	.w7(32'h39379bc8),
	.w8(32'hb9906766),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67376f3),
	.w1(32'h38e2664e),
	.w2(32'hbaa08bf2),
	.w3(32'hba049161),
	.w4(32'h3a027054),
	.w5(32'hba0c5600),
	.w6(32'hb906d615),
	.w7(32'hba63e4bf),
	.w8(32'hbb0f6cab),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb222b5a),
	.w1(32'hb9c58a52),
	.w2(32'hb9bfdd8d),
	.w3(32'hba73e1a2),
	.w4(32'hb9b2be2a),
	.w5(32'hba33703f),
	.w6(32'hba34fe84),
	.w7(32'hba24a0c4),
	.w8(32'hba6936c7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4714),
	.w1(32'h3996a457),
	.w2(32'h3a50c12f),
	.w3(32'hba32d1c4),
	.w4(32'hb9ce2b79),
	.w5(32'h3924b8e0),
	.w6(32'h397878dd),
	.w7(32'h3908348c),
	.w8(32'hb9ac01d6),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c38da2),
	.w1(32'hb918e848),
	.w2(32'hba35c3e7),
	.w3(32'h397babcd),
	.w4(32'h390913a5),
	.w5(32'hb98d8fad),
	.w6(32'hb9ceb87d),
	.w7(32'hba435bcd),
	.w8(32'hba9f23c9),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e995f),
	.w1(32'hba2499dc),
	.w2(32'hbad3d247),
	.w3(32'hb9d5e1c9),
	.w4(32'h39e54be0),
	.w5(32'hba7af24b),
	.w6(32'h3a7a3ee8),
	.w7(32'hbb022423),
	.w8(32'hba515dcc),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac818d2),
	.w1(32'h3a2d96c6),
	.w2(32'hba804220),
	.w3(32'h393cc71e),
	.w4(32'h399c773c),
	.w5(32'hba9a9cc1),
	.w6(32'h39ed9485),
	.w7(32'h383abe4f),
	.w8(32'hba7ab386),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b765),
	.w1(32'hba1b4f37),
	.w2(32'hb98b1ea1),
	.w3(32'hba1bf39c),
	.w4(32'hba04487c),
	.w5(32'h3a02ca84),
	.w6(32'hba3cbd7f),
	.w7(32'hb95d5efd),
	.w8(32'h38e924c2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f76d8),
	.w1(32'hbb113f3c),
	.w2(32'hbaaea80a),
	.w3(32'hba039bd5),
	.w4(32'hbb151639),
	.w5(32'hbb013e9b),
	.w6(32'hbb676f32),
	.w7(32'hbaa7797d),
	.w8(32'hbada7f37),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0be32),
	.w1(32'hbaf060fd),
	.w2(32'hb987abdc),
	.w3(32'hbaf45840),
	.w4(32'hbb3f7215),
	.w5(32'hbb18389f),
	.w6(32'hbb2f070f),
	.w7(32'hbad2d51b),
	.w8(32'hba87537c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902891a),
	.w1(32'h3984e1a4),
	.w2(32'hba7d1193),
	.w3(32'hbaac53d5),
	.w4(32'hbaa025f1),
	.w5(32'hbb064220),
	.w6(32'hb9d28998),
	.w7(32'hba8e79f9),
	.w8(32'hba32fcd4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9589ff),
	.w1(32'h3a70f165),
	.w2(32'hba18c752),
	.w3(32'hbb07593b),
	.w4(32'h3a0f48fa),
	.w5(32'hb981474f),
	.w6(32'h3ac8c3ac),
	.w7(32'h3a269f50),
	.w8(32'h38ccd139),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7005de),
	.w1(32'h3abb2aa0),
	.w2(32'h3ac13477),
	.w3(32'h3a6af2d2),
	.w4(32'h3a6d3702),
	.w5(32'h3a33d639),
	.w6(32'h3a8e1841),
	.w7(32'h38fedf45),
	.w8(32'hb9f7ebad),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd180c),
	.w1(32'hb99903fd),
	.w2(32'h383b83db),
	.w3(32'hba46b6ad),
	.w4(32'hba687172),
	.w5(32'hb910f813),
	.w6(32'hb9f5ba01),
	.w7(32'hb9f7a68b),
	.w8(32'hb967a204),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9245cdc),
	.w1(32'hb9ce033f),
	.w2(32'h3801cae3),
	.w3(32'hb9ad4ae9),
	.w4(32'hba845d48),
	.w5(32'hba20e570),
	.w6(32'hba1a344d),
	.w7(32'hba58c4b1),
	.w8(32'hbaa528db),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba681041),
	.w1(32'hbab700f3),
	.w2(32'hba852df7),
	.w3(32'hba75167e),
	.w4(32'hbb1a3e02),
	.w5(32'hbb032272),
	.w6(32'hbb3d1662),
	.w7(32'hbb0b2591),
	.w8(32'hbb1cd3e3),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef7b78),
	.w1(32'h3b3f9b16),
	.w2(32'hbb7139dc),
	.w3(32'hbafaaaa6),
	.w4(32'h3a821605),
	.w5(32'hbb549fee),
	.w6(32'h3a94ea43),
	.w7(32'h397dd6aa),
	.w8(32'hbac92a21),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15c5fc),
	.w1(32'h3b0efd6c),
	.w2(32'h3b814fea),
	.w3(32'hba8da97b),
	.w4(32'h3b061d37),
	.w5(32'h3b222a1c),
	.w6(32'h3aafefac),
	.w7(32'h3ad14638),
	.w8(32'h3a506833),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a23d831),
	.w1(32'h3afbb5d0),
	.w2(32'hba2edf1e),
	.w3(32'h3ac55264),
	.w4(32'h3b086d33),
	.w5(32'hb908761f),
	.w6(32'h3b17445a),
	.w7(32'h3a71ef59),
	.w8(32'h3a503cad),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a985148),
	.w1(32'hb7e86713),
	.w2(32'hb9c26ce9),
	.w3(32'h3aba1042),
	.w4(32'h3a8e09cb),
	.w5(32'h3a0c322a),
	.w6(32'h3a046883),
	.w7(32'h3a4a1503),
	.w8(32'h3a317858),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f19b1b),
	.w1(32'hb985a876),
	.w2(32'hb9b4705e),
	.w3(32'hb9482437),
	.w4(32'h3a7ba96d),
	.w5(32'h3a144f8d),
	.w6(32'h39df484c),
	.w7(32'hba456b8e),
	.w8(32'hbab21418),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b530),
	.w1(32'hbab0ebaa),
	.w2(32'h3900ef83),
	.w3(32'h3940b405),
	.w4(32'h396e3fab),
	.w5(32'hb72a2410),
	.w6(32'hba61ccc5),
	.w7(32'hb9863e61),
	.w8(32'h39dd99b5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32d0ac),
	.w1(32'h3b836c7c),
	.w2(32'hbb2fe9c0),
	.w3(32'hb9bfe5a8),
	.w4(32'h3b184032),
	.w5(32'hba3448fa),
	.w6(32'h3b22f048),
	.w7(32'hb9bee2af),
	.w8(32'hba4c6655),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09f87f),
	.w1(32'hba05b9ea),
	.w2(32'hba2856f5),
	.w3(32'hb9b42c26),
	.w4(32'hb8e8b816),
	.w5(32'hba6a241b),
	.w6(32'hba893f44),
	.w7(32'hba8ef8c7),
	.w8(32'hbad3f350),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaac9f28),
	.w1(32'hba465d2e),
	.w2(32'hb9627b58),
	.w3(32'hbad6f3c8),
	.w4(32'hbabf3a07),
	.w5(32'hba2dde43),
	.w6(32'h3866a17f),
	.w7(32'hba723734),
	.w8(32'hbade2b40),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0332ea),
	.w1(32'hb9f49fc2),
	.w2(32'hb8ee7e71),
	.w3(32'h37896583),
	.w4(32'h38ccf437),
	.w5(32'h39829640),
	.w6(32'hba1ca8b6),
	.w7(32'hba2fe1fc),
	.w8(32'h3914a0b9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba973aa4),
	.w1(32'h3a266e55),
	.w2(32'h3a3ad4c0),
	.w3(32'hb9c3af72),
	.w4(32'hb9b8362e),
	.w5(32'hb9e390b9),
	.w6(32'h39a18ba1),
	.w7(32'hba3f52c9),
	.w8(32'hbad6baa2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac8272),
	.w1(32'h3ae7f0cb),
	.w2(32'hbb21a643),
	.w3(32'hb9ee7738),
	.w4(32'h39440575),
	.w5(32'hbace7558),
	.w6(32'h3aafc2fa),
	.w7(32'hbab89439),
	.w8(32'h39a38ef9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cd5ca),
	.w1(32'hbabd2598),
	.w2(32'hba90e0c4),
	.w3(32'h3a7f6b3f),
	.w4(32'hbacc305c),
	.w5(32'hbab65ab3),
	.w6(32'hbb120e83),
	.w7(32'hba5687d2),
	.w8(32'hba8ec160),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa013ee),
	.w1(32'hba3dfe06),
	.w2(32'h399e1f94),
	.w3(32'hbab1c815),
	.w4(32'hbaa2ab74),
	.w5(32'h37d5200c),
	.w6(32'hba2ad224),
	.w7(32'hb888f8cd),
	.w8(32'hb8ecdeff),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9db5922),
	.w1(32'h3b1d7fe3),
	.w2(32'hbb086b18),
	.w3(32'hba45450f),
	.w4(32'h3aa5e73b),
	.w5(32'hb9007592),
	.w6(32'h3adf511e),
	.w7(32'hb972fde6),
	.w8(32'h3a2fcacc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e9913),
	.w1(32'hb868d2fb),
	.w2(32'hb9b7d399),
	.w3(32'h3914feb7),
	.w4(32'h3a89de45),
	.w5(32'h39bc8881),
	.w6(32'h39e7f4a6),
	.w7(32'hba676995),
	.w8(32'hb8a1d401),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6441e8),
	.w1(32'hba96fb76),
	.w2(32'hbafeedcc),
	.w3(32'h39ea997b),
	.w4(32'h3a00acbf),
	.w5(32'hb9f88b2f),
	.w6(32'hb9eefd69),
	.w7(32'hbb06afe3),
	.w8(32'h38106d6c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae635e6),
	.w1(32'h3a474d1a),
	.w2(32'h3af267dd),
	.w3(32'h3a04cd92),
	.w4(32'h3a1379e3),
	.w5(32'h39ebf097),
	.w6(32'h3a416d3d),
	.w7(32'h3a838631),
	.w8(32'hb8bc63f8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c6d22a),
	.w1(32'hba84bc89),
	.w2(32'hbb120e90),
	.w3(32'h391adf1d),
	.w4(32'hbb6100c7),
	.w5(32'hbb165ab7),
	.w6(32'hbb04e8e3),
	.w7(32'hbb17f9c5),
	.w8(32'hbad0424b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba972586),
	.w1(32'hba77fc56),
	.w2(32'hba718479),
	.w3(32'hbb04c1d3),
	.w4(32'hb9b72ee9),
	.w5(32'hb9fb0e2a),
	.w6(32'hba6b226d),
	.w7(32'hba289336),
	.w8(32'hba67a252),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba601b37),
	.w1(32'h39fac348),
	.w2(32'h3a525c24),
	.w3(32'hba0f57bf),
	.w4(32'h38dfea74),
	.w5(32'h39842f5f),
	.w6(32'h3a189708),
	.w7(32'h3947aaeb),
	.w8(32'h38e91701),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e457d),
	.w1(32'h39a10701),
	.w2(32'h3a3aa8c6),
	.w3(32'h38a3da52),
	.w4(32'hb9915e0a),
	.w5(32'h39517640),
	.w6(32'h3a2e95cf),
	.w7(32'h3a1ca3d2),
	.w8(32'hb93cd3df),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6de478b),
	.w1(32'hb9c74f00),
	.w2(32'h399fffe1),
	.w3(32'h38f67e6f),
	.w4(32'hba8087df),
	.w5(32'hba35c827),
	.w6(32'hba1a4fa4),
	.w7(32'hb9ddd6ef),
	.w8(32'hba6c3a5c),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4c86),
	.w1(32'hb991b706),
	.w2(32'hba0e6f9e),
	.w3(32'hba7d5eb0),
	.w4(32'hba0668cd),
	.w5(32'hba2afcae),
	.w6(32'hb9c50d13),
	.w7(32'hba35feae),
	.w8(32'hbac5488e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8f21c),
	.w1(32'h3b0b11f5),
	.w2(32'hbb0728ab),
	.w3(32'hba45b45f),
	.w4(32'hb9ebdc12),
	.w5(32'hba384aaa),
	.w6(32'h3b13f3de),
	.w7(32'h39c67064),
	.w8(32'h39370b40),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de2416),
	.w1(32'h3a0205b2),
	.w2(32'h3a87684d),
	.w3(32'hba136487),
	.w4(32'hb87f5e0b),
	.w5(32'h3a35ff9e),
	.w6(32'h38fd58a9),
	.w7(32'hb8c262f6),
	.w8(32'h38e23eb4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d5fcc),
	.w1(32'hb98edddf),
	.w2(32'hbacc3cd8),
	.w3(32'h3886aade),
	.w4(32'hba5150c0),
	.w5(32'hbabb71ff),
	.w6(32'hb916a3a1),
	.w7(32'hbac8c912),
	.w8(32'hba641ef5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac5982),
	.w1(32'hb9940758),
	.w2(32'hb9d6760c),
	.w3(32'h3998b3b8),
	.w4(32'h3b1aff87),
	.w5(32'h3b4c20e8),
	.w6(32'h3a6d8cdc),
	.w7(32'h3b0c3225),
	.w8(32'h3b5bc228),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af78ecd),
	.w1(32'hba04b58c),
	.w2(32'hba394a6a),
	.w3(32'h3aad2ff9),
	.w4(32'hba19fe54),
	.w5(32'hba48d255),
	.w6(32'hba506628),
	.w7(32'hbac8d6fa),
	.w8(32'hba8ce17e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce0be4),
	.w1(32'hba3483be),
	.w2(32'hba8435c0),
	.w3(32'hba18473f),
	.w4(32'h383887fb),
	.w5(32'hba07c334),
	.w6(32'hba64a129),
	.w7(32'hbb062937),
	.w8(32'hba20596d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1ede5),
	.w1(32'hb964dcbb),
	.w2(32'hba11e3d5),
	.w3(32'h39b6a79a),
	.w4(32'h396c619f),
	.w5(32'hbaa0981b),
	.w6(32'hba16528d),
	.w7(32'hbaac0dde),
	.w8(32'hbb0fbe20),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbb98),
	.w1(32'h3aaa7bd4),
	.w2(32'h3a6cde85),
	.w3(32'hbaa46d58),
	.w4(32'h3a95cbe9),
	.w5(32'h39906bc5),
	.w6(32'h3a9aa5fd),
	.w7(32'h3a66c682),
	.w8(32'h399c96db),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395e9274),
	.w1(32'hba4d5c78),
	.w2(32'hb9d70d98),
	.w3(32'h39c37a88),
	.w4(32'hb9e18f04),
	.w5(32'hba4a812b),
	.w6(32'hba36c5f3),
	.w7(32'hba8f315d),
	.w8(32'hba7ba48a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad01367),
	.w1(32'hbaef80bb),
	.w2(32'hba69213f),
	.w3(32'hba9b50ed),
	.w4(32'hba157899),
	.w5(32'hba9ee846),
	.w6(32'h39ae75d0),
	.w7(32'hbb2c0914),
	.w8(32'hbac6d7a1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6debd1),
	.w1(32'h3986c6c9),
	.w2(32'h38f05f98),
	.w3(32'hba656b56),
	.w4(32'h3aa01cb2),
	.w5(32'h3a190eba),
	.w6(32'h3946e780),
	.w7(32'hb9595d0e),
	.w8(32'h3885e618),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75e194),
	.w1(32'hbad1e339),
	.w2(32'hbac2c96b),
	.w3(32'hb7598b66),
	.w4(32'hbb080ff5),
	.w5(32'hbaa6c5f0),
	.w6(32'hbabeaa8b),
	.w7(32'hbb087bfb),
	.w8(32'hbaa4471c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc6644),
	.w1(32'hb93c1fbf),
	.w2(32'h3928a168),
	.w3(32'hba80ee28),
	.w4(32'hb99a4803),
	.w5(32'hb99bf400),
	.w6(32'hba0f99b5),
	.w7(32'hba4198d3),
	.w8(32'hba3cb4d4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba124f9a),
	.w1(32'h3870cceb),
	.w2(32'hb90f8ca4),
	.w3(32'hba0dbbff),
	.w4(32'h3a1710dc),
	.w5(32'hb8f03bb2),
	.w6(32'h38899ff4),
	.w7(32'h39824011),
	.w8(32'hb8c39151),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f6c73),
	.w1(32'hba8b1a49),
	.w2(32'h3897e286),
	.w3(32'hb9756c09),
	.w4(32'hbaa89a81),
	.w5(32'hba817ec0),
	.w6(32'hba93e5ac),
	.w7(32'hbabae5ee),
	.w8(32'hbab3ab70),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba933655),
	.w1(32'hbac1f301),
	.w2(32'hba8e48ec),
	.w3(32'hbab47bbf),
	.w4(32'hbb021e57),
	.w5(32'hbac2073e),
	.w6(32'hba32ce7e),
	.w7(32'hbb06065b),
	.w8(32'hbb1db30d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc3eeb),
	.w1(32'hbb04e834),
	.w2(32'hbab2f513),
	.w3(32'hbae02d4c),
	.w4(32'hbb3fbaed),
	.w5(32'hbb3668fc),
	.w6(32'hbb222155),
	.w7(32'hbb062463),
	.w8(32'hbb07f68d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabefc45),
	.w1(32'h39bbb4ef),
	.w2(32'hba25ff09),
	.w3(32'hbab879a7),
	.w4(32'h3a69789f),
	.w5(32'h39a059f5),
	.w6(32'hb8372907),
	.w7(32'hb9ffbe7e),
	.w8(32'hb9b6ff6b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48aa5f),
	.w1(32'h39222ee2),
	.w2(32'h3982ee38),
	.w3(32'hb923a43d),
	.w4(32'h3a9086f0),
	.w5(32'h3a53be86),
	.w6(32'hb9a901e2),
	.w7(32'hba0597a2),
	.w8(32'hb4a476b8),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ca1d6),
	.w1(32'hba882a0a),
	.w2(32'hb8eb0111),
	.w3(32'h39ed1ff4),
	.w4(32'hb90dac1f),
	.w5(32'hba154feb),
	.w6(32'hb9ad9038),
	.w7(32'hb9e53ddd),
	.w8(32'hba5b85bc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2068db),
	.w1(32'h39bf518a),
	.w2(32'h3a416640),
	.w3(32'hb9743a8a),
	.w4(32'h3a591a1d),
	.w5(32'h3a910ecc),
	.w6(32'h38a599ce),
	.w7(32'hba89b7ae),
	.w8(32'h39db42fb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a961253),
	.w1(32'hba00795f),
	.w2(32'hba982a95),
	.w3(32'hba540dea),
	.w4(32'h3a534f48),
	.w5(32'h39d85ef1),
	.w6(32'h3a36a555),
	.w7(32'hba41019a),
	.w8(32'h3af9f31c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab84ead),
	.w1(32'h3b3667d8),
	.w2(32'hb91500c2),
	.w3(32'h3b7442f8),
	.w4(32'h3aeb0d53),
	.w5(32'h3aad7deb),
	.w6(32'h3aa45a4d),
	.w7(32'h3985bb71),
	.w8(32'h3aa01144),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa72f45),
	.w1(32'hba2bb029),
	.w2(32'hba22fea0),
	.w3(32'h3a9eb659),
	.w4(32'hb94d5934),
	.w5(32'hba6b5bef),
	.w6(32'hba3c8614),
	.w7(32'hba6e0118),
	.w8(32'hbad5ded9),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c193),
	.w1(32'h3a828819),
	.w2(32'h39af02a5),
	.w3(32'hba744f11),
	.w4(32'h3a264d1c),
	.w5(32'h39c686bb),
	.w6(32'h39ef1190),
	.w7(32'h39689535),
	.w8(32'hba464b0d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96d737),
	.w1(32'h3b85accc),
	.w2(32'hbb330e18),
	.w3(32'h3a3c447e),
	.w4(32'h3b558ac5),
	.w5(32'hb9d138d8),
	.w6(32'h3b583302),
	.w7(32'h3a193090),
	.w8(32'h3aba0186),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02035b),
	.w1(32'h3b262f3a),
	.w2(32'hbb20751f),
	.w3(32'hb92624e8),
	.w4(32'h3ac475ff),
	.w5(32'h38f82aee),
	.w6(32'h3b3ca200),
	.w7(32'h38c1c207),
	.w8(32'h3a3807ef),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49c4e1),
	.w1(32'hba3f2ac9),
	.w2(32'h3a98c3c2),
	.w3(32'hbafd2b8f),
	.w4(32'hbb005bce),
	.w5(32'hba4c72e9),
	.w6(32'hb887b43d),
	.w7(32'hbaa23efc),
	.w8(32'hbb02d7ca),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398aa342),
	.w1(32'h3a7c42a0),
	.w2(32'h3a7751cd),
	.w3(32'h36c709c0),
	.w4(32'h39c90301),
	.w5(32'h395f4fc8),
	.w6(32'h3a8cac27),
	.w7(32'h395d7c8e),
	.w8(32'h38c9557b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a331828),
	.w1(32'h39dbf088),
	.w2(32'h3a400f46),
	.w3(32'h3a1211a0),
	.w4(32'hb8f2c53c),
	.w5(32'h39ae0a77),
	.w6(32'h391a891f),
	.w7(32'hb7c4bcb3),
	.w8(32'hb9480c93),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380365af),
	.w1(32'h3a66fe6c),
	.w2(32'h3a693290),
	.w3(32'hb95d1428),
	.w4(32'hb97879c9),
	.w5(32'h38b8be11),
	.w6(32'h3a196022),
	.w7(32'h39643b47),
	.w8(32'hb9ab37ae),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed8f1b),
	.w1(32'hba7db5ab),
	.w2(32'hb9bbee18),
	.w3(32'h398b69e2),
	.w4(32'hba590db0),
	.w5(32'hba73bdcc),
	.w6(32'hba2b8391),
	.w7(32'hba9e9dbc),
	.w8(32'hbae41696),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86b879),
	.w1(32'hba1a9338),
	.w2(32'hb9808b48),
	.w3(32'hba35f625),
	.w4(32'hba270611),
	.w5(32'hba1f86d1),
	.w6(32'hba83c7c6),
	.w7(32'hbab39bba),
	.w8(32'hbaa9d52f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf954d),
	.w1(32'h39d7ec2c),
	.w2(32'h3a53a477),
	.w3(32'hba9b8f82),
	.w4(32'hb93a48d5),
	.w5(32'h3987d817),
	.w6(32'h38fc33c2),
	.w7(32'hb8734cae),
	.w8(32'hb997f867),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3916e4cb),
	.w1(32'hbb41f364),
	.w2(32'hbb1c279d),
	.w3(32'hb768e4cf),
	.w4(32'hbb81cf2f),
	.w5(32'hbb1dbb0b),
	.w6(32'hbb2691f1),
	.w7(32'hbb0ba135),
	.w8(32'hbb0cd868),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa06ab5),
	.w1(32'h3a974317),
	.w2(32'h3a45d591),
	.w3(32'hbaacb942),
	.w4(32'h38a36590),
	.w5(32'hb815cc94),
	.w6(32'h3a582fe0),
	.w7(32'h3a66cfaf),
	.w8(32'hb9a8394d),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba127115),
	.w1(32'h3acfb635),
	.w2(32'hbb2620b8),
	.w3(32'h389cd432),
	.w4(32'hb8fe9f76),
	.w5(32'hba9b82e3),
	.w6(32'h3a5311ca),
	.w7(32'hbaa55041),
	.w8(32'hbac670c5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a4dd6),
	.w1(32'h3a0d533b),
	.w2(32'h3aa49283),
	.w3(32'hba979a79),
	.w4(32'hb9cb0cef),
	.w5(32'hb958daac),
	.w6(32'h3a2bb16d),
	.w7(32'h3a4b0790),
	.w8(32'hb93859fb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f6f0f7),
	.w1(32'hba988ea3),
	.w2(32'hbb088cfa),
	.w3(32'h39800c02),
	.w4(32'hba8b5b84),
	.w5(32'hbada71e3),
	.w6(32'hbae311f0),
	.w7(32'hbabecac7),
	.w8(32'hbb1f3384),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0d5c0),
	.w1(32'h3a97f316),
	.w2(32'h3a758fa2),
	.w3(32'hba6cbf36),
	.w4(32'h39d0e4d4),
	.w5(32'h3a36ec10),
	.w6(32'h39dcef3f),
	.w7(32'hb8d2a500),
	.w8(32'hba956cfa),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39545465),
	.w1(32'h3a19bc72),
	.w2(32'h3a969474),
	.w3(32'hb9a04ef3),
	.w4(32'hb966138f),
	.w5(32'h39e2f9aa),
	.w6(32'h39380360),
	.w7(32'hb88082a1),
	.w8(32'hb9a7cfd1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a275e7),
	.w1(32'h3a12b2d3),
	.w2(32'h3a04ce43),
	.w3(32'h38b1743a),
	.w4(32'h3982dd32),
	.w5(32'h39edc0d6),
	.w6(32'h39d87104),
	.w7(32'hb7f26a4a),
	.w8(32'hb9586feb),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391ec02c),
	.w1(32'h3a4cbbb7),
	.w2(32'h3a28ff18),
	.w3(32'h3924982c),
	.w4(32'h39e08005),
	.w5(32'h3a2a8141),
	.w6(32'h3a002daa),
	.w7(32'h38cf3488),
	.w8(32'h37fd5dd3),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3909fdeb),
	.w1(32'h3a9311bd),
	.w2(32'h3a891e2a),
	.w3(32'h39862285),
	.w4(32'hb8dcde66),
	.w5(32'hba0bff77),
	.w6(32'h3a5116ea),
	.w7(32'h39b06069),
	.w8(32'hb9ac435e),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0bb9b),
	.w1(32'h3ad92a51),
	.w2(32'h39cb3616),
	.w3(32'h39035ba2),
	.w4(32'h3a7029bf),
	.w5(32'h3a850f0d),
	.w6(32'h3a16b105),
	.w7(32'h3a83cab7),
	.w8(32'hb94c0abf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5fdcba),
	.w1(32'h3a1f2def),
	.w2(32'h3ad7cdc8),
	.w3(32'hb8b9aca2),
	.w4(32'h3909acef),
	.w5(32'hb8dd6720),
	.w6(32'h3a3dc3da),
	.w7(32'h3a4f97c4),
	.w8(32'hb934e413),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d6827),
	.w1(32'h3a5d1c8f),
	.w2(32'h3aadaeb8),
	.w3(32'hb92570b7),
	.w4(32'h39b62d88),
	.w5(32'h39edba61),
	.w6(32'hb887e8aa),
	.w7(32'h3a014af2),
	.w8(32'h38187a5d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3628796a),
	.w1(32'h38b0aee4),
	.w2(32'h3a087440),
	.w3(32'h3a0ffdad),
	.w4(32'hb9ee55fd),
	.w5(32'h37f71bf6),
	.w6(32'h3894a392),
	.w7(32'hb98fd808),
	.w8(32'hba53cd22),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3f1e2),
	.w1(32'h3a6ee7c2),
	.w2(32'h3a11688f),
	.w3(32'hb9f3a08e),
	.w4(32'h39679ce0),
	.w5(32'hb975af04),
	.w6(32'h3a9ac0ff),
	.w7(32'h3aabf7c2),
	.w8(32'h3ad5036b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a945f61),
	.w1(32'h3af6f01d),
	.w2(32'h3b5b1ff2),
	.w3(32'hba5c9efc),
	.w4(32'h3b2dcac4),
	.w5(32'h3b4b16f5),
	.w6(32'h3a9b3d16),
	.w7(32'h3a55c233),
	.w8(32'h3a808358),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a8630),
	.w1(32'hb9bec678),
	.w2(32'hb9851030),
	.w3(32'h3af01ae6),
	.w4(32'hbaa5c54d),
	.w5(32'hba92146b),
	.w6(32'hba8754e1),
	.w7(32'hbae2ef10),
	.w8(32'hbaacf40a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88959a),
	.w1(32'h3a5951fc),
	.w2(32'hbad65176),
	.w3(32'hba8ff258),
	.w4(32'hb9ba9783),
	.w5(32'hba22520a),
	.w6(32'hba515034),
	.w7(32'h38f94f51),
	.w8(32'hba08d15c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b523ec),
	.w1(32'hbabbdf35),
	.w2(32'hbb0477ab),
	.w3(32'h38c16c20),
	.w4(32'hb9f4bf3d),
	.w5(32'hba887677),
	.w6(32'hb92f05e9),
	.w7(32'hba15328a),
	.w8(32'hba0c1136),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule