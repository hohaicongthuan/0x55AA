module layer_10_featuremap_169(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc264fec),
	.w1(32'hbc156ed6),
	.w2(32'hbbe91e28),
	.w3(32'hbbb4a18d),
	.w4(32'hbc59830e),
	.w5(32'hbc3f5c59),
	.w6(32'hbc237739),
	.w7(32'hbc3148b7),
	.w8(32'hbb9614de),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9961d66),
	.w1(32'h3ae4511e),
	.w2(32'h3bed2f9f),
	.w3(32'hbc275b8f),
	.w4(32'hb9c76953),
	.w5(32'h3b3e1dae),
	.w6(32'hbb08eff2),
	.w7(32'h3b1410dd),
	.w8(32'h39a36384),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89a67c),
	.w1(32'hbaa034b3),
	.w2(32'h3b8f1122),
	.w3(32'h39adb3d2),
	.w4(32'hbb9c7c02),
	.w5(32'hbb8f52e2),
	.w6(32'hbb396c3b),
	.w7(32'h3a5b5506),
	.w8(32'h39e5827c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4474c0),
	.w1(32'hbb676c38),
	.w2(32'hbbed2a54),
	.w3(32'hbbd48c44),
	.w4(32'h3b9d06b1),
	.w5(32'h3bb35b52),
	.w6(32'hbb257b4e),
	.w7(32'hbb22f795),
	.w8(32'hbb1cc45a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2ba0c),
	.w1(32'hbb91d6f0),
	.w2(32'h3aee9913),
	.w3(32'h3c38de94),
	.w4(32'hbb85b581),
	.w5(32'h3af4e905),
	.w6(32'hbbcfe695),
	.w7(32'hbb7358ad),
	.w8(32'hbbc0cf0e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb955507),
	.w1(32'hbc89c0c1),
	.w2(32'hbc9d3475),
	.w3(32'hbbaad03f),
	.w4(32'hbc39f39c),
	.w5(32'hbc6a9136),
	.w6(32'hbc9d37cc),
	.w7(32'hbca6052a),
	.w8(32'hbc8a89d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ba058),
	.w1(32'hbaace47a),
	.w2(32'h3b902f42),
	.w3(32'hbc404d80),
	.w4(32'hbb776347),
	.w5(32'h3a7fe13c),
	.w6(32'hbba54d5f),
	.w7(32'hb8bfb5bb),
	.w8(32'hba990dd9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7eada1),
	.w1(32'h3b3c9b38),
	.w2(32'h38012f4b),
	.w3(32'hb88729db),
	.w4(32'h3bfeef99),
	.w5(32'h3ba53edc),
	.w6(32'h3ba1e3ac),
	.w7(32'h3b662ce0),
	.w8(32'h3bac0e07),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ded68),
	.w1(32'hbb77e5cb),
	.w2(32'hbb806db9),
	.w3(32'h3be09d87),
	.w4(32'hbb278a1a),
	.w5(32'hbb2cefa9),
	.w6(32'hbb7e04dc),
	.w7(32'hbb8b7f39),
	.w8(32'hbb3f0d2b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c0290),
	.w1(32'h3a1b20bc),
	.w2(32'h3bf07156),
	.w3(32'hbb0804ad),
	.w4(32'hbba1ac60),
	.w5(32'hb9c09406),
	.w6(32'hbb0f1a9b),
	.w7(32'h3a19fb62),
	.w8(32'hbb42fb47),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888396),
	.w1(32'hbb9a96ec),
	.w2(32'hbbf21c56),
	.w3(32'hbbaad791),
	.w4(32'hbb48289e),
	.w5(32'hbb1c39ab),
	.w6(32'hbb63d8f7),
	.w7(32'hbb725fcd),
	.w8(32'h39ac8b45),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1df3ca),
	.w1(32'hbc0e66d1),
	.w2(32'hbc111802),
	.w3(32'hbb25b2a5),
	.w4(32'hbba35d45),
	.w5(32'h3adf9bfd),
	.w6(32'hbc0b9b9b),
	.w7(32'hbc291785),
	.w8(32'hbbb4e8fe),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8043f3),
	.w1(32'hb9f3a4d5),
	.w2(32'h39ab4ec4),
	.w3(32'h3b7fc121),
	.w4(32'h3b1e3f0a),
	.w5(32'h3b29091c),
	.w6(32'h3b00da85),
	.w7(32'h3b04c2dd),
	.w8(32'h3b8ad5c1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c47f4),
	.w1(32'hbc1e128c),
	.w2(32'hbc12858c),
	.w3(32'h3b6c31a7),
	.w4(32'hbb8c82d0),
	.w5(32'hbb636f3e),
	.w6(32'hbbe8a6bd),
	.w7(32'hbc080a48),
	.w8(32'h39827ac8),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba872300),
	.w1(32'hba6711b8),
	.w2(32'hbb73de15),
	.w3(32'h3aee7029),
	.w4(32'h394c4619),
	.w5(32'h3c573e75),
	.w6(32'hbb5daaf4),
	.w7(32'hbb552a1c),
	.w8(32'hb9ff4a1a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa7bc5),
	.w1(32'hbbdc405b),
	.w2(32'hbb80e69e),
	.w3(32'h3b975ec7),
	.w4(32'hbb9f48f0),
	.w5(32'hbb10f810),
	.w6(32'hbbee6096),
	.w7(32'hbbddf928),
	.w8(32'hbb82516e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdbf96f),
	.w1(32'hbb294311),
	.w2(32'hbafd5cdd),
	.w3(32'hbb996c99),
	.w4(32'hba8e26f3),
	.w5(32'hba40ab59),
	.w6(32'hbaea19fc),
	.w7(32'hbaf4863b),
	.w8(32'h398dfbbe),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafbc3f),
	.w1(32'h3b998e19),
	.w2(32'h3c43b0c1),
	.w3(32'hba812edf),
	.w4(32'h3a4c2157),
	.w5(32'h3bbe9390),
	.w6(32'h3b53fc1f),
	.w7(32'h3c04e7a5),
	.w8(32'h3b8bd0b7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17982),
	.w1(32'hbacaaf3f),
	.w2(32'h3b844dcb),
	.w3(32'h3af20c05),
	.w4(32'hbab5646f),
	.w5(32'h3aea45cf),
	.w6(32'hbab5ff7b),
	.w7(32'h3aa37292),
	.w8(32'hb7cd6337),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba036e0f),
	.w1(32'hbb806e65),
	.w2(32'hbb5b7f3a),
	.w3(32'hba85a183),
	.w4(32'hbb3f4875),
	.w5(32'hbb32baec),
	.w6(32'hbb90e5da),
	.w7(32'hbb7e7042),
	.w8(32'hbb81bcc9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833567),
	.w1(32'h3b48e717),
	.w2(32'h3b3c5385),
	.w3(32'hbb25093e),
	.w4(32'h3bb82d4a),
	.w5(32'h3bb499ff),
	.w6(32'h3b853e5e),
	.w7(32'h3b3a31cf),
	.w8(32'h3b645b4d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2601cd),
	.w1(32'hbba12c09),
	.w2(32'h3b38446f),
	.w3(32'h3ba3c146),
	.w4(32'hbb5e673f),
	.w5(32'hbbc7b424),
	.w6(32'hbc45be23),
	.w7(32'hbb96d811),
	.w8(32'hbba22ffd),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f35e7a),
	.w1(32'h39b1bce7),
	.w2(32'h3ac0dd2b),
	.w3(32'hbb619b4e),
	.w4(32'hb8ec20be),
	.w5(32'hb8883ca3),
	.w6(32'h3b1f4137),
	.w7(32'h3b8e9a69),
	.w8(32'h3b290cff),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad30024),
	.w1(32'hbb2053c0),
	.w2(32'hbb67a396),
	.w3(32'h3aecbb64),
	.w4(32'h3b226cf0),
	.w5(32'h3b179e09),
	.w6(32'hbb142b94),
	.w7(32'hbb1e78f5),
	.w8(32'h3b3387c2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06b7d9),
	.w1(32'h3af1678a),
	.w2(32'hb9be8c77),
	.w3(32'h3ba19799),
	.w4(32'h3aa494b3),
	.w5(32'hba0f8410),
	.w6(32'hba0a76ed),
	.w7(32'h3ae08d0e),
	.w8(32'hbb10fa84),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb987e2c),
	.w1(32'hbb3bf54c),
	.w2(32'hbb35200a),
	.w3(32'hbb84140d),
	.w4(32'hba3fe46d),
	.w5(32'hbb73643c),
	.w6(32'h3964b0ef),
	.w7(32'h396bd794),
	.w8(32'h3a8803ff),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb077815),
	.w1(32'hbb491f34),
	.w2(32'hbad12ec1),
	.w3(32'hbbad9333),
	.w4(32'hbaa25919),
	.w5(32'hb9e28cd0),
	.w6(32'hbb695629),
	.w7(32'hbb293dd6),
	.w8(32'hbabca8a6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dfe5b),
	.w1(32'hbb91c232),
	.w2(32'hbb9f7d28),
	.w3(32'hbb47d742),
	.w4(32'hbb8f15d1),
	.w5(32'hbbd372c8),
	.w6(32'hbc16e511),
	.w7(32'hbbb2d04b),
	.w8(32'hbbf93e16),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc389fef),
	.w1(32'h3c061aa9),
	.w2(32'h3b145266),
	.w3(32'hbc07db82),
	.w4(32'h3bc8fc97),
	.w5(32'h39fad1fb),
	.w6(32'h3bdc7218),
	.w7(32'h3a9acb1d),
	.w8(32'h3a95e843),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e63bc),
	.w1(32'hbab628a2),
	.w2(32'hbb9e1d98),
	.w3(32'hbb5dd3e3),
	.w4(32'h3948eae8),
	.w5(32'hba46c933),
	.w6(32'hbb48baaa),
	.w7(32'hbb4e43b6),
	.w8(32'hbaddc044),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c5cf8),
	.w1(32'hba128fef),
	.w2(32'h38a3aa58),
	.w3(32'hbac6eb79),
	.w4(32'h398c8958),
	.w5(32'h39f70284),
	.w6(32'h38fa135d),
	.w7(32'h397be6d5),
	.w8(32'h39835e52),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce8557),
	.w1(32'hbabfda84),
	.w2(32'hbae76899),
	.w3(32'h38d22cc9),
	.w4(32'hb9016784),
	.w5(32'hb9db2783),
	.w6(32'hbaab1c41),
	.w7(32'hbabe731d),
	.w8(32'hba3f2cf2),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac95dfe),
	.w1(32'hbbbd886f),
	.w2(32'hbaf595e3),
	.w3(32'hb9996001),
	.w4(32'hbb74d9b1),
	.w5(32'hbae4d675),
	.w6(32'hbb79f6a9),
	.w7(32'h3a8211fa),
	.w8(32'h3b39425c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42bd17),
	.w1(32'hbb90781c),
	.w2(32'hbbb5fd6a),
	.w3(32'hbb84a536),
	.w4(32'hbbaacce6),
	.w5(32'hbb9f8ccd),
	.w6(32'hbb2a955f),
	.w7(32'hbb1ffee0),
	.w8(32'hbafe30dd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ed1ac),
	.w1(32'hbb911107),
	.w2(32'h3ba108f2),
	.w3(32'hbb00b9df),
	.w4(32'hbbf4099f),
	.w5(32'hbb3f2308),
	.w6(32'hbbc3c779),
	.w7(32'hbaa3122d),
	.w8(32'hbb8d56a2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39282db1),
	.w1(32'hbb7b1396),
	.w2(32'hbb90fad8),
	.w3(32'hbb6552d0),
	.w4(32'hbb0b2489),
	.w5(32'hbb494c43),
	.w6(32'hbb27baea),
	.w7(32'hbb3c6b06),
	.w8(32'hbb12a851),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a78a8),
	.w1(32'hbb0ccf16),
	.w2(32'hbb84180a),
	.w3(32'hbad00c14),
	.w4(32'hbb529a1c),
	.w5(32'hbba51256),
	.w6(32'hbb9229f8),
	.w7(32'hbb53e0ae),
	.w8(32'hbc01aa5d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a0ebc),
	.w1(32'h3b2597ad),
	.w2(32'h3bd60f5a),
	.w3(32'hbb8c5303),
	.w4(32'hbad9ee31),
	.w5(32'h3a83ff69),
	.w6(32'hbbbbc3be),
	.w7(32'h3a8e9d5c),
	.w8(32'hbabe5cfd),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4d6b11),
	.w1(32'hbbaea975),
	.w2(32'hbbd12977),
	.w3(32'hbad509aa),
	.w4(32'hba92d379),
	.w5(32'hbaa23151),
	.w6(32'hbc2ebaa3),
	.w7(32'hbbedba95),
	.w8(32'hbb453546),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9154af),
	.w1(32'hba8f1dd3),
	.w2(32'h3b23a388),
	.w3(32'hb9d551d6),
	.w4(32'hbb7cbde2),
	.w5(32'h3a93f670),
	.w6(32'hbacacb61),
	.w7(32'h3ad68193),
	.w8(32'h3a04a20b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcb8d5),
	.w1(32'hbb79838a),
	.w2(32'hbb51bed1),
	.w3(32'h3a922690),
	.w4(32'hbb2bcc9f),
	.w5(32'hba9ad0d5),
	.w6(32'hbaf91614),
	.w7(32'hbb06967d),
	.w8(32'hbabf3084),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a30b6),
	.w1(32'h3a9179a1),
	.w2(32'h3b665ae0),
	.w3(32'hb98d00ba),
	.w4(32'hba8cc7cd),
	.w5(32'h3b26ad14),
	.w6(32'h3af6488d),
	.w7(32'h3b7373e0),
	.w8(32'h3b3651b3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba28d9b),
	.w1(32'hb929fdd2),
	.w2(32'hba285964),
	.w3(32'h3a26c580),
	.w4(32'h3ab73d06),
	.w5(32'h3aa4ab88),
	.w6(32'h39df3ba9),
	.w7(32'h3a35141b),
	.w8(32'h3b334c9c),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaece326),
	.w1(32'h3a958baa),
	.w2(32'h3c3d4fe3),
	.w3(32'h3a9850bc),
	.w4(32'hba9290d0),
	.w5(32'h3bc6f4e5),
	.w6(32'hb98874d2),
	.w7(32'h3b3faa10),
	.w8(32'h3b8f099c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a37ff),
	.w1(32'h3b4d35a0),
	.w2(32'h3c13d7fc),
	.w3(32'h3b44b17e),
	.w4(32'hbb8c7234),
	.w5(32'hbb98b8c7),
	.w6(32'h3ba4689c),
	.w7(32'h3c2d66b1),
	.w8(32'h3bd31fe3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c405365),
	.w1(32'h3a1b1b36),
	.w2(32'h3baaa92b),
	.w3(32'hbaf10fcc),
	.w4(32'hbbce1d47),
	.w5(32'hbbef27da),
	.w6(32'hbbf25e98),
	.w7(32'h39704391),
	.w8(32'hbbfad94b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe41795),
	.w1(32'hbb358ded),
	.w2(32'hbb433b34),
	.w3(32'hbc2eb7b1),
	.w4(32'h3b537d06),
	.w5(32'h3c8e3214),
	.w6(32'hbbb530f9),
	.w7(32'hbbb37be9),
	.w8(32'hbb85be41),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf1f85),
	.w1(32'h396c0081),
	.w2(32'hb9c5c3e0),
	.w3(32'h3c67eb42),
	.w4(32'h39e94e55),
	.w5(32'hba982ed3),
	.w6(32'h3b8bca16),
	.w7(32'hb8d64915),
	.w8(32'h3a5fdefc),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a1c09),
	.w1(32'hbb35e8f2),
	.w2(32'hbb1efdae),
	.w3(32'hbb4f56de),
	.w4(32'hba866a14),
	.w5(32'hba71399b),
	.w6(32'hbb301def),
	.w7(32'hbb2f88ce),
	.w8(32'hba7b68e3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a266),
	.w1(32'h3b1566c6),
	.w2(32'hb8b1f90f),
	.w3(32'hba3c4c61),
	.w4(32'h3bce7eb7),
	.w5(32'h3b9a83fb),
	.w6(32'h3b84b1fe),
	.w7(32'h3b278962),
	.w8(32'h3bba424b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b630b3e),
	.w1(32'h3ba94f23),
	.w2(32'h3c08a828),
	.w3(32'h3bd71ea0),
	.w4(32'hba6db565),
	.w5(32'h391ca21d),
	.w6(32'h3ba904b8),
	.w7(32'h3b847141),
	.w8(32'hbaa3e3d7),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacee0e8),
	.w1(32'hbc821f55),
	.w2(32'hbc622573),
	.w3(32'hbbdba41e),
	.w4(32'hbc2e6e3c),
	.w5(32'hbb2dfa4c),
	.w6(32'hbc5439b5),
	.w7(32'hbc296ecb),
	.w8(32'hbb885f15),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1312a8),
	.w1(32'hbca191de),
	.w2(32'hbc9089f3),
	.w3(32'h3c58381b),
	.w4(32'hbc8fbd24),
	.w5(32'hbc88392c),
	.w6(32'hbca6c87d),
	.w7(32'hbc9ed384),
	.w8(32'hbca11a33),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3905d),
	.w1(32'hbc838231),
	.w2(32'hbc018ae1),
	.w3(32'hbc92e248),
	.w4(32'hbc701bea),
	.w5(32'hbc1db4d6),
	.w6(32'hbc8c463b),
	.w7(32'hbc2bf310),
	.w8(32'hbbae9664),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd94ec3),
	.w1(32'h3b4dee1e),
	.w2(32'h3bc6cead),
	.w3(32'hbc18053e),
	.w4(32'h3b40063f),
	.w5(32'h3b810600),
	.w6(32'h3b644111),
	.w7(32'h3b869c02),
	.w8(32'h3b3ebb1f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae39a26),
	.w1(32'hbb143459),
	.w2(32'h39e72238),
	.w3(32'h3ac168b7),
	.w4(32'h39475176),
	.w5(32'h3ae94cbc),
	.w6(32'hbaf7d70b),
	.w7(32'hba9e34a7),
	.w8(32'hbb195980),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3e599),
	.w1(32'h3bbfd642),
	.w2(32'h3c67aada),
	.w3(32'hb9e17797),
	.w4(32'h39476b1d),
	.w5(32'h3b51e9c0),
	.w6(32'h3ba0daa5),
	.w7(32'h3c2d443a),
	.w8(32'h3bd54e0c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d1cfa),
	.w1(32'h3b8dd206),
	.w2(32'h3bbfd8b4),
	.w3(32'h3b0a0539),
	.w4(32'h3b06f65e),
	.w5(32'h3b1b06ce),
	.w6(32'hbaf89600),
	.w7(32'h3a6c0183),
	.w8(32'hbb56c230),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3497),
	.w1(32'hba11cd0d),
	.w2(32'h3b77e1aa),
	.w3(32'hbbc41883),
	.w4(32'hbaf029ba),
	.w5(32'h3a5df1e8),
	.w6(32'hba3a49b8),
	.w7(32'h3abac5ad),
	.w8(32'hbabf7a01),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c441e),
	.w1(32'hbbe57e35),
	.w2(32'hbbe3ace7),
	.w3(32'h39a2aabe),
	.w4(32'hbb36bf36),
	.w5(32'hbb0e443e),
	.w6(32'hbbd54f3a),
	.w7(32'hbbceeff1),
	.w8(32'hbacef93d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c4493),
	.w1(32'hba9cfbd3),
	.w2(32'h3b86ddc0),
	.w3(32'h3a3c5c76),
	.w4(32'hbb08bcdd),
	.w5(32'h3b054497),
	.w6(32'hbb296b58),
	.w7(32'h3a2b5ea7),
	.w8(32'hb993cd5a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981e578),
	.w1(32'hbb90a501),
	.w2(32'hbac914c9),
	.w3(32'hbb6650d7),
	.w4(32'hbaa37912),
	.w5(32'h3a553d67),
	.w6(32'hbac839ae),
	.w7(32'h3a38f7ab),
	.w8(32'h3bdb4fd2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b72eba1),
	.w1(32'hbb42e2db),
	.w2(32'h3b5d0038),
	.w3(32'h3b404f08),
	.w4(32'hbbbdeabe),
	.w5(32'hbb0f43f4),
	.w6(32'h3b53af9f),
	.w7(32'h3c0cff04),
	.w8(32'hba843ad3),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093d7b),
	.w1(32'h3a0fcaf4),
	.w2(32'h3bab6326),
	.w3(32'hbbb91965),
	.w4(32'hbb126a3c),
	.w5(32'h3a210047),
	.w6(32'hbb23997c),
	.w7(32'hb8ee71e0),
	.w8(32'hbac4ba56),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8387ea),
	.w1(32'h39ea225b),
	.w2(32'h391c99e2),
	.w3(32'hb9656704),
	.w4(32'hba7eff8d),
	.w5(32'hb9b6ae0c),
	.w6(32'hbb016748),
	.w7(32'h37aee320),
	.w8(32'hbb0e0142),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb812c4c),
	.w1(32'hbb24921f),
	.w2(32'hbb107cce),
	.w3(32'hbbb89dc8),
	.w4(32'hbb2d1dbf),
	.w5(32'hbbbc2d4e),
	.w6(32'hbbbe02e3),
	.w7(32'hbba0b614),
	.w8(32'hbbc554ee),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe851e),
	.w1(32'hbc120e78),
	.w2(32'hbb13c2f9),
	.w3(32'hbbaf9e2a),
	.w4(32'hbbc9fb9c),
	.w5(32'hbac935d0),
	.w6(32'hbbbcd3cb),
	.w7(32'hbbb9a043),
	.w8(32'hba3a81cb),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d18ae),
	.w1(32'hb9a91699),
	.w2(32'h3a23e229),
	.w3(32'hbb13b4a8),
	.w4(32'h3b2722c1),
	.w5(32'h3b1c88bc),
	.w6(32'h3a8b7f4f),
	.w7(32'h3b6ff90b),
	.w8(32'h3bab6c3e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba309986),
	.w1(32'hbc06a872),
	.w2(32'hbbaa7a40),
	.w3(32'h3ad1b059),
	.w4(32'hbbc5e9c0),
	.w5(32'hbb6047ff),
	.w6(32'hbc1319c1),
	.w7(32'hbc0601a2),
	.w8(32'hbb95addf),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac41a),
	.w1(32'h3c1979f5),
	.w2(32'h3bebf633),
	.w3(32'hbb9f6bf7),
	.w4(32'h3a16d381),
	.w5(32'hbb7c7767),
	.w6(32'h39f3dc5a),
	.w7(32'h3b7b41dd),
	.w8(32'hbbb80fc2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d07a8),
	.w1(32'hbac5c635),
	.w2(32'h3b6da65d),
	.w3(32'hbc575b77),
	.w4(32'hbb5821ac),
	.w5(32'hb8276cf9),
	.w6(32'hbb80a6c6),
	.w7(32'hba26da64),
	.w8(32'hbb186f27),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f55d3),
	.w1(32'hbb855ef2),
	.w2(32'hbb993141),
	.w3(32'hb9b4a227),
	.w4(32'hba0b6f28),
	.w5(32'hbb028c20),
	.w6(32'hbb7f0cc6),
	.w7(32'hbb97077d),
	.w8(32'hbb73ab1e),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98cb04),
	.w1(32'hbbed5f6f),
	.w2(32'hbbf57f8c),
	.w3(32'hbab232b6),
	.w4(32'hbb58f929),
	.w5(32'hbb383607),
	.w6(32'hbbf1c9ef),
	.w7(32'hbbeee95d),
	.w8(32'hbb747971),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d353e),
	.w1(32'hbb82e017),
	.w2(32'hbb60928b),
	.w3(32'hb8289e67),
	.w4(32'hbb03bdad),
	.w5(32'hbad90d85),
	.w6(32'hbb479f62),
	.w7(32'hbb42a373),
	.w8(32'hbaee600e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b5241),
	.w1(32'hbad054a2),
	.w2(32'h39f54fa3),
	.w3(32'hbb030b3a),
	.w4(32'hbb2a1d54),
	.w5(32'h39a66fb9),
	.w6(32'hba8847e9),
	.w7(32'hbaa549e9),
	.w8(32'hbb37d46f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a105096),
	.w1(32'hbba16018),
	.w2(32'hbbbd5cd1),
	.w3(32'hbab10b70),
	.w4(32'hb99464a4),
	.w5(32'h3c37d223),
	.w6(32'h3b3350b3),
	.w7(32'h3b25f12f),
	.w8(32'h3b8cefc5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c085f1a),
	.w1(32'hba0bb20a),
	.w2(32'hbbb823d4),
	.w3(32'h3c4c5891),
	.w4(32'h3bc87577),
	.w5(32'h3a2cbbfa),
	.w6(32'h3b03ba4f),
	.w7(32'hba7f07ec),
	.w8(32'h3b659e6a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bd3b56),
	.w1(32'hba17d8ea),
	.w2(32'h3b7645ef),
	.w3(32'h3bab908f),
	.w4(32'hb89ac13d),
	.w5(32'h3ace043a),
	.w6(32'hbab95ac6),
	.w7(32'h3b1a5c67),
	.w8(32'hbaf4950f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0d19b),
	.w1(32'h3bb5813c),
	.w2(32'h3bb9b7ed),
	.w3(32'hbae11864),
	.w4(32'h3b80f553),
	.w5(32'h3b74f2bf),
	.w6(32'h3ba543bb),
	.w7(32'h3b755c75),
	.w8(32'h3b8b21c1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aed2704),
	.w1(32'h3a390b7a),
	.w2(32'h3a852994),
	.w3(32'hba670806),
	.w4(32'h3b491868),
	.w5(32'h3b11d3a2),
	.w6(32'h3b1bb2a8),
	.w7(32'h3a0e19e2),
	.w8(32'h3ad90db3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25c8eb),
	.w1(32'h3b0f3d73),
	.w2(32'h3b8a78b0),
	.w3(32'h3ac2473d),
	.w4(32'h3ae6656f),
	.w5(32'h3b55a058),
	.w6(32'h3b21705a),
	.w7(32'h3b3520c4),
	.w8(32'h3b5acd46),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8d90),
	.w1(32'h3b067edd),
	.w2(32'h3c044065),
	.w3(32'h3b4348f5),
	.w4(32'h394ba6bd),
	.w5(32'h3ba3c0bb),
	.w6(32'h3b025a71),
	.w7(32'h3bb1cf62),
	.w8(32'h3c0230b8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c352ce6),
	.w1(32'hba87c247),
	.w2(32'hb9129736),
	.w3(32'h3bde0d8a),
	.w4(32'hbab2c69a),
	.w5(32'hba6f463a),
	.w6(32'hba898f7d),
	.w7(32'hb9b22e7b),
	.w8(32'hbae1ce8a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8dc69),
	.w1(32'hb9ce17e2),
	.w2(32'h3b38255d),
	.w3(32'hbb044016),
	.w4(32'hbaf49b90),
	.w5(32'h38aeef47),
	.w6(32'hbb07474b),
	.w7(32'h37d2ab44),
	.w8(32'hba775ded),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8029b4),
	.w1(32'h38e926b7),
	.w2(32'h39f06c1c),
	.w3(32'h3a163e4e),
	.w4(32'h39901566),
	.w5(32'hb924c56c),
	.w6(32'h3b80daf9),
	.w7(32'h3a0e48eb),
	.w8(32'h3b53ecca),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1d598),
	.w1(32'h3c0f9076),
	.w2(32'h3c687dbe),
	.w3(32'h3af1a2e1),
	.w4(32'h3bddf984),
	.w5(32'h3c2070d3),
	.w6(32'h3bc2ff8d),
	.w7(32'h3c1b40fb),
	.w8(32'h3c246372),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6bfb5a),
	.w1(32'hbc17f9a6),
	.w2(32'hbba19f51),
	.w3(32'h3c1b6f73),
	.w4(32'hbc02d369),
	.w5(32'hbbbc73fa),
	.w6(32'hbbd34553),
	.w7(32'hbb8b8470),
	.w8(32'hbbaced2f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba533a2c),
	.w1(32'hba35b20f),
	.w2(32'hba1a74f6),
	.w3(32'hbbb66e90),
	.w4(32'h3941ec24),
	.w5(32'h39626294),
	.w6(32'h399e653c),
	.w7(32'hb834bffc),
	.w8(32'h3808d744),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f6fe7),
	.w1(32'h3b6c17db),
	.w2(32'h3bcc9d42),
	.w3(32'h39d5c49a),
	.w4(32'h3b1c99a2),
	.w5(32'h3b7672e4),
	.w6(32'h3b03ba2c),
	.w7(32'h3b93db04),
	.w8(32'h3b65dd98),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c4e26),
	.w1(32'h3aa5230c),
	.w2(32'h3b523a76),
	.w3(32'h3ad7b1c9),
	.w4(32'h3b5aa39e),
	.w5(32'h3baa546d),
	.w6(32'h3b2e70f6),
	.w7(32'h3b26112c),
	.w8(32'h3b771c8a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15ac06),
	.w1(32'hbac8efcb),
	.w2(32'hbb24bd0a),
	.w3(32'h3b85746f),
	.w4(32'hb9ade126),
	.w5(32'hba8fd452),
	.w6(32'hba9cae82),
	.w7(32'hba4b61bc),
	.w8(32'hb8322ce2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2fb34),
	.w1(32'h3c0544b8),
	.w2(32'h3c6fd2c5),
	.w3(32'hba9e8773),
	.w4(32'h3b0e7a95),
	.w5(32'h3bba1bc8),
	.w6(32'h3bcc6925),
	.w7(32'h3c0d734d),
	.w8(32'h3b8f6eda),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f9255),
	.w1(32'hbb8e4df9),
	.w2(32'hbb09f344),
	.w3(32'h3ae5a18a),
	.w4(32'hbbaa4d9e),
	.w5(32'hbb65955c),
	.w6(32'hbbd600e0),
	.w7(32'hbb92ab18),
	.w8(32'hbbb38922),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc13b),
	.w1(32'h3bb02651),
	.w2(32'h3c14d62f),
	.w3(32'hbbe061bd),
	.w4(32'h3b7aeae7),
	.w5(32'h3bfa6eb1),
	.w6(32'h3b948b4f),
	.w7(32'h3bb862db),
	.w8(32'h3b9e9369),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b196874),
	.w1(32'hbab9e678),
	.w2(32'h3ae9e2bd),
	.w3(32'h3a6f9019),
	.w4(32'hbb77158c),
	.w5(32'hbb5cb2b5),
	.w6(32'hbb8436e8),
	.w7(32'hbb36fad5),
	.w8(32'hbb5222bf),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31e64d),
	.w1(32'hbc6436ce),
	.w2(32'hbc44b409),
	.w3(32'hbbaea08a),
	.w4(32'hbc367f61),
	.w5(32'hbc3d4c6f),
	.w6(32'hbcc0c901),
	.w7(32'hbc8f0470),
	.w8(32'hbc85bc59),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6dfff1),
	.w1(32'hb9d125c6),
	.w2(32'h378d5f02),
	.w3(32'hbc56ca3f),
	.w4(32'hbac0cc2d),
	.w5(32'hbb102a73),
	.w6(32'h3aed56a2),
	.w7(32'h3b599e4e),
	.w8(32'h3b39442a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b546e82),
	.w1(32'h39fdd852),
	.w2(32'hbb475cdd),
	.w3(32'h3ba06057),
	.w4(32'h3b1dd016),
	.w5(32'hb834586a),
	.w6(32'h39c1a9a0),
	.w7(32'hbaf4ee65),
	.w8(32'hbb14bf74),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4af8aa),
	.w1(32'hba20581a),
	.w2(32'h3bd8015e),
	.w3(32'hbacb3c86),
	.w4(32'hbae6c9d5),
	.w5(32'h3b51a9ea),
	.w6(32'h3aff9cda),
	.w7(32'h3bb8e4c4),
	.w8(32'h3b8521d6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f930),
	.w1(32'hbbc060e1),
	.w2(32'hbc4180e5),
	.w3(32'h3b7eea4c),
	.w4(32'hbbf8cd24),
	.w5(32'hbc54df64),
	.w6(32'hbc0cf567),
	.w7(32'hbc2897fc),
	.w8(32'hbc739a7a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4845ff),
	.w1(32'h3b9303a8),
	.w2(32'h3a3c56f4),
	.w3(32'hbc26d0ae),
	.w4(32'h381c4871),
	.w5(32'hbb981fed),
	.w6(32'hba950e36),
	.w7(32'h3b79e406),
	.w8(32'h3a4eab51),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6ae30),
	.w1(32'h385ac1ea),
	.w2(32'h3c0040e2),
	.w3(32'hbbd4b569),
	.w4(32'hbb087761),
	.w5(32'hbb23eb2f),
	.w6(32'hbbd7c8fd),
	.w7(32'h3bce292d),
	.w8(32'hbabb5953),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93aa5a6),
	.w1(32'h37a24721),
	.w2(32'hbc11114d),
	.w3(32'hbbaa8a10),
	.w4(32'h3c08b6bf),
	.w5(32'hb907463d),
	.w6(32'h3b181532),
	.w7(32'hbb72c675),
	.w8(32'h3b93a65b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9576b2),
	.w1(32'hbb5d0ce0),
	.w2(32'hbb8c7b84),
	.w3(32'h3c0ddb4e),
	.w4(32'h3aa58ac6),
	.w5(32'hb9dd6383),
	.w6(32'hbb8d79d0),
	.w7(32'hbbb30533),
	.w8(32'hbb6df9ed),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72f31),
	.w1(32'h3b01feff),
	.w2(32'hbbd0ea6a),
	.w3(32'hbb0e1a12),
	.w4(32'h3b8bb9c4),
	.w5(32'hbb15d4dd),
	.w6(32'h3adac3d6),
	.w7(32'hbaeabf40),
	.w8(32'hba0d6d02),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d6e34),
	.w1(32'hbb220c56),
	.w2(32'hbb0aae60),
	.w3(32'h3ba8ce07),
	.w4(32'h39191099),
	.w5(32'hba189392),
	.w6(32'hbaf27e93),
	.w7(32'hbaacab55),
	.w8(32'hb9b18642),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391c112d),
	.w1(32'hba52f54f),
	.w2(32'h3b26c63c),
	.w3(32'h3a9f5ea4),
	.w4(32'hbb88c79c),
	.w5(32'hbb99e218),
	.w6(32'hbaa25535),
	.w7(32'hba175c6d),
	.w8(32'hbb09a8d0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c464),
	.w1(32'hbb0d5fb5),
	.w2(32'hbabb06b8),
	.w3(32'hbbaa8a8e),
	.w4(32'hb9165c21),
	.w5(32'h39891687),
	.w6(32'h390f7f1d),
	.w7(32'hb96e0bb0),
	.w8(32'h3a8e79bc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab550ab),
	.w1(32'hba0bd434),
	.w2(32'hbb6a44d9),
	.w3(32'h3980b211),
	.w4(32'h3b99cb32),
	.w5(32'h3ad6a6f8),
	.w6(32'h3ad6ccf6),
	.w7(32'hba4a526c),
	.w8(32'h3b84c9fb),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961c95d),
	.w1(32'hbaf1faaf),
	.w2(32'h3b3b9299),
	.w3(32'h3b81ca01),
	.w4(32'hbbcf9d8b),
	.w5(32'hbb46dc1e),
	.w6(32'hbb0bb521),
	.w7(32'h3936ee9f),
	.w8(32'hbb15d138),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e67b9),
	.w1(32'hbc0b7ef0),
	.w2(32'hbc12a276),
	.w3(32'hbbbfa577),
	.w4(32'hbbd22edb),
	.w5(32'hbbaac436),
	.w6(32'hbc3133e0),
	.w7(32'hbc1e8874),
	.w8(32'hbbfb8559),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3b7cd),
	.w1(32'hbc792352),
	.w2(32'hbbd434c1),
	.w3(32'hbb04b12a),
	.w4(32'hbc367274),
	.w5(32'hbbd4fe31),
	.w6(32'hbbf83398),
	.w7(32'hbb0f2c42),
	.w8(32'h3c17d10e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e8d1e),
	.w1(32'hbc2d33ff),
	.w2(32'hbc47dd85),
	.w3(32'h3c139b6a),
	.w4(32'hbc071fa9),
	.w5(32'hbc10bde3),
	.w6(32'hbc381d2f),
	.w7(32'hbc3adfc1),
	.w8(32'hbc2f0360),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c9aab),
	.w1(32'hbb0233e4),
	.w2(32'h3b990527),
	.w3(32'hbc134c27),
	.w4(32'hbb8a3068),
	.w5(32'h3ab70406),
	.w6(32'hba94a5f8),
	.w7(32'hba2db705),
	.w8(32'hba875fef),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9deed51),
	.w1(32'hba812504),
	.w2(32'h3b384300),
	.w3(32'hbb9674df),
	.w4(32'h3ad2bf8d),
	.w5(32'h3b8753f0),
	.w6(32'h3af3715f),
	.w7(32'h3b692ef2),
	.w8(32'h3bf94f2a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10b478),
	.w1(32'h387d2476),
	.w2(32'hbbb59ec2),
	.w3(32'h3bd6427f),
	.w4(32'h3be27c0c),
	.w5(32'h3aba43d1),
	.w6(32'h3ac9dc26),
	.w7(32'hbb081721),
	.w8(32'h3b88390a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58719f),
	.w1(32'hbadd36c6),
	.w2(32'hbb71a564),
	.w3(32'h3bcb0e55),
	.w4(32'h3b822229),
	.w5(32'h3b11a1b2),
	.w6(32'hbb0ed644),
	.w7(32'hbb540477),
	.w8(32'h3a4c1fa7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3e60e4),
	.w1(32'hbb319a35),
	.w2(32'hbba5f44c),
	.w3(32'h3b6eba36),
	.w4(32'h3b5aa066),
	.w5(32'h3aa4b885),
	.w6(32'hbb3509cb),
	.w7(32'hbb9784d5),
	.w8(32'h39b5c1a2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac23bcd),
	.w1(32'hbbf89c8b),
	.w2(32'hbb2930c5),
	.w3(32'h3b561e92),
	.w4(32'hbc0b5ccf),
	.w5(32'hbc180723),
	.w6(32'hbc04ba08),
	.w7(32'hbaf85b64),
	.w8(32'h3b028e2f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a487d79),
	.w1(32'hbb09bf48),
	.w2(32'hba42a363),
	.w3(32'hbbc5001c),
	.w4(32'hbba239d3),
	.w5(32'hbbd67c31),
	.w6(32'hbbc9d28b),
	.w7(32'hbb87e81b),
	.w8(32'hbbb931b5),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc059fa8),
	.w1(32'hbc210b0c),
	.w2(32'hbc0ec0ac),
	.w3(32'hbc16a916),
	.w4(32'hbbf6fbd4),
	.w5(32'hbc0487f5),
	.w6(32'hbc39f3cb),
	.w7(32'hbc251edf),
	.w8(32'hbc23574a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21c3c9),
	.w1(32'hbc45bb03),
	.w2(32'hbc28ee85),
	.w3(32'hbc13a113),
	.w4(32'hbc2d9cdb),
	.w5(32'hbc27980e),
	.w6(32'hbc42236b),
	.w7(32'hbc35b4ea),
	.w8(32'hbc3760d4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41f6e5),
	.w1(32'hbb0b5671),
	.w2(32'hbb8338ae),
	.w3(32'hbc2c83d2),
	.w4(32'h3af97ddb),
	.w5(32'h3a9597e6),
	.w6(32'hbb8443d0),
	.w7(32'hbb3ce6b4),
	.w8(32'h3af097d2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a9d75),
	.w1(32'hba0bba63),
	.w2(32'h3bbc453c),
	.w3(32'h3b671471),
	.w4(32'hbbf42c24),
	.w5(32'hbc1bb197),
	.w6(32'hbbb55100),
	.w7(32'h3b4b91ad),
	.w8(32'hba41c19a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fae4bb),
	.w1(32'hbcd46083),
	.w2(32'hbcc499c8),
	.w3(32'hbbea3c61),
	.w4(32'hbcc144c3),
	.w5(32'hbcbd18be),
	.w6(32'hbce083b5),
	.w7(32'hbcdb7351),
	.w8(32'hbcddda6f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd689fc),
	.w1(32'hbb9ccd04),
	.w2(32'hbbabbdb9),
	.w3(32'hbccde396),
	.w4(32'hbb598ce1),
	.w5(32'hbb8577fd),
	.w6(32'hbb6d1b61),
	.w7(32'hbb99f4af),
	.w8(32'hbb8d44c0),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb50c65),
	.w1(32'h37b0457d),
	.w2(32'h380590df),
	.w3(32'hbb8d6699),
	.w4(32'hb73f6548),
	.w5(32'h376ee243),
	.w6(32'hb88c2063),
	.w7(32'hb61b4895),
	.w8(32'h37e48a19),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b021936),
	.w1(32'h39a57119),
	.w2(32'hba7479c9),
	.w3(32'h3b3c9ce3),
	.w4(32'h3a6c1c65),
	.w5(32'h3aa553bd),
	.w6(32'hb9ab9380),
	.w7(32'h3a2b94f1),
	.w8(32'h3a9c7d3b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd60e1),
	.w1(32'hba9f4bfa),
	.w2(32'h3a525b5d),
	.w3(32'hba152a8b),
	.w4(32'hba4e4bbc),
	.w5(32'h3a85989e),
	.w6(32'hb9326265),
	.w7(32'h3808e339),
	.w8(32'h3abdeca5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dea5f5),
	.w1(32'hb93a5171),
	.w2(32'h38417a42),
	.w3(32'hb938c3df),
	.w4(32'hb941674c),
	.w5(32'h38a0726f),
	.w6(32'hb8cc4095),
	.w7(32'hb8fb546d),
	.w8(32'h37f9e9d7),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec4289),
	.w1(32'h3976c621),
	.w2(32'h39d10d45),
	.w3(32'hb8958597),
	.w4(32'h391e369e),
	.w5(32'h393e7858),
	.w6(32'hb9903b12),
	.w7(32'h39ad2c08),
	.w8(32'h39ad0745),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d73173),
	.w1(32'h3902c83f),
	.w2(32'hb8af5d7f),
	.w3(32'hb928d6e5),
	.w4(32'h391ec316),
	.w5(32'hb8b00d2f),
	.w6(32'hb936648c),
	.w7(32'hb7f40634),
	.w8(32'hb8bc0882),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9687fae),
	.w1(32'h389d6cf2),
	.w2(32'h3a669486),
	.w3(32'hb9a58d2e),
	.w4(32'h378af0ef),
	.w5(32'h3a4c6000),
	.w6(32'hb964d663),
	.w7(32'h396f0a0d),
	.w8(32'h3a1559a8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f63f68),
	.w1(32'h39a2a808),
	.w2(32'h3abc1305),
	.w3(32'hba9b3f50),
	.w4(32'hb9686c48),
	.w5(32'h3a5338a4),
	.w6(32'hba8f448a),
	.w7(32'hba24628c),
	.w8(32'h3911b629),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cfe38),
	.w1(32'hbad0295a),
	.w2(32'h3993fae0),
	.w3(32'hb9816c9c),
	.w4(32'hba0e8450),
	.w5(32'h3a2ee283),
	.w6(32'h3a11ed03),
	.w7(32'h388b7b21),
	.w8(32'h3ad15944),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a60bdb),
	.w1(32'h3a0c0811),
	.w2(32'hb9319167),
	.w3(32'hb9b86041),
	.w4(32'h39cb9b77),
	.w5(32'hb8086431),
	.w6(32'hba068230),
	.w7(32'h395b83f3),
	.w8(32'hb8f4c29f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37aa7e14),
	.w1(32'hb9250246),
	.w2(32'h3a0625e0),
	.w3(32'h391477d1),
	.w4(32'h38e67a29),
	.w5(32'h3a2503e7),
	.w6(32'hb9ec481a),
	.w7(32'hb93b9673),
	.w8(32'h39a640a4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3680c2ad),
	.w1(32'hba62b0c9),
	.w2(32'hb932b99d),
	.w3(32'hb7eb6d00),
	.w4(32'hba05b0b0),
	.w5(32'h38ffcfb9),
	.w6(32'h38b2054a),
	.w7(32'hb8d7ef76),
	.w8(32'h3a302bed),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921742c),
	.w1(32'h39fe8214),
	.w2(32'hba2e8fcf),
	.w3(32'h389cc17b),
	.w4(32'h3950e874),
	.w5(32'hba2b6619),
	.w6(32'hba0c073f),
	.w7(32'h388dde64),
	.w8(32'hb9f3a776),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cb1d54),
	.w1(32'hb9be532e),
	.w2(32'h39d601ba),
	.w3(32'hb9a28013),
	.w4(32'hb9c6ded3),
	.w5(32'h396e282b),
	.w6(32'h38d9b261),
	.w7(32'h38c8facf),
	.w8(32'h3a09a9da),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8008b93),
	.w1(32'h388c33f2),
	.w2(32'h377c1a78),
	.w3(32'h37f5f68b),
	.w4(32'h38d63c29),
	.w5(32'h38a9482c),
	.w6(32'hb811dfcf),
	.w7(32'h38b9ae1b),
	.w8(32'h38c78104),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54d33a),
	.w1(32'h3a5afc07),
	.w2(32'hb881f829),
	.w3(32'hbae346d6),
	.w4(32'h3ae93f2d),
	.w5(32'h3a85e5ec),
	.w6(32'hbb120a58),
	.w7(32'h3aaad980),
	.w8(32'h3a678352),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94971a4),
	.w1(32'h393bf0f2),
	.w2(32'h3a01f4f3),
	.w3(32'hb946cc60),
	.w4(32'hb92b0259),
	.w5(32'h39b8ee66),
	.w6(32'hb91ff4d5),
	.w7(32'h39ceb888),
	.w8(32'h399d0345),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885b105),
	.w1(32'hb636ae02),
	.w2(32'h3880ffbc),
	.w3(32'hb70c1d2a),
	.w4(32'hb581eab4),
	.w5(32'h38a6e358),
	.w6(32'hb84e5b1a),
	.w7(32'h382c3410),
	.w8(32'h38e2f2a1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8232068),
	.w1(32'hb818f1bf),
	.w2(32'hb8917b4a),
	.w3(32'h3519f68a),
	.w4(32'hb7c7cfb7),
	.w5(32'hb7fc4e4a),
	.w6(32'hb5c2bea0),
	.w7(32'h36e50a98),
	.w8(32'hb6ebee40),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932b29a),
	.w1(32'hb9cf09f5),
	.w2(32'hba2bdf9d),
	.w3(32'hb8306629),
	.w4(32'hb9493325),
	.w5(32'hba2832e3),
	.w6(32'h36d4a39c),
	.w7(32'hb8e19aa4),
	.w8(32'hb9e25a83),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3912a41e),
	.w1(32'h39f1c211),
	.w2(32'hb9d9a470),
	.w3(32'hba1b08a2),
	.w4(32'hb6b1e0ca),
	.w5(32'hba1abf5e),
	.w6(32'hb95703fa),
	.w7(32'h39b96192),
	.w8(32'hb9a9af0d),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994c2e6),
	.w1(32'hb9a4c53f),
	.w2(32'h37e439d9),
	.w3(32'hb8136061),
	.w4(32'h37fc769f),
	.w5(32'h39c8849d),
	.w6(32'hb8ec71e4),
	.w7(32'h39558473),
	.w8(32'h3a04a844),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367861dd),
	.w1(32'h37416ff9),
	.w2(32'h3682eba9),
	.w3(32'h35d4d333),
	.w4(32'h3622372f),
	.w5(32'hb728041b),
	.w6(32'h374e0c68),
	.w7(32'h36ebd38d),
	.w8(32'h361229c2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9151fb4),
	.w1(32'hb9f01aab),
	.w2(32'h39f68fdb),
	.w3(32'hb9c0e01a),
	.w4(32'hb9a2cacb),
	.w5(32'h3a22ff84),
	.w6(32'h39705ca0),
	.w7(32'h39e1c7b4),
	.w8(32'h3a5fedde),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90331c6),
	.w1(32'h39901c2d),
	.w2(32'h39f81e54),
	.w3(32'hb7758752),
	.w4(32'h39ef2d9e),
	.w5(32'h39f46b66),
	.w6(32'h384d48d6),
	.w7(32'h39c78a12),
	.w8(32'h3a09c7db),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a166a2f),
	.w1(32'hba2b1942),
	.w2(32'hba43c7ed),
	.w3(32'h390d58ea),
	.w4(32'hb9fb1953),
	.w5(32'hb9874140),
	.w6(32'h386d4db4),
	.w7(32'hb9817ef0),
	.w8(32'h391fde62),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb409f67),
	.w1(32'h3a3636a6),
	.w2(32'h3ac90d9d),
	.w3(32'hbb25fc69),
	.w4(32'hb8d4670f),
	.w5(32'h39b8a6b4),
	.w6(32'hbb164388),
	.w7(32'hb9cd0dd8),
	.w8(32'h3afa60d2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b29914),
	.w1(32'h392e9740),
	.w2(32'h39cfac07),
	.w3(32'hb99a2acb),
	.w4(32'h3908720e),
	.w5(32'h3a04deec),
	.w6(32'hba1dcc27),
	.w7(32'h38722f51),
	.w8(32'h39caaa9a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983d60b),
	.w1(32'hb981d898),
	.w2(32'h390d0dbd),
	.w3(32'hb90e9cba),
	.w4(32'h38f8149d),
	.w5(32'hb75ddbc9),
	.w6(32'hb906d190),
	.w7(32'hb952b410),
	.w8(32'hb8fcd58d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e7ef4c),
	.w1(32'h390561b9),
	.w2(32'hb827f0f3),
	.w3(32'h3987f0f4),
	.w4(32'h39e5b117),
	.w5(32'hb92c756b),
	.w6(32'h37d9ddab),
	.w7(32'h39e34a51),
	.w8(32'h38cf2d3f),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb9a61),
	.w1(32'h3979ac50),
	.w2(32'hb9287f51),
	.w3(32'hba144476),
	.w4(32'hb8feeee5),
	.w5(32'hb96a9a37),
	.w6(32'hba1586d5),
	.w7(32'hb95ad451),
	.w8(32'hb9825695),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a853d6),
	.w1(32'h3982daf9),
	.w2(32'hb923a0e9),
	.w3(32'hb9b8f659),
	.w4(32'h391b91bb),
	.w5(32'hb947ffc8),
	.w6(32'hb9d78dcd),
	.w7(32'h38a93d5b),
	.w8(32'hb9514c50),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb889b8c4),
	.w1(32'hb99d1d32),
	.w2(32'hb9cdb326),
	.w3(32'h378d7178),
	.w4(32'hb96a8dc2),
	.w5(32'hb9549177),
	.w6(32'hb78173bb),
	.w7(32'hb8aca7c4),
	.w8(32'hb910d792),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3744be7c),
	.w1(32'h382f1962),
	.w2(32'h381ec6dc),
	.w3(32'h37ebf00c),
	.w4(32'h388f5f2d),
	.w5(32'h38198bf3),
	.w6(32'hb6ad423d),
	.w7(32'h3884b3d2),
	.w8(32'h37fdcf88),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84f5163),
	.w1(32'hb9ed79b5),
	.w2(32'h39630b33),
	.w3(32'hb9443f64),
	.w4(32'hb98f09cb),
	.w5(32'h39f7dc57),
	.w6(32'hb9763c17),
	.w7(32'h386f8928),
	.w8(32'h3a235ca7),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c15b25),
	.w1(32'hb9d4619f),
	.w2(32'hba440cc2),
	.w3(32'h39893551),
	.w4(32'hb9c7f0af),
	.w5(32'hb9a3f0b5),
	.w6(32'hb64da442),
	.w7(32'hb9aff2cf),
	.w8(32'hb9322187),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60c237),
	.w1(32'h37b76dac),
	.w2(32'h3a62c8a1),
	.w3(32'hb97e7a66),
	.w4(32'h398398bb),
	.w5(32'h3a4ea0c0),
	.w6(32'hbaa1f1f7),
	.w7(32'h3961e594),
	.w8(32'h3a2c3025),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38895953),
	.w1(32'hb902e314),
	.w2(32'hb722d243),
	.w3(32'hb8193aa2),
	.w4(32'hb945100e),
	.w5(32'h3881f69f),
	.w6(32'hb66993b6),
	.w7(32'hb8f2a8a6),
	.w8(32'h3809e970),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e2f6b),
	.w1(32'hba8b2ab6),
	.w2(32'hb9dbe316),
	.w3(32'h3a029885),
	.w4(32'h375918e2),
	.w5(32'h3a5b09de),
	.w6(32'h3a05ea6d),
	.w7(32'h3a0c57cc),
	.w8(32'h3aa13f04),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb708a6e7),
	.w1(32'hb77d13dc),
	.w2(32'hb719e2ba),
	.w3(32'hb7394671),
	.w4(32'hb83e5eb0),
	.w5(32'hb80ac4ca),
	.w6(32'hb8a9c40a),
	.w7(32'hb8b27b81),
	.w8(32'hb864df71),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3815dadc),
	.w1(32'h370c6b73),
	.w2(32'h37ba42ae),
	.w3(32'h36173286),
	.w4(32'hb6e97f58),
	.w5(32'hb72e1b1a),
	.w6(32'hb818d8a5),
	.w7(32'h36b7d553),
	.w8(32'h377c13fd),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb943800a),
	.w1(32'h390cf35f),
	.w2(32'h38b3586b),
	.w3(32'hb9056019),
	.w4(32'h38f4593a),
	.w5(32'h3958be55),
	.w6(32'hb9c1b81f),
	.w7(32'hb8d57054),
	.w8(32'h387d07d5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b5187),
	.w1(32'hba5f09e2),
	.w2(32'hbafd9567),
	.w3(32'h3ab4a0d9),
	.w4(32'h37b19b50),
	.w5(32'hba9de1b4),
	.w6(32'h3a172bd0),
	.w7(32'h3a2f6914),
	.w8(32'h39219ce9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cc6348),
	.w1(32'hb8b04303),
	.w2(32'h38bd7a58),
	.w3(32'hba1d11c6),
	.w4(32'hb978436d),
	.w5(32'hb8c0c29a),
	.w6(32'hba0d84ca),
	.w7(32'hb94d988a),
	.w8(32'hb8906573),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d303c3),
	.w1(32'h39976794),
	.w2(32'h392c56df),
	.w3(32'hb9984628),
	.w4(32'h39c74f5b),
	.w5(32'h39d47a34),
	.w6(32'hba546355),
	.w7(32'hb8fdf425),
	.w8(32'hb914b9b4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0aa3a2),
	.w1(32'hb8d7bf94),
	.w2(32'h38e62494),
	.w3(32'hba89da50),
	.w4(32'hba361211),
	.w5(32'hb911560f),
	.w6(32'hba587202),
	.w7(32'hba2cb16d),
	.w8(32'hb82780d5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07c85d),
	.w1(32'hbaa7e80d),
	.w2(32'h3a1d8592),
	.w3(32'hba41b47a),
	.w4(32'h39107e08),
	.w5(32'h3ac67b1e),
	.w6(32'h3919ac9b),
	.w7(32'hb9ac3b35),
	.w8(32'h3ae1f8b7),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba211f7e),
	.w1(32'h38814bb0),
	.w2(32'h3a633cf3),
	.w3(32'hbaa0c3fe),
	.w4(32'h3941d10d),
	.w5(32'h3a89f760),
	.w6(32'hba7219b8),
	.w7(32'hb95eaa12),
	.w8(32'h3a145a00),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bf633),
	.w1(32'hba7c2583),
	.w2(32'h3a1e3136),
	.w3(32'hb9779467),
	.w4(32'hb9b04a84),
	.w5(32'h3a77fe68),
	.w6(32'h3906c04c),
	.w7(32'h39cb0be3),
	.w8(32'h3aaab7ec),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9180f37),
	.w1(32'hb93da67a),
	.w2(32'h387fcffc),
	.w3(32'hb94d6101),
	.w4(32'hb976c486),
	.w5(32'h38277587),
	.w6(32'hb97d016c),
	.w7(32'hb993d03b),
	.w8(32'h37f8ea7c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fcb8ae),
	.w1(32'h395ab1c6),
	.w2(32'h3ab85e6a),
	.w3(32'hba0d44a6),
	.w4(32'h383195b1),
	.w5(32'h3a993da7),
	.w6(32'hb9c66d3a),
	.w7(32'hb7a4fe2b),
	.w8(32'h3a470147),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365fc29e),
	.w1(32'hb7104541),
	.w2(32'hb70f2518),
	.w3(32'h34b88c15),
	.w4(32'hb6c94999),
	.w5(32'hb71e0016),
	.w6(32'h37024d3b),
	.w7(32'h36404ad3),
	.w8(32'hb6a29775),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906acf3),
	.w1(32'hb9487ad5),
	.w2(32'hb8fba6a9),
	.w3(32'hb8af1630),
	.w4(32'hb8e4fc0c),
	.w5(32'hb78e8dd9),
	.w6(32'h35dc9e74),
	.w7(32'hb8d8e9bb),
	.w8(32'hb8309999),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ced8d),
	.w1(32'h3895b855),
	.w2(32'h37ea634a),
	.w3(32'hb89e1805),
	.w4(32'h3811b940),
	.w5(32'hb7be0508),
	.w6(32'hb959fdd9),
	.w7(32'hb3be5484),
	.w8(32'hb7616e1f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56a389),
	.w1(32'hb9aa48cb),
	.w2(32'h3af4aa7e),
	.w3(32'hba9e450f),
	.w4(32'hb959021b),
	.w5(32'h3ad23a04),
	.w6(32'hb9ffbbb0),
	.w7(32'hb989b0f4),
	.w8(32'h3ac101c7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369699f8),
	.w1(32'h36a9133a),
	.w2(32'hb5b540d0),
	.w3(32'h368f4281),
	.w4(32'h36182537),
	.w5(32'hb7193d9b),
	.w6(32'h359b0527),
	.w7(32'h3623a022),
	.w8(32'hb72d198c),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb857e9b3),
	.w1(32'hb810db17),
	.w2(32'h3814d0f1),
	.w3(32'hb7b4c563),
	.w4(32'h379c8060),
	.w5(32'h388b2516),
	.w6(32'hb7321197),
	.w7(32'h37d671a4),
	.w8(32'h3858ec9d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ac748),
	.w1(32'hb8dbee96),
	.w2(32'h39e6613e),
	.w3(32'hb9c4c899),
	.w4(32'hb92cc47b),
	.w5(32'h375332e6),
	.w6(32'hba4669ea),
	.w7(32'hb9ecd521),
	.w8(32'h38f8be17),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915ef51),
	.w1(32'h3949edf3),
	.w2(32'h38f4cba8),
	.w3(32'hba819e42),
	.w4(32'h38242f46),
	.w5(32'hb9e9ff1b),
	.w6(32'hb9fe56dc),
	.w7(32'hba9344b3),
	.w8(32'hba55156d),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa95069),
	.w1(32'h3a1bb5e5),
	.w2(32'hbb0b4e28),
	.w3(32'h399ee52e),
	.w4(32'h391da82d),
	.w5(32'hbb23bbe8),
	.w6(32'hb8eb7b38),
	.w7(32'hb9e66538),
	.w8(32'hbb19a703),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f2416),
	.w1(32'hb7b988f2),
	.w2(32'hb91c8ef3),
	.w3(32'hb7c576d8),
	.w4(32'hb8eaed92),
	.w5(32'hb8abd473),
	.w6(32'hb8b33665),
	.w7(32'hb8cf5c71),
	.w8(32'hb8f591f2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac95833),
	.w1(32'hbad2b6a3),
	.w2(32'h3a8ee0ae),
	.w3(32'hb8b69c9e),
	.w4(32'hb9e26bb7),
	.w5(32'h3b024665),
	.w6(32'hb961d853),
	.w7(32'h39bed659),
	.w8(32'h3b31af15),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccc787),
	.w1(32'hb93c8279),
	.w2(32'h3a680884),
	.w3(32'hbb51b5a7),
	.w4(32'hbaf0765a),
	.w5(32'h390c250e),
	.w6(32'hba90cbe9),
	.w7(32'hba637327),
	.w8(32'h3aeaadc0),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a336322),
	.w1(32'hb9aa0f05),
	.w2(32'hba845626),
	.w3(32'h3957f9a5),
	.w4(32'hb9825684),
	.w5(32'hb990884b),
	.w6(32'h39c27344),
	.w7(32'hb92eb09c),
	.w8(32'hb90c5bd5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374fc995),
	.w1(32'h37141f8e),
	.w2(32'h369116f8),
	.w3(32'h3712b94d),
	.w4(32'h367193a0),
	.w5(32'h36b4b72a),
	.w6(32'h3760a9bc),
	.w7(32'h3732c3b6),
	.w8(32'hb62dcc58),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8903ae1),
	.w1(32'h37cd2cad),
	.w2(32'h392455d0),
	.w3(32'h38d7b4e3),
	.w4(32'h3904e8d6),
	.w5(32'h3950b585),
	.w6(32'h390e29fd),
	.w7(32'h3906856c),
	.w8(32'h390abe4f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34557e67),
	.w1(32'hb61d516b),
	.w2(32'hb6faf435),
	.w3(32'h3781bfb0),
	.w4(32'h371759e9),
	.w5(32'hb6812edb),
	.w6(32'h36cd01d8),
	.w7(32'h3530a6f9),
	.w8(32'hb6ad51ce),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e9517),
	.w1(32'hba267b7f),
	.w2(32'hba993cc3),
	.w3(32'h3a3a8aae),
	.w4(32'h390395bf),
	.w5(32'hb98b4cfb),
	.w6(32'h3a0b4f5d),
	.w7(32'hb8f95369),
	.w8(32'h39651eb6),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8bf06),
	.w1(32'hb9eef977),
	.w2(32'hb92872f5),
	.w3(32'hb986145d),
	.w4(32'hb9299964),
	.w5(32'h389a3c0b),
	.w6(32'hb9e53828),
	.w7(32'hb78747ba),
	.w8(32'h38cd414d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39796180),
	.w1(32'h3a640f74),
	.w2(32'h397afafe),
	.w3(32'hb930fd89),
	.w4(32'h3a74d8f8),
	.w5(32'h396df841),
	.w6(32'hba2a54f7),
	.w7(32'h395fd9a0),
	.w8(32'hb9d34200),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376192b0),
	.w1(32'h3794c242),
	.w2(32'h38a382c8),
	.w3(32'h378ad896),
	.w4(32'h37afe0c9),
	.w5(32'h37e7ba9d),
	.w6(32'hb92ca23f),
	.w7(32'h37ef1203),
	.w8(32'h38a60473),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca0ef4),
	.w1(32'hba7e08be),
	.w2(32'h3910ecac),
	.w3(32'h382fa053),
	.w4(32'hb82181da),
	.w5(32'h3a4cc809),
	.w6(32'h3988b0fa),
	.w7(32'h398e248a),
	.w8(32'h3a92d7dc),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39486ffe),
	.w1(32'h39b5a5c6),
	.w2(32'hba27a2ca),
	.w3(32'h39c5eecf),
	.w4(32'h39ca60fe),
	.w5(32'hba4e28c9),
	.w6(32'hb9f3dd21),
	.w7(32'hb9bf9c2f),
	.w8(32'hba174e78),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f303e5),
	.w1(32'hb6661fdc),
	.w2(32'hb75928c0),
	.w3(32'h3680b7d1),
	.w4(32'hb6993edc),
	.w5(32'hb7602d4f),
	.w6(32'h366364e7),
	.w7(32'hb68d2674),
	.w8(32'hb751b4c6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6821d2),
	.w1(32'h395eec70),
	.w2(32'h3a8ee104),
	.w3(32'hb99fb6dc),
	.w4(32'h3a5fd800),
	.w5(32'h3a993b0c),
	.w6(32'hb79f8af8),
	.w7(32'h3a82118b),
	.w8(32'h3a863bf2),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375e29dd),
	.w1(32'h3621ee98),
	.w2(32'hb7b8049f),
	.w3(32'h37493b44),
	.w4(32'hb6865f23),
	.w5(32'hb7f77ac0),
	.w6(32'h378b2b33),
	.w7(32'h35d08e13),
	.w8(32'hb7c61770),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a850d6),
	.w1(32'hb9cb73e6),
	.w2(32'h37f2b4d0),
	.w3(32'hb94213b0),
	.w4(32'hb89f532b),
	.w5(32'h39bedf8d),
	.w6(32'hb99a5581),
	.w7(32'hb9043c32),
	.w8(32'h39bb6bb3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a57702),
	.w1(32'h3a1d5108),
	.w2(32'h39fffd57),
	.w3(32'hb9e1687b),
	.w4(32'hb8800418),
	.w5(32'hb83b1beb),
	.w6(32'hba664735),
	.w7(32'hb93aad35),
	.w8(32'h38938de5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961566e),
	.w1(32'h39885f18),
	.w2(32'h3915d232),
	.w3(32'hb933bbfa),
	.w4(32'h391f49e1),
	.w5(32'h3907cee3),
	.w6(32'hb9ebdb79),
	.w7(32'hb7061b91),
	.w8(32'h370667d8),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876316b),
	.w1(32'hb7cee329),
	.w2(32'h37697626),
	.w3(32'hb89e65e3),
	.w4(32'hb81143e7),
	.w5(32'h376ba117),
	.w6(32'hb88181ec),
	.w7(32'hb81325fe),
	.w8(32'h3624fbb5),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1cc923),
	.w1(32'h3a132a02),
	.w2(32'h39f74359),
	.w3(32'hba6cd088),
	.w4(32'h36fb8b43),
	.w5(32'h399a6fac),
	.w6(32'hba9a79b7),
	.w7(32'hb9f579d2),
	.w8(32'h385f2128),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a62e2b),
	.w1(32'hb9df2a59),
	.w2(32'h3a5014f1),
	.w3(32'hb9b1596c),
	.w4(32'hb874bdd4),
	.w5(32'h3a416f53),
	.w6(32'hb8c6e2ef),
	.w7(32'hb90ef41c),
	.w8(32'h3a20bf9a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9941dbe),
	.w1(32'hba016b01),
	.w2(32'hb929e1c5),
	.w3(32'hb9556a16),
	.w4(32'hb9106a09),
	.w5(32'h398f5f2d),
	.w6(32'hb9a28aa9),
	.w7(32'hb89a0231),
	.w8(32'h39d12b25),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4433c78),
	.w1(32'h371d0b90),
	.w2(32'h37732e0a),
	.w3(32'hb68ff046),
	.w4(32'hb5373494),
	.w5(32'h372f32f1),
	.w6(32'hb68ea5b9),
	.w7(32'h37847aa2),
	.w8(32'h37a8bc77),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369f7906),
	.w1(32'hb79e3c45),
	.w2(32'hb7b3b592),
	.w3(32'hb7124958),
	.w4(32'hb723d8f3),
	.w5(32'hb832070b),
	.w6(32'hb6c886a9),
	.w7(32'hb7bb68c3),
	.w8(32'hb7c74f1a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4e902),
	.w1(32'hba310d79),
	.w2(32'hba8639bf),
	.w3(32'h3ab13e76),
	.w4(32'h3a541b89),
	.w5(32'hb4cf85e0),
	.w6(32'hba530f87),
	.w7(32'h38911df8),
	.w8(32'h3a06dff4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23b321),
	.w1(32'hb950335a),
	.w2(32'h390223c0),
	.w3(32'h389e6e68),
	.w4(32'h39920d4b),
	.w5(32'h39a0866c),
	.w6(32'hba6bc84a),
	.w7(32'h39bb30d4),
	.w8(32'h3a85e459),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3862ca98),
	.w1(32'h39a74311),
	.w2(32'h39a25ba0),
	.w3(32'h385b00f8),
	.w4(32'h39602904),
	.w5(32'h39dceacc),
	.w6(32'hba1bb6d2),
	.w7(32'h39369563),
	.w8(32'h3961a143),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0af644),
	.w1(32'hbad8bde1),
	.w2(32'hba3dacdf),
	.w3(32'hbaa3aba7),
	.w4(32'hba8339ee),
	.w5(32'hba53b86d),
	.w6(32'h3a08ab1d),
	.w7(32'hba9faecd),
	.w8(32'h397f10cc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9d361),
	.w1(32'hb6080507),
	.w2(32'h39917177),
	.w3(32'hb88dde54),
	.w4(32'h3765e433),
	.w5(32'h39c03435),
	.w6(32'hb9410ace),
	.w7(32'h38a79331),
	.w8(32'h39f44f9d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f1c00c),
	.w1(32'hb87346c8),
	.w2(32'h3a0eb3bc),
	.w3(32'hb95fc804),
	.w4(32'h38282959),
	.w5(32'h39ba1fee),
	.w6(32'hb958e7f9),
	.w7(32'h397d4dbd),
	.w8(32'h39954c38),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa2666),
	.w1(32'hbafe63ef),
	.w2(32'hbbc5a0eb),
	.w3(32'h3b362355),
	.w4(32'hbad5c815),
	.w5(32'hbb78fc4d),
	.w6(32'h38f664d2),
	.w7(32'hbb055b50),
	.w8(32'hbb18587b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7c74e),
	.w1(32'hba91ab6f),
	.w2(32'h3a0be485),
	.w3(32'h38079492),
	.w4(32'hba0ce0d9),
	.w5(32'h3a5be208),
	.w6(32'hb7d38dce),
	.w7(32'h39be5f5e),
	.w8(32'h3ae33864),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8daf71),
	.w1(32'h3873d61a),
	.w2(32'hbab1e5ba),
	.w3(32'h3a324155),
	.w4(32'hb9a824cd),
	.w5(32'hbaaf9560),
	.w6(32'h39822205),
	.w7(32'hb921a428),
	.w8(32'hba0f6a2f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c9f38),
	.w1(32'h39ba1a6b),
	.w2(32'h37e28381),
	.w3(32'hb9e5eb7d),
	.w4(32'h39d11928),
	.w5(32'hb817848a),
	.w6(32'hba718aee),
	.w7(32'h39124697),
	.w8(32'h383376b6),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe64cf),
	.w1(32'h3a3eb5f6),
	.w2(32'h3a16c317),
	.w3(32'hba3cdda4),
	.w4(32'h39324ca7),
	.w5(32'h398eba04),
	.w6(32'hba67928a),
	.w7(32'hb8020c83),
	.w8(32'h3997a08e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6033844),
	.w1(32'hb6800922),
	.w2(32'hb6f22c70),
	.w3(32'hb66171c0),
	.w4(32'hb6c69cd4),
	.w5(32'hb706f04e),
	.w6(32'hb6885d91),
	.w7(32'hb6d12dce),
	.w8(32'hb6f2a032),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365afdff),
	.w1(32'h34b2d6d5),
	.w2(32'hb62bc2e8),
	.w3(32'h36360276),
	.w4(32'hb4c49590),
	.w5(32'hb6b60944),
	.w6(32'h36177d77),
	.w7(32'h358636c8),
	.w8(32'hb669f7c0),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d5e462),
	.w1(32'hb9cf20fe),
	.w2(32'hb858f976),
	.w3(32'h39036d5a),
	.w4(32'h39344bd7),
	.w5(32'h3a2cde47),
	.w6(32'hb86d42ca),
	.w7(32'h393ef530),
	.w8(32'h3a284f5e),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h368be92d),
	.w1(32'hb69d36cd),
	.w2(32'hb720c8c9),
	.w3(32'h36b2e1d5),
	.w4(32'hb65ba6e9),
	.w5(32'hb70b9594),
	.w6(32'h36e67f42),
	.w7(32'hb5ad926e),
	.w8(32'hb6701e90),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a460edd),
	.w1(32'h37ff7a68),
	.w2(32'hb99c0006),
	.w3(32'h39e8aefd),
	.w4(32'h3949dfdd),
	.w5(32'h3992110a),
	.w6(32'h39795387),
	.w7(32'hb9108901),
	.w8(32'h3788d2f4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c576f6),
	.w1(32'h3a402e6a),
	.w2(32'h3a4b98a6),
	.w3(32'h3a3e9e3e),
	.w4(32'h39d9fc55),
	.w5(32'h39a0d94a),
	.w6(32'hba56144a),
	.w7(32'h3a341161),
	.w8(32'h3aba194d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8324327),
	.w1(32'h3902ce9d),
	.w2(32'hb6cb5de9),
	.w3(32'h37b88e4a),
	.w4(32'h39210f5a),
	.w5(32'h37f4e2cd),
	.w6(32'hb906a428),
	.w7(32'h38dce4eb),
	.w8(32'h390eff70),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36aa40f3),
	.w1(32'hb52d4302),
	.w2(32'hb687b5b1),
	.w3(32'h355f66a9),
	.w4(32'h365eadf0),
	.w5(32'hb6196e4b),
	.w6(32'hb6ae8613),
	.w7(32'h3551581e),
	.w8(32'hb68ec525),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a74e8),
	.w1(32'hb9a4f6b5),
	.w2(32'hbab13193),
	.w3(32'h3a86fb8b),
	.w4(32'h39735b1f),
	.w5(32'hbab457bd),
	.w6(32'h39f35834),
	.w7(32'hba0fc880),
	.w8(32'hb999267b),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ac802),
	.w1(32'hba2e3753),
	.w2(32'h38d0c589),
	.w3(32'hb801ea71),
	.w4(32'hb996cbc4),
	.w5(32'h39669c06),
	.w6(32'h381f6ef0),
	.w7(32'h388e2a56),
	.w8(32'h3a3a40e9),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h367c6562),
	.w1(32'hb5dd0049),
	.w2(32'h37149e7b),
	.w3(32'h3651f63e),
	.w4(32'hb683f2a2),
	.w5(32'h36a15a83),
	.w6(32'h370707f8),
	.w7(32'h35d94beb),
	.w8(32'h37042d6d),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b6ff5),
	.w1(32'hba7dcdd6),
	.w2(32'hba1ea8d0),
	.w3(32'hb808f253),
	.w4(32'hba35a820),
	.w5(32'hb946f14f),
	.w6(32'h394fc212),
	.w7(32'h37818bea),
	.w8(32'h3a181c62),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f38a8e),
	.w1(32'hb7d9150c),
	.w2(32'hb5f4899f),
	.w3(32'hb7cfacf3),
	.w4(32'hb7ef7086),
	.w5(32'h367d0a99),
	.w6(32'hb7e4c69b),
	.w7(32'hb78efa46),
	.w8(32'h376bd097),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74b0318),
	.w1(32'hb6117ddc),
	.w2(32'h38991939),
	.w3(32'hb8ae9969),
	.w4(32'hb835a02a),
	.w5(32'h371efa91),
	.w6(32'hb82a2ea0),
	.w7(32'h381d4a1a),
	.w8(32'h38ec064d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37af1aab),
	.w1(32'h37027044),
	.w2(32'hb70e33a5),
	.w3(32'h3651b72d),
	.w4(32'hb6f33a09),
	.w5(32'hb7694080),
	.w6(32'h36e9f54c),
	.w7(32'hb6ee53a6),
	.w8(32'hb7fc9b7f),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7405ec8),
	.w1(32'hb7501ba8),
	.w2(32'hb6f4125f),
	.w3(32'hb665bcfd),
	.w4(32'hb7898c86),
	.w5(32'hb742cdcd),
	.w6(32'hb740baaa),
	.w7(32'hb76afd7b),
	.w8(32'hb66c6737),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a93b),
	.w1(32'h36a7f706),
	.w2(32'hb9df31d1),
	.w3(32'h38a8d86a),
	.w4(32'h3932ee86),
	.w5(32'hb8b9317c),
	.w6(32'hb900a57c),
	.w7(32'h38f15e9f),
	.w8(32'hb920f8d6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04547a),
	.w1(32'hba956a8b),
	.w2(32'h3ab08ff0),
	.w3(32'hba73dcd7),
	.w4(32'hba403f06),
	.w5(32'h3ad49e33),
	.w6(32'hb8fcb312),
	.w7(32'hba78e670),
	.w8(32'h3ac190ec),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910928c),
	.w1(32'hba31cc11),
	.w2(32'h398144d3),
	.w3(32'h373d8a40),
	.w4(32'hb9881abf),
	.w5(32'h3a05a9d4),
	.w6(32'h3927f8fa),
	.w7(32'h39a90c5b),
	.w8(32'h3a839543),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10775c),
	.w1(32'hbaa68613),
	.w2(32'h39a4818d),
	.w3(32'hba4ca29b),
	.w4(32'hba07f4c4),
	.w5(32'h3a7d748d),
	.w6(32'h385ebf5f),
	.w7(32'hb9db9e22),
	.w8(32'h3a981cb8),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83430d2),
	.w1(32'hb82ccc1e),
	.w2(32'h3754dd38),
	.w3(32'hb82723d0),
	.w4(32'hb82204e1),
	.w5(32'hb6966db8),
	.w6(32'hb7b4ac2b),
	.w7(32'hb7dff306),
	.w8(32'hb6c8b63a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38def35a),
	.w1(32'h39036a64),
	.w2(32'h399f46d8),
	.w3(32'hb8c922b8),
	.w4(32'hb7e3aa73),
	.w5(32'h392f2780),
	.w6(32'h389f7a2d),
	.w7(32'h38940589),
	.w8(32'h390e63e4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374fc830),
	.w1(32'h36a4bd58),
	.w2(32'hb7fa83b3),
	.w3(32'h36b24f0b),
	.w4(32'hb794372d),
	.w5(32'hb834ebee),
	.w6(32'h372aa873),
	.w7(32'hb69f7eb6),
	.w8(32'hb79ddfd4),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ab603d),
	.w1(32'h36a79df0),
	.w2(32'h36bc0ebc),
	.w3(32'hb6b04148),
	.w4(32'hb70a8398),
	.w5(32'hb70757ef),
	.w6(32'h360ee8fb),
	.w7(32'h351ec384),
	.w8(32'h363c8c28),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31e902),
	.w1(32'h391adaab),
	.w2(32'h3b0a0311),
	.w3(32'hba05dc6a),
	.w4(32'hb7b35900),
	.w5(32'h3aea54a2),
	.w6(32'hb9c29c1c),
	.w7(32'h39dcc37b),
	.w8(32'h3abd4785),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fa9e47),
	.w1(32'h3814f283),
	.w2(32'h3924996c),
	.w3(32'h38f6bfa4),
	.w4(32'h39241763),
	.w5(32'h394f0034),
	.w6(32'h3908f487),
	.w7(32'h391823bb),
	.w8(32'h390892f1),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f7711),
	.w1(32'hb804c38f),
	.w2(32'h38c57f7f),
	.w3(32'hb966e5ff),
	.w4(32'hb8a120f1),
	.w5(32'h37a6caa6),
	.w6(32'hb9397f92),
	.w7(32'hb88c8bce),
	.w8(32'hb78548aa),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da3965),
	.w1(32'h39313a06),
	.w2(32'h39dd5aea),
	.w3(32'hb9a6b4c9),
	.w4(32'hb7f0b70b),
	.w5(32'h39b424ea),
	.w6(32'hb9dc1c85),
	.w7(32'hb937724d),
	.w8(32'h3807d03c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787beea),
	.w1(32'h37b8567f),
	.w2(32'h384d4a54),
	.w3(32'hb6a77227),
	.w4(32'h3819905d),
	.w5(32'h37e33ec5),
	.w6(32'h380e84aa),
	.w7(32'h3833974b),
	.w8(32'h381c96b3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923e644),
	.w1(32'hb9876a97),
	.w2(32'h38687f33),
	.w3(32'hb88087e5),
	.w4(32'hb8c767c8),
	.w5(32'h394b3db3),
	.w6(32'h368a129c),
	.w7(32'h383fe8dc),
	.w8(32'h39ae0722),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb807b0ab),
	.w1(32'h37bd5ff3),
	.w2(32'h391ff764),
	.w3(32'hb8124b6f),
	.w4(32'h3904aff0),
	.w5(32'h3915a181),
	.w6(32'h37a4f96d),
	.w7(32'h38cb3933),
	.w8(32'h390e3fd2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2c87b),
	.w1(32'hba02c247),
	.w2(32'h3b7c672d),
	.w3(32'hbada0ac7),
	.w4(32'hb7ffdb42),
	.w5(32'h3b80e24b),
	.w6(32'hba8a792c),
	.w7(32'hb9fcc219),
	.w8(32'h3b44ec3c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7803a4a),
	.w1(32'h3a299418),
	.w2(32'hb985fabe),
	.w3(32'hb4f4b87f),
	.w4(32'h39ab314c),
	.w5(32'hba7b3d74),
	.w6(32'h3ac83a85),
	.w7(32'hb7beac2d),
	.w8(32'h391c2166),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e7a59),
	.w1(32'h3986fce2),
	.w2(32'hba28ba2d),
	.w3(32'h3a57d843),
	.w4(32'hb8ac5c5f),
	.w5(32'hbabad943),
	.w6(32'h395eabfe),
	.w7(32'h3a19cc1f),
	.w8(32'hb9b66c5a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule