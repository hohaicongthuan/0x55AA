module layer_10_featuremap_458(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c1f161),
	.w1(32'h3a85354b),
	.w2(32'h3a5bdae7),
	.w3(32'h3a798a7d),
	.w4(32'h3aabb085),
	.w5(32'h3a0f8aa0),
	.w6(32'h3aba78e9),
	.w7(32'h3aad51dd),
	.w8(32'h3a94438d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7d6800),
	.w1(32'hba961b15),
	.w2(32'h381fd1ac),
	.w3(32'h3aa5ad55),
	.w4(32'hbb0b299b),
	.w5(32'hb911796c),
	.w6(32'h3a1ea494),
	.w7(32'hbb0e82a3),
	.w8(32'hb9e57e0a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e0fb4),
	.w1(32'hb86424dd),
	.w2(32'hbaa8f972),
	.w3(32'hba8a3e15),
	.w4(32'hba862b8b),
	.w5(32'hbb3586ce),
	.w6(32'hba116ff4),
	.w7(32'hba648af7),
	.w8(32'hba8c4aaf),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8699280),
	.w1(32'h3aaaf530),
	.w2(32'h39a26e9d),
	.w3(32'hbaea8f31),
	.w4(32'h3a0165ec),
	.w5(32'h3a10ac76),
	.w6(32'hba5f22ae),
	.w7(32'h3a02b376),
	.w8(32'hba463bd3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394212dd),
	.w1(32'hba6ea7d9),
	.w2(32'hba486641),
	.w3(32'hba515699),
	.w4(32'hb92b6eb3),
	.w5(32'h39157c4e),
	.w6(32'hba81ce3a),
	.w7(32'h38fdc986),
	.w8(32'h3a0f6df2),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998aad5),
	.w1(32'h390ebada),
	.w2(32'h3ae68865),
	.w3(32'h3a32a530),
	.w4(32'h3a327772),
	.w5(32'h3b4fda72),
	.w6(32'h39f3b894),
	.w7(32'h39ae29d4),
	.w8(32'h3b44d361),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772d767),
	.w1(32'hb90f6b79),
	.w2(32'hb8e7a2c7),
	.w3(32'h3a8a44c5),
	.w4(32'hbac3d342),
	.w5(32'h3853f9d8),
	.w6(32'h39f79975),
	.w7(32'hbaa2266f),
	.w8(32'h39a0cbdd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7338),
	.w1(32'h3af4587b),
	.w2(32'h3b0f7ccc),
	.w3(32'h3affdf43),
	.w4(32'h3aa72948),
	.w5(32'h3acc40e1),
	.w6(32'h3adba710),
	.w7(32'h3ac6d709),
	.w8(32'h3b15fa04),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8058e0),
	.w1(32'h39b29c5f),
	.w2(32'hb72d0eef),
	.w3(32'h39b94d9e),
	.w4(32'hb855fe50),
	.w5(32'hba41a2f7),
	.w6(32'hba6deca4),
	.w7(32'h3a1cce17),
	.w8(32'h398499dc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393dc01c),
	.w1(32'h3bbcaa72),
	.w2(32'h3bc0b933),
	.w3(32'hbaa342d0),
	.w4(32'h3b76fe82),
	.w5(32'h3ba39f45),
	.w6(32'hba78487f),
	.w7(32'h3b41b847),
	.w8(32'h3bad172b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d1aaa),
	.w1(32'hba1466ad),
	.w2(32'hbb24df6d),
	.w3(32'hb9670983),
	.w4(32'h39e7f458),
	.w5(32'hba1dafcb),
	.w6(32'h3a60a350),
	.w7(32'h3a698c16),
	.w8(32'h384a42aa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42866c),
	.w1(32'hbb65cd0e),
	.w2(32'hbae77e1e),
	.w3(32'hbafc3792),
	.w4(32'hbb889a69),
	.w5(32'hbad896fa),
	.w6(32'hba7fc842),
	.w7(32'hbb6b4a6b),
	.w8(32'hbb25b034),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43a35),
	.w1(32'h3b918369),
	.w2(32'h3b584e66),
	.w3(32'h3ae264ad),
	.w4(32'h3b5c6c93),
	.w5(32'h3b8e46bd),
	.w6(32'h38d23adf),
	.w7(32'h3b616ef4),
	.w8(32'h3b5814fc),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74faddd),
	.w1(32'hb94d5ad8),
	.w2(32'h351f7cca),
	.w3(32'hba7df15e),
	.w4(32'hb980bad3),
	.w5(32'h399bbaa5),
	.w6(32'hb94a2b91),
	.w7(32'h394ee0ae),
	.w8(32'h3a9faf7e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6dc7594),
	.w1(32'hb98d2c19),
	.w2(32'hb91720bc),
	.w3(32'hb95dafe7),
	.w4(32'hbb020b06),
	.w5(32'hba7249ed),
	.w6(32'h395c6246),
	.w7(32'hbafaad93),
	.w8(32'hb979824c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b991b),
	.w1(32'h3af517a7),
	.w2(32'h3b5632f1),
	.w3(32'hb9ece367),
	.w4(32'h39de001f),
	.w5(32'h3b21378a),
	.w6(32'hba54413f),
	.w7(32'h3a46b680),
	.w8(32'h3b2ad225),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00d042),
	.w1(32'hb92804f5),
	.w2(32'hba74862d),
	.w3(32'h39b7ace6),
	.w4(32'hb8e6bd4e),
	.w5(32'hba2b4bc7),
	.w6(32'h3a507e20),
	.w7(32'hb7a8f213),
	.w8(32'hb9ffdb4a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac21bce),
	.w1(32'h3b6c5b1f),
	.w2(32'h3b893336),
	.w3(32'h3a397791),
	.w4(32'h3b74cf60),
	.w5(32'h3b693669),
	.w6(32'h3ac9677f),
	.w7(32'h3b890316),
	.w8(32'h3b6508fb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a461b0d),
	.w1(32'h3b1b8351),
	.w2(32'h3ae16835),
	.w3(32'h3a7727f4),
	.w4(32'h3ad136e5),
	.w5(32'h3b668f64),
	.w6(32'h3ad2d569),
	.w7(32'h3ac06e2a),
	.w8(32'h3b517292),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950c1b2),
	.w1(32'h3904afd9),
	.w2(32'hbaf7e0ef),
	.w3(32'hb98d2ce4),
	.w4(32'h38c95d8b),
	.w5(32'hba166073),
	.w6(32'hb9a7fb51),
	.w7(32'hb99e01a1),
	.w8(32'hbb138454),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bb08b),
	.w1(32'hba2b3e45),
	.w2(32'h39fc81b2),
	.w3(32'hbb357ca9),
	.w4(32'h39e982cc),
	.w5(32'h3b145c03),
	.w6(32'hbaded8a8),
	.w7(32'h39aa555b),
	.w8(32'h3ad86098),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bee9de),
	.w1(32'hba9055d1),
	.w2(32'hba7c981b),
	.w3(32'h3a09ac56),
	.w4(32'hbac1484b),
	.w5(32'hbae89769),
	.w6(32'h3927e267),
	.w7(32'hbb00a53c),
	.w8(32'hbb1a5f69),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51a745),
	.w1(32'h39d60674),
	.w2(32'h3b8ca2ff),
	.w3(32'hbbbc881e),
	.w4(32'hbb022b4d),
	.w5(32'h3bd006fc),
	.w6(32'hbb6a8ebb),
	.w7(32'hbb6eb4b2),
	.w8(32'h3b98f72b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43846a),
	.w1(32'h3b055687),
	.w2(32'h3ada3f1c),
	.w3(32'hba20805a),
	.w4(32'hba6f9b3a),
	.w5(32'h39ccf6c1),
	.w6(32'hba82c944),
	.w7(32'hba84bd4c),
	.w8(32'h3a73913b),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a8d2a),
	.w1(32'h3a335f29),
	.w2(32'h3b60718b),
	.w3(32'hba0908cc),
	.w4(32'hb9653333),
	.w5(32'h3b298443),
	.w6(32'hba4b6086),
	.w7(32'hb966e612),
	.w8(32'h3ac4b013),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba353456),
	.w1(32'h398b9382),
	.w2(32'hb996500e),
	.w3(32'hbaddcbd7),
	.w4(32'hb99aa59a),
	.w5(32'hbb2c9ea4),
	.w6(32'hbab38cc1),
	.w7(32'hba14bb6f),
	.w8(32'hba1f7875),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba60d9f6),
	.w1(32'hba3ed1eb),
	.w2(32'hba96698e),
	.w3(32'hb995cff7),
	.w4(32'hbb0fbcae),
	.w5(32'hba82dbbc),
	.w6(32'hba0410fa),
	.w7(32'hbb21fcde),
	.w8(32'hb98c55b1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83933b),
	.w1(32'h39a97914),
	.w2(32'hb94eba09),
	.w3(32'hba52380f),
	.w4(32'h3a053a03),
	.w5(32'h388551bd),
	.w6(32'h38ff7699),
	.w7(32'h391b6477),
	.w8(32'hb9e7e5cb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb427),
	.w1(32'hbb369830),
	.w2(32'hba1b0679),
	.w3(32'hbb18ad3e),
	.w4(32'hbb75f72c),
	.w5(32'hba38aa30),
	.w6(32'hbb2e7b94),
	.w7(32'hbb7f660a),
	.w8(32'hbb0f0739),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb882c586),
	.w1(32'h3b57a68f),
	.w2(32'h3b945d93),
	.w3(32'hb9af3f02),
	.w4(32'h3b2b9d1f),
	.w5(32'h3b621412),
	.w6(32'h3a932f20),
	.w7(32'h3ad21276),
	.w8(32'h3b228884),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a9462),
	.w1(32'h3a5df2e3),
	.w2(32'h3a352dd9),
	.w3(32'h3a62130a),
	.w4(32'h390814ee),
	.w5(32'h3abfbfdc),
	.w6(32'h39ab587e),
	.w7(32'hb98d72e6),
	.w8(32'hb9c8aa30),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a147ea9),
	.w1(32'hb927badd),
	.w2(32'hbaa34f44),
	.w3(32'h3aa97810),
	.w4(32'hba6ba1a6),
	.w5(32'hba3ad726),
	.w6(32'h3a9dbddf),
	.w7(32'hba954f53),
	.w8(32'hb7e53152),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85f42e),
	.w1(32'h3ab9c8f6),
	.w2(32'h3ad72ebe),
	.w3(32'hb983a83d),
	.w4(32'h3a38f273),
	.w5(32'h3a37184a),
	.w6(32'hba663802),
	.w7(32'hb9dbc4b0),
	.w8(32'h3afd2171),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390cbccf),
	.w1(32'h39f00f74),
	.w2(32'h3a9be601),
	.w3(32'hba8229d4),
	.w4(32'h39d2f05e),
	.w5(32'h3af3d25f),
	.w6(32'h362fe6fa),
	.w7(32'hb967caa6),
	.w8(32'h3ac81e41),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81921f0),
	.w1(32'h3a143be3),
	.w2(32'h39f84ddc),
	.w3(32'hba09f080),
	.w4(32'hba007b4f),
	.w5(32'h38073233),
	.w6(32'hb984f665),
	.w7(32'h3a3c90fe),
	.w8(32'h39a5d0c3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395c5b72),
	.w1(32'h3a5d2522),
	.w2(32'h3ac85ba9),
	.w3(32'h399adf5f),
	.w4(32'h39aa3a87),
	.w5(32'h3a922eae),
	.w6(32'h38be95f7),
	.w7(32'h3a2de76e),
	.w8(32'h3a981ee9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0b263),
	.w1(32'h3b194f21),
	.w2(32'h3aed0ec5),
	.w3(32'hba829b49),
	.w4(32'h39cfd576),
	.w5(32'h3add0967),
	.w6(32'hb9f10357),
	.w7(32'hba7396cb),
	.w8(32'h3a9ca4e9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14fc58),
	.w1(32'hbb6ce99f),
	.w2(32'hbae900fd),
	.w3(32'hba60e78d),
	.w4(32'hbbb18111),
	.w5(32'hbb39e93d),
	.w6(32'hb9e30ea9),
	.w7(32'hbbc2bcf9),
	.w8(32'hbb609ad9),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a3a7d),
	.w1(32'hbbc26989),
	.w2(32'hbb66522d),
	.w3(32'hbb5c1a63),
	.w4(32'hbb95373f),
	.w5(32'hbaf10cc5),
	.w6(32'hbb337f60),
	.w7(32'hbb9fb80f),
	.w8(32'hbb6d8942),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871226),
	.w1(32'h3a371382),
	.w2(32'hb94cba3c),
	.w3(32'h3aaa0a45),
	.w4(32'h3ae71092),
	.w5(32'h3a92ea15),
	.w6(32'h3aa64935),
	.w7(32'h3afe3f15),
	.w8(32'h3ad6c719),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d86e8),
	.w1(32'hba7b480a),
	.w2(32'hba75ef39),
	.w3(32'h3a8ff570),
	.w4(32'hb9effc2c),
	.w5(32'hbab029a2),
	.w6(32'h39b45a79),
	.w7(32'hb9828ea6),
	.w8(32'hba80d1e5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad240f9),
	.w1(32'hbaba13f6),
	.w2(32'hbae76dad),
	.w3(32'hba74a1c1),
	.w4(32'hbaa19edc),
	.w5(32'h3985f88f),
	.w6(32'hbacbf08f),
	.w7(32'hba766047),
	.w8(32'hb95eb207),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cc245),
	.w1(32'h3aae49b5),
	.w2(32'h3a61a62c),
	.w3(32'h37783e85),
	.w4(32'h39605117),
	.w5(32'h3a2803bc),
	.w6(32'hba32d04f),
	.w7(32'h390f866c),
	.w8(32'hb891e4da),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93ba68),
	.w1(32'h3bbd24ee),
	.w2(32'h3b6beed2),
	.w3(32'h3b06dd79),
	.w4(32'h3ba73854),
	.w5(32'h3b86a332),
	.w6(32'h3a90397c),
	.w7(32'h3b986aca),
	.w8(32'h3b92eef4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02c886),
	.w1(32'h3ab696be),
	.w2(32'h3b06ff2b),
	.w3(32'h381991f1),
	.w4(32'hbaa7bef3),
	.w5(32'h3a958813),
	.w6(32'hbad087db),
	.w7(32'hbb18971a),
	.w8(32'h3a5133c2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a933bf8),
	.w1(32'h3a1b634a),
	.w2(32'h3b19ae9a),
	.w3(32'hbaa395ef),
	.w4(32'hbb2e3055),
	.w5(32'h3a5e598c),
	.w6(32'hbaec52a5),
	.w7(32'hbaf2e6b7),
	.w8(32'h3aafd323),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae90351),
	.w1(32'h3b5a9e63),
	.w2(32'h3b9ae310),
	.w3(32'h3a36df5e),
	.w4(32'h3af1f60a),
	.w5(32'h3b886b98),
	.w6(32'hba80c2cc),
	.w7(32'h39cbd41d),
	.w8(32'h3b5b7cff),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5ab8a),
	.w1(32'h3b24b891),
	.w2(32'h3b5b0908),
	.w3(32'h3b86a389),
	.w4(32'h3b96f762),
	.w5(32'h3bdd50e6),
	.w6(32'h3bc2b223),
	.w7(32'h3ba39010),
	.w8(32'h3bc7fefb),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a5ae1),
	.w1(32'hba202576),
	.w2(32'h3ac6cc32),
	.w3(32'hba495f72),
	.w4(32'hb6872468),
	.w5(32'h3b061221),
	.w6(32'hb9d3667f),
	.w7(32'h398c46d3),
	.w8(32'h3b186ddc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb742905b),
	.w1(32'hb98fdf56),
	.w2(32'h3b1fd1d0),
	.w3(32'h3a304a65),
	.w4(32'h3a0ab48c),
	.w5(32'h3b424228),
	.w6(32'h39c689c9),
	.w7(32'h3a229519),
	.w8(32'h3b7e7685),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a512d10),
	.w1(32'hba28d97b),
	.w2(32'hba48b2d5),
	.w3(32'h3a0a3501),
	.w4(32'hbb0e8d27),
	.w5(32'hb9925f14),
	.w6(32'hba145562),
	.w7(32'hbaaccea6),
	.w8(32'hba5be14b),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3955cbfb),
	.w1(32'hba3347b9),
	.w2(32'h3a2467fb),
	.w3(32'hba2e8a82),
	.w4(32'hbaf48561),
	.w5(32'hb9d01a03),
	.w6(32'hba4799ab),
	.w7(32'hba4a189c),
	.w8(32'h397e2039),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf78bcf),
	.w1(32'h39739642),
	.w2(32'h3afa4235),
	.w3(32'hbaa91efa),
	.w4(32'h3a3799ab),
	.w5(32'h3b22d0f3),
	.w6(32'hbb0a0c30),
	.w7(32'h39b60e85),
	.w8(32'h3b2aaf51),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871573),
	.w1(32'h3a8d921e),
	.w2(32'h3b070b73),
	.w3(32'h39157d49),
	.w4(32'h39e9561b),
	.w5(32'h3afc39d7),
	.w6(32'h3a0d2994),
	.w7(32'h3ab83905),
	.w8(32'h3b6796b8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbadf0),
	.w1(32'h3a981bac),
	.w2(32'hba144158),
	.w3(32'hba216e97),
	.w4(32'h3a55dbef),
	.w5(32'h38a0dd63),
	.w6(32'h3a141a41),
	.w7(32'hb893a666),
	.w8(32'hb9af8c3e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2097db),
	.w1(32'hbad5fa28),
	.w2(32'hba8dd181),
	.w3(32'hba9a0e26),
	.w4(32'hba96c651),
	.w5(32'hb9b09423),
	.w6(32'hbab8ad64),
	.w7(32'hba2547da),
	.w8(32'h3a52881d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1096f8),
	.w1(32'hb9383c2e),
	.w2(32'hb9a1df47),
	.w3(32'hbac2cb9d),
	.w4(32'h38c8f2f5),
	.w5(32'hb90067e7),
	.w6(32'hb9f415ad),
	.w7(32'h391fb4ad),
	.w8(32'hb8082efd),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379f30cd),
	.w1(32'hba62f42f),
	.w2(32'hbacac424),
	.w3(32'hb9a3db96),
	.w4(32'hba6ef5cb),
	.w5(32'hba324fb5),
	.w6(32'h3868ac17),
	.w7(32'hba2f8d61),
	.w8(32'hb9c5d4fb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ef941),
	.w1(32'h3a4c74d7),
	.w2(32'hba867876),
	.w3(32'hb90521b6),
	.w4(32'h3a68e52c),
	.w5(32'hba84ae63),
	.w6(32'hb9c7361f),
	.w7(32'h3a7a373a),
	.w8(32'hba940411),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed5de),
	.w1(32'hb9c1b1f5),
	.w2(32'hb921f1fe),
	.w3(32'hb74b6260),
	.w4(32'hb912e8e7),
	.w5(32'hbac9175a),
	.w6(32'h3978acce),
	.w7(32'h3a0c9e45),
	.w8(32'hbadb9064),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2ff9b),
	.w1(32'h3b04244c),
	.w2(32'h3b1643b4),
	.w3(32'h3ab08877),
	.w4(32'h3a8efd78),
	.w5(32'h3b4e0ddf),
	.w6(32'h39392200),
	.w7(32'h3ab4de03),
	.w8(32'h3b41a51b),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acba207),
	.w1(32'h37587bcc),
	.w2(32'hba8c627e),
	.w3(32'h3b1b4f0d),
	.w4(32'hb9de92b9),
	.w5(32'h3929e6c4),
	.w6(32'h3ab45b65),
	.w7(32'hba8cbfa4),
	.w8(32'h3957caf2),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980505a),
	.w1(32'h3adfdb09),
	.w2(32'hb9ef1e95),
	.w3(32'hba4c1f76),
	.w4(32'h3a6584d2),
	.w5(32'hba7daeac),
	.w6(32'hba6f0d82),
	.w7(32'h3ad097b4),
	.w8(32'hbaa0886f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96efc7),
	.w1(32'hba140356),
	.w2(32'hb9df82fd),
	.w3(32'hbae8bf05),
	.w4(32'hbab2e462),
	.w5(32'hba800536),
	.w6(32'hba538ad6),
	.w7(32'hba55b12a),
	.w8(32'hbab85170),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8c9c7),
	.w1(32'h3abeb51b),
	.w2(32'h3b0d96a2),
	.w3(32'hba9923c5),
	.w4(32'h3ad95bbe),
	.w5(32'h3aa4f4e4),
	.w6(32'hb982386f),
	.w7(32'h3ae47d9b),
	.w8(32'h3af4f97b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28646f),
	.w1(32'h39a57835),
	.w2(32'hb93a027e),
	.w3(32'h3b0e396d),
	.w4(32'h3a0ef78b),
	.w5(32'h3a5da796),
	.w6(32'h3af51342),
	.w7(32'h3a935d1b),
	.w8(32'h3ac84aca),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e0d2d),
	.w1(32'h3ae688a1),
	.w2(32'h3b008d71),
	.w3(32'h3b245698),
	.w4(32'h3a3a75f7),
	.w5(32'h3ad168c2),
	.w6(32'h3b1c732e),
	.w7(32'h3a9ed924),
	.w8(32'h3b029cc7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9e8bb),
	.w1(32'h3a26109d),
	.w2(32'h3b3502ba),
	.w3(32'hbb12e653),
	.w4(32'hba8e3fa0),
	.w5(32'h3b1b4dd5),
	.w6(32'hbb251d0a),
	.w7(32'hbb225b74),
	.w8(32'h3a299590),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e367e),
	.w1(32'hba181737),
	.w2(32'h3a2d430b),
	.w3(32'hbac611ef),
	.w4(32'hbb42df60),
	.w5(32'hba01b2c1),
	.w6(32'hbb61b059),
	.w7(32'hbb843b89),
	.w8(32'hbad306e4),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae10952),
	.w1(32'hbc30ad59),
	.w2(32'h3b4ab0ac),
	.w3(32'hbb492d31),
	.w4(32'hbc422c9e),
	.w5(32'h3c11090c),
	.w6(32'hbb87c74d),
	.w7(32'hbc43ad90),
	.w8(32'h3af907eb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1222a6),
	.w1(32'hbb1029d1),
	.w2(32'h3a768ea7),
	.w3(32'hbaac3882),
	.w4(32'hbb608d0a),
	.w5(32'h3a010834),
	.w6(32'hbb6121be),
	.w7(32'hbb322fb8),
	.w8(32'h39d1caf6),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f5d2c),
	.w1(32'h3bfce92a),
	.w2(32'hbae38350),
	.w3(32'h3b94e101),
	.w4(32'h3b03bb34),
	.w5(32'hbb859f36),
	.w6(32'h3b80277b),
	.w7(32'h3af6e602),
	.w8(32'h3a394f2f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8a04d),
	.w1(32'h3ba7caf3),
	.w2(32'h3b81a787),
	.w3(32'hbb098921),
	.w4(32'h3a23b34d),
	.w5(32'h3a7beef8),
	.w6(32'h3b9ffd35),
	.w7(32'hba6c51be),
	.w8(32'h3b31a02f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af97b6f),
	.w1(32'h3babbe0e),
	.w2(32'h3c223a6f),
	.w3(32'h3a33a882),
	.w4(32'h3b8bc15c),
	.w5(32'h3bea2292),
	.w6(32'h39b63c11),
	.w7(32'h3c0302e3),
	.w8(32'h3c2b41c1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5d365),
	.w1(32'h3c37693b),
	.w2(32'h3c1ab234),
	.w3(32'h3bc79dfe),
	.w4(32'h3b183b7e),
	.w5(32'hba88971d),
	.w6(32'h3bd09ca7),
	.w7(32'h3b885b40),
	.w8(32'h3bbf55e1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b479c84),
	.w1(32'h3c1d5f4c),
	.w2(32'h39db8778),
	.w3(32'hbbe84068),
	.w4(32'h3c020688),
	.w5(32'hbadb1a87),
	.w6(32'h3ada507f),
	.w7(32'h3b8d7c36),
	.w8(32'h3b6c134c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb8a51),
	.w1(32'h3bed587f),
	.w2(32'h3bab6cf3),
	.w3(32'hbb407d30),
	.w4(32'h3bded87d),
	.w5(32'h3a06f493),
	.w6(32'hbb3ac216),
	.w7(32'h3c2d39b2),
	.w8(32'h3b9a38b6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a500ab7),
	.w1(32'h3b255e83),
	.w2(32'hb9e8889f),
	.w3(32'h3a4eaa79),
	.w4(32'hbbede76d),
	.w5(32'hbbe0549c),
	.w6(32'h388b5dfa),
	.w7(32'hbb534c50),
	.w8(32'hbbe8647e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1758da),
	.w1(32'hbc18428d),
	.w2(32'hbb9c1e0e),
	.w3(32'hbbc8caaf),
	.w4(32'hbc81d979),
	.w5(32'hbc600e72),
	.w6(32'hbc103843),
	.w7(32'hbc65b9a0),
	.w8(32'hbbbb5382),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99130e1),
	.w1(32'hb93df665),
	.w2(32'hba9f6a38),
	.w3(32'hbbefc80f),
	.w4(32'h3a646cfd),
	.w5(32'hba86605c),
	.w6(32'hbbc8e3ee),
	.w7(32'h3ad95a85),
	.w8(32'h3982abe7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6bc5d),
	.w1(32'h3bfd84ea),
	.w2(32'hbb53d3da),
	.w3(32'hbb965a83),
	.w4(32'h3c12a96d),
	.w5(32'hbbab7601),
	.w6(32'hbb26838d),
	.w7(32'h3b93ff09),
	.w8(32'hbb8de197),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd963c),
	.w1(32'h3916f42c),
	.w2(32'h39a899ad),
	.w3(32'h3b2ab25a),
	.w4(32'h3aa644b5),
	.w5(32'h3a801424),
	.w6(32'hba3ef81f),
	.w7(32'h3a1e4aa6),
	.w8(32'hbaa0384e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23c856),
	.w1(32'h3c30da29),
	.w2(32'h3bb879a4),
	.w3(32'h39dfd73c),
	.w4(32'h3c72a4d1),
	.w5(32'h3b99c61f),
	.w6(32'hbb8518d2),
	.w7(32'h3bd9df0d),
	.w8(32'hbad8b6c7),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fd478),
	.w1(32'h3bb64052),
	.w2(32'h3b2d8625),
	.w3(32'h3afb7f56),
	.w4(32'h3bce9ecd),
	.w5(32'h3a322aa9),
	.w6(32'h39d1c92f),
	.w7(32'hba57d1c9),
	.w8(32'hbb1defec),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f10a1),
	.w1(32'h3994d98d),
	.w2(32'h3c165339),
	.w3(32'h3b0078e9),
	.w4(32'hba65de31),
	.w5(32'h3b871462),
	.w6(32'h3a8857e7),
	.w7(32'hbb4e3271),
	.w8(32'h3bf051c8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1958c5),
	.w1(32'hbb9d9711),
	.w2(32'hbabf7081),
	.w3(32'h3baf8ce0),
	.w4(32'h3a8af796),
	.w5(32'hbb1712ec),
	.w6(32'h3b97d66e),
	.w7(32'h3a2f6495),
	.w8(32'hbb150e0f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e1d57),
	.w1(32'hbc7941dd),
	.w2(32'hbbe4683c),
	.w3(32'hbb7877ec),
	.w4(32'hbc42c67b),
	.w5(32'hbbf89dbb),
	.w6(32'hbae99306),
	.w7(32'hbbc42994),
	.w8(32'hbbca9a37),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b2c17),
	.w1(32'hbb2adca3),
	.w2(32'hba6600e1),
	.w3(32'hbc0a611d),
	.w4(32'h3aba6d26),
	.w5(32'h3b0230c0),
	.w6(32'hbc123599),
	.w7(32'h3bef114c),
	.w8(32'h3a5caea0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40bb73),
	.w1(32'hbae43fd4),
	.w2(32'hb6d5936a),
	.w3(32'hbb6c5601),
	.w4(32'h3b883879),
	.w5(32'h3a939b26),
	.w6(32'hba251425),
	.w7(32'h3ae37a4d),
	.w8(32'h3b79a048),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06641e),
	.w1(32'hbb86138b),
	.w2(32'hbb024b23),
	.w3(32'hbbab9e1e),
	.w4(32'hbb5af9d1),
	.w5(32'h38b28b48),
	.w6(32'hbadaf429),
	.w7(32'hbb1a9540),
	.w8(32'h3a571d3f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba36ef8),
	.w1(32'hbbbbd2b5),
	.w2(32'h3ba017fc),
	.w3(32'hbbc7c55b),
	.w4(32'hbb5e197e),
	.w5(32'h3b3b57cc),
	.w6(32'hbbf506e3),
	.w7(32'hbbff066f),
	.w8(32'h3acc7866),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95a759),
	.w1(32'hba812af5),
	.w2(32'h3b8f7ab8),
	.w3(32'h3bb945ae),
	.w4(32'hb983fe9d),
	.w5(32'h3ac503e0),
	.w6(32'hba8ac108),
	.w7(32'hbb276e5a),
	.w8(32'h39b77d14),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95ac7b),
	.w1(32'hbb7d68a3),
	.w2(32'hbb593aae),
	.w3(32'hbb32cdd9),
	.w4(32'hba0bf4ce),
	.w5(32'hba99881b),
	.w6(32'hb93fb266),
	.w7(32'hbb9c1164),
	.w8(32'hbbacea0c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caed0c),
	.w1(32'hbb182837),
	.w2(32'hb9f178af),
	.w3(32'h3a8ab2e3),
	.w4(32'h3aa5da43),
	.w5(32'h3ad4b26e),
	.w6(32'hbb30d0ba),
	.w7(32'h3b167079),
	.w8(32'h3b81f226),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fe0dd),
	.w1(32'hbba90c12),
	.w2(32'hbba75f13),
	.w3(32'h3bcb28ff),
	.w4(32'hbb69e06e),
	.w5(32'hbbcf753b),
	.w6(32'h3b754895),
	.w7(32'h3a3499b0),
	.w8(32'h3b36c266),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef16cd),
	.w1(32'hbabcd068),
	.w2(32'h3b8dcc90),
	.w3(32'hbc35239c),
	.w4(32'h3aa0a58a),
	.w5(32'h3ca0bf25),
	.w6(32'h3b1961eb),
	.w7(32'hbb0a7d18),
	.w8(32'h3c49dd5e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f1e89),
	.w1(32'hbb22ad78),
	.w2(32'h3ad80864),
	.w3(32'h3bf65e5e),
	.w4(32'hba1faa67),
	.w5(32'h39ffcead),
	.w6(32'h3ba7f8f1),
	.w7(32'h3b54bd45),
	.w8(32'h3c08d511),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08a9cd),
	.w1(32'hbb17b3f3),
	.w2(32'hbaa4d67e),
	.w3(32'h3a955553),
	.w4(32'hbb93448d),
	.w5(32'hbb73dd66),
	.w6(32'h3be685ab),
	.w7(32'hbb738236),
	.w8(32'hb9f3610b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baac60d),
	.w1(32'hbc124035),
	.w2(32'hba54a2c3),
	.w3(32'h3b85d835),
	.w4(32'hbc2b844c),
	.w5(32'hbb673b0a),
	.w6(32'hba0c0390),
	.w7(32'hbb953d15),
	.w8(32'h3ad7c4f8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6a95c),
	.w1(32'hbbbefae3),
	.w2(32'hb94215cc),
	.w3(32'hbc043c25),
	.w4(32'hbbe8dfa9),
	.w5(32'hb96ba0fa),
	.w6(32'hbb6de9a7),
	.w7(32'hbb813e55),
	.w8(32'h3b5d16f6),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2d87c),
	.w1(32'h3ad29dce),
	.w2(32'h3b42ea98),
	.w3(32'h3b6e0cc3),
	.w4(32'hb7484d7d),
	.w5(32'h3ab3bb82),
	.w6(32'h3a81709d),
	.w7(32'hba06e5bb),
	.w8(32'h3b595543),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20d636),
	.w1(32'h3bb88fc7),
	.w2(32'h3c8b9a09),
	.w3(32'h3bd830d6),
	.w4(32'h3c3fb230),
	.w5(32'h3ccddac3),
	.w6(32'h3c0004df),
	.w7(32'h393f80de),
	.w8(32'h3c864858),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e58fd),
	.w1(32'hbc0e27d1),
	.w2(32'hbc86696e),
	.w3(32'h3c857dc0),
	.w4(32'hbb3630ca),
	.w5(32'hbbbec3da),
	.w6(32'h3c5a6538),
	.w7(32'hbbb68479),
	.w8(32'hbc153ae0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a8ecd),
	.w1(32'hbb989a73),
	.w2(32'h3bdd5c65),
	.w3(32'hbbe5cf1f),
	.w4(32'hbab1f21f),
	.w5(32'h3b0d74c6),
	.w6(32'hbc3c39d7),
	.w7(32'hbb7953b1),
	.w8(32'h3bbf04e2),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b13c2),
	.w1(32'hbb1eaa88),
	.w2(32'hbb0b04f8),
	.w3(32'hbbd0d340),
	.w4(32'h3a095365),
	.w5(32'hbae0ea18),
	.w6(32'hbc0e3835),
	.w7(32'hbb0a29f3),
	.w8(32'h3b78a34a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d3aaf),
	.w1(32'h3b07dce5),
	.w2(32'h3be38fc4),
	.w3(32'h3b62035e),
	.w4(32'h3bb777f6),
	.w5(32'h3badd97b),
	.w6(32'h3b425186),
	.w7(32'h3be2a03f),
	.w8(32'h3c14bf1c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb433d),
	.w1(32'h3b927bd4),
	.w2(32'hbaceacc9),
	.w3(32'h3b8094c9),
	.w4(32'h3b3076df),
	.w5(32'hbba31c19),
	.w6(32'h3b88002a),
	.w7(32'hbba39caf),
	.w8(32'hbbf39ebf),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf3f44),
	.w1(32'hbafaa5f7),
	.w2(32'h3bc05260),
	.w3(32'h3bbe943e),
	.w4(32'hbbf37d2d),
	.w5(32'h3c350eb3),
	.w6(32'h3b0e7080),
	.w7(32'hbc329811),
	.w8(32'h3c0a834c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1306bd),
	.w1(32'h3bcf24e3),
	.w2(32'h3b2a37b5),
	.w3(32'h3bd8fe6c),
	.w4(32'h3be545c4),
	.w5(32'h3b3712a0),
	.w6(32'h3bb2bcb7),
	.w7(32'h3ba20aa1),
	.w8(32'h3bd3138b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34d1da),
	.w1(32'h3bd66fb2),
	.w2(32'h3ba5bc29),
	.w3(32'hbaa2c82f),
	.w4(32'h3b7c6702),
	.w5(32'h3bda197f),
	.w6(32'h3afa034a),
	.w7(32'hbc2d78ab),
	.w8(32'hbb3f4646),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46649a),
	.w1(32'h3bdd2f04),
	.w2(32'h3bad7c2e),
	.w3(32'hba584eb4),
	.w4(32'hb92c0039),
	.w5(32'hba8674eb),
	.w6(32'hb9c5bcf3),
	.w7(32'hbb1e715f),
	.w8(32'hbb971b78),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61b7c8),
	.w1(32'h3b226ee6),
	.w2(32'h3a8037d5),
	.w3(32'hbbb0414f),
	.w4(32'hb7fa4264),
	.w5(32'h3ae9a0d8),
	.w6(32'hbbcfbc9a),
	.w7(32'h3b9b6c35),
	.w8(32'h3b901778),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b018e),
	.w1(32'hbb5b7838),
	.w2(32'h3ad95296),
	.w3(32'hbaa8d076),
	.w4(32'h3b13fa9f),
	.w5(32'h3c1625a9),
	.w6(32'h3a6ffb51),
	.w7(32'h3a128688),
	.w8(32'h3bb84522),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4ce98),
	.w1(32'h3c86d976),
	.w2(32'hbbc84ce1),
	.w3(32'h3bd89f8c),
	.w4(32'h3d001bed),
	.w5(32'hbc3336c6),
	.w6(32'h3b7650a0),
	.w7(32'h3c7e46b3),
	.w8(32'hbbd89081),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3666b),
	.w1(32'hbbc98eee),
	.w2(32'hbbaa129a),
	.w3(32'hbca4a781),
	.w4(32'hbc0e7258),
	.w5(32'hbbe57c55),
	.w6(32'hbca6b4a0),
	.w7(32'hbba43ea4),
	.w8(32'hbbbf53e9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab2dc4),
	.w1(32'h3ad8ba49),
	.w2(32'h3a52b6b2),
	.w3(32'hbc2fd5e5),
	.w4(32'hbb45777d),
	.w5(32'h3b7463eb),
	.w6(32'hbc14adb9),
	.w7(32'h3890146f),
	.w8(32'h3bc0906f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49c805),
	.w1(32'hbb77193b),
	.w2(32'h3acf5c7d),
	.w3(32'h3b5c0bfe),
	.w4(32'hb8aa193b),
	.w5(32'h3bd1fb58),
	.w6(32'h3b483375),
	.w7(32'hbb62c0fa),
	.w8(32'hb9964b67),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba192fec),
	.w1(32'hbc68e9d9),
	.w2(32'hbbf9dcef),
	.w3(32'h3a16f52d),
	.w4(32'hbc686222),
	.w5(32'hbbe4ee0f),
	.w6(32'h3aaa32f2),
	.w7(32'hbbaf75ef),
	.w8(32'h3b678888),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0fe908),
	.w1(32'hbb785d54),
	.w2(32'hbac69ff1),
	.w3(32'h3ba27ab2),
	.w4(32'hbac6f4e7),
	.w5(32'h3ae5852c),
	.w6(32'h3b6038dc),
	.w7(32'h3809840a),
	.w8(32'h3b15e39e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eeb94),
	.w1(32'h3b2e9333),
	.w2(32'hbc31ed35),
	.w3(32'h3ab327e4),
	.w4(32'h3c0a3ae7),
	.w5(32'hbb221a16),
	.w6(32'h3a1ec05e),
	.w7(32'h3b68b031),
	.w8(32'hbc0fc224),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8366ec),
	.w1(32'h3c141c27),
	.w2(32'h3b5b4241),
	.w3(32'hb93f9273),
	.w4(32'h3c5c5680),
	.w5(32'h3b165747),
	.w6(32'hbacfb99e),
	.w7(32'h3bdee42e),
	.w8(32'h3b5840f6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883c575),
	.w1(32'hbbafa277),
	.w2(32'hbad67cd5),
	.w3(32'h3b19eee9),
	.w4(32'hbb31a24f),
	.w5(32'h3afa7dd9),
	.w6(32'hbb166c6c),
	.w7(32'hbb9f5e90),
	.w8(32'h3c236699),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11e4c7),
	.w1(32'hbbeceaab),
	.w2(32'hbb965608),
	.w3(32'h3a8af620),
	.w4(32'hb8eda63c),
	.w5(32'h3b85e1f3),
	.w6(32'hb920172e),
	.w7(32'hbad51678),
	.w8(32'h3b5c264e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac48a1c),
	.w1(32'hba812253),
	.w2(32'h3ba0ecc0),
	.w3(32'h3bb9f94c),
	.w4(32'h3b402db8),
	.w5(32'h3c22b30f),
	.w6(32'h3bd2c2e9),
	.w7(32'h3b0f0386),
	.w8(32'h3bda052c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d92e),
	.w1(32'hbb560730),
	.w2(32'hbb5070ee),
	.w3(32'h3b57a1cf),
	.w4(32'hbafab536),
	.w5(32'hbbd106e9),
	.w6(32'h3b167ac2),
	.w7(32'hbbf3b1c2),
	.w8(32'hbb6895bc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc43ae),
	.w1(32'hbbca5b6d),
	.w2(32'hbbf04dc2),
	.w3(32'hbb964b14),
	.w4(32'hbbdd20a9),
	.w5(32'hbbd11316),
	.w6(32'hb8a86838),
	.w7(32'hbbcc7ac5),
	.w8(32'h3b529e8b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc75e5fa),
	.w1(32'hbbf8b747),
	.w2(32'h3b52cb7b),
	.w3(32'hbc94082a),
	.w4(32'hbc2a2827),
	.w5(32'h3aca2975),
	.w6(32'hbc7106a3),
	.w7(32'hbab33fce),
	.w8(32'h3b031c9e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39877985),
	.w1(32'hbbaa2c04),
	.w2(32'hbabec044),
	.w3(32'hb93bc491),
	.w4(32'hbb62e6b1),
	.w5(32'hba8e2c72),
	.w6(32'h3bbc388d),
	.w7(32'h3a799846),
	.w8(32'h3abf1408),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd4ee8),
	.w1(32'hbb569cde),
	.w2(32'hbb6eb6a8),
	.w3(32'hbc093f81),
	.w4(32'hbb26799e),
	.w5(32'hbb8f54b3),
	.w6(32'hbbbab605),
	.w7(32'h3a8e0d37),
	.w8(32'hba56c303),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a08d2),
	.w1(32'hbbb2c9c4),
	.w2(32'hbc10529c),
	.w3(32'hbbfd681e),
	.w4(32'hbbb5a86d),
	.w5(32'hbb908ca1),
	.w6(32'hbb9a4898),
	.w7(32'hbb7503f5),
	.w8(32'hbbdea3ca),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3db445),
	.w1(32'hba2acb92),
	.w2(32'h38ab3086),
	.w3(32'hbc53dcca),
	.w4(32'h3b9ed127),
	.w5(32'hbb0cc6f3),
	.w6(32'hbc5e1d63),
	.w7(32'h3ad0c318),
	.w8(32'h3850cb03),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1379f8),
	.w1(32'hbc0bdc4d),
	.w2(32'hbba5bc0e),
	.w3(32'h3c2a9f5c),
	.w4(32'hbc01174f),
	.w5(32'hbb8c2ac1),
	.w6(32'h3bf2b3b1),
	.w7(32'hbc16f268),
	.w8(32'h3b0e1f5a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f156b),
	.w1(32'h3b8b614f),
	.w2(32'h3be3f59d),
	.w3(32'hbbb938ec),
	.w4(32'h3b9975f4),
	.w5(32'h3c2bfcd8),
	.w6(32'hbb818ab3),
	.w7(32'h3afb5fd2),
	.w8(32'h3c12b7b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24cf97),
	.w1(32'h3b2d16ad),
	.w2(32'h3b994097),
	.w3(32'h3c04ddcc),
	.w4(32'h3b9e6073),
	.w5(32'h3bb92977),
	.w6(32'h3c0e8cfd),
	.w7(32'h3bfac630),
	.w8(32'h3c14d541),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99eb0b),
	.w1(32'h3bc0afae),
	.w2(32'h3bb14af1),
	.w3(32'h3b82aab7),
	.w4(32'h3bb71955),
	.w5(32'h3b024b4b),
	.w6(32'h3bbe6b63),
	.w7(32'h3c4367e2),
	.w8(32'h3bca6ffa),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9458fd),
	.w1(32'hbbdc7307),
	.w2(32'hbbd166ad),
	.w3(32'hb9831816),
	.w4(32'h3b39ae4d),
	.w5(32'h3b76c2bb),
	.w6(32'h3b3ba404),
	.w7(32'h3b8631cc),
	.w8(32'h3ba934ca),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e553d),
	.w1(32'hbb9fb3fb),
	.w2(32'h3c7dd9fb),
	.w3(32'h3b05b56f),
	.w4(32'hbbf448ff),
	.w5(32'h3c164871),
	.w6(32'hbb38a3f6),
	.w7(32'hbb86b51d),
	.w8(32'h3c8e17c3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c554d28),
	.w1(32'h3bb322fb),
	.w2(32'h3b78ba23),
	.w3(32'h3c142189),
	.w4(32'h3b36ee74),
	.w5(32'hba507d9c),
	.w6(32'h3b643348),
	.w7(32'h3a9f066f),
	.w8(32'h3bbc1fdc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98d573),
	.w1(32'hb9e80b28),
	.w2(32'hbb1d3111),
	.w3(32'h3b52419e),
	.w4(32'hbb2e2d41),
	.w5(32'hbb203a3b),
	.w6(32'h3c133f9e),
	.w7(32'hbba99bd6),
	.w8(32'hb8e1dd37),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d3e93),
	.w1(32'h3c252a70),
	.w2(32'h3be9cb42),
	.w3(32'hbb8266d3),
	.w4(32'h3c51d23e),
	.w5(32'h3b1a2fd8),
	.w6(32'h3b0710e9),
	.w7(32'h3c260fd0),
	.w8(32'h3aa0a81c),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba707a73),
	.w1(32'hbb4f9bf7),
	.w2(32'hbba579cc),
	.w3(32'hbab8965a),
	.w4(32'hbb460d4c),
	.w5(32'hbb8e8fb7),
	.w6(32'hbb799f97),
	.w7(32'hbbd47c6f),
	.w8(32'h3a6a96ef),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0c239),
	.w1(32'h3b995184),
	.w2(32'h3c0617f2),
	.w3(32'hbb8b18d5),
	.w4(32'h3beeeeb7),
	.w5(32'h3c240fc7),
	.w6(32'hbbbd27e6),
	.w7(32'h3b29ff83),
	.w8(32'h3bbe060e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4cc1),
	.w1(32'hbc0c181c),
	.w2(32'h39efcdb9),
	.w3(32'h3bbcf848),
	.w4(32'hbbb75532),
	.w5(32'h3bacd187),
	.w6(32'h3bc744ea),
	.w7(32'hbc041d03),
	.w8(32'h38b8effd),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f719),
	.w1(32'h3af6e851),
	.w2(32'hbb04f87c),
	.w3(32'h3bf1f205),
	.w4(32'hba3933f6),
	.w5(32'hbb4b3e3d),
	.w6(32'h3b8a114b),
	.w7(32'hbb4ea072),
	.w8(32'hbbfa838f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4eb95c),
	.w1(32'h3b84324d),
	.w2(32'h3ba520ed),
	.w3(32'hbb3082b2),
	.w4(32'hbb147ad9),
	.w5(32'hb9148bc8),
	.w6(32'hbc099417),
	.w7(32'hbab8b5c3),
	.w8(32'hba3bad8b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c1e04),
	.w1(32'hbbe63213),
	.w2(32'hbbebb268),
	.w3(32'h3b28dfbf),
	.w4(32'hbbabf39a),
	.w5(32'hbbcafb3d),
	.w6(32'hbad9e21d),
	.w7(32'hbb6f16f9),
	.w8(32'hba7b04f2),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56e520),
	.w1(32'hbbbcc9f8),
	.w2(32'h3aa9db93),
	.w3(32'hbc016681),
	.w4(32'hbc0c57bd),
	.w5(32'hbbd023f1),
	.w6(32'hbb7284ea),
	.w7(32'hbbf4259c),
	.w8(32'hba67ffcd),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bab88),
	.w1(32'h3c2b6901),
	.w2(32'h3b884570),
	.w3(32'h3b133c8b),
	.w4(32'h3c5a84b2),
	.w5(32'h3ba7b3b8),
	.w6(32'h3aa1182d),
	.w7(32'h3c0d2f54),
	.w8(32'h3ba69be8),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13df2a),
	.w1(32'h3b8ba2cb),
	.w2(32'h3b003e86),
	.w3(32'h3b06e1d3),
	.w4(32'h3c2877b7),
	.w5(32'hba9c4935),
	.w6(32'hbb273c67),
	.w7(32'h3bf0b7f6),
	.w8(32'hb8ffce10),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadca29b),
	.w1(32'h399df254),
	.w2(32'h3bfe0a16),
	.w3(32'hbb80e027),
	.w4(32'h3bbbaffd),
	.w5(32'h3c26820e),
	.w6(32'hbb7a4187),
	.w7(32'hba8eeb63),
	.w8(32'h3bb5d1d6),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb00033),
	.w1(32'hbadbcbf7),
	.w2(32'hbb161f8b),
	.w3(32'hbbc72a29),
	.w4(32'hbbb9777d),
	.w5(32'h3a571ecc),
	.w6(32'hbbca9cf2),
	.w7(32'hbb06d52b),
	.w8(32'h3b2e215d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ba4b7),
	.w1(32'h3c3ef48e),
	.w2(32'h3b4f689f),
	.w3(32'hbacb25d9),
	.w4(32'h3b8ad675),
	.w5(32'hbaa76ba2),
	.w6(32'h3bbb4c1f),
	.w7(32'h3adf5da7),
	.w8(32'hbbb26b07),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc85196),
	.w1(32'hba8b272e),
	.w2(32'hba321751),
	.w3(32'h3af83a41),
	.w4(32'hbb11a17e),
	.w5(32'hbb176d08),
	.w6(32'hb7732086),
	.w7(32'h3b15c526),
	.w8(32'hb9e7974c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd46ae),
	.w1(32'hbb9dc2f9),
	.w2(32'hba0b1a64),
	.w3(32'h3ac43bd5),
	.w4(32'hbb03f9f0),
	.w5(32'hb9431855),
	.w6(32'hb945b54c),
	.w7(32'hbb82732c),
	.w8(32'hba8b7cdf),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61b1d0),
	.w1(32'h3bac4099),
	.w2(32'h3c20da1d),
	.w3(32'h3b4675c1),
	.w4(32'hb88ff9c1),
	.w5(32'h3b7e83ff),
	.w6(32'hba0cc42c),
	.w7(32'h3b586504),
	.w8(32'h3b9d227f),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5053c9),
	.w1(32'hba891d37),
	.w2(32'hbae6b8ab),
	.w3(32'h3c1b10f5),
	.w4(32'h38e736f5),
	.w5(32'hba428b75),
	.w6(32'h3bb389a3),
	.w7(32'hba9c32a8),
	.w8(32'h3a4dcf0c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf3d27),
	.w1(32'h3b90ce6a),
	.w2(32'h3a3237ed),
	.w3(32'hbbcdc79b),
	.w4(32'hbad90592),
	.w5(32'hbb3aa26f),
	.w6(32'hbbbeb3ba),
	.w7(32'h39ea6070),
	.w8(32'hbb033272),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbe9f9),
	.w1(32'hbb6a9ebb),
	.w2(32'h3aef7962),
	.w3(32'hbb84cc34),
	.w4(32'hba7e33f2),
	.w5(32'hbb601f63),
	.w6(32'h3ba644ae),
	.w7(32'hbb06df39),
	.w8(32'hbb47468f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2656ff),
	.w1(32'h3b1ac04b),
	.w2(32'h3b7cf312),
	.w3(32'h39e4f2a8),
	.w4(32'h3be806e1),
	.w5(32'h3ae39baa),
	.w6(32'hba72b332),
	.w7(32'h3b7453e7),
	.w8(32'h3a40bfd5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42f07d),
	.w1(32'h3c6cf718),
	.w2(32'hbb995f85),
	.w3(32'h3941140b),
	.w4(32'h3cb60a69),
	.w5(32'h3b876ae8),
	.w6(32'hbb276dab),
	.w7(32'h3c875e4c),
	.w8(32'h3b8e0b87),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea71a1),
	.w1(32'hbb35a664),
	.w2(32'hbb316542),
	.w3(32'h3b3d12d9),
	.w4(32'hbb503e83),
	.w5(32'hbbcdd94c),
	.w6(32'h3acf90cd),
	.w7(32'h3b5330de),
	.w8(32'h39862e87),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc54037),
	.w1(32'hbb8a012c),
	.w2(32'h3a4352b8),
	.w3(32'hbbb55baf),
	.w4(32'hbb30bfab),
	.w5(32'h3a488d50),
	.w6(32'hbb937062),
	.w7(32'h3a7bb7a4),
	.w8(32'h3bc337b4),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1d597),
	.w1(32'h3ba3ca11),
	.w2(32'h3b6febd5),
	.w3(32'h3b390c33),
	.w4(32'h3c6b46bb),
	.w5(32'h3c388a7a),
	.w6(32'hb9401cdf),
	.w7(32'h3be814b1),
	.w8(32'h3b02b52c),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb909f757),
	.w1(32'hbb8f743a),
	.w2(32'hbc176b0e),
	.w3(32'h3bcd6e49),
	.w4(32'hbc2a02c6),
	.w5(32'hbc8bf821),
	.w6(32'hbb0615d6),
	.w7(32'hbc1f76a4),
	.w8(32'hbc25c7a9),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1cb9d3),
	.w1(32'hbbc3713b),
	.w2(32'hbbb1de22),
	.w3(32'hbc777519),
	.w4(32'hbba6959d),
	.w5(32'hbc175908),
	.w6(32'hbc537bd7),
	.w7(32'hbb13e494),
	.w8(32'hbb9a9571),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be4f7),
	.w1(32'h3bb4ad4d),
	.w2(32'hbbceeda4),
	.w3(32'hbc31799d),
	.w4(32'h3a6fd7ce),
	.w5(32'hbc050743),
	.w6(32'hbbece9bf),
	.w7(32'h3b9edb4d),
	.w8(32'hbb96e88a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb963a11),
	.w1(32'hbb7e5a3b),
	.w2(32'h3b0b1530),
	.w3(32'hbbceeb2d),
	.w4(32'hbbcad617),
	.w5(32'h3c0ee0b3),
	.w6(32'hbbf91b58),
	.w7(32'hbc0d264d),
	.w8(32'h39853e11),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca7c4),
	.w1(32'hbb0e163b),
	.w2(32'hbb7a2815),
	.w3(32'h3b997420),
	.w4(32'hbb4775d7),
	.w5(32'hbbbfef41),
	.w6(32'h3b033d9c),
	.w7(32'hbb8db9b5),
	.w8(32'hbb699cb2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c9741),
	.w1(32'hb9dc8959),
	.w2(32'h3bff41c2),
	.w3(32'hbb191aa6),
	.w4(32'hbb34bcd1),
	.w5(32'h3c40620c),
	.w6(32'hbbfe8fe5),
	.w7(32'hbb89c6cc),
	.w8(32'h3bb1c90e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6812),
	.w1(32'hbc319c3d),
	.w2(32'hbb8338c4),
	.w3(32'h3b28a431),
	.w4(32'hbb3922fc),
	.w5(32'h3bac4631),
	.w6(32'h3bc4f20a),
	.w7(32'hbc0b0a60),
	.w8(32'h3a37becf),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4ae3),
	.w1(32'hbc2919b9),
	.w2(32'hbbc1a69c),
	.w3(32'h3c8d710a),
	.w4(32'hbc3a291d),
	.w5(32'hbb10e725),
	.w6(32'h3c513a35),
	.w7(32'hbc1a55ab),
	.w8(32'h3ac64e0e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b8325),
	.w1(32'hbb662404),
	.w2(32'hbb3d41a9),
	.w3(32'hbc02ac1f),
	.w4(32'hb9fe4e04),
	.w5(32'hbbaf4008),
	.w6(32'hbb945496),
	.w7(32'hba06b6f1),
	.w8(32'hbbb3d2bd),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadbfd0),
	.w1(32'h3b620fc2),
	.w2(32'h3b49217e),
	.w3(32'h3b53d212),
	.w4(32'hb995cba1),
	.w5(32'h3add0d2e),
	.w6(32'h3b3311f0),
	.w7(32'hbb134a6a),
	.w8(32'h3b390f81),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b678c50),
	.w1(32'hba0b0b65),
	.w2(32'hb963942a),
	.w3(32'hba9d4832),
	.w4(32'hbb1b61b0),
	.w5(32'h3adb897a),
	.w6(32'hbade67fa),
	.w7(32'hbba210c4),
	.w8(32'hbb1df346),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f9a629),
	.w1(32'hbb59b2d7),
	.w2(32'hbb3cc01f),
	.w3(32'hbb7883e6),
	.w4(32'hbb9baba2),
	.w5(32'hbbdbc336),
	.w6(32'hbb81b63c),
	.w7(32'hbc3b56b8),
	.w8(32'hbbe16523),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb273656),
	.w1(32'h3b11f12c),
	.w2(32'h3859cfba),
	.w3(32'hbb0e6fb0),
	.w4(32'hbb40b5f9),
	.w5(32'hbb8ec59b),
	.w6(32'hbc025e13),
	.w7(32'h3b43188d),
	.w8(32'hbb7edd16),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d8888),
	.w1(32'hbb040672),
	.w2(32'h3ba11125),
	.w3(32'h3bae094b),
	.w4(32'hbaf21aad),
	.w5(32'hbb057fbb),
	.w6(32'h3bb9ad7a),
	.w7(32'hbb48a6c0),
	.w8(32'h3ae400ab),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0ffe3),
	.w1(32'h3c156d5a),
	.w2(32'h3a330ce2),
	.w3(32'hbbba077f),
	.w4(32'h3c799f65),
	.w5(32'h3b5054d8),
	.w6(32'hbbcce274),
	.w7(32'h3c399aa6),
	.w8(32'h390a53ae),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c62a7),
	.w1(32'h3bc3de7d),
	.w2(32'h3b61dcc1),
	.w3(32'h3b612aca),
	.w4(32'h3b2c7a28),
	.w5(32'h3b474b38),
	.w6(32'h3a8d2b04),
	.w7(32'h3bc218f3),
	.w8(32'h3b8c0643),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49d416),
	.w1(32'h3b76b96c),
	.w2(32'h3ad3cc9b),
	.w3(32'h3b27ab04),
	.w4(32'h3b19b83a),
	.w5(32'hbb321310),
	.w6(32'h3b97aee2),
	.w7(32'h3b3fa4aa),
	.w8(32'hbaffd37b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c6b24),
	.w1(32'hbadbc3ee),
	.w2(32'h3b7d0f2b),
	.w3(32'h3baab271),
	.w4(32'hba91efda),
	.w5(32'h3bb622d4),
	.w6(32'h3b69b8f2),
	.w7(32'h3a55098b),
	.w8(32'h3b798228),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3d01),
	.w1(32'hbbc99a5e),
	.w2(32'hbc17f15d),
	.w3(32'h3c233efa),
	.w4(32'hbbc5c047),
	.w5(32'hbc2d5217),
	.w6(32'h3bc4a0ae),
	.w7(32'hbc233160),
	.w8(32'hbc290753),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9593f),
	.w1(32'h3a7b29ba),
	.w2(32'hba9aee03),
	.w3(32'hbbc83156),
	.w4(32'h3b0584b8),
	.w5(32'h39b574a6),
	.w6(32'hbc150e76),
	.w7(32'h3b40b52f),
	.w8(32'h3ba505c1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d4c3),
	.w1(32'hbc50b77d),
	.w2(32'h39a476da),
	.w3(32'h3ae4b5b1),
	.w4(32'hbc5635aa),
	.w5(32'h3a860cbd),
	.w6(32'h3b079a64),
	.w7(32'hbcad55b8),
	.w8(32'hbb5c8bb7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cb1b0),
	.w1(32'hba4504c1),
	.w2(32'hba71c365),
	.w3(32'hbc6d727d),
	.w4(32'hbb7476e5),
	.w5(32'hbb387429),
	.w6(32'hbc9f1204),
	.w7(32'hbb41d756),
	.w8(32'hbb2516ed),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b464b42),
	.w1(32'h3a2ad410),
	.w2(32'hba1ab741),
	.w3(32'h39f74576),
	.w4(32'h3ab7961b),
	.w5(32'hbaf102dd),
	.w6(32'h39787886),
	.w7(32'hbaa1bf25),
	.w8(32'hbab4e506),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf26388),
	.w1(32'hbbaa61da),
	.w2(32'hbc3b4c2b),
	.w3(32'hbbbf55e1),
	.w4(32'hbb5d408c),
	.w5(32'hbc31b16e),
	.w6(32'hbc072166),
	.w7(32'hbb9df63d),
	.w8(32'hbc115d49),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3364c8),
	.w1(32'h3ac216ca),
	.w2(32'h3b1629e2),
	.w3(32'hbb703005),
	.w4(32'hb74c68ef),
	.w5(32'h3bafa371),
	.w6(32'hbbcd32b0),
	.w7(32'h3b3d8ff5),
	.w8(32'h3bc20931),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac0589),
	.w1(32'h3a2083e9),
	.w2(32'h3bcaf0e1),
	.w3(32'h39b4e97f),
	.w4(32'hbbbbbcd8),
	.w5(32'h3a31df7a),
	.w6(32'hb94b1ea9),
	.w7(32'hbbf8d0e7),
	.w8(32'hbb8b2635),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b276119),
	.w1(32'hbc18ec6e),
	.w2(32'hbc0be4b6),
	.w3(32'h3bbe0ec1),
	.w4(32'hbb926954),
	.w5(32'hb9801aad),
	.w6(32'h3aa362d9),
	.w7(32'hbc141033),
	.w8(32'hbb621c3f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e59ef),
	.w1(32'h3bea514a),
	.w2(32'hbc16fc07),
	.w3(32'hbb461a79),
	.w4(32'h3b6e7ffb),
	.w5(32'hbbedd9c3),
	.w6(32'hbb91d9f2),
	.w7(32'h3b869829),
	.w8(32'hbbd9a37b),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb5b29),
	.w1(32'h3af991d5),
	.w2(32'h3aa88f5f),
	.w3(32'h3b33882f),
	.w4(32'h38bf3cf9),
	.w5(32'h3a09addc),
	.w6(32'h3b44ded2),
	.w7(32'h3b18e8df),
	.w8(32'h3bb1fe2c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaabca6),
	.w1(32'h3b89b59a),
	.w2(32'hba1f555a),
	.w3(32'hba6e1b88),
	.w4(32'h3aa9c306),
	.w5(32'hbbdfbbf9),
	.w6(32'h3a49d690),
	.w7(32'h3a57c06e),
	.w8(32'hbb3ac4ee),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59cc74),
	.w1(32'h3ad2ddd6),
	.w2(32'h3b876217),
	.w3(32'h3b5315b9),
	.w4(32'h3bc7fa87),
	.w5(32'h3c1fb177),
	.w6(32'h3b0199d2),
	.w7(32'hba7f6397),
	.w8(32'h3b61075b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d60e3),
	.w1(32'hbbded306),
	.w2(32'hbbd7dcdc),
	.w3(32'h3bb7d671),
	.w4(32'hbbe48823),
	.w5(32'hbbc4b51e),
	.w6(32'h3bfc9b6c),
	.w7(32'hbb128645),
	.w8(32'h3a55b596),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d2eac),
	.w1(32'h3b5f4f53),
	.w2(32'h3c137e2f),
	.w3(32'hbc3d66e1),
	.w4(32'h3a24d16e),
	.w5(32'h3b26741e),
	.w6(32'hbbf93d56),
	.w7(32'h3bea8b71),
	.w8(32'h3bf96263),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a7b3),
	.w1(32'h38ede719),
	.w2(32'hbc03d905),
	.w3(32'hb9dd9506),
	.w4(32'hbb99e043),
	.w5(32'hbc065a57),
	.w6(32'hbaec112c),
	.w7(32'h39ea6b9f),
	.w8(32'hbc0cff96),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3b95e),
	.w1(32'h3b050cbc),
	.w2(32'h3bcc1c04),
	.w3(32'hbc45aa73),
	.w4(32'h3b27807c),
	.w5(32'h3c277b40),
	.w6(32'hbbcf172c),
	.w7(32'h3b060042),
	.w8(32'h3c168736),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e988de),
	.w1(32'hba7c8807),
	.w2(32'hbac097f1),
	.w3(32'h39887071),
	.w4(32'hba9d4b87),
	.w5(32'hbb3515a2),
	.w6(32'h3b2e2a5c),
	.w7(32'hbafa59f4),
	.w8(32'hbaa6139f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9723e),
	.w1(32'h3a8f9b72),
	.w2(32'h39593ce6),
	.w3(32'hbb87cfe3),
	.w4(32'hb95e8524),
	.w5(32'h39dcb955),
	.w6(32'hbb3c5375),
	.w7(32'hba82780c),
	.w8(32'h3990d635),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b432e91),
	.w1(32'hbb63bdaa),
	.w2(32'hba007db5),
	.w3(32'h3b1f8ded),
	.w4(32'hba82f7f2),
	.w5(32'h3b7cf623),
	.w6(32'h3b20f4e9),
	.w7(32'hbb2cf859),
	.w8(32'h3a9d65df),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5b22d),
	.w1(32'hba2cc9fb),
	.w2(32'h397899e8),
	.w3(32'hb9b4a1e7),
	.w4(32'hba2fa905),
	.w5(32'hbb01132f),
	.w6(32'h39d7af27),
	.w7(32'hbad33238),
	.w8(32'hbafece9d),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae10a55),
	.w1(32'hb9a4774d),
	.w2(32'h3ad9cd86),
	.w3(32'hbb10f6db),
	.w4(32'hbaa3cae6),
	.w5(32'h3adf75c0),
	.w6(32'hbadf25fd),
	.w7(32'hbb1e34b1),
	.w8(32'h3a9fdc72),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3479d1),
	.w1(32'h3908858e),
	.w2(32'h3b11a870),
	.w3(32'h3ad01094),
	.w4(32'h397f3aec),
	.w5(32'hbaafe5b3),
	.w6(32'hba62afcd),
	.w7(32'hba36f19d),
	.w8(32'h3a1bee58),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63b691),
	.w1(32'hbb0a8aae),
	.w2(32'hba8ad2ac),
	.w3(32'hba8489d1),
	.w4(32'hbb0c266b),
	.w5(32'hbb3f102b),
	.w6(32'hba132eea),
	.w7(32'hbb3c5ee0),
	.w8(32'hbab65faa),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3bf27),
	.w1(32'hbb2d438e),
	.w2(32'hbb4869f3),
	.w3(32'hba817589),
	.w4(32'hbaf75db5),
	.w5(32'h39b44b31),
	.w6(32'hb8afdfcc),
	.w7(32'hbb5c08d3),
	.w8(32'hbb88cfa2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdd72f),
	.w1(32'h3ae13889),
	.w2(32'h3ad9aa80),
	.w3(32'hba926bb2),
	.w4(32'h3a2187e4),
	.w5(32'h3b23bf00),
	.w6(32'hbbc10b31),
	.w7(32'h3a6fc492),
	.w8(32'h3a920fea),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b162c08),
	.w1(32'h3a930a3a),
	.w2(32'hba1d223e),
	.w3(32'hb925a509),
	.w4(32'h3ab004c9),
	.w5(32'h3a00ef11),
	.w6(32'h39da5847),
	.w7(32'hb8445ab2),
	.w8(32'h3aa0744d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b491a05),
	.w1(32'h3c1c4988),
	.w2(32'h3c3b69b6),
	.w3(32'h3bc337bd),
	.w4(32'h3c23c38d),
	.w5(32'h3bb93ad3),
	.w6(32'h3acea658),
	.w7(32'h3c4ce123),
	.w8(32'h3c2f2d05),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb49a1),
	.w1(32'h3ac57b45),
	.w2(32'h3afb32af),
	.w3(32'h3bb90e71),
	.w4(32'h373bf843),
	.w5(32'h3a5e4d7f),
	.w6(32'h3c1a29f5),
	.w7(32'hb82aab32),
	.w8(32'hb91b0511),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cc220d),
	.w1(32'hba2edaaf),
	.w2(32'hb9f5ecff),
	.w3(32'hbb12bb1d),
	.w4(32'hb8a0d86b),
	.w5(32'hba827a4f),
	.w6(32'hbac45b1b),
	.w7(32'h3a5f03aa),
	.w8(32'hba06009c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad956b7),
	.w1(32'hb8c648be),
	.w2(32'h3b815f05),
	.w3(32'hb9a1789a),
	.w4(32'h3b4fbbbb),
	.w5(32'h3bd34c43),
	.w6(32'h398f79ad),
	.w7(32'h3b035f18),
	.w8(32'h3b851a00),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c171),
	.w1(32'hbafe56e1),
	.w2(32'h3b4998c3),
	.w3(32'hb91b9e8b),
	.w4(32'hbb2a7bbf),
	.w5(32'h3b47378f),
	.w6(32'hbaf17036),
	.w7(32'hbb4ab0fd),
	.w8(32'h3b228f98),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea3247),
	.w1(32'hbb312a99),
	.w2(32'hba3fd5e7),
	.w3(32'hbb44c610),
	.w4(32'hbae15de1),
	.w5(32'h3a3fb0f6),
	.w6(32'hba7e4ff2),
	.w7(32'h3a9bc4b3),
	.w8(32'h3b18a6ea),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22c411),
	.w1(32'hbac95c7b),
	.w2(32'hba825310),
	.w3(32'hbabd2694),
	.w4(32'h3a7407a2),
	.w5(32'h3b1830cf),
	.w6(32'hbaf3f4c2),
	.w7(32'h3b5440b0),
	.w8(32'h39cbe943),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdc839),
	.w1(32'hbb3d58a0),
	.w2(32'hbb5588ed),
	.w3(32'h3a2e0739),
	.w4(32'hb9d94a85),
	.w5(32'hbac6b5a1),
	.w6(32'h3a24fda5),
	.w7(32'hba65bd21),
	.w8(32'hba0d96fa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61a458),
	.w1(32'h3b4c1ed6),
	.w2(32'h3b711811),
	.w3(32'hbb05bfab),
	.w4(32'h3b248bd9),
	.w5(32'h3b2c19ef),
	.w6(32'hba628d3a),
	.w7(32'h3a9c2fb2),
	.w8(32'h3b5925cb),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00f36e),
	.w1(32'hb8eefafb),
	.w2(32'hb9241c05),
	.w3(32'h3ac5fa25),
	.w4(32'hba9962f7),
	.w5(32'h3aff8d8b),
	.w6(32'h3b26739d),
	.w7(32'hbaa1f1f4),
	.w8(32'hbaf64ca8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33c372),
	.w1(32'h3b4be919),
	.w2(32'h3b956b4d),
	.w3(32'h38740963),
	.w4(32'h3b5cb7e0),
	.w5(32'h3b3a5d65),
	.w6(32'hbb2e347a),
	.w7(32'h3b18151f),
	.w8(32'h3a854dab),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd8759),
	.w1(32'h3b8243e8),
	.w2(32'h3bb76fe6),
	.w3(32'h3ad083e9),
	.w4(32'h3ba5b96d),
	.w5(32'h3be2f86e),
	.w6(32'h3b27e907),
	.w7(32'h3b9f2c45),
	.w8(32'h3bdb8bbd),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943f16),
	.w1(32'hba89dbb2),
	.w2(32'h3aa00bdc),
	.w3(32'h3b85d5ba),
	.w4(32'hbaa6911b),
	.w5(32'hbaa78142),
	.w6(32'h3bb4239b),
	.w7(32'h3a176bb3),
	.w8(32'h3b18d87f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92beea),
	.w1(32'h3ae82fd2),
	.w2(32'h3b992a96),
	.w3(32'h3a23a5b5),
	.w4(32'h3ac4e7ea),
	.w5(32'h3b49f914),
	.w6(32'h3ac0198d),
	.w7(32'h3a95ffd7),
	.w8(32'h3b2f341f),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a2f17),
	.w1(32'h3a90e22b),
	.w2(32'h3b3f9a9b),
	.w3(32'h3a8662a5),
	.w4(32'h3b4e222e),
	.w5(32'h3b0a7ad0),
	.w6(32'h3b4db13d),
	.w7(32'h3b03c2a3),
	.w8(32'h3b50a7d5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be5f6),
	.w1(32'h3aa6b5a5),
	.w2(32'hba5d8463),
	.w3(32'h3b221a9d),
	.w4(32'hbb3988f7),
	.w5(32'hbb32f346),
	.w6(32'h3b4c2b11),
	.w7(32'hbb74184b),
	.w8(32'hbb1db2ca),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85b390),
	.w1(32'hba1caa5c),
	.w2(32'hb9244ba6),
	.w3(32'hbb8d5261),
	.w4(32'h3976e1e7),
	.w5(32'h3ab75e44),
	.w6(32'hb8df400f),
	.w7(32'hba4a1e10),
	.w8(32'h39b0b125),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5ee3b),
	.w1(32'h3b123fff),
	.w2(32'hbac027c3),
	.w3(32'hba540797),
	.w4(32'h3ae7609e),
	.w5(32'hbae58cfe),
	.w6(32'h39af883f),
	.w7(32'h3b6ce433),
	.w8(32'hba0d69a8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054b8a),
	.w1(32'hb93d122b),
	.w2(32'hba829244),
	.w3(32'hbb7a417c),
	.w4(32'hb89220fc),
	.w5(32'hbbaa4521),
	.w6(32'hbbb9ca8e),
	.w7(32'hba8011b6),
	.w8(32'hbb985eee),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389272dc),
	.w1(32'h3b9bab02),
	.w2(32'h3bb1bf4e),
	.w3(32'hbb49263b),
	.w4(32'h3b192600),
	.w5(32'h3bc4979c),
	.w6(32'hbb5ff158),
	.w7(32'h39abb33f),
	.w8(32'h3b143c86),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88064a),
	.w1(32'h378dade3),
	.w2(32'h3aef4d6d),
	.w3(32'h3b931be9),
	.w4(32'h3b0792c9),
	.w5(32'h39d996cf),
	.w6(32'h3a9ed2a9),
	.w7(32'h38e7711e),
	.w8(32'h3a95d138),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a565b6b),
	.w1(32'hbb2be402),
	.w2(32'hbac1afcb),
	.w3(32'h3962282f),
	.w4(32'hbb7a9e5a),
	.w5(32'hba834155),
	.w6(32'h3a3235d2),
	.w7(32'hbb3d4f95),
	.w8(32'hbb633dbd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb801d9b),
	.w1(32'hba3659d1),
	.w2(32'h3a9986e0),
	.w3(32'hbbb0f515),
	.w4(32'h386c85a5),
	.w5(32'h3b161ead),
	.w6(32'hbb398f55),
	.w7(32'hb9f86dc0),
	.w8(32'h3b61059a),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9013ab),
	.w1(32'hba6049ef),
	.w2(32'h3b72e05a),
	.w3(32'h3ba8d29d),
	.w4(32'hbb541eb0),
	.w5(32'h3b008858),
	.w6(32'h3b526fbc),
	.w7(32'hba6fb851),
	.w8(32'hbab1eca8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ba6a7),
	.w1(32'h3aca0a4d),
	.w2(32'h38d2d408),
	.w3(32'hbb2f1ee7),
	.w4(32'h3b0a48b9),
	.w5(32'hba9eecef),
	.w6(32'hb7927b64),
	.w7(32'h3a84d88e),
	.w8(32'h3b1521ce),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8101ca),
	.w1(32'h3b0909e2),
	.w2(32'h3b505d5e),
	.w3(32'hba6aa216),
	.w4(32'h3b03efbb),
	.w5(32'h3ac9a2f7),
	.w6(32'hb8af5682),
	.w7(32'h3aee6ff1),
	.w8(32'h3b0f6ff7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa80b83),
	.w1(32'h3b1f4e79),
	.w2(32'h3ab2a6c4),
	.w3(32'h3a444f0f),
	.w4(32'h38655fc0),
	.w5(32'hba3ae859),
	.w6(32'h3a2ecd90),
	.w7(32'h3a77623a),
	.w8(32'hb9dda4a7),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af978a7),
	.w1(32'h3a46b935),
	.w2(32'h3779bee5),
	.w3(32'hbb0208e0),
	.w4(32'h3af78085),
	.w5(32'h381919e7),
	.w6(32'hba1025aa),
	.w7(32'h3b08d671),
	.w8(32'h39242e64),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3fcd2),
	.w1(32'hbb278b58),
	.w2(32'hb962e8b9),
	.w3(32'h3b1858a6),
	.w4(32'hbaf5568d),
	.w5(32'hbae80912),
	.w6(32'h3aa76a3f),
	.w7(32'hba8b21d5),
	.w8(32'h3a391fe1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8cfc4),
	.w1(32'h3acff16a),
	.w2(32'h3b69e6c9),
	.w3(32'hba82c6b2),
	.w4(32'hba8ac665),
	.w5(32'h3a24e5df),
	.w6(32'hbac5109b),
	.w7(32'h39dba8a4),
	.w8(32'h3a90026e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a281),
	.w1(32'hb959c204),
	.w2(32'hb975ab63),
	.w3(32'hbb0a2710),
	.w4(32'h39e88c67),
	.w5(32'h3a67fd8c),
	.w6(32'hbb3d3e73),
	.w7(32'h3aa08249),
	.w8(32'h393b2a66),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cb295),
	.w1(32'h3af5e874),
	.w2(32'h3b102b97),
	.w3(32'h3a589ecf),
	.w4(32'hbabf8207),
	.w5(32'h3a04de7e),
	.w6(32'h3ad1e3fe),
	.w7(32'h3a97bce0),
	.w8(32'h39b2bf2f),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa47e4a),
	.w1(32'hb914a4af),
	.w2(32'h3a928b53),
	.w3(32'hbb36069b),
	.w4(32'hb9dfc8b4),
	.w5(32'h3ab7cb17),
	.w6(32'hbb8c5a46),
	.w7(32'hba8b5dfd),
	.w8(32'h3956e2cf),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad91b6),
	.w1(32'h3b30e05a),
	.w2(32'h3b753982),
	.w3(32'h3adaa497),
	.w4(32'hbac05bff),
	.w5(32'hba3e035f),
	.w6(32'h39dff7c5),
	.w7(32'h3b46a01e),
	.w8(32'h3ba4c57c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11ea38),
	.w1(32'hbad44b59),
	.w2(32'h39c1428e),
	.w3(32'h3a2960f4),
	.w4(32'hbaa73fb1),
	.w5(32'h3b31c9f5),
	.w6(32'h391af5ed),
	.w7(32'h3a3ad6c8),
	.w8(32'h3b40525e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a453f68),
	.w1(32'hbab654a3),
	.w2(32'hbb25a20f),
	.w3(32'h3a396441),
	.w4(32'hbafe9358),
	.w5(32'hbb57e2a1),
	.w6(32'h3b348694),
	.w7(32'hbb6dbce4),
	.w8(32'hbb83f302),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014f65),
	.w1(32'h3a8fb547),
	.w2(32'h3b39bbd2),
	.w3(32'hbb102831),
	.w4(32'h3aa10de6),
	.w5(32'h3b5b042c),
	.w6(32'hbaea694e),
	.w7(32'hbaae61c4),
	.w8(32'hb82aa54a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac018c7),
	.w1(32'h3a642227),
	.w2(32'h3b2c2dea),
	.w3(32'hb9736abe),
	.w4(32'h3a8e14aa),
	.w5(32'h3a32b7cb),
	.w6(32'hba006ce2),
	.w7(32'h3b585f89),
	.w8(32'h3ac5d06c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a976e),
	.w1(32'hbb4eea07),
	.w2(32'hbb33e010),
	.w3(32'hba64320a),
	.w4(32'hbb7698a5),
	.w5(32'hbb1c351f),
	.w6(32'hb923a0c7),
	.w7(32'hbba66aa4),
	.w8(32'hbb0a5023),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacdb8d2),
	.w1(32'hba9b124c),
	.w2(32'h3a6f0198),
	.w3(32'hbb0a8b3f),
	.w4(32'hb9b0cb8a),
	.w5(32'h3b31153e),
	.w6(32'hbb5ed722),
	.w7(32'h384a3ce9),
	.w8(32'h3b67092b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb18bde),
	.w1(32'h39e4a2b4),
	.w2(32'h3b07aa52),
	.w3(32'h3bc38b18),
	.w4(32'h3a71a65f),
	.w5(32'hb9b506aa),
	.w6(32'h3bc27436),
	.w7(32'hba82ad3f),
	.w8(32'hb99bb1f4),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ce501),
	.w1(32'h3b612171),
	.w2(32'h3a503423),
	.w3(32'h3b1699d6),
	.w4(32'h3acd9fed),
	.w5(32'hbb45d8a7),
	.w6(32'h3b8a70f4),
	.w7(32'hba9bee99),
	.w8(32'h3a7b4bc6),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa0a4d9),
	.w1(32'h3af7ab47),
	.w2(32'h3a29a8c8),
	.w3(32'h3b4ae149),
	.w4(32'h3b0d09a4),
	.w5(32'hb9dc51f0),
	.w6(32'h3b5fdc16),
	.w7(32'h3a9278f3),
	.w8(32'h3a4c3942),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f4785),
	.w1(32'h3bc20ea7),
	.w2(32'h3c02c3d4),
	.w3(32'h3a2eacba),
	.w4(32'h3b9ed3fa),
	.w5(32'h3b9c25d7),
	.w6(32'h3b244f6f),
	.w7(32'h3bb1b776),
	.w8(32'h3bb143b2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86597c),
	.w1(32'h39037b73),
	.w2(32'h3b428e2a),
	.w3(32'h3b2bb405),
	.w4(32'hb9b96b2f),
	.w5(32'hb995c83e),
	.w6(32'h3ba5997e),
	.w7(32'hba624b42),
	.w8(32'h3b23ea02),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22ecde),
	.w1(32'h3b19f43a),
	.w2(32'h3ae23792),
	.w3(32'hba53457b),
	.w4(32'h37b24f49),
	.w5(32'h3a42f260),
	.w6(32'h3aa9fd4c),
	.w7(32'hba1dd074),
	.w8(32'h3a7d78a0),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9467b1a),
	.w1(32'hbaef3d7d),
	.w2(32'hbadd044e),
	.w3(32'hba569786),
	.w4(32'hbb2547ca),
	.w5(32'hbaf43e8c),
	.w6(32'hba2a7882),
	.w7(32'h3aa4e2e8),
	.w8(32'h3af554de),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ec6f1),
	.w1(32'hbb52f8f6),
	.w2(32'hbbb905e8),
	.w3(32'hba897718),
	.w4(32'hbad532fe),
	.w5(32'hbb8aa900),
	.w6(32'h3ae156c9),
	.w7(32'hbb76afba),
	.w8(32'hbb65c1b0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule