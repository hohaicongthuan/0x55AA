module layer_10_featuremap_295(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bf7e7),
	.w1(32'h39725e60),
	.w2(32'hb97ed448),
	.w3(32'h390e5331),
	.w4(32'hb9c6413d),
	.w5(32'h3a0c30e4),
	.w6(32'h3942bdc8),
	.w7(32'hb9b56e6f),
	.w8(32'h388e5ca8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39823802),
	.w1(32'h390b34f9),
	.w2(32'h39005e71),
	.w3(32'h39bc4bc3),
	.w4(32'h39a69d89),
	.w5(32'hba7e57d5),
	.w6(32'h3980ac1f),
	.w7(32'h3914e73c),
	.w8(32'hb9071cbb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a9e0f),
	.w1(32'hb91ef654),
	.w2(32'hb922ec38),
	.w3(32'hba616000),
	.w4(32'hba0cead7),
	.w5(32'h38ab635c),
	.w6(32'h39b56e16),
	.w7(32'h3896d2ba),
	.w8(32'h399608f3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f58f68),
	.w1(32'h39bd5584),
	.w2(32'h3a3a7b01),
	.w3(32'h391df923),
	.w4(32'h3a200dea),
	.w5(32'h3981777b),
	.w6(32'h39fe4ca7),
	.w7(32'h3a271dcc),
	.w8(32'hb98f0eae),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a007a26),
	.w1(32'h39b2cec1),
	.w2(32'h395e9ac5),
	.w3(32'h395ddaf9),
	.w4(32'h39719f01),
	.w5(32'hb7594674),
	.w6(32'hba992c72),
	.w7(32'hba5d7d44),
	.w8(32'h393b5d9e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cfbf6),
	.w1(32'h3984acc9),
	.w2(32'h39788fe8),
	.w3(32'h39792ba2),
	.w4(32'h39a13eab),
	.w5(32'h3a104fc0),
	.w6(32'h390a22f0),
	.w7(32'h36a35aaa),
	.w8(32'h39d2b31b),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35d8bb),
	.w1(32'h39ced3a4),
	.w2(32'h3a03a478),
	.w3(32'h3a244c7d),
	.w4(32'h3a2281fe),
	.w5(32'h39a20b7d),
	.w6(32'h39ca04c4),
	.w7(32'h39c08850),
	.w8(32'h39d62055),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fe6bea),
	.w1(32'h3969f2e8),
	.w2(32'h3a3b675c),
	.w3(32'h3901bfdb),
	.w4(32'h3a06bcb2),
	.w5(32'h38d49690),
	.w6(32'h39acaca7),
	.w7(32'h3a819e84),
	.w8(32'h397f615a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9be70),
	.w1(32'h39825908),
	.w2(32'h38da4704),
	.w3(32'h395c1a05),
	.w4(32'h39bd6efa),
	.w5(32'h393507ad),
	.w6(32'h38eceedb),
	.w7(32'h3985ec55),
	.w8(32'h39aed7a4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fef922),
	.w1(32'h397e5660),
	.w2(32'h392505e0),
	.w3(32'h39cfbb5e),
	.w4(32'h39ff9abb),
	.w5(32'hb97b10f3),
	.w6(32'h398e4406),
	.w7(32'h397c636a),
	.w8(32'h392ba5f8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a57fd),
	.w1(32'h39c8ce2c),
	.w2(32'h39feb0c1),
	.w3(32'hb8f02f40),
	.w4(32'h3950059d),
	.w5(32'hb9740f79),
	.w6(32'h38f4b953),
	.w7(32'h398afdfc),
	.w8(32'h39abf9fc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d88d3d),
	.w1(32'hba5ac827),
	.w2(32'hbaa19c54),
	.w3(32'hb99b22b0),
	.w4(32'hb83f86e9),
	.w5(32'hba6b58f2),
	.w6(32'h3a2bf338),
	.w7(32'h39276b83),
	.w8(32'hba8610d9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab16cdc),
	.w1(32'hbae0bb51),
	.w2(32'hbaad478d),
	.w3(32'hba7c38b5),
	.w4(32'hbaabcec6),
	.w5(32'h385aa44a),
	.w6(32'hbab151cd),
	.w7(32'hbaa9f1c9),
	.w8(32'h39ab6894),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a37e8),
	.w1(32'hb9baaeb9),
	.w2(32'hba2eb82a),
	.w3(32'hba4f68d6),
	.w4(32'hba76eacf),
	.w5(32'hba18cc23),
	.w6(32'hba7b65fd),
	.w7(32'hba9c65c6),
	.w8(32'hb9ca82f1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91581b2),
	.w1(32'hb883ee4c),
	.w2(32'h38dd0d10),
	.w3(32'hb92a0990),
	.w4(32'h3a0d8c0e),
	.w5(32'hb777cb55),
	.w6(32'hb7994882),
	.w7(32'h388d7cb0),
	.w8(32'h39073f16),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27ca7a),
	.w1(32'h39e58bee),
	.w2(32'h38bfeee9),
	.w3(32'h378f28e2),
	.w4(32'hb9816d55),
	.w5(32'h39b37571),
	.w6(32'h39d1a266),
	.w7(32'h3969ecfa),
	.w8(32'h38b54614),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3961a062),
	.w1(32'h3a08b55c),
	.w2(32'h3a0895d3),
	.w3(32'h39d80121),
	.w4(32'h39c2d178),
	.w5(32'hb9fbf0e3),
	.w6(32'h3a21f1bb),
	.w7(32'h3a0d9a67),
	.w8(32'hba4bf911),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fbe8d),
	.w1(32'hba6b2991),
	.w2(32'hb9faa8ef),
	.w3(32'hba0853a1),
	.w4(32'hba00f0a5),
	.w5(32'hba517424),
	.w6(32'hb9d2894e),
	.w7(32'hba30ffe8),
	.w8(32'hba47a442),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6007a9),
	.w1(32'hba419c2e),
	.w2(32'hb93711f7),
	.w3(32'hba1d6ecd),
	.w4(32'hba4ce683),
	.w5(32'hb9ab37f2),
	.w6(32'hba7b22ca),
	.w7(32'hba362d64),
	.w8(32'hba20bed0),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aec60a),
	.w1(32'h39478558),
	.w2(32'hb991c744),
	.w3(32'hb941e0f7),
	.w4(32'hb8dfe8d9),
	.w5(32'hb8f4313d),
	.w6(32'hba2326c2),
	.w7(32'hb9d4f98e),
	.w8(32'h396530e3),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72de2c),
	.w1(32'h39b87632),
	.w2(32'hb87611a1),
	.w3(32'hb97861e0),
	.w4(32'hb95a036d),
	.w5(32'h3a5c9b2d),
	.w6(32'hb943f32e),
	.w7(32'h391a113a),
	.w8(32'h3a85dcd1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa75118),
	.w1(32'h3aa6dd02),
	.w2(32'h3ac5b5bf),
	.w3(32'h3a9169ad),
	.w4(32'h3ac52639),
	.w5(32'h391171eb),
	.w6(32'h3a865766),
	.w7(32'h3acac992),
	.w8(32'h37eab165),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba253977),
	.w1(32'hba6d186b),
	.w2(32'hba748bae),
	.w3(32'hb9110f75),
	.w4(32'hb95fcb8c),
	.w5(32'h39472e88),
	.w6(32'h39180ae7),
	.w7(32'hb9ea6908),
	.w8(32'h39d51bf9),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ae85e),
	.w1(32'hba03a933),
	.w2(32'hba4eb7bc),
	.w3(32'h37ddcba8),
	.w4(32'hb90871f1),
	.w5(32'hb9b82000),
	.w6(32'h398ff292),
	.w7(32'h393aa62d),
	.w8(32'hba7dcfd4),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb8966),
	.w1(32'hb9823e2d),
	.w2(32'hb9849d13),
	.w3(32'hb9655291),
	.w4(32'hb9cfb6ae),
	.w5(32'h390a44c5),
	.w6(32'hba0bb220),
	.w7(32'hb98f7d6b),
	.w8(32'h39a3707e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3995155e),
	.w1(32'h3a617779),
	.w2(32'h3a1f05ff),
	.w3(32'h3a35deda),
	.w4(32'h3a402523),
	.w5(32'hb88c6aaa),
	.w6(32'h3a51a9b1),
	.w7(32'h3a828769),
	.w8(32'h39578e6b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901260f),
	.w1(32'h3a3dd7bd),
	.w2(32'h399484bf),
	.w3(32'h39ee575d),
	.w4(32'h394675db),
	.w5(32'h39a87807),
	.w6(32'h3a85ef48),
	.w7(32'h3a17a454),
	.w8(32'h39cf0cf6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a478645),
	.w1(32'h39f2c298),
	.w2(32'hb9a50eae),
	.w3(32'h39c5918d),
	.w4(32'h38a5bd92),
	.w5(32'h399aa7ad),
	.w6(32'h39010d02),
	.w7(32'hb9aa83c1),
	.w8(32'hb721450a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02143f),
	.w1(32'h3a32d1c2),
	.w2(32'h39ae7f1a),
	.w3(32'h39a8d2ff),
	.w4(32'h39dba05f),
	.w5(32'hba08247d),
	.w6(32'hb86a1f6a),
	.w7(32'h38f1edeb),
	.w8(32'hb9a136f9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b232a4),
	.w1(32'h39c38ae6),
	.w2(32'h39bcb074),
	.w3(32'h399ddc0d),
	.w4(32'h391b6f26),
	.w5(32'hba20d003),
	.w6(32'h3a09b989),
	.w7(32'h396985dd),
	.w8(32'hba400ba6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c184a7),
	.w1(32'hb89bf255),
	.w2(32'hb935fc27),
	.w3(32'h38c53903),
	.w4(32'h3a1bbdca),
	.w5(32'hba36de8d),
	.w6(32'hb873ceac),
	.w7(32'hb972f85e),
	.w8(32'h3a068c49),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbc05d),
	.w1(32'h3952b385),
	.w2(32'h3a43d3a8),
	.w3(32'hba5646d1),
	.w4(32'hb9076a68),
	.w5(32'hba1e03ed),
	.w6(32'h3a155ae0),
	.w7(32'h3a386f58),
	.w8(32'hb9fc5c2f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38868f44),
	.w1(32'h39e254da),
	.w2(32'h3967ab12),
	.w3(32'hb949f6ca),
	.w4(32'hba15957f),
	.w5(32'hb9e95a03),
	.w6(32'hb9d08f7a),
	.w7(32'h39c442b2),
	.w8(32'hba9d4771),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa73098),
	.w1(32'hba96f19e),
	.w2(32'hba80464f),
	.w3(32'hba0e7cec),
	.w4(32'hba26b681),
	.w5(32'hb9f17a05),
	.w6(32'hba69020d),
	.w7(32'hba9e2750),
	.w8(32'hb9a3ddfb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f0a68),
	.w1(32'hb991e6a1),
	.w2(32'hb9162e94),
	.w3(32'hb9d2a2e5),
	.w4(32'hba0b51b5),
	.w5(32'hba15a928),
	.w6(32'hba404c2a),
	.w7(32'hb9fd798d),
	.w8(32'hba8623e2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f76c95),
	.w1(32'hb9fa1763),
	.w2(32'hb980cec8),
	.w3(32'hba1b61cb),
	.w4(32'hb9ee6ff1),
	.w5(32'h38027d45),
	.w6(32'hba0390b5),
	.w7(32'hba1c0641),
	.w8(32'hba346e04),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399138c0),
	.w1(32'h3a7df064),
	.w2(32'h3a136927),
	.w3(32'hb91f6961),
	.w4(32'hb9c50dbf),
	.w5(32'hb926e7d3),
	.w6(32'h39eb40d7),
	.w7(32'h3a631782),
	.w8(32'h39d5082e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38843d10),
	.w1(32'h3a009822),
	.w2(32'h3a08395c),
	.w3(32'h396a8c14),
	.w4(32'h3950c93a),
	.w5(32'hba0575be),
	.w6(32'h399dd3d7),
	.w7(32'h374f9ed0),
	.w8(32'hba83ca37),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88deb0b),
	.w1(32'h37b6a716),
	.w2(32'hba09160e),
	.w3(32'hb9954b51),
	.w4(32'h3998fa11),
	.w5(32'h39eedd3e),
	.w6(32'hba82f739),
	.w7(32'hbaa4e830),
	.w8(32'h39d0c5c6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eeddd6),
	.w1(32'hb9822ae5),
	.w2(32'hb7330bda),
	.w3(32'h39ac2978),
	.w4(32'h39bc1c50),
	.w5(32'h3894a4e7),
	.w6(32'hba840c9e),
	.w7(32'h39b58702),
	.w8(32'h383b3ed0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953fefb),
	.w1(32'hb9e4b213),
	.w2(32'hb9943010),
	.w3(32'hb9b4336f),
	.w4(32'hba27d175),
	.w5(32'h3a822b63),
	.w6(32'hb9c351ff),
	.w7(32'hba13ca27),
	.w8(32'h3aa26f38),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e3f1b),
	.w1(32'h3ac70f3b),
	.w2(32'h3aa0f9ba),
	.w3(32'h3aadf09f),
	.w4(32'h3ad02b21),
	.w5(32'hba336781),
	.w6(32'h3ac55d2d),
	.w7(32'h3ad7d044),
	.w8(32'hb9e0d898),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba944d6a),
	.w1(32'hba84d79d),
	.w2(32'hba819284),
	.w3(32'hba94badc),
	.w4(32'hba88b2d9),
	.w5(32'hbaca2b2d),
	.w6(32'hba25eabc),
	.w7(32'hba82da72),
	.w8(32'hbaa78ca7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae9aa0),
	.w1(32'hba632842),
	.w2(32'hba3c5d70),
	.w3(32'hbaa9e1af),
	.w4(32'hba8cfc93),
	.w5(32'hb9de4e31),
	.w6(32'hb9d873a6),
	.w7(32'hba607ec9),
	.w8(32'h3854dea0),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7241d),
	.w1(32'hb8543fb2),
	.w2(32'hb953a9fd),
	.w3(32'hba48633e),
	.w4(32'hba4c311b),
	.w5(32'h3aa13a61),
	.w6(32'hb9defae2),
	.w7(32'hb91c26b1),
	.w8(32'h3a9265cd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa98caf),
	.w1(32'h3a810b83),
	.w2(32'h3a92cbfa),
	.w3(32'h3ab88715),
	.w4(32'h3a6444ab),
	.w5(32'h38f187b8),
	.w6(32'h3a73b4b5),
	.w7(32'h3aa49e4e),
	.w8(32'h3a6c4060),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa45456),
	.w1(32'h3aaccdd2),
	.w2(32'h3a54ec00),
	.w3(32'h3a1a6c79),
	.w4(32'h39816f72),
	.w5(32'h3a172b7c),
	.w6(32'h3a692572),
	.w7(32'h3a713d2d),
	.w8(32'h3a2b92f6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a947ef6),
	.w1(32'h3abcd38f),
	.w2(32'h3ac32089),
	.w3(32'h3aa53dcc),
	.w4(32'h3adf13f7),
	.w5(32'hbac5b680),
	.w6(32'h3aa18843),
	.w7(32'h3acbc664),
	.w8(32'hbab7c8d6),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeef31c),
	.w1(32'hbb01bdbe),
	.w2(32'hbac7280f),
	.w3(32'hbacf7d74),
	.w4(32'hbab98c94),
	.w5(32'h3a7fae8c),
	.w6(32'hbaca65af),
	.w7(32'hbaecf46f),
	.w8(32'h3a89b3fa),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8cfed),
	.w1(32'h3aa7a204),
	.w2(32'h3ac32e6a),
	.w3(32'h3aa2cf46),
	.w4(32'h3abed65b),
	.w5(32'hba727c14),
	.w6(32'h3a92e959),
	.w7(32'h3aad1eeb),
	.w8(32'hbab66eaf),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c8260),
	.w1(32'hb8cace0b),
	.w2(32'hb8b94770),
	.w3(32'hb9a34946),
	.w4(32'hba4f7dae),
	.w5(32'hb85963fd),
	.w6(32'hba7509c2),
	.w7(32'hba50d0ce),
	.w8(32'hb9d881e9),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4919b7),
	.w1(32'hba6a84b7),
	.w2(32'hb9b1397e),
	.w3(32'hba467c3c),
	.w4(32'hb91fcac7),
	.w5(32'hba83b9a3),
	.w6(32'hba09e802),
	.w7(32'hba03ce64),
	.w8(32'hb8b94f1e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395965f6),
	.w1(32'hb95f8baa),
	.w2(32'hb9751180),
	.w3(32'hb9cab093),
	.w4(32'hb9f48f4f),
	.w5(32'h39d4f63e),
	.w6(32'h37dd97f3),
	.w7(32'hb9bea5c8),
	.w8(32'h399c4ff6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39538447),
	.w1(32'h3a64d5dd),
	.w2(32'hb971cf60),
	.w3(32'h3a407017),
	.w4(32'hb9d34563),
	.w5(32'h38e2adcf),
	.w6(32'h3a916d55),
	.w7(32'h39d398a0),
	.w8(32'hb8069867),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac7ec2),
	.w1(32'h392cc8a4),
	.w2(32'hb719cb5b),
	.w3(32'hb862887c),
	.w4(32'h38dd936e),
	.w5(32'hb9b5a6c6),
	.w6(32'hb9d6fb66),
	.w7(32'hb8920502),
	.w8(32'hb9cffac6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37540e23),
	.w1(32'hb8a1a999),
	.w2(32'h393b1926),
	.w3(32'hba0a0166),
	.w4(32'hb9085d4a),
	.w5(32'h38abf48e),
	.w6(32'hba84007a),
	.w7(32'hba2263b0),
	.w8(32'hb78078e5),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a0edf5),
	.w1(32'h37667456),
	.w2(32'h37b5876a),
	.w3(32'hb91496e8),
	.w4(32'hb83d2693),
	.w5(32'h3679e2c0),
	.w6(32'hba019272),
	.w7(32'hb9524d35),
	.w8(32'h39de8f59),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a535e48),
	.w1(32'h3a9f69f2),
	.w2(32'h38a2c70e),
	.w3(32'h3a3ccb8b),
	.w4(32'hb790d05a),
	.w5(32'h3a7ba0b8),
	.w6(32'h3a99cb51),
	.w7(32'hb9d653fe),
	.w8(32'h3a7a757c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a968d47),
	.w1(32'h3a873084),
	.w2(32'h3a9615bc),
	.w3(32'h3a9a1bca),
	.w4(32'h3aaac81a),
	.w5(32'h396f4dec),
	.w6(32'h3a85ac95),
	.w7(32'h3a9291f3),
	.w8(32'h3a54f30f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cea58),
	.w1(32'h3ac3218a),
	.w2(32'h3aba0e98),
	.w3(32'h3a970139),
	.w4(32'h3aaa45fe),
	.w5(32'hb9b75c31),
	.w6(32'h3a809e11),
	.w7(32'h3a9f239e),
	.w8(32'hba21da2e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b019f),
	.w1(32'h397c364c),
	.w2(32'hb91492d1),
	.w3(32'hb9c4a21e),
	.w4(32'h38b97491),
	.w5(32'h3a6dbd03),
	.w6(32'hb9f33369),
	.w7(32'hba263910),
	.w8(32'h3a3247c1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9504f3),
	.w1(32'h3a9915a8),
	.w2(32'h3aa2a56a),
	.w3(32'h3a9fb83a),
	.w4(32'h3aaaa142),
	.w5(32'hb9d60037),
	.w6(32'h3aaaba39),
	.w7(32'h3ac8ba32),
	.w8(32'hba3c3bc3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e7549),
	.w1(32'hba0386a4),
	.w2(32'hb9a6ac03),
	.w3(32'hb9cc401f),
	.w4(32'h38e27614),
	.w5(32'hb9a8a48c),
	.w6(32'hba807ad6),
	.w7(32'hb9e88704),
	.w8(32'hba4923fe),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba458a3d),
	.w1(32'hba0f1e3a),
	.w2(32'hba02fc3c),
	.w3(32'hba008df8),
	.w4(32'hba0a3e04),
	.w5(32'hba838b42),
	.w6(32'hba88313a),
	.w7(32'hba6b3d8a),
	.w8(32'hba261c27),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba188ce9),
	.w1(32'h390e2010),
	.w2(32'hb9d9c0fb),
	.w3(32'hba51a50a),
	.w4(32'hba858fe3),
	.w5(32'hb9bd7763),
	.w6(32'hba810ece),
	.w7(32'hbaa94160),
	.w8(32'hba0dc882),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39011bfc),
	.w1(32'hb891bf6d),
	.w2(32'hb99759b6),
	.w3(32'hb928588f),
	.w4(32'h39e3988a),
	.w5(32'h396332b3),
	.w6(32'hb9fe1db1),
	.w7(32'hb9eb0645),
	.w8(32'hb8805424),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39956719),
	.w1(32'h3994bbd4),
	.w2(32'h3a0815ff),
	.w3(32'h39e164eb),
	.w4(32'h397d9a32),
	.w5(32'hbaabd128),
	.w6(32'h387963f6),
	.w7(32'h39428e63),
	.w8(32'hbaa586be),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba781699),
	.w1(32'hb689e672),
	.w2(32'hb9c2a347),
	.w3(32'hba0f6b7e),
	.w4(32'hb9ca6f4b),
	.w5(32'hb8bc8109),
	.w6(32'h39a38c60),
	.w7(32'h36fac513),
	.w8(32'hb8098ca2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a717b7),
	.w1(32'h39fb34a1),
	.w2(32'hb9588084),
	.w3(32'hb822b169),
	.w4(32'hba004d0e),
	.w5(32'hba575d74),
	.w6(32'hb9165b7f),
	.w7(32'hb9cf0fc1),
	.w8(32'hba957701),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaca38e),
	.w1(32'hbb0ad922),
	.w2(32'hbaa096bb),
	.w3(32'hbab35a7a),
	.w4(32'hba708045),
	.w5(32'hba418e29),
	.w6(32'hbad1cc37),
	.w7(32'hbad1a0a3),
	.w8(32'hb9d14da4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca33c5),
	.w1(32'hb8e34f7f),
	.w2(32'hb86ee2df),
	.w3(32'hba108815),
	.w4(32'hb9cf3483),
	.w5(32'h399c8d25),
	.w6(32'h396e7929),
	.w7(32'h397c3666),
	.w8(32'h39555628),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2550d8),
	.w1(32'hb95e4d6d),
	.w2(32'h391e0a20),
	.w3(32'h3872d394),
	.w4(32'h39c22d0b),
	.w5(32'h398dba03),
	.w6(32'h3a306035),
	.w7(32'h399a61e2),
	.w8(32'hb98f945d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba04f71d),
	.w1(32'hb4459bd3),
	.w2(32'hba565308),
	.w3(32'h3a463264),
	.w4(32'h3a5fa34f),
	.w5(32'h37e8d754),
	.w6(32'h3a411bb0),
	.w7(32'hb91a2072),
	.w8(32'hba4fb0af),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba624613),
	.w1(32'hba31afc9),
	.w2(32'hba266a99),
	.w3(32'hb9a92030),
	.w4(32'h39107b53),
	.w5(32'hb9143392),
	.w6(32'hba8e8718),
	.w7(32'hb98dc394),
	.w8(32'hb843c8a1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38630d12),
	.w1(32'h39208a60),
	.w2(32'hb95f9767),
	.w3(32'hb9cc889c),
	.w4(32'hba81ab29),
	.w5(32'hbabf184a),
	.w6(32'hb9abd3a3),
	.w7(32'hba14151f),
	.w8(32'hbacc3341),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7bcf0),
	.w1(32'hbb0c31d7),
	.w2(32'hbae91c37),
	.w3(32'hbae740d5),
	.w4(32'hbacc8783),
	.w5(32'h39dbe5d6),
	.w6(32'hbb0cfc40),
	.w7(32'hbb00bbb7),
	.w8(32'h36f161c2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a95a0),
	.w1(32'hb9f5a209),
	.w2(32'hb985d420),
	.w3(32'h399b060f),
	.w4(32'h3940ff83),
	.w5(32'hb9ef300a),
	.w6(32'hb837c343),
	.w7(32'hba0a4a1a),
	.w8(32'hba95be50),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65fff5),
	.w1(32'hbabcdb84),
	.w2(32'hbaa4559c),
	.w3(32'hba69da35),
	.w4(32'hba8dcb34),
	.w5(32'hb9e7b0c2),
	.w6(32'hbab34f38),
	.w7(32'hbad8aa49),
	.w8(32'hb9f3732a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d23a9),
	.w1(32'hba1f4fc5),
	.w2(32'hb985d227),
	.w3(32'hb9997b68),
	.w4(32'hb976f6d4),
	.w5(32'h39128353),
	.w6(32'hb9da25db),
	.w7(32'hb94a8d0b),
	.w8(32'hb9a87fea),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de476d),
	.w1(32'h396ea602),
	.w2(32'h3977f156),
	.w3(32'h39c7c3e1),
	.w4(32'h39d4de3b),
	.w5(32'hba353e5d),
	.w6(32'h39062048),
	.w7(32'hb85e6bf6),
	.w8(32'hba1256cc),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba749e02),
	.w1(32'hbad6618d),
	.w2(32'hbaae9be1),
	.w3(32'hba9ef7c3),
	.w4(32'hba228734),
	.w5(32'hba1a73b5),
	.w6(32'hbad7d065),
	.w7(32'hb9d82b34),
	.w8(32'hba6b55d9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba939949),
	.w1(32'hba99ee75),
	.w2(32'hba7be21d),
	.w3(32'hba58871d),
	.w4(32'hba20a80a),
	.w5(32'h39899e76),
	.w6(32'hba8345d5),
	.w7(32'hba92dc2c),
	.w8(32'hb6cf7914),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1971a8),
	.w1(32'hb98fdf16),
	.w2(32'hba2b6ae3),
	.w3(32'hb82cf0bf),
	.w4(32'hba0c7b90),
	.w5(32'hba939ef6),
	.w6(32'hb8cc3034),
	.w7(32'hb9ec057b),
	.w8(32'hba7600e6),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36475d),
	.w1(32'hb8953fd1),
	.w2(32'hb7d2b79a),
	.w3(32'hba23e6db),
	.w4(32'hb9c5b732),
	.w5(32'hb95e2b0b),
	.w6(32'hb9335276),
	.w7(32'h398e6c70),
	.w8(32'hba2a71de),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54cf29),
	.w1(32'hba57fec7),
	.w2(32'hba74f5f3),
	.w3(32'hba45d565),
	.w4(32'hba5b1f2f),
	.w5(32'hb869028c),
	.w6(32'hba3f421f),
	.w7(32'hba1188f1),
	.w8(32'h38e42c70),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d28f),
	.w1(32'h3a1a646d),
	.w2(32'h3a53fc8a),
	.w3(32'h3a000fb7),
	.w4(32'h39d21992),
	.w5(32'h396ec98a),
	.w6(32'h39194d64),
	.w7(32'hb849f1ec),
	.w8(32'h3a0d7c65),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394614f4),
	.w1(32'h3a01e2d4),
	.w2(32'hba7e6153),
	.w3(32'h3a338df3),
	.w4(32'hb9ac2886),
	.w5(32'h3a27a1af),
	.w6(32'h3ab64678),
	.w7(32'hba0e4089),
	.w8(32'hb9a95019),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39030e97),
	.w1(32'hb9597d06),
	.w2(32'hb94663f4),
	.w3(32'h3a1e0d47),
	.w4(32'h3a1ce488),
	.w5(32'h3903a1df),
	.w6(32'hb9ddb244),
	.w7(32'hb9a44fbd),
	.w8(32'hb8c63745),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39418c64),
	.w1(32'h3957a448),
	.w2(32'h399feac8),
	.w3(32'h39eeff69),
	.w4(32'h3a0b92aa),
	.w5(32'hb95fbfc7),
	.w6(32'h39aff03d),
	.w7(32'h39622568),
	.w8(32'hb944c0b0),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d20a13),
	.w1(32'hba0bdd7a),
	.w2(32'h399c5559),
	.w3(32'hba277fe2),
	.w4(32'hb8e94552),
	.w5(32'h39e26e4e),
	.w6(32'hba518126),
	.w7(32'hb927172c),
	.w8(32'hb8fe58ec),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ff569),
	.w1(32'hba537f38),
	.w2(32'hb9931814),
	.w3(32'hb9292a4a),
	.w4(32'hb78f0ec7),
	.w5(32'hba72e1ab),
	.w6(32'hb9f546b2),
	.w7(32'hb9857905),
	.w8(32'hba24c4a5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0beb83),
	.w1(32'h39993f43),
	.w2(32'h38dffbdf),
	.w3(32'h38b2783d),
	.w4(32'hba1f56b2),
	.w5(32'hb98e9773),
	.w6(32'h390f8d86),
	.w7(32'hb8c85300),
	.w8(32'hb9efc337),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c4ade7),
	.w1(32'hb9197f01),
	.w2(32'h397ee585),
	.w3(32'hba2f145a),
	.w4(32'hba16b2d5),
	.w5(32'hb993873f),
	.w6(32'hb9c405d8),
	.w7(32'hb9a5af72),
	.w8(32'hb95a0678),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d45e35),
	.w1(32'h398f2250),
	.w2(32'hb966d7c1),
	.w3(32'h3953d406),
	.w4(32'hb8dae9ec),
	.w5(32'h3905ce85),
	.w6(32'h392d35d8),
	.w7(32'hb994c7a7),
	.w8(32'h392f5824),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d78914),
	.w1(32'h391ee714),
	.w2(32'h39a2dca3),
	.w3(32'h3939827a),
	.w4(32'h394b0c20),
	.w5(32'hb9a61e41),
	.w6(32'h38a26a4e),
	.w7(32'h3832bcf4),
	.w8(32'h3a2745ca),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81d5da),
	.w1(32'hba314a27),
	.w2(32'hb9ad286f),
	.w3(32'hb94613e6),
	.w4(32'hb9d8f8b2),
	.w5(32'hb98ce8ab),
	.w6(32'h3aa06894),
	.w7(32'h393c79ef),
	.w8(32'hb9069829),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8fca0),
	.w1(32'hb92509df),
	.w2(32'hba0a435c),
	.w3(32'hb966ae1c),
	.w4(32'h37bb2c73),
	.w5(32'h3a52c167),
	.w6(32'hba61f481),
	.w7(32'hb9020e07),
	.w8(32'h3a4fb035),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17b7c8),
	.w1(32'hb8590cb8),
	.w2(32'h3982eb6a),
	.w3(32'h39bb8acb),
	.w4(32'h39327dde),
	.w5(32'h3c01de62),
	.w6(32'hb8d4c6cd),
	.w7(32'h39f6dfa1),
	.w8(32'h399c05e5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf1435),
	.w1(32'hbbd77872),
	.w2(32'hbb47a356),
	.w3(32'h3bd50682),
	.w4(32'h3b38d4cf),
	.w5(32'hbc0d7051),
	.w6(32'hbb92a058),
	.w7(32'hbaf76766),
	.w8(32'h3ad1a76d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b194b4e),
	.w1(32'h3c2a60e0),
	.w2(32'hb9c7f43b),
	.w3(32'hbb9af904),
	.w4(32'hbbcd3137),
	.w5(32'h3abc40de),
	.w6(32'h3b8c07ec),
	.w7(32'h3ab9cbda),
	.w8(32'hbc3a514f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c5e98),
	.w1(32'h3a0245a5),
	.w2(32'h3a325e3f),
	.w3(32'h3aa6c3dc),
	.w4(32'h3b68b95b),
	.w5(32'h3a0c7b86),
	.w6(32'hbc81c46b),
	.w7(32'hbbe80eb5),
	.w8(32'h3cb26b2f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c12fc68),
	.w1(32'h3bf6bc86),
	.w2(32'h3c4a1f04),
	.w3(32'h3a003f4f),
	.w4(32'h3c0a6bc8),
	.w5(32'h3b8bb14a),
	.w6(32'h3d0b0344),
	.w7(32'h3d09907e),
	.w8(32'hbc20b21d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3a63),
	.w1(32'hba87437c),
	.w2(32'hbaaf0300),
	.w3(32'hbb58db94),
	.w4(32'hbc03f88b),
	.w5(32'hbc66a888),
	.w6(32'hbc1f89c4),
	.w7(32'hbb8c102c),
	.w8(32'h3b8f2e13),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd63077),
	.w1(32'h3c550955),
	.w2(32'hbb0371db),
	.w3(32'hbc198531),
	.w4(32'hbc3abbca),
	.w5(32'hbb00e3f5),
	.w6(32'h3c0e4579),
	.w7(32'hbbe8ab3b),
	.w8(32'hbbcaf57c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b821200),
	.w1(32'h3b44a5de),
	.w2(32'h3b641140),
	.w3(32'hbc2e6493),
	.w4(32'hba5f6598),
	.w5(32'hbb8f239a),
	.w6(32'h3b40a655),
	.w7(32'h3b1f6b82),
	.w8(32'hbc241f67),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e9442),
	.w1(32'h3bcbd77a),
	.w2(32'hbb818dee),
	.w3(32'hb97e9cca),
	.w4(32'h3aa90f40),
	.w5(32'hbb89a39f),
	.w6(32'hbc73098f),
	.w7(32'hbbd07f89),
	.w8(32'h3a69e07b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3426dd),
	.w1(32'hbb4397bf),
	.w2(32'hbb936d61),
	.w3(32'hbb0fc020),
	.w4(32'hbc375fbb),
	.w5(32'hbb7ccd92),
	.w6(32'hba9d6455),
	.w7(32'h3adffb19),
	.w8(32'hbbea4565),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b365),
	.w1(32'h3ba9ddc1),
	.w2(32'hbb888f20),
	.w3(32'h3b07bdaa),
	.w4(32'h39986882),
	.w5(32'hbab88328),
	.w6(32'hbbd14277),
	.w7(32'hbbc2e6eb),
	.w8(32'hbbb93a96),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ec7d),
	.w1(32'hbc1bc2c0),
	.w2(32'hbb5afeda),
	.w3(32'h3b5a405d),
	.w4(32'hbb7d0790),
	.w5(32'h3aabd516),
	.w6(32'hbbe25702),
	.w7(32'h3a293081),
	.w8(32'h39a93b99),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9d837),
	.w1(32'h3a17c2d1),
	.w2(32'hba90c31b),
	.w3(32'hb9bb60da),
	.w4(32'hba3a02f8),
	.w5(32'hb68fcd37),
	.w6(32'hbb5f4c18),
	.w7(32'hbb27c11c),
	.w8(32'hbaa5b1ae),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf3942),
	.w1(32'hb9bc0ff8),
	.w2(32'hbb683ad2),
	.w3(32'hbc084188),
	.w4(32'hbb97cee2),
	.w5(32'hbc2ab219),
	.w6(32'hbb3f585b),
	.w7(32'hbb07506f),
	.w8(32'hbc47c592),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ec523),
	.w1(32'hbbd7694b),
	.w2(32'hbc19da4f),
	.w3(32'hbb767b8d),
	.w4(32'h3b7f32d8),
	.w5(32'hbb418d41),
	.w6(32'hbb9863e5),
	.w7(32'hbc8bfac9),
	.w8(32'hb921308c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba353971),
	.w1(32'h3ae4129d),
	.w2(32'h3b15455f),
	.w3(32'hbb95e2bb),
	.w4(32'hbb2847e4),
	.w5(32'h3be42172),
	.w6(32'hbbb19b4c),
	.w7(32'h3b1cc89f),
	.w8(32'hbba03e7c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6392d),
	.w1(32'h3b250eae),
	.w2(32'h3c0c098e),
	.w3(32'h3c89fc33),
	.w4(32'h3c5ea838),
	.w5(32'h3b8dad2b),
	.w6(32'hbc046320),
	.w7(32'hbb98d186),
	.w8(32'h3c37869f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e95fe),
	.w1(32'h3b464b9d),
	.w2(32'h3b0e097e),
	.w3(32'h3b9acc9a),
	.w4(32'h3b92f602),
	.w5(32'hbb937682),
	.w6(32'h3b66a0ae),
	.w7(32'h3ae4dd99),
	.w8(32'h3c794f75),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab51c2a),
	.w1(32'h3b9c2869),
	.w2(32'hbb80daf4),
	.w3(32'h3b645ca9),
	.w4(32'h3cd55436),
	.w5(32'hbac99e82),
	.w6(32'h3cb7b487),
	.w7(32'h3c3a7a93),
	.w8(32'hbbbbcc46),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8fecc),
	.w1(32'hbba507ab),
	.w2(32'hbb20e693),
	.w3(32'hbb0018aa),
	.w4(32'h3b8021fd),
	.w5(32'h3b3ab397),
	.w6(32'hbc19f426),
	.w7(32'hbb811207),
	.w8(32'h3b3bc363),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb879540),
	.w1(32'hbab553bc),
	.w2(32'h3bae2a8e),
	.w3(32'hbc5be4fa),
	.w4(32'hbc360d39),
	.w5(32'h3be0b1ab),
	.w6(32'h3c84e265),
	.w7(32'h3c3ba99e),
	.w8(32'hbb897788),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b507d29),
	.w1(32'h3b357754),
	.w2(32'h3bb4e774),
	.w3(32'h3c8463de),
	.w4(32'h3c203dc7),
	.w5(32'hbae2ec38),
	.w6(32'hbb3d0718),
	.w7(32'h3a47cf00),
	.w8(32'hbb6a697d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25b67),
	.w1(32'hbbb9d3e1),
	.w2(32'h3bc5534d),
	.w3(32'h3c3ecd6e),
	.w4(32'hbbf4bd50),
	.w5(32'hbaf805bb),
	.w6(32'h3a3d75f7),
	.w7(32'h3bd801b4),
	.w8(32'h3c3b5fc2),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20815f),
	.w1(32'h39665720),
	.w2(32'h3b2a9c9f),
	.w3(32'hbb7075e5),
	.w4(32'hbaabf34d),
	.w5(32'hbb811d7f),
	.w6(32'h3c5b475f),
	.w7(32'hbb1723a0),
	.w8(32'hbb6c6421),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb220fd),
	.w1(32'h3b4c8a42),
	.w2(32'h3bda2a0a),
	.w3(32'hbbe8f7e3),
	.w4(32'hbc7f9c5e),
	.w5(32'hbc4c5ec5),
	.w6(32'h3b85304f),
	.w7(32'hbb0176b6),
	.w8(32'hbc74dac2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21bba5),
	.w1(32'hba7e3731),
	.w2(32'hbc1b7741),
	.w3(32'hbc28bdb9),
	.w4(32'hbc5203b2),
	.w5(32'hb93a5e96),
	.w6(32'h3c3760e3),
	.w7(32'hbc1c6b90),
	.w8(32'h3c2068d7),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c0677),
	.w1(32'h3baf105a),
	.w2(32'h3b860837),
	.w3(32'hbc0e432f),
	.w4(32'hbb9a1052),
	.w5(32'hbbf9fa8e),
	.w6(32'h3c66b708),
	.w7(32'hbafad5db),
	.w8(32'h39c4f7f8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b838d),
	.w1(32'hbb1921ca),
	.w2(32'hbb1e587c),
	.w3(32'hbb02fefb),
	.w4(32'hbb61740b),
	.w5(32'hbb1757c0),
	.w6(32'h3c5d8c99),
	.w7(32'hbb9f7948),
	.w8(32'h3b46d3c5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf686db),
	.w1(32'hbc5c1f0b),
	.w2(32'hbc351472),
	.w3(32'h3b8922be),
	.w4(32'hbbc0b7be),
	.w5(32'h3bb9ae4c),
	.w6(32'h3d0ceeac),
	.w7(32'h3b748815),
	.w8(32'h3b62b11f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34b0ef),
	.w1(32'h3b7d030d),
	.w2(32'hb9b1cab3),
	.w3(32'h3a60bccc),
	.w4(32'h3b8cba51),
	.w5(32'h3bcd8489),
	.w6(32'h3b30537d),
	.w7(32'hbad16568),
	.w8(32'hbbb645da),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e282),
	.w1(32'hbb7e2332),
	.w2(32'hba16589b),
	.w3(32'h3c3d8cdf),
	.w4(32'hb85a8933),
	.w5(32'hbb4d14c4),
	.w6(32'hbb75bef8),
	.w7(32'hbb998eae),
	.w8(32'hbb01b013),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba904785),
	.w1(32'hbc0368a9),
	.w2(32'hbc17b3e7),
	.w3(32'hbb361e0d),
	.w4(32'hbbbb1646),
	.w5(32'hbbad2596),
	.w6(32'hbba0bd02),
	.w7(32'hbbdc42db),
	.w8(32'h391d4d2a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b590f74),
	.w1(32'h3bcd7979),
	.w2(32'hbb00a12c),
	.w3(32'hb9abd366),
	.w4(32'hbb6de215),
	.w5(32'hbc27affd),
	.w6(32'h3a43377f),
	.w7(32'h3a731f08),
	.w8(32'h3c0e1b6c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f2b51),
	.w1(32'h3b9adf24),
	.w2(32'hbc63e5ea),
	.w3(32'hbca28df5),
	.w4(32'hbbb37336),
	.w5(32'h3aba7993),
	.w6(32'h3c500efa),
	.w7(32'h3a5ce816),
	.w8(32'hbb25f2d7),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0ef39),
	.w1(32'h3b2a650b),
	.w2(32'hbbd8c1ba),
	.w3(32'hbb880997),
	.w4(32'hbb7d8cd5),
	.w5(32'hbbddda6c),
	.w6(32'h3ad191cc),
	.w7(32'hbbcf8707),
	.w8(32'h3a1c9461),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fb7d8),
	.w1(32'hba12e049),
	.w2(32'hbbaceb1f),
	.w3(32'hbc28b3c1),
	.w4(32'hbbc9dfa5),
	.w5(32'h3b744e55),
	.w6(32'h3c38f89e),
	.w7(32'hba8fceaa),
	.w8(32'h3a982b5a),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba96a7b),
	.w1(32'h3c036860),
	.w2(32'h3b71c1ab),
	.w3(32'h397f6b0a),
	.w4(32'h3a123e97),
	.w5(32'hbb723cc4),
	.w6(32'h3b4436c9),
	.w7(32'h3b1f0d83),
	.w8(32'h3aacc845),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b4765),
	.w1(32'h3b72f794),
	.w2(32'h3b91c51c),
	.w3(32'hba8a1936),
	.w4(32'h3b4348f3),
	.w5(32'hbc105e83),
	.w6(32'h3b7fe064),
	.w7(32'h3bbe011f),
	.w8(32'hbc3fc2de),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc38b3),
	.w1(32'hbb91ed05),
	.w2(32'h3971a836),
	.w3(32'hbc2fb72f),
	.w4(32'hbc05afa2),
	.w5(32'hb9e42df1),
	.w6(32'hbc43ee41),
	.w7(32'hbbebd527),
	.w8(32'hbb2d7e89),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa87a0c),
	.w1(32'hba36f779),
	.w2(32'h3a35d869),
	.w3(32'hba0edec5),
	.w4(32'h3b5e8bd0),
	.w5(32'h3b84927f),
	.w6(32'hbc02fd23),
	.w7(32'h3b0c71f8),
	.w8(32'h39dc28a9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9aeb09),
	.w1(32'h3bf43aa8),
	.w2(32'h3b5413e1),
	.w3(32'hb976a2e7),
	.w4(32'h3a2900d2),
	.w5(32'h3b83f23b),
	.w6(32'h3b404672),
	.w7(32'hb854fb31),
	.w8(32'hbbc97b86),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315b4c),
	.w1(32'h3bfd4f7a),
	.w2(32'h3b17d820),
	.w3(32'h3b76dfc5),
	.w4(32'hba97c724),
	.w5(32'h3aa83829),
	.w6(32'h3a0cc7d0),
	.w7(32'hba82ba02),
	.w8(32'hbc45f632),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07d24e),
	.w1(32'h3c10a61a),
	.w2(32'h3c3d4890),
	.w3(32'h3c943c52),
	.w4(32'h3a08d2cc),
	.w5(32'hbc250798),
	.w6(32'hbc15db12),
	.w7(32'hbbd70f16),
	.w8(32'hba87db44),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0c68),
	.w1(32'h3c3921a0),
	.w2(32'hb8624f33),
	.w3(32'hbc625ae5),
	.w4(32'hbb91e8d0),
	.w5(32'hbc1aa9b3),
	.w6(32'hbb3aa644),
	.w7(32'hbc1bc271),
	.w8(32'hbc859dd8),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17ca5b),
	.w1(32'hbc4bf3b7),
	.w2(32'hbbe9e887),
	.w3(32'hbbb04910),
	.w4(32'hbc257c50),
	.w5(32'h3b8002fa),
	.w6(32'h3bdf74b4),
	.w7(32'h3aca5a8f),
	.w8(32'hba27c982),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaf983),
	.w1(32'hbb14793f),
	.w2(32'h3aa25e4c),
	.w3(32'h3b07cb50),
	.w4(32'hba3a50f9),
	.w5(32'hba054248),
	.w6(32'h3b2f04be),
	.w7(32'h3b2e08f1),
	.w8(32'hbb204040),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982189c),
	.w1(32'hbb85f83d),
	.w2(32'hbb1af645),
	.w3(32'h3b107439),
	.w4(32'hbc05f283),
	.w5(32'hbc0dc990),
	.w6(32'h3be3d274),
	.w7(32'hbb7e12f8),
	.w8(32'hbbc3a07a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0b2c6),
	.w1(32'hbb42bfaa),
	.w2(32'h39f4d5dd),
	.w3(32'hbc1fdbba),
	.w4(32'hbbc98be9),
	.w5(32'hbb691759),
	.w6(32'hbc099cd3),
	.w7(32'h38d34d8b),
	.w8(32'hbaa2f015),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31e9cc),
	.w1(32'h3a8f851c),
	.w2(32'hb9eee4a9),
	.w3(32'hbbc58e2b),
	.w4(32'hbc0860eb),
	.w5(32'hbb7036a3),
	.w6(32'hba7b3add),
	.w7(32'hb9c93940),
	.w8(32'h3b2facf6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb406a3),
	.w1(32'h3b42869c),
	.w2(32'hbbba9953),
	.w3(32'hbbcf86e4),
	.w4(32'hb9d390cb),
	.w5(32'hbc867451),
	.w6(32'h3b5791d3),
	.w7(32'h3b839b17),
	.w8(32'h3bc67f7b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90b4b9),
	.w1(32'hbb32ccb7),
	.w2(32'hbc85cb42),
	.w3(32'hbbfa6ceb),
	.w4(32'h3c9e3b4a),
	.w5(32'hbbd23bb4),
	.w6(32'hbca7a04b),
	.w7(32'hbc86d67c),
	.w8(32'hba8cd9d5),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30e6c3),
	.w1(32'hbb5a6dd9),
	.w2(32'hba575eea),
	.w3(32'hbaf8f61d),
	.w4(32'hbb84438f),
	.w5(32'hbac430e6),
	.w6(32'h39cf9ef9),
	.w7(32'h3aaa7e26),
	.w8(32'hbbef782c),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb683d2c),
	.w1(32'hbbc2166b),
	.w2(32'hbb0b772c),
	.w3(32'hbb0b8602),
	.w4(32'h3ab93301),
	.w5(32'h3c17f8b0),
	.w6(32'hbc277634),
	.w7(32'hbb8aeffa),
	.w8(32'hbbbed977),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81d904),
	.w1(32'hbbd80e83),
	.w2(32'h3b00855a),
	.w3(32'h3be1bd34),
	.w4(32'hbac59e72),
	.w5(32'hbb0fa60c),
	.w6(32'hbc52cb4f),
	.w7(32'hb9d66042),
	.w8(32'hbbe687a6),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aaddbf),
	.w1(32'hbbaeb3f2),
	.w2(32'hbbf928d5),
	.w3(32'hbc8f894d),
	.w4(32'hbc9b4023),
	.w5(32'h3cd04e0c),
	.w6(32'hbb23c2e1),
	.w7(32'hbb936260),
	.w8(32'h3ccd7ddb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f89e7),
	.w1(32'hbc0bf7cb),
	.w2(32'h3bf29478),
	.w3(32'h3cafa6c0),
	.w4(32'h3d06a78c),
	.w5(32'hb911da65),
	.w6(32'h3c136e0a),
	.w7(32'h3d05a591),
	.w8(32'h3a3c4614),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba65200),
	.w1(32'hbb82a3a1),
	.w2(32'hb9c39a67),
	.w3(32'hbb054c16),
	.w4(32'hbaccd20f),
	.w5(32'hbb102e61),
	.w6(32'hbb9b7c24),
	.w7(32'hbb445ce9),
	.w8(32'h3ae7c87b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8918a0),
	.w1(32'hba20766b),
	.w2(32'h3bb4770b),
	.w3(32'hbc0980d6),
	.w4(32'hbb46366f),
	.w5(32'h393285ae),
	.w6(32'hbbb3fd04),
	.w7(32'hba43b94a),
	.w8(32'hbb6aacac),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99ab04),
	.w1(32'hbbb257db),
	.w2(32'hbbb582d4),
	.w3(32'h3a118a2c),
	.w4(32'hbad1db8a),
	.w5(32'h3cb33e40),
	.w6(32'hbbddffcd),
	.w7(32'hbb2d7a57),
	.w8(32'h3c1411bf),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5ddee3),
	.w1(32'h3c4e6937),
	.w2(32'h3c85bea3),
	.w3(32'h3d0b25f8),
	.w4(32'hbbdca202),
	.w5(32'hbc211636),
	.w6(32'h3d1889ae),
	.w7(32'h3c9fe229),
	.w8(32'hbb6434a8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38012a),
	.w1(32'hbb5996a8),
	.w2(32'hbb65af66),
	.w3(32'hbc8f7e3a),
	.w4(32'h3a9a0590),
	.w5(32'hbc0597da),
	.w6(32'hba0638cf),
	.w7(32'h3aea907f),
	.w8(32'hbad13b5e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f0c8a),
	.w1(32'hbafa4b15),
	.w2(32'hbbf3507f),
	.w3(32'hbc453599),
	.w4(32'hbc47fa43),
	.w5(32'hbc054951),
	.w6(32'h3c18c187),
	.w7(32'hbbbe435b),
	.w8(32'h3acae1ca),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3750c5),
	.w1(32'hba7df36f),
	.w2(32'hbc079a98),
	.w3(32'hbb24e02f),
	.w4(32'hbbfcc375),
	.w5(32'h3ad975bc),
	.w6(32'h3c53e3c2),
	.w7(32'hbb91f994),
	.w8(32'h3cca6fb7),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04961f),
	.w1(32'hb9926515),
	.w2(32'hbc0eaafe),
	.w3(32'h3cb1abbb),
	.w4(32'h3c91cac4),
	.w5(32'h3ad4ed3e),
	.w6(32'h3bf1a333),
	.w7(32'hbb9cdc41),
	.w8(32'hb8ad7d63),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9950a5),
	.w1(32'hbac80807),
	.w2(32'h3acfe878),
	.w3(32'h3af858f1),
	.w4(32'hbc54b87a),
	.w5(32'h3ceaa57f),
	.w6(32'h3bd6e778),
	.w7(32'h3af7ba66),
	.w8(32'hbb275c43),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855970),
	.w1(32'h3b9ea286),
	.w2(32'h3c49fd7b),
	.w3(32'h3cc75687),
	.w4(32'hbbb3adde),
	.w5(32'hbbb5085b),
	.w6(32'hbad72fe2),
	.w7(32'h3ca51fc6),
	.w8(32'h3c798559),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b4c07),
	.w1(32'h3bb761df),
	.w2(32'h3b9fbcc8),
	.w3(32'hbc3ed4d0),
	.w4(32'h3b232fcd),
	.w5(32'h3c63a160),
	.w6(32'h3c41df51),
	.w7(32'h3c6c0cad),
	.w8(32'hb9357cbc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabee81b),
	.w1(32'hbbd121f4),
	.w2(32'h3bcb51ff),
	.w3(32'h3c853aa6),
	.w4(32'h3bf35f0e),
	.w5(32'h3b4b2804),
	.w6(32'h3c34d510),
	.w7(32'h3c15f38b),
	.w8(32'hbba52c9a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8de3f),
	.w1(32'h3bc40ce7),
	.w2(32'h3c402aab),
	.w3(32'hbb799050),
	.w4(32'hb91e55a3),
	.w5(32'hbb254c42),
	.w6(32'hbbd02ad0),
	.w7(32'h3aa40aa9),
	.w8(32'hba2ee1f9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2449d7),
	.w1(32'h3a8c66f4),
	.w2(32'h3b44cc3b),
	.w3(32'hbc0d3e02),
	.w4(32'hbc26ce7f),
	.w5(32'hbbec49c5),
	.w6(32'h3c54676e),
	.w7(32'h3b94417f),
	.w8(32'hbc240e0f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b5a30),
	.w1(32'hbb82d773),
	.w2(32'hbaa1841f),
	.w3(32'hbb256364),
	.w4(32'hbb30b76a),
	.w5(32'h3c40767c),
	.w6(32'hbbd4b4ba),
	.w7(32'hbbf842dc),
	.w8(32'hbc304b0b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2532a),
	.w1(32'h3ce511ef),
	.w2(32'h3c8e3757),
	.w3(32'h3d0ad38a),
	.w4(32'h3b2b0f91),
	.w5(32'h3ada69e1),
	.w6(32'h3b939e43),
	.w7(32'h3c999e65),
	.w8(32'h3a935d60),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe265a),
	.w1(32'h3b482e07),
	.w2(32'h3aa58e87),
	.w3(32'hbad5dec8),
	.w4(32'hb982b7d4),
	.w5(32'hba3ea482),
	.w6(32'hbb7ed9cd),
	.w7(32'hba9c6c53),
	.w8(32'hbb75428d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37e2db),
	.w1(32'h3c3013bb),
	.w2(32'h3ba53ac8),
	.w3(32'hbbb02f28),
	.w4(32'h3b5d567f),
	.w5(32'h3a9bc8a8),
	.w6(32'hbb69d6a5),
	.w7(32'h3bb9a84c),
	.w8(32'hbb02db0b),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f9b0f),
	.w1(32'h3b8a1a38),
	.w2(32'hb999d05e),
	.w3(32'hbbda499e),
	.w4(32'hbbb9ae8d),
	.w5(32'hbb9f0185),
	.w6(32'h3bfc35fb),
	.w7(32'h3a33fff7),
	.w8(32'hbb617ff7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82764b),
	.w1(32'hb8b3689c),
	.w2(32'hbc02b1f1),
	.w3(32'hbb87a2fd),
	.w4(32'hbbd9ca69),
	.w5(32'hbaeda087),
	.w6(32'hbc03d6c9),
	.w7(32'hbbd5944c),
	.w8(32'hbb7f99d1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc4af7),
	.w1(32'hbb24b29b),
	.w2(32'hbb133b1b),
	.w3(32'hbbdf9b69),
	.w4(32'hbb6d30b4),
	.w5(32'h3b299835),
	.w6(32'hbc492594),
	.w7(32'hbbd083b7),
	.w8(32'h3af1fcb1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b7a60),
	.w1(32'hba2c6134),
	.w2(32'h3b8a743a),
	.w3(32'h3bb51236),
	.w4(32'h3ba28b69),
	.w5(32'hbaddb206),
	.w6(32'hbc0ba69b),
	.w7(32'hbac479ab),
	.w8(32'hbb9ca909),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b973040),
	.w1(32'h3acac128),
	.w2(32'h3be57f4c),
	.w3(32'hbb0423a3),
	.w4(32'hbabb2d2b),
	.w5(32'hb95e8cb1),
	.w6(32'hbbe3d53a),
	.w7(32'h39ef7e89),
	.w8(32'h3c0feaed),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf96da),
	.w1(32'h3b9cb0b1),
	.w2(32'h3b04a09c),
	.w3(32'hbc182475),
	.w4(32'hbae8a902),
	.w5(32'hbb9ef061),
	.w6(32'h3b4eff5e),
	.w7(32'hb9fe2024),
	.w8(32'hbc21d47b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99c830),
	.w1(32'hbbf53183),
	.w2(32'hbb97aa8a),
	.w3(32'hbbc1ce31),
	.w4(32'hbb850b21),
	.w5(32'hbc249828),
	.w6(32'hbc8525c7),
	.w7(32'hbc21dbf9),
	.w8(32'h3c891e9d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42caa1),
	.w1(32'hbae137b0),
	.w2(32'hb9f767f5),
	.w3(32'hbc010329),
	.w4(32'h3b8c8b75),
	.w5(32'hbba70740),
	.w6(32'h3c845cc7),
	.w7(32'h3c857fbb),
	.w8(32'h3b5c1705),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0be6b9),
	.w1(32'h3b82be94),
	.w2(32'h3b5a62da),
	.w3(32'hbc37fc44),
	.w4(32'h3aa72b61),
	.w5(32'h3b066dfc),
	.w6(32'hbb856e57),
	.w7(32'hbbc5447a),
	.w8(32'hbc59ee4e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799b30),
	.w1(32'h3978e6b2),
	.w2(32'hbb8be537),
	.w3(32'hba982b20),
	.w4(32'hbc470905),
	.w5(32'hb9d09948),
	.w6(32'hbc8d01fa),
	.w7(32'hbc7dce9c),
	.w8(32'hbb0e2ea0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39023a88),
	.w1(32'hbad08c73),
	.w2(32'h3b94a89b),
	.w3(32'h3bfcbd72),
	.w4(32'hbbcedb80),
	.w5(32'hbbaacda7),
	.w6(32'hba2b0c6f),
	.w7(32'h3bcb5091),
	.w8(32'hbb20df80),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce09a54),
	.w1(32'h3bcc0314),
	.w2(32'hbb2b69bd),
	.w3(32'h3bd56b91),
	.w4(32'h3d02d4c2),
	.w5(32'h3c00a103),
	.w6(32'hbcdb4ec7),
	.w7(32'hbc77feff),
	.w8(32'h3c2bebae),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76ea36),
	.w1(32'h3c9c19f0),
	.w2(32'h3c9646f9),
	.w3(32'h3bb8651b),
	.w4(32'hbbf65c80),
	.w5(32'h3c306684),
	.w6(32'h3ccc9df6),
	.w7(32'h3c9e978f),
	.w8(32'hbaa8d86a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6186f),
	.w1(32'h3accf8cc),
	.w2(32'h3c1e8281),
	.w3(32'h3c7e2c22),
	.w4(32'hbae717c5),
	.w5(32'hbbda90b4),
	.w6(32'h3c335f81),
	.w7(32'h3c5f38b0),
	.w8(32'hbbd0d61f),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11acaa),
	.w1(32'hba80c885),
	.w2(32'hba9c94ce),
	.w3(32'h38ffb815),
	.w4(32'hb9b0f0bc),
	.w5(32'hbb86f582),
	.w6(32'hb9dcbb0d),
	.w7(32'h39e179db),
	.w8(32'hbbdb685d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d5e95),
	.w1(32'hbbc71f43),
	.w2(32'hbb1e71b7),
	.w3(32'hbbc9c1d0),
	.w4(32'hbba64342),
	.w5(32'h3b315d9d),
	.w6(32'hbc58f925),
	.w7(32'hbbbfdaf4),
	.w8(32'h3b0744d0),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201d3c),
	.w1(32'hbb2e9aa6),
	.w2(32'h3ba53a98),
	.w3(32'h3aba0da1),
	.w4(32'h3b853c08),
	.w5(32'hbb03f214),
	.w6(32'hbba95831),
	.w7(32'h3b9b0519),
	.w8(32'h3b8dc540),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e0d4a),
	.w1(32'h3b593184),
	.w2(32'h3a87b66e),
	.w3(32'hba98a24f),
	.w4(32'hbb41fb46),
	.w5(32'hbb671f48),
	.w6(32'h3b832742),
	.w7(32'hbb943872),
	.w8(32'hba280202),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b871432),
	.w1(32'h3a714f65),
	.w2(32'hbaa2e03b),
	.w3(32'hbbcc9a11),
	.w4(32'hbb97d9d8),
	.w5(32'hb9147195),
	.w6(32'h3ad24344),
	.w7(32'hbbfdaecc),
	.w8(32'h3b51ab17),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecc8c9),
	.w1(32'h3b434272),
	.w2(32'hbb7c2ea5),
	.w3(32'h3990fbc0),
	.w4(32'hbb556d43),
	.w5(32'h3c86105a),
	.w6(32'h3cc519c2),
	.w7(32'h3b900f60),
	.w8(32'hbba4c6fb),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b60a9),
	.w1(32'h3b93fce9),
	.w2(32'h3c36d49d),
	.w3(32'h3cd5e4d1),
	.w4(32'h3a682c36),
	.w5(32'hbbddc12b),
	.w6(32'h3b8f1482),
	.w7(32'h3cae8f28),
	.w8(32'hbbe9e834),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9722628),
	.w1(32'hba3257d9),
	.w2(32'hbb941687),
	.w3(32'hbc0225d9),
	.w4(32'h3bb65e76),
	.w5(32'h3c006d79),
	.w6(32'h3c013baa),
	.w7(32'hbc007eab),
	.w8(32'hbc9653b2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a48fa),
	.w1(32'h3b695509),
	.w2(32'h3aa0274b),
	.w3(32'h3c5dcbce),
	.w4(32'h3c7faf86),
	.w5(32'hb9e69734),
	.w6(32'hbbbe993b),
	.w7(32'hbc9927bd),
	.w8(32'hbbac3403),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61f901),
	.w1(32'hbb0851aa),
	.w2(32'h3a834116),
	.w3(32'hbb95de3f),
	.w4(32'hbbbe2d67),
	.w5(32'hbb136a48),
	.w6(32'hbb3247bb),
	.w7(32'hbb149c91),
	.w8(32'hbad0ea5e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65404b),
	.w1(32'hba942e8a),
	.w2(32'hbabf9aa8),
	.w3(32'h3957e7b4),
	.w4(32'h3c85e2b0),
	.w5(32'hbc1124c2),
	.w6(32'h3a804755),
	.w7(32'h3b2ed929),
	.w8(32'h3c49729c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec5db7),
	.w1(32'hbc361b60),
	.w2(32'hbbc72983),
	.w3(32'h3c34966e),
	.w4(32'h3ccc0979),
	.w5(32'h3b1d9cbe),
	.w6(32'h3b407f87),
	.w7(32'hbc1ef72f),
	.w8(32'hbb5b9dce),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d1aea),
	.w1(32'h3ba6e031),
	.w2(32'hbb028f8e),
	.w3(32'h3a92cc6f),
	.w4(32'h3a6039c6),
	.w5(32'hb87c8525),
	.w6(32'hbc94f06b),
	.w7(32'h3b90691d),
	.w8(32'h3a2a73c8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa207f6),
	.w1(32'h39c46145),
	.w2(32'h3bd26cb0),
	.w3(32'hbae62d2a),
	.w4(32'h3b947a38),
	.w5(32'hbc14d69a),
	.w6(32'hbbafc92c),
	.w7(32'h393a52bf),
	.w8(32'hbace3af7),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab91fd3),
	.w1(32'hb9b6e523),
	.w2(32'hbb41146c),
	.w3(32'hbc32d87d),
	.w4(32'hbc53b845),
	.w5(32'hbc13a8d1),
	.w6(32'hbb9f621d),
	.w7(32'hbbade008),
	.w8(32'h3bdbc315),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbfbe6),
	.w1(32'h3bb6b8a9),
	.w2(32'h3b96ea82),
	.w3(32'hbc741577),
	.w4(32'hbc841ff6),
	.w5(32'hbad750e2),
	.w6(32'h3c6f0b78),
	.w7(32'h3ade8b97),
	.w8(32'h3c02e10d),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b405be4),
	.w1(32'h3b3aa932),
	.w2(32'hba027c73),
	.w3(32'hbb89818d),
	.w4(32'h3a7428e7),
	.w5(32'h3c010c27),
	.w6(32'h3b93f46b),
	.w7(32'hbae26018),
	.w8(32'h3b3d1bda),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3dd54),
	.w1(32'h3bf334f3),
	.w2(32'h3a923ee4),
	.w3(32'h3b0e1864),
	.w4(32'hbbd23eee),
	.w5(32'hbc16e87b),
	.w6(32'h3b415392),
	.w7(32'hb82d81ea),
	.w8(32'h3ad63d9a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d12c),
	.w1(32'h3bef84d2),
	.w2(32'h3ba202c7),
	.w3(32'hbc4bd837),
	.w4(32'hbc33e8c9),
	.w5(32'h3b828d51),
	.w6(32'h3bb7c4c5),
	.w7(32'h3b5bd548),
	.w8(32'hbc3ec90b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27eddc),
	.w1(32'h3c5e8172),
	.w2(32'h3bd119c4),
	.w3(32'h3bea1da0),
	.w4(32'hba8ff092),
	.w5(32'hbb44930a),
	.w6(32'hbc4f9e2a),
	.w7(32'hbb98ed9c),
	.w8(32'hbb4c743b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f60f7),
	.w1(32'h3ad38f6a),
	.w2(32'h3b8182a6),
	.w3(32'hbb1b391c),
	.w4(32'hbb95521f),
	.w5(32'hbbd75b3e),
	.w6(32'h3bbc2d04),
	.w7(32'hbb908a8e),
	.w8(32'hbb427b5b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77d82),
	.w1(32'h3a8d674c),
	.w2(32'hbbb9742c),
	.w3(32'hbbec60e1),
	.w4(32'hbbe4c498),
	.w5(32'h3a9897df),
	.w6(32'h3b3c1dd5),
	.w7(32'hbbcc69d4),
	.w8(32'h3be54e72),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87aaa1),
	.w1(32'h3a735f47),
	.w2(32'hbaacc73e),
	.w3(32'hbb71fc63),
	.w4(32'hbbb98060),
	.w5(32'hbacbda42),
	.w6(32'h3c3263bc),
	.w7(32'h3b3144d0),
	.w8(32'hbb8565b7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c075),
	.w1(32'h3b9def51),
	.w2(32'h3ad6d1bd),
	.w3(32'hbb56e1da),
	.w4(32'h3bb1bf12),
	.w5(32'hbb9087f2),
	.w6(32'hbc11a07c),
	.w7(32'hbbe134d6),
	.w8(32'h3b8f9d2d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab27dd7),
	.w1(32'h3b88979c),
	.w2(32'hbb89c23a),
	.w3(32'hbc30163e),
	.w4(32'hba755c75),
	.w5(32'hbc190a1b),
	.w6(32'h3b56ca00),
	.w7(32'hb632cf44),
	.w8(32'h3b75ba74),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb190f),
	.w1(32'h3b06f343),
	.w2(32'hba12ef9c),
	.w3(32'hbbdcb8a2),
	.w4(32'hbaea260c),
	.w5(32'h3a666b20),
	.w6(32'h3bc1f68f),
	.w7(32'hbc039ead),
	.w8(32'hbb962cd6),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1bf42),
	.w1(32'h3b835028),
	.w2(32'h3b32651c),
	.w3(32'hbbab1f6e),
	.w4(32'h39e55cba),
	.w5(32'hbb42a04b),
	.w6(32'hbb1ec30d),
	.w7(32'h39f654da),
	.w8(32'h3bd4346b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70a5f8),
	.w1(32'hbc367765),
	.w2(32'hbc07d94e),
	.w3(32'hbbb8a052),
	.w4(32'h3b2ecf96),
	.w5(32'hbb8a7cf0),
	.w6(32'h3bbd3dae),
	.w7(32'hbabe67e3),
	.w8(32'hbc0bc85f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b544c3),
	.w1(32'hbb6431ee),
	.w2(32'hbacab9b8),
	.w3(32'hbba1675c),
	.w4(32'hbbd3418d),
	.w5(32'hbc179983),
	.w6(32'hbb93f4b5),
	.w7(32'hbc50b803),
	.w8(32'hbb6562a8),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5933bf),
	.w1(32'hbbd9256f),
	.w2(32'hbc1a0658),
	.w3(32'hbc4b8c39),
	.w4(32'hbb780c3e),
	.w5(32'hbc5c8c96),
	.w6(32'hbb8573f2),
	.w7(32'hbc6a6f69),
	.w8(32'h3bf13304),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8678c9),
	.w1(32'hba853bf0),
	.w2(32'hbb898c07),
	.w3(32'hbb95f5cb),
	.w4(32'hba5a87ce),
	.w5(32'hba331b4a),
	.w6(32'h3c95a197),
	.w7(32'h38380aac),
	.w8(32'h3b0e14e1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951dd9),
	.w1(32'h3ba018ed),
	.w2(32'h3bbb34ef),
	.w3(32'hb9ca8929),
	.w4(32'h3aa439b7),
	.w5(32'hbbdacd91),
	.w6(32'h3a54f6d1),
	.w7(32'h3b285196),
	.w8(32'h3a31aa37),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5abd48),
	.w1(32'h3b1cbe1c),
	.w2(32'hbc001590),
	.w3(32'hbc3a9823),
	.w4(32'hbc91b0ef),
	.w5(32'hba7d93d5),
	.w6(32'hbbaeb428),
	.w7(32'hbc0445b5),
	.w8(32'h3b73e1c0),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abcf5df),
	.w1(32'hba511d37),
	.w2(32'hbb831e2e),
	.w3(32'hbbb0d523),
	.w4(32'hbbe2c81c),
	.w5(32'hbc0e5b5c),
	.w6(32'hba916690),
	.w7(32'hbbcfd4e1),
	.w8(32'h3aeb7abb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a115648),
	.w1(32'h3becc8e4),
	.w2(32'hbab566d8),
	.w3(32'hbc47e354),
	.w4(32'hbac2fa11),
	.w5(32'hbba5052e),
	.w6(32'h3bd2c712),
	.w7(32'hbaa8977e),
	.w8(32'h3a268f11),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0eaec),
	.w1(32'hbb73f68a),
	.w2(32'hbbdc35f5),
	.w3(32'hbbfd7dbc),
	.w4(32'hbc88c9ab),
	.w5(32'hbbe46301),
	.w6(32'h3c800ae7),
	.w7(32'h39e307dc),
	.w8(32'h3c121881),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f3908),
	.w1(32'h3b63af09),
	.w2(32'h3c101bbd),
	.w3(32'hbc31ad5b),
	.w4(32'hbb15f377),
	.w5(32'hbac0ae46),
	.w6(32'h3c93ebda),
	.w7(32'h3c50d7f7),
	.w8(32'h3a98368e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d455c),
	.w1(32'hbb8fe8cb),
	.w2(32'hbb8d717e),
	.w3(32'hb9fecbbf),
	.w4(32'hbb76e75e),
	.w5(32'h38cdccd1),
	.w6(32'hbb409f20),
	.w7(32'h39302317),
	.w8(32'hbaff5ec0),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf12b5),
	.w1(32'hbb806617),
	.w2(32'hbbc74101),
	.w3(32'hbaea54f5),
	.w4(32'hbb8951a1),
	.w5(32'hba61e379),
	.w6(32'h3c209f76),
	.w7(32'h38a6c74c),
	.w8(32'h3b106757),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccd9a3),
	.w1(32'h3ba33afa),
	.w2(32'h39933e0f),
	.w3(32'h39eb3d91),
	.w4(32'hbb3b4d3b),
	.w5(32'hbc14aaa2),
	.w6(32'h3bf0e819),
	.w7(32'hb9ef8326),
	.w8(32'hbc34ae36),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba3b05),
	.w1(32'h3a8c4aac),
	.w2(32'hbbc17519),
	.w3(32'hbc8aaae5),
	.w4(32'hbc9f84df),
	.w5(32'hb975d3e2),
	.w6(32'hbc5c6a47),
	.w7(32'hbc238ac6),
	.w8(32'hb999e4f0),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2d428),
	.w1(32'hb974315b),
	.w2(32'hba984b47),
	.w3(32'hb91b18cc),
	.w4(32'hba44256a),
	.w5(32'h39f5fdfb),
	.w6(32'hb959592a),
	.w7(32'hba6fbcd7),
	.w8(32'hb89260b8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28fb57),
	.w1(32'h3a79eab6),
	.w2(32'h399f481e),
	.w3(32'h39bba0c3),
	.w4(32'h39320048),
	.w5(32'hbad52832),
	.w6(32'h3a042882),
	.w7(32'h39b239ad),
	.w8(32'hba62f3c2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad546a3),
	.w1(32'hba49a3a5),
	.w2(32'hbabc88ba),
	.w3(32'hba5d557a),
	.w4(32'hbaa90888),
	.w5(32'hb9d6fb40),
	.w6(32'hb953f023),
	.w7(32'hba46f772),
	.w8(32'hba893ac2),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fdc536),
	.w1(32'h3a463203),
	.w2(32'h3a8b382a),
	.w3(32'hba17281d),
	.w4(32'h38f74238),
	.w5(32'hb8ece090),
	.w6(32'hba188002),
	.w7(32'h39389658),
	.w8(32'hb95f49ee),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d1443),
	.w1(32'h3994a01d),
	.w2(32'hb993d65b),
	.w3(32'h38b4bf43),
	.w4(32'hb92adf92),
	.w5(32'hbb46fc07),
	.w6(32'h3987e361),
	.w7(32'h372a5372),
	.w8(32'hbb7efe0c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70636a),
	.w1(32'hbb8af056),
	.w2(32'hbb561caa),
	.w3(32'hbb2d9f00),
	.w4(32'hbafa297b),
	.w5(32'h3a90ae5f),
	.w6(32'hbb623fc5),
	.w7(32'hbb2b613a),
	.w8(32'h3ae0dba4),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8be74),
	.w1(32'h3a230f23),
	.w2(32'hb8eeb617),
	.w3(32'h383e5c86),
	.w4(32'hba9581f9),
	.w5(32'h3a38fa5a),
	.w6(32'h39d1c3c8),
	.w7(32'hb9c56c9c),
	.w8(32'h39d34ede),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3976e8eb),
	.w1(32'hba19d563),
	.w2(32'hb8482484),
	.w3(32'h393ade40),
	.w4(32'hb8a865c7),
	.w5(32'h3a150d7b),
	.w6(32'h38f19ac7),
	.w7(32'hb8a38ef2),
	.w8(32'h3af06f5f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ff77f),
	.w1(32'h3a747d2e),
	.w2(32'hb808b2e1),
	.w3(32'h3a671ae5),
	.w4(32'hb8a942e2),
	.w5(32'hb9cefaa2),
	.w6(32'h3ac4cc4a),
	.w7(32'h36ec112a),
	.w8(32'hb9ae1b5d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba093b8e),
	.w1(32'hb9eb4b54),
	.w2(32'hb9a339bf),
	.w3(32'hb9e85979),
	.w4(32'hb96e403c),
	.w5(32'h3a8a3aa3),
	.w6(32'hba12c90c),
	.w7(32'hb98bb96e),
	.w8(32'h3a8118d4),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a708293),
	.w1(32'h39963f57),
	.w2(32'hba893473),
	.w3(32'h3a115ce5),
	.w4(32'hb98acc60),
	.w5(32'hb98ca475),
	.w6(32'h3a0ab710),
	.w7(32'hba0d3c99),
	.w8(32'hb8e35fb9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cef1e9),
	.w1(32'h3a4f6fc8),
	.w2(32'h3a3e3df4),
	.w3(32'h38f66c23),
	.w4(32'h3980ac6c),
	.w5(32'h391f6984),
	.w6(32'h3908981a),
	.w7(32'h39bd3fb9),
	.w8(32'hb94f5d9f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fbc8df),
	.w1(32'hb8fb9963),
	.w2(32'hb79d0873),
	.w3(32'hb9bae0f9),
	.w4(32'hb8084ce1),
	.w5(32'hba98a80b),
	.w6(32'hba9e8b4f),
	.w7(32'hba0f5da9),
	.w8(32'hba23ae80),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9547e9c),
	.w1(32'h3940ef54),
	.w2(32'h38cfc473),
	.w3(32'hba39d320),
	.w4(32'hb9bbdf89),
	.w5(32'h3b59eb01),
	.w6(32'hb9cd81d9),
	.w7(32'hb7b0fbf4),
	.w8(32'h3b6b792e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b663c4b),
	.w1(32'h3b71b593),
	.w2(32'h3b58a518),
	.w3(32'h3b60d0b5),
	.w4(32'h3b4b9db7),
	.w5(32'hb9c26395),
	.w6(32'h3b4adb19),
	.w7(32'h3b2bf088),
	.w8(32'hba169572),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbcae6),
	.w1(32'hba5ae9ff),
	.w2(32'hbac29885),
	.w3(32'hb939a103),
	.w4(32'hb9a14c5b),
	.w5(32'hba817bcf),
	.w6(32'hb99eb594),
	.w7(32'hba490eab),
	.w8(32'hba6caa2b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa671a4),
	.w1(32'hbacf7ae2),
	.w2(32'hba830cd0),
	.w3(32'hba9cc648),
	.w4(32'hbaafdc05),
	.w5(32'hba675f88),
	.w6(32'hba00e4e2),
	.w7(32'hba943ae0),
	.w8(32'hba76cea3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93078e0),
	.w1(32'h3996bc6c),
	.w2(32'h3a141afa),
	.w3(32'hba5ce0d4),
	.w4(32'hb9b64b9b),
	.w5(32'h3a7af1d1),
	.w6(32'hba5799b3),
	.w7(32'h38277325),
	.w8(32'h3a9b906f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4d979),
	.w1(32'h3aca6245),
	.w2(32'h3acc7452),
	.w3(32'h3a9097e8),
	.w4(32'h3a9b0793),
	.w5(32'hba4a235a),
	.w6(32'h3ac6a9ec),
	.w7(32'h3ac1ff92),
	.w8(32'hba580bdf),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf89a5a),
	.w1(32'hbaabd8c6),
	.w2(32'hbad41b6e),
	.w3(32'hba4f9c08),
	.w4(32'hbae82843),
	.w5(32'hba687920),
	.w6(32'hba8c1d08),
	.w7(32'hbab00f5c),
	.w8(32'hbabe7d53),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac915e9),
	.w1(32'hb9dc831b),
	.w2(32'hba88938a),
	.w3(32'hb9c6b562),
	.w4(32'hba16ebca),
	.w5(32'hbb80cbd6),
	.w6(32'hba197622),
	.w7(32'hba80d652),
	.w8(32'hbb8bb3cf),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80d60a),
	.w1(32'hbb7c54e7),
	.w2(32'hbb85aa04),
	.w3(32'hbb4a51e2),
	.w4(32'hbb224c48),
	.w5(32'hb910c0f3),
	.w6(32'hbb61c0db),
	.w7(32'hbb5d6ba2),
	.w8(32'hb9b70f4f),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08a5e8),
	.w1(32'hba14c141),
	.w2(32'h38f2678b),
	.w3(32'hb9d1313b),
	.w4(32'h389a56b9),
	.w5(32'h3b2064a0),
	.w6(32'hba1c013c),
	.w7(32'hb9cb2775),
	.w8(32'h3b1b0145),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae43792),
	.w1(32'h3ac19ef7),
	.w2(32'h3ab3806a),
	.w3(32'h3b035701),
	.w4(32'h3aaa6777),
	.w5(32'h3b1b1a33),
	.w6(32'h3aea5ffd),
	.w7(32'h3ab60322),
	.w8(32'h3af1c90e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb3f7f),
	.w1(32'h3aab49f7),
	.w2(32'h3ac471d7),
	.w3(32'h3b1172f0),
	.w4(32'h3b4d5648),
	.w5(32'h3ad268b1),
	.w6(32'h3ae77eb4),
	.w7(32'h3b1a4098),
	.w8(32'h3b09b9bd),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa367c),
	.w1(32'h3ae54b4f),
	.w2(32'h3ae85c2a),
	.w3(32'h3ab0a84e),
	.w4(32'h3a72ab53),
	.w5(32'h3b1e43a5),
	.w6(32'h3a8f0e6f),
	.w7(32'h3aa9070a),
	.w8(32'h3ab6830d),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa8f40),
	.w1(32'h3aaf69a0),
	.w2(32'h3af23abe),
	.w3(32'h3b2f8a5c),
	.w4(32'h3b32b8da),
	.w5(32'hb9dbbd22),
	.w6(32'h3aa03889),
	.w7(32'h3b104cc5),
	.w8(32'hb9dc5159),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad8517),
	.w1(32'h39b1028d),
	.w2(32'h39c387f3),
	.w3(32'hb9b44c2a),
	.w4(32'hb9060a16),
	.w5(32'hb9e228fe),
	.w6(32'hba35d628),
	.w7(32'hb9a2ceb6),
	.w8(32'hb98ad1b6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956cde2),
	.w1(32'h3954501e),
	.w2(32'h39372a48),
	.w3(32'hb9422489),
	.w4(32'h39c28cb8),
	.w5(32'hb91099d3),
	.w6(32'hba25e0ad),
	.w7(32'h381a8c70),
	.w8(32'hb82168f5),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb924922d),
	.w1(32'h37b933f9),
	.w2(32'hb94814c9),
	.w3(32'hb90cd6e6),
	.w4(32'hb9ac7f99),
	.w5(32'h3aa13a47),
	.w6(32'h393e55d5),
	.w7(32'hb9c83ba8),
	.w8(32'h3ac0a895),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule