module layer_10_featuremap_506(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57894e5),
	.w1(32'hb44b1caf),
	.w2(32'hb5c79862),
	.w3(32'hb5b86234),
	.w4(32'hb417430b),
	.w5(32'hb5dbf301),
	.w6(32'hb5b476ed),
	.w7(32'h34375e00),
	.w8(32'hb55a1e1f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a89563),
	.w1(32'h398de9ed),
	.w2(32'h39886299),
	.w3(32'h39c55b17),
	.w4(32'h392e3d4d),
	.w5(32'h396a3dc5),
	.w6(32'h3a074f34),
	.w7(32'h39987298),
	.w8(32'h39a6565e),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb55f4917),
	.w1(32'h3445f1fa),
	.w2(32'hb51db845),
	.w3(32'hb45e66a8),
	.w4(32'h35684888),
	.w5(32'h3482fae7),
	.w6(32'h34a986ee),
	.w7(32'h3570db98),
	.w8(32'hb499390f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8753332),
	.w1(32'hb8f577a4),
	.w2(32'hb8b3e0bf),
	.w3(32'hb75d3d8f),
	.w4(32'hb8645d4e),
	.w5(32'hb7c5daff),
	.w6(32'hb572aa50),
	.w7(32'hb893d1e3),
	.w8(32'hb81e39ae),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb663e2a1),
	.w1(32'hb5f0bfb3),
	.w2(32'hb6208efa),
	.w3(32'hb6726f45),
	.w4(32'hb600e85d),
	.w5(32'hb62c612c),
	.w6(32'hb6503f1e),
	.w7(32'hb5cd9dce),
	.w8(32'hb637580e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f97dc0),
	.w1(32'hb58cf83b),
	.w2(32'hb5be1868),
	.w3(32'hb43dac79),
	.w4(32'h334bb5e9),
	.w5(32'hb59ba201),
	.w6(32'hb4812a11),
	.w7(32'hb4a600b1),
	.w8(32'hb4cf9dc0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb911b4f0),
	.w1(32'h39118125),
	.w2(32'h39a0d840),
	.w3(32'hb9209159),
	.w4(32'h39b3105d),
	.w5(32'h39d96b15),
	.w6(32'hba1eb257),
	.w7(32'hb91a79e7),
	.w8(32'h397158a4),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07c8f),
	.w1(32'h3a64a808),
	.w2(32'h39465d51),
	.w3(32'h3a5cfb70),
	.w4(32'h39d28f6d),
	.w5(32'h3989eb0a),
	.w6(32'h3922ca60),
	.w7(32'hb8731ff0),
	.w8(32'hb80ddb6e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359ddad8),
	.w1(32'hb69e31a2),
	.w2(32'hb7472114),
	.w3(32'h371c5f0a),
	.w4(32'h361794e8),
	.w5(32'hb6fe031b),
	.w6(32'h37404fbd),
	.w7(32'h36ca5b26),
	.w8(32'hb6f7a427),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3930d5ca),
	.w1(32'h378815e1),
	.w2(32'h39bd3d83),
	.w3(32'h3977aaa5),
	.w4(32'h38ad9743),
	.w5(32'h3997bf85),
	.w6(32'hb80edeb0),
	.w7(32'hb8e6bc71),
	.w8(32'h39328fe2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3599f9ca),
	.w1(32'h36bb5a72),
	.w2(32'h36875995),
	.w3(32'hb5bb733b),
	.w4(32'h35aa7317),
	.w5(32'hb681a278),
	.w6(32'h3650371b),
	.w7(32'hb6551fc3),
	.w8(32'hb59dc7ab),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995c958),
	.w1(32'hb97d51fa),
	.w2(32'h38ec4fa4),
	.w3(32'hb9adbd79),
	.w4(32'hb7e6560a),
	.w5(32'h3991d23b),
	.w6(32'hba3691cc),
	.w7(32'hb9cc2f1f),
	.w8(32'h38d89bba),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7cf05),
	.w1(32'hb7eeb2ae),
	.w2(32'h39a317ce),
	.w3(32'hb875eb42),
	.w4(32'hb8d823c1),
	.w5(32'h392ca342),
	.w6(32'hb9b9e933),
	.w7(32'hb9b73569),
	.w8(32'hb7fd24fe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39273844),
	.w1(32'h39cd1bbd),
	.w2(32'h39ab9c09),
	.w3(32'h391251cf),
	.w4(32'h3989c38d),
	.w5(32'h396da2f9),
	.w6(32'hb81b59ec),
	.w7(32'h39181b4d),
	.w8(32'h38f09918),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391f6b9d),
	.w1(32'h36c77b9c),
	.w2(32'h38cb57e8),
	.w3(32'h3947a9ff),
	.w4(32'hb6a03d15),
	.w5(32'h38a2d020),
	.w6(32'h39968c9e),
	.w7(32'h38b7829e),
	.w8(32'h392a99cf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b76c0),
	.w1(32'h3a35aa54),
	.w2(32'h3a3f3af1),
	.w3(32'h3a627ff3),
	.w4(32'h3a007d99),
	.w5(32'h398923dd),
	.w6(32'h3a431e0f),
	.w7(32'h39b48888),
	.w8(32'h394b8b83),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357dfcfd),
	.w1(32'hb58cbb99),
	.w2(32'hb6399fc2),
	.w3(32'hb5c590a3),
	.w4(32'hb60483dc),
	.w5(32'hb6d08522),
	.w6(32'h3650ceb3),
	.w7(32'h346861f7),
	.w8(32'hb6b55b81),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bfa8a),
	.w1(32'h39aa13b0),
	.w2(32'h39f4c0eb),
	.w3(32'h398d7d12),
	.w4(32'h38f0ff22),
	.w5(32'h3973e80c),
	.w6(32'hb9ac2460),
	.w7(32'hb9ee3004),
	.w8(32'h36ceadda),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954c7f1),
	.w1(32'h374bf111),
	.w2(32'h39309560),
	.w3(32'hb6cc9f6f),
	.w4(32'hb8cde2df),
	.w5(32'h3814bd32),
	.w6(32'hb99b9b15),
	.w7(32'hb9ac3e5d),
	.w8(32'hb89466b2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37174bd9),
	.w1(32'hb6b45af6),
	.w2(32'h36664ef3),
	.w3(32'h362a205b),
	.w4(32'hb765e3da),
	.w5(32'h35e221ac),
	.w6(32'h36fff310),
	.w7(32'hb71f258f),
	.w8(32'h364ef34a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb603bbe9),
	.w1(32'h3723b627),
	.w2(32'h372c311e),
	.w3(32'h31867b57),
	.w4(32'h36d4d21a),
	.w5(32'h3691a4c0),
	.w6(32'hb65c1583),
	.w7(32'h34d6641a),
	.w8(32'hb4b87168),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34bdae3f),
	.w1(32'hb89d191b),
	.w2(32'hb6492caa),
	.w3(32'h385b4009),
	.w4(32'hb8803d9a),
	.w5(32'h3801c606),
	.w6(32'h38d973e5),
	.w7(32'h36545317),
	.w8(32'h3844f3fa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cdaf3),
	.w1(32'h3a10d4f8),
	.w2(32'h3a52d05b),
	.w3(32'h39cb7647),
	.w4(32'hb843463f),
	.w5(32'h39ce0532),
	.w6(32'h38f2d112),
	.w7(32'hb97c7f5e),
	.w8(32'h39c9b8d2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac8ca1),
	.w1(32'hb85add69),
	.w2(32'h3982530e),
	.w3(32'h38cab8b5),
	.w4(32'hb8899469),
	.w5(32'h392e55b0),
	.w6(32'h38ad881b),
	.w7(32'hb88b5bfc),
	.w8(32'h39379ed2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a05ffa),
	.w1(32'hb87ef5cb),
	.w2(32'h39949b1f),
	.w3(32'h39ea5542),
	.w4(32'hb8fc1298),
	.w5(32'h3953904b),
	.w6(32'h3a650b09),
	.w7(32'h3974854b),
	.w8(32'h39f3961f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c1af61),
	.w1(32'h378d34cb),
	.w2(32'h37721bd2),
	.w3(32'h346200e4),
	.w4(32'h37acbdc6),
	.w5(32'h379f3167),
	.w6(32'h366925c0),
	.w7(32'h37a6c5a2),
	.w8(32'h37961f95),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c24211),
	.w1(32'hb6a00fa2),
	.w2(32'hb6ca15ef),
	.w3(32'hb6937185),
	.w4(32'hb675ed64),
	.w5(32'hb6c1d53f),
	.w6(32'h344178e1),
	.w7(32'hb5f46919),
	.w8(32'hb68b4316),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7fb8345),
	.w1(32'hba1b05ab),
	.w2(32'hb90f5b81),
	.w3(32'h39db64c4),
	.w4(32'hb9da84a1),
	.w5(32'hb99337eb),
	.w6(32'h390535e9),
	.w7(32'hba01c323),
	.w8(32'hb9d2e75e),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37797430),
	.w1(32'hb74f5977),
	.w2(32'hb7c1bc92),
	.w3(32'h378e6618),
	.w4(32'hb78c98a7),
	.w5(32'hb7d652a3),
	.w6(32'h37d014af),
	.w7(32'hb7042f50),
	.w8(32'hb7b696a2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c2aa4),
	.w1(32'hba1d10bf),
	.w2(32'hb9805e84),
	.w3(32'h391bcfcc),
	.w4(32'hb9a2c661),
	.w5(32'hb8107b66),
	.w6(32'h39c64dfb),
	.w7(32'h3808d50a),
	.w8(32'h391ed5e3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f03f1e),
	.w1(32'hb5a77c6c),
	.w2(32'hb593a784),
	.w3(32'hb5a6c3b9),
	.w4(32'hb58efd76),
	.w5(32'hb59539c2),
	.w6(32'hb53098e2),
	.w7(32'hb496ef24),
	.w8(32'h353709c3),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65c6584),
	.w1(32'hb5bcf09b),
	.w2(32'hb606bb5f),
	.w3(32'h351ef601),
	.w4(32'hb53e80bd),
	.w5(32'hb5a2125f),
	.w6(32'h358922f6),
	.w7(32'h34aef0ca),
	.w8(32'hb4dc847c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388b6e29),
	.w1(32'h38239215),
	.w2(32'h393e0cdd),
	.w3(32'h38203480),
	.w4(32'h37b1d328),
	.w5(32'h38dab2c1),
	.w6(32'hb8cdf837),
	.w7(32'hb8b42d12),
	.w8(32'h3824bf59),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fa7cf),
	.w1(32'h394e30c7),
	.w2(32'h39122cf8),
	.w3(32'h395bc938),
	.w4(32'h3902df40),
	.w5(32'h38d1a88b),
	.w6(32'h39995de6),
	.w7(32'h3948a9d5),
	.w8(32'h392c860c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a4d255),
	.w1(32'hb75bae7a),
	.w2(32'h371dafe2),
	.w3(32'h385a0631),
	.w4(32'h388643ea),
	.w5(32'h3818d25d),
	.w6(32'hb7abbdb6),
	.w7(32'hb6495075),
	.w8(32'h36b47912),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e47edd),
	.w1(32'h38deda21),
	.w2(32'h391d1b9c),
	.w3(32'hb9672599),
	.w4(32'hb7f0a284),
	.w5(32'h38c5e725),
	.w6(32'hb9b9690d),
	.w7(32'hb99243b3),
	.w8(32'hb8a0292a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b989a),
	.w1(32'h398fbde5),
	.w2(32'hb7dcc454),
	.w3(32'h39f7c1ae),
	.w4(32'hb9044a6b),
	.w5(32'h38ab6bca),
	.w6(32'h38849341),
	.w7(32'hba3b9ebf),
	.w8(32'h398068b6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dd3cb7),
	.w1(32'hb9ffb5d6),
	.w2(32'h39845b75),
	.w3(32'h3a00c985),
	.w4(32'hb9ff7588),
	.w5(32'h39166080),
	.w6(32'h3a8d3316),
	.w7(32'h393bfc20),
	.w8(32'h39e983c4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9deb77a),
	.w1(32'hba455fc8),
	.w2(32'h38e9ee3e),
	.w3(32'hb894474b),
	.w4(32'hba2b6d0a),
	.w5(32'h38364393),
	.w6(32'h394072af),
	.w7(32'hb92d7003),
	.w8(32'h397322ef),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378ead56),
	.w1(32'hb8bddaa9),
	.w2(32'hb80d7a6d),
	.w3(32'h3891a2f8),
	.w4(32'hb8d3e9ab),
	.w5(32'hb8208b15),
	.w6(32'h3928d99d),
	.w7(32'hb729790f),
	.w8(32'h37ad936a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63fbaa5),
	.w1(32'hb5e76a53),
	.w2(32'hb695023f),
	.w3(32'hb55080e3),
	.w4(32'h356dae01),
	.w5(32'hb627b27b),
	.w6(32'hb5c1996c),
	.w7(32'hb5348fa9),
	.w8(32'hb64186be),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b4ed87),
	.w1(32'hb698ac2f),
	.w2(32'hb6aa25e2),
	.w3(32'hb61221c7),
	.w4(32'hb65cda07),
	.w5(32'hb6b101ee),
	.w6(32'h3659ed91),
	.w7(32'h35b3d68b),
	.w8(32'hb5447f25),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ddf40d),
	.w1(32'hb6b96cc0),
	.w2(32'h36e5e297),
	.w3(32'h37e206f6),
	.w4(32'hb6670f38),
	.w5(32'h37443c7f),
	.w6(32'h37a2403e),
	.w7(32'h37409baf),
	.w8(32'h3750c2d3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f02215),
	.w1(32'h3908ce79),
	.w2(32'h3a1fa68d),
	.w3(32'h39760a8c),
	.w4(32'hb946382c),
	.w5(32'h389c91f8),
	.w6(32'hb9296bc5),
	.w7(32'hb9e5a3c6),
	.w8(32'hb882814a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390fae02),
	.w1(32'hb89c4d40),
	.w2(32'h39681a5d),
	.w3(32'h39577e06),
	.w4(32'hb8def1dd),
	.w5(32'h3919eb66),
	.w6(32'h39cc941f),
	.w7(32'h38c812bc),
	.w8(32'h39b241fe),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a53388),
	.w1(32'h3896aa4c),
	.w2(32'h39765936),
	.w3(32'h379c287c),
	.w4(32'hb919383d),
	.w5(32'h38813d0f),
	.w6(32'h3991f7e6),
	.w7(32'hb82be526),
	.w8(32'h3979f213),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dc09b),
	.w1(32'h38c6f69f),
	.w2(32'h39a27d8c),
	.w3(32'h39aebc8f),
	.w4(32'h38349f53),
	.w5(32'h395ce662),
	.w6(32'h399d86b7),
	.w7(32'h38c1899b),
	.w8(32'h3956ea30),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de1e55),
	.w1(32'h392e8870),
	.w2(32'h39fe78e4),
	.w3(32'h37dae2ae),
	.w4(32'hb867df72),
	.w5(32'h398637e0),
	.w6(32'hba2cd490),
	.w7(32'hba2c7b8c),
	.w8(32'hb89ed34c),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35677846),
	.w1(32'h358a8e99),
	.w2(32'hb65b0c51),
	.w3(32'h35fa65ec),
	.w4(32'h361d4725),
	.w5(32'hb58fddb9),
	.w6(32'h345debd1),
	.w7(32'h35209f16),
	.w8(32'hb507396b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7372446),
	.w1(32'hb6e12c3a),
	.w2(32'hb799d557),
	.w3(32'hb683ea19),
	.w4(32'hb6ff1a69),
	.w5(32'hb78607d9),
	.w6(32'hb50a40e5),
	.w7(32'hb5858f25),
	.w8(32'hb6a57007),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36562cee),
	.w1(32'h36b073e9),
	.w2(32'h3363b536),
	.w3(32'h36d38e66),
	.w4(32'h36d5f4f0),
	.w5(32'h35d6831c),
	.w6(32'h36b3d189),
	.w7(32'h369911fc),
	.w8(32'h36311531),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7ed7d),
	.w1(32'h39099224),
	.w2(32'h39954f4e),
	.w3(32'h3961d14e),
	.w4(32'h38918575),
	.w5(32'h395a027e),
	.w6(32'h39644669),
	.w7(32'h3775c711),
	.w8(32'h3912f9be),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925a9ea),
	.w1(32'h38dea9d4),
	.w2(32'h372508a9),
	.w3(32'h38bbe165),
	.w4(32'h38847241),
	.w5(32'hb7256635),
	.w6(32'h37e76e07),
	.w7(32'h35bbf945),
	.w8(32'hb7bf6ddb),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d9f2c7),
	.w1(32'h394c77c2),
	.w2(32'h3a093fe7),
	.w3(32'h398468fb),
	.w4(32'h38e4301b),
	.w5(32'h39a87336),
	.w6(32'hb9c1e893),
	.w7(32'hb9a1bdf4),
	.w8(32'h38def302),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390dbf3e),
	.w1(32'hb67eb84a),
	.w2(32'h38e5f201),
	.w3(32'h3844499a),
	.w4(32'hb7b950af),
	.w5(32'h388ae814),
	.w6(32'h36754d63),
	.w7(32'hb8948c94),
	.w8(32'h382b974b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb505f4d3),
	.w1(32'hb709158a),
	.w2(32'hb723cc64),
	.w3(32'h368fd424),
	.w4(32'hb7719f24),
	.w5(32'hb727ee31),
	.w6(32'h37c4eb56),
	.w7(32'h36d448b7),
	.w8(32'h36656786),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35b29011),
	.w1(32'h3472235b),
	.w2(32'hb5221534),
	.w3(32'h35ba8af5),
	.w4(32'hb4424368),
	.w5(32'h34b4fdbc),
	.w6(32'h3685694a),
	.w7(32'h362720c0),
	.w8(32'h36281e44),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb816ee76),
	.w1(32'hb875cf71),
	.w2(32'hb68f1899),
	.w3(32'hb7ae69ef),
	.w4(32'hb82a3258),
	.w5(32'hb6457dba),
	.w6(32'hb6d229a2),
	.w7(32'hb7619cc5),
	.w8(32'h37a50e04),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7352d2b),
	.w1(32'hb82970f1),
	.w2(32'hb7f3b746),
	.w3(32'h363ab0c2),
	.w4(32'hb82a9814),
	.w5(32'hb7f5eed8),
	.w6(32'h37638471),
	.w7(32'hb7984f96),
	.w8(32'hb781716e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70017fa),
	.w1(32'hb77b786b),
	.w2(32'hb71bf503),
	.w3(32'h3609c342),
	.w4(32'h36d2ae93),
	.w5(32'h376aee0d),
	.w6(32'hb70aff48),
	.w7(32'hb502a3f3),
	.w8(32'h37a2a0ab),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398827ae),
	.w1(32'h39107db5),
	.w2(32'h391f5771),
	.w3(32'h39098d40),
	.w4(32'h378aeb27),
	.w5(32'h3884d456),
	.w6(32'hb8acd6ea),
	.w7(32'hb91879fb),
	.w8(32'hb616519d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24c30e),
	.w1(32'h39364a00),
	.w2(32'h3a0c9f95),
	.w3(32'h39fe3077),
	.w4(32'h38e00b72),
	.w5(32'h39991400),
	.w6(32'h396aebd4),
	.w7(32'hb8b33042),
	.w8(32'h39370100),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61d8c5c),
	.w1(32'hb6365c47),
	.w2(32'hb693c55d),
	.w3(32'hb5470330),
	.w4(32'hb5462351),
	.w5(32'hb6648f87),
	.w6(32'h342fcab6),
	.w7(32'h34f926cc),
	.w8(32'hb62fe3f6),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63f2e80),
	.w1(32'hb643cea2),
	.w2(32'hb60b6c30),
	.w3(32'hb5de6d98),
	.w4(32'hb5fda49e),
	.w5(32'hb5e41ccf),
	.w6(32'hb41401cf),
	.w7(32'hb5143a0f),
	.w8(32'hb5c3833e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6257c02),
	.w1(32'hb56a3736),
	.w2(32'hb62f36a7),
	.w3(32'hb598528a),
	.w4(32'hb4969553),
	.w5(32'hb5acb788),
	.w6(32'hb61f91ab),
	.w7(32'hb3e8d3d8),
	.w8(32'hb5d7f08b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68220d7),
	.w1(32'hb6021be5),
	.w2(32'hb61ef0eb),
	.w3(32'hb6537d7e),
	.w4(32'hb61c9b84),
	.w5(32'hb6447633),
	.w6(32'hb6324269),
	.w7(32'hb4ace8ff),
	.w8(32'hb61cb621),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2a7bf),
	.w1(32'h39bd2a6e),
	.w2(32'h3a4c83dc),
	.w3(32'h3a889382),
	.w4(32'h3a2430a7),
	.w5(32'h3a08ee55),
	.w6(32'h391abe45),
	.w7(32'h399acb6f),
	.w8(32'h393646b7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a255e0e),
	.w1(32'h3a227c7d),
	.w2(32'h3a1e9b4a),
	.w3(32'h37db760f),
	.w4(32'h3972fc1c),
	.w5(32'h39d44057),
	.w6(32'h39784e52),
	.w7(32'h38b84b8c),
	.w8(32'h3988f31f),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2db10c),
	.w1(32'h39c80c6a),
	.w2(32'h3a261b1b),
	.w3(32'h3983e49f),
	.w4(32'h3910fbbd),
	.w5(32'h39ac7dad),
	.w6(32'h39049fe1),
	.w7(32'hb8e5f168),
	.w8(32'h3974c50f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4747e),
	.w1(32'hbae28922),
	.w2(32'hbc0f9f47),
	.w3(32'h3995e3d5),
	.w4(32'h3b0324f1),
	.w5(32'hbb01ba65),
	.w6(32'h3a870d53),
	.w7(32'hbbc32180),
	.w8(32'hbbd4c4ac),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80688a),
	.w1(32'h3ae87389),
	.w2(32'h3bb706dc),
	.w3(32'hbbe07c7d),
	.w4(32'h3ac05681),
	.w5(32'hbbc73ab8),
	.w6(32'hbb40a8fe),
	.w7(32'h3b2c1fe7),
	.w8(32'h3a2047b5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d529),
	.w1(32'hbb6995b7),
	.w2(32'hbbb5d115),
	.w3(32'hb7c301eb),
	.w4(32'hbbaf8d96),
	.w5(32'hbbe8ef41),
	.w6(32'hbac7a2ac),
	.w7(32'hbb5588be),
	.w8(32'hbbcbd9f8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9564b1),
	.w1(32'hba3ea961),
	.w2(32'hbb11bab1),
	.w3(32'hbb3cf2f2),
	.w4(32'hbb1dc154),
	.w5(32'h3b36e935),
	.w6(32'hbc1acd3d),
	.w7(32'hbbfca976),
	.w8(32'hbb9dcaed),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91e7c3),
	.w1(32'hbad9193f),
	.w2(32'hba914880),
	.w3(32'hbc2d23c2),
	.w4(32'hba4ddb85),
	.w5(32'h3c1ab56e),
	.w6(32'hbbfb32fa),
	.w7(32'hba264b15),
	.w8(32'h3aefe410),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3073bc),
	.w1(32'h3b7ecf13),
	.w2(32'h3b465946),
	.w3(32'h3b8bcb62),
	.w4(32'h3a4b270c),
	.w5(32'h3c491f80),
	.w6(32'hbb451b8a),
	.w7(32'hbbacfe29),
	.w8(32'h3b904878),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7d6db),
	.w1(32'h3b9fbb06),
	.w2(32'h3b2038f7),
	.w3(32'h3c0fb1df),
	.w4(32'h3b4c51fd),
	.w5(32'h3c144896),
	.w6(32'h3c279281),
	.w7(32'h3c023f40),
	.w8(32'h3c2b91dc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecdcce),
	.w1(32'hbc061900),
	.w2(32'hbc5359b4),
	.w3(32'h3bee640c),
	.w4(32'hbc3193b1),
	.w5(32'hbb512dd3),
	.w6(32'h3b7a6b14),
	.w7(32'hbc2b7c10),
	.w8(32'hbc430b33),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6af0be),
	.w1(32'h3bc9c4bf),
	.w2(32'hbb29c83c),
	.w3(32'hbc5d4ea2),
	.w4(32'hbb5b1139),
	.w5(32'hbc69731b),
	.w6(32'hbc11133e),
	.w7(32'h3b7a3149),
	.w8(32'h3bd36f59),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4fa5e),
	.w1(32'hbb1b05df),
	.w2(32'hbadd9f86),
	.w3(32'h3b63c031),
	.w4(32'h3bb0144e),
	.w5(32'h3bde987f),
	.w6(32'h3c019fbe),
	.w7(32'h3b97bc19),
	.w8(32'h3b4c9b5f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96a0747),
	.w1(32'hbbf671b2),
	.w2(32'h3bb275d4),
	.w3(32'h3ad5710c),
	.w4(32'hbc1de66e),
	.w5(32'hb98f5104),
	.w6(32'h3bb2639e),
	.w7(32'hbbbaaf6b),
	.w8(32'hbb937711),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd9532),
	.w1(32'hbbc76ca1),
	.w2(32'hbb731d3d),
	.w3(32'hbb6a64f6),
	.w4(32'hbbe62082),
	.w5(32'hbc1486df),
	.w6(32'hbb5876ad),
	.w7(32'hbba1fa01),
	.w8(32'hbba6e305),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca9679),
	.w1(32'h3b072321),
	.w2(32'h3b2abacd),
	.w3(32'hbc32bc5b),
	.w4(32'h3b669321),
	.w5(32'hbb1892e3),
	.w6(32'hbc371113),
	.w7(32'hbaf45214),
	.w8(32'hbb912be7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac700f0),
	.w1(32'h3bc677a0),
	.w2(32'h3baa11c1),
	.w3(32'hbbafe276),
	.w4(32'h3bb0a0ab),
	.w5(32'h3b9420ea),
	.w6(32'hba952db1),
	.w7(32'h3babfab2),
	.w8(32'hbac235da),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0662b),
	.w1(32'hbb7aebda),
	.w2(32'hbc219634),
	.w3(32'hba9b9353),
	.w4(32'hbbc07266),
	.w5(32'hbb6f87b9),
	.w6(32'hbb0d724d),
	.w7(32'h3b10eb04),
	.w8(32'hba3eaf8f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d90322),
	.w1(32'h3b7e174e),
	.w2(32'h3a9a60e6),
	.w3(32'hbbc7e21c),
	.w4(32'hbad3e711),
	.w5(32'hbb722d08),
	.w6(32'hba970146),
	.w7(32'hbb89ab58),
	.w8(32'h3ab1f74a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d823f),
	.w1(32'hbc28ba9b),
	.w2(32'h3bfe138a),
	.w3(32'hbb872c46),
	.w4(32'h3c14a09a),
	.w5(32'h3bc2fecd),
	.w6(32'h3b07fc49),
	.w7(32'hbc10021b),
	.w8(32'hbbb7a6c9),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b54a65),
	.w1(32'h3b1b6185),
	.w2(32'hbb5f11de),
	.w3(32'hbb7c131b),
	.w4(32'h3ab6a789),
	.w5(32'hbc9863dd),
	.w6(32'h3a7adab6),
	.w7(32'hbb37a49d),
	.w8(32'hbb87ed8b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacaeb6),
	.w1(32'h3b0d0f60),
	.w2(32'h3b24fd93),
	.w3(32'hbc038f36),
	.w4(32'h3c217259),
	.w5(32'h3aaf8f04),
	.w6(32'hbbd15a33),
	.w7(32'hbadf46ff),
	.w8(32'h3b813a3c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b2b6f),
	.w1(32'hbbffc171),
	.w2(32'hbb83bbfe),
	.w3(32'hbba1ee3a),
	.w4(32'hbb7d0a99),
	.w5(32'hbabff11a),
	.w6(32'hbbeb6ffd),
	.w7(32'hbc207696),
	.w8(32'hbc1f1049),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a713e),
	.w1(32'h3b0d7476),
	.w2(32'h3b2a3a18),
	.w3(32'hbb87fddf),
	.w4(32'h3abe9e89),
	.w5(32'hbb95d787),
	.w6(32'hbae7d47d),
	.w7(32'hb9c76417),
	.w8(32'hbb890d60),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bd81e),
	.w1(32'h3b988ee9),
	.w2(32'hbac4b473),
	.w3(32'hbb2ffbf4),
	.w4(32'hbad1a6d7),
	.w5(32'h3bb8a308),
	.w6(32'h3b207f81),
	.w7(32'hbb01cad5),
	.w8(32'hbb1a0da7),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d305),
	.w1(32'hbb0f8d0a),
	.w2(32'hbbb30c4b),
	.w3(32'h3bc2388e),
	.w4(32'h3ace97cd),
	.w5(32'h3ad78ea8),
	.w6(32'hbb2a2c92),
	.w7(32'hbb6594ad),
	.w8(32'h3a8eb824),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e009f),
	.w1(32'h3b5f4265),
	.w2(32'h3b9a2860),
	.w3(32'h36bc9bd1),
	.w4(32'h3bfac9d6),
	.w5(32'h3c3293e6),
	.w6(32'hbab74ba1),
	.w7(32'h3be53ebc),
	.w8(32'hbb80cafa),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f4f29),
	.w1(32'h3b166f7e),
	.w2(32'h3be3fdc9),
	.w3(32'h3ba4d4f6),
	.w4(32'h3bff180a),
	.w5(32'h3b9b22dc),
	.w6(32'hbafbe7f4),
	.w7(32'h3b84f9ab),
	.w8(32'h390c8e02),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba986dc1),
	.w1(32'hbadd6938),
	.w2(32'hbbc0d775),
	.w3(32'h3b09c5b4),
	.w4(32'hbc09d83b),
	.w5(32'hbb16fd52),
	.w6(32'hbb133c80),
	.w7(32'hba88e4fa),
	.w8(32'hbbf2e5b6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaca3dc),
	.w1(32'hb98d721f),
	.w2(32'hbc111128),
	.w3(32'h3afcf26f),
	.w4(32'hbbad89b0),
	.w5(32'h3b7e5243),
	.w6(32'hbb868d39),
	.w7(32'h3ac6235d),
	.w8(32'h3bfe3b13),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83fa0a9),
	.w1(32'hbb02cd3d),
	.w2(32'h3badb7de),
	.w3(32'h3bea2e11),
	.w4(32'h3b23a702),
	.w5(32'h3b26d9fc),
	.w6(32'h3aa17230),
	.w7(32'hbac7ffc7),
	.w8(32'hbb2e45c7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bc6b2),
	.w1(32'hbbc57ebb),
	.w2(32'hbc186fb0),
	.w3(32'hb9c9a783),
	.w4(32'hbb35a595),
	.w5(32'hbb0bfa11),
	.w6(32'hbb65b87e),
	.w7(32'hbbfa531f),
	.w8(32'hbc0aa5da),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828563),
	.w1(32'h3bc2a21a),
	.w2(32'h3bf009ae),
	.w3(32'hbbd08c37),
	.w4(32'h3c08ab3d),
	.w5(32'hbb457058),
	.w6(32'h38362829),
	.w7(32'hbb3c756e),
	.w8(32'h3b47836e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10976e),
	.w1(32'h3beec0fe),
	.w2(32'hbad89b63),
	.w3(32'hba75cf77),
	.w4(32'hba935c5b),
	.w5(32'h3c385a92),
	.w6(32'hbb3d7557),
	.w7(32'h3aa2a10a),
	.w8(32'h3b254571),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74b9f1),
	.w1(32'h3a966719),
	.w2(32'hba0c0ff7),
	.w3(32'hbbf60d0b),
	.w4(32'hba954ce5),
	.w5(32'h3a111239),
	.w6(32'h3bc7b7aa),
	.w7(32'hbada4d47),
	.w8(32'hbbe757a7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba303982),
	.w1(32'hba2f0807),
	.w2(32'h3a4ad3a6),
	.w3(32'h3b8fc194),
	.w4(32'h3b99048f),
	.w5(32'h3bbd28dd),
	.w6(32'hbb3eef4b),
	.w7(32'h3a9655d9),
	.w8(32'h3b1175f2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dbd84d),
	.w1(32'hba8b2c84),
	.w2(32'hbaadd44d),
	.w3(32'hbbfdf0fc),
	.w4(32'h3a2f21ae),
	.w5(32'h3b5ae1e9),
	.w6(32'hba644f57),
	.w7(32'hbb46cb75),
	.w8(32'h3bdac9e9),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e0e5f),
	.w1(32'h3b17a677),
	.w2(32'hbae4b9a0),
	.w3(32'hbb999525),
	.w4(32'h3b90e81c),
	.w5(32'h389af1ee),
	.w6(32'h3a9a4fdb),
	.w7(32'h3b20f5f8),
	.w8(32'h3a29080c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b483074),
	.w1(32'h3b79c7ea),
	.w2(32'h3c145c29),
	.w3(32'hbbcf72fe),
	.w4(32'h3c009bf6),
	.w5(32'h3baa785a),
	.w6(32'h3aeda9ba),
	.w7(32'h3bd82d9c),
	.w8(32'hba923a21),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccdc2b),
	.w1(32'h3be9627e),
	.w2(32'h3c47dd28),
	.w3(32'h3b89c69c),
	.w4(32'h3c47646b),
	.w5(32'h3be08eab),
	.w6(32'h3bd0053e),
	.w7(32'h3b925f1a),
	.w8(32'hba94c3d4),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba594d3),
	.w1(32'h3bb97dc3),
	.w2(32'h3b91bf98),
	.w3(32'h3a82442a),
	.w4(32'h3b8d3612),
	.w5(32'hbb341273),
	.w6(32'h3b16f5a8),
	.w7(32'h3c0cadfc),
	.w8(32'h3ae772bc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b255efa),
	.w1(32'h3a524a78),
	.w2(32'hbc12a2c2),
	.w3(32'h389b77f4),
	.w4(32'h3b3d5e0e),
	.w5(32'hbc39e5d8),
	.w6(32'h3a362c33),
	.w7(32'hba34fe0a),
	.w8(32'hbc08d845),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc3aa8),
	.w1(32'h3c08ce11),
	.w2(32'h3ab6c56e),
	.w3(32'hba0a9de8),
	.w4(32'h3b18076d),
	.w5(32'h3afe8d2a),
	.w6(32'h3b4e27be),
	.w7(32'h3b1ec954),
	.w8(32'h3baad01d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920d4d),
	.w1(32'h3a9bf432),
	.w2(32'hbaa4eb4d),
	.w3(32'hb9b56eb0),
	.w4(32'hbb17984d),
	.w5(32'hbc48f8bd),
	.w6(32'h3992a374),
	.w7(32'hbae93a7f),
	.w8(32'hbbecbac6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2576f),
	.w1(32'hbc8eb3fe),
	.w2(32'hbc2d93fb),
	.w3(32'hb9db1852),
	.w4(32'hbc0fb3e9),
	.w5(32'hbba7ea32),
	.w6(32'h3afa3eb8),
	.w7(32'hbbd64670),
	.w8(32'h3b7114ba),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75a62),
	.w1(32'hbc1142da),
	.w2(32'hbbdb04d5),
	.w3(32'hbc0ff40e),
	.w4(32'hbbed0b3b),
	.w5(32'hbc161210),
	.w6(32'hbc1fd7de),
	.w7(32'h3936b241),
	.w8(32'hbbb717f9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e233f8),
	.w1(32'hbb1b97eb),
	.w2(32'h3ad82c35),
	.w3(32'hbb493f10),
	.w4(32'h3a3599a0),
	.w5(32'h3c844543),
	.w6(32'hbb154b69),
	.w7(32'hbb0b8668),
	.w8(32'h3bbdc0a7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fa83a),
	.w1(32'h3bb7e19b),
	.w2(32'h3c119d1e),
	.w3(32'h3ae964ff),
	.w4(32'hba27582a),
	.w5(32'h3c6d86ac),
	.w6(32'h3a6cb0a4),
	.w7(32'h3ba16354),
	.w8(32'hbad58d1b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf2c11),
	.w1(32'hbb7a1a36),
	.w2(32'h3c1151a3),
	.w3(32'hba547612),
	.w4(32'hba13de7f),
	.w5(32'h3cc9f343),
	.w6(32'hbaa568fb),
	.w7(32'h3a379760),
	.w8(32'hbc10d462),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b5344),
	.w1(32'hbc021ecc),
	.w2(32'hbbe87fcc),
	.w3(32'hbaca2bd0),
	.w4(32'hbb9f084c),
	.w5(32'hbc210677),
	.w6(32'hbbd3b284),
	.w7(32'hbb8aca52),
	.w8(32'hbbaefc1f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0bd3),
	.w1(32'h3bb89874),
	.w2(32'h3b2fd397),
	.w3(32'hbbd07561),
	.w4(32'h3b2ba7e4),
	.w5(32'h3ce0eee5),
	.w6(32'hbbdbe260),
	.w7(32'h3bc98301),
	.w8(32'h3bd67719),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951364f),
	.w1(32'h3b159ec8),
	.w2(32'h3c0a92ec),
	.w3(32'h3bd1fc82),
	.w4(32'h39ea9989),
	.w5(32'h3bf79b78),
	.w6(32'h3c1e4099),
	.w7(32'h3a15afde),
	.w8(32'hbba6ac1b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3de05f),
	.w1(32'hbb49e5da),
	.w2(32'hbb35fd76),
	.w3(32'h3a5f6ab2),
	.w4(32'h3b09a120),
	.w5(32'h3a9dabd2),
	.w6(32'hbb95ee71),
	.w7(32'h3b54a46f),
	.w8(32'hb9f58e86),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa69ee2),
	.w1(32'hbb357d4e),
	.w2(32'hbb86a57f),
	.w3(32'h3aa49eff),
	.w4(32'hbb4147cd),
	.w5(32'hbbe9b149),
	.w6(32'hbae41075),
	.w7(32'hbacab5e9),
	.w8(32'h3a91604d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d601f1),
	.w1(32'hbbc0125f),
	.w2(32'hbc4a6f2a),
	.w3(32'h3af71a73),
	.w4(32'hbc131603),
	.w5(32'hbbdd7c37),
	.w6(32'h3ae5ac36),
	.w7(32'hbc1f9fbe),
	.w8(32'hbbc93aec),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc64871),
	.w1(32'hbb9957ea),
	.w2(32'hbbd582ca),
	.w3(32'hbc235909),
	.w4(32'hbbe53387),
	.w5(32'hbc124d76),
	.w6(32'hbb86bc36),
	.w7(32'hbbe5ac50),
	.w8(32'hba4b2ff3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb250ae),
	.w1(32'h39efa709),
	.w2(32'h3b591840),
	.w3(32'hbb90889e),
	.w4(32'hbb76ab93),
	.w5(32'hbc0a3afd),
	.w6(32'hbb5b31ea),
	.w7(32'hb9e5e447),
	.w8(32'h3b35911d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2a8de),
	.w1(32'hbc01a1ee),
	.w2(32'hba876700),
	.w3(32'hbbbfff6a),
	.w4(32'h3b3aed36),
	.w5(32'hb9da18d8),
	.w6(32'hbb787d02),
	.w7(32'hbba3e4cb),
	.w8(32'hbb376d4a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45a227),
	.w1(32'h3c1565d0),
	.w2(32'hbbe07af9),
	.w3(32'h3b191327),
	.w4(32'hbbae6354),
	.w5(32'hbc712eaf),
	.w6(32'hbb1a2fcb),
	.w7(32'hb97e0db1),
	.w8(32'hbb9f5bfd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46b979),
	.w1(32'hbbdb86ba),
	.w2(32'hba1378a1),
	.w3(32'hb9e9946a),
	.w4(32'hb93465c4),
	.w5(32'h3c4deca0),
	.w6(32'hb9a7607c),
	.w7(32'hbb22b93f),
	.w8(32'hbb1697a3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2dfda),
	.w1(32'h3c238de5),
	.w2(32'h3c818497),
	.w3(32'hba4d8f0a),
	.w4(32'h3c874223),
	.w5(32'h3c637014),
	.w6(32'hbb009c7c),
	.w7(32'h3c518aa0),
	.w8(32'h3ca1d501),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af93007),
	.w1(32'h380438da),
	.w2(32'hba9eaf1c),
	.w3(32'h3c1572db),
	.w4(32'hbb67c2ed),
	.w5(32'hbac27ab6),
	.w6(32'h3c3c5188),
	.w7(32'hbb8e149d),
	.w8(32'hbbe432a6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03ceef),
	.w1(32'hbbd46250),
	.w2(32'hbc02e79d),
	.w3(32'hbbe69fde),
	.w4(32'hbbed7f1d),
	.w5(32'hbbce6e91),
	.w6(32'hbc0a4fdf),
	.w7(32'hbb5809df),
	.w8(32'hba286f49),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd2bac),
	.w1(32'hbbf02e88),
	.w2(32'hb9df9ea8),
	.w3(32'hbbf88070),
	.w4(32'hbbad2164),
	.w5(32'h3b98ed2a),
	.w6(32'hb9dfe25f),
	.w7(32'hbbd73a9b),
	.w8(32'hbbcecc09),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe26bfd),
	.w1(32'h3ac57b52),
	.w2(32'hba991211),
	.w3(32'hbc377073),
	.w4(32'h3b39e78c),
	.w5(32'hbbd57632),
	.w6(32'hbc0a947b),
	.w7(32'hb9af3e27),
	.w8(32'hbbb40091),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08f06b),
	.w1(32'hbb232cce),
	.w2(32'hbb299435),
	.w3(32'h3bd9ca97),
	.w4(32'hbb2434fc),
	.w5(32'hb994be97),
	.w6(32'h3b2fd5fa),
	.w7(32'h3b3e80fb),
	.w8(32'hbb06754d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8df306),
	.w1(32'hbb388ac4),
	.w2(32'hbb5f5039),
	.w3(32'h3a99f783),
	.w4(32'hbbac189a),
	.w5(32'hba795114),
	.w6(32'hbb79f62b),
	.w7(32'hbbba4d31),
	.w8(32'h3b007566),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1ffd8),
	.w1(32'h3afe21f6),
	.w2(32'hbb3381de),
	.w3(32'hbb7f4f49),
	.w4(32'h3baf7e3f),
	.w5(32'h3d0f41fb),
	.w6(32'hba9b15e9),
	.w7(32'h3b20e7ee),
	.w8(32'hbb047d6a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7fbb7),
	.w1(32'hba6f81f1),
	.w2(32'hbb915334),
	.w3(32'hba46ee24),
	.w4(32'h3a62159f),
	.w5(32'hbb61d00b),
	.w6(32'h3a086158),
	.w7(32'h3b8f94b5),
	.w8(32'h3c011adb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae95f47),
	.w1(32'h3b1d7c11),
	.w2(32'h3b12c8c2),
	.w3(32'h3a3a13ba),
	.w4(32'h3c0fdbbb),
	.w5(32'h3bdea0d8),
	.w6(32'h395a864a),
	.w7(32'h3b826e69),
	.w8(32'h3b5ffaec),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991f91e),
	.w1(32'h3a74e62e),
	.w2(32'h3ba44d3a),
	.w3(32'h3c084d3b),
	.w4(32'h3b652ebf),
	.w5(32'h3c0ed36d),
	.w6(32'hbbbaf22b),
	.w7(32'h3b0c25ef),
	.w8(32'hbb88d4c1),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ac0b),
	.w1(32'hbafebc0d),
	.w2(32'hb9c05efb),
	.w3(32'h3a539d74),
	.w4(32'hbb107fef),
	.w5(32'h3b3c7541),
	.w6(32'hbb39c496),
	.w7(32'h3a9268d5),
	.w8(32'hbc001315),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd929e),
	.w1(32'h3a1d6a42),
	.w2(32'hbb4af4a2),
	.w3(32'hbbe221b7),
	.w4(32'hb795410a),
	.w5(32'h3c39f027),
	.w6(32'hbc6222e9),
	.w7(32'hbad91d18),
	.w8(32'h3b635795),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c6105),
	.w1(32'hbb54466f),
	.w2(32'hbc0a16dc),
	.w3(32'h3b0e1bd2),
	.w4(32'hbb9768c8),
	.w5(32'hbb66c0f8),
	.w6(32'h3b28fb03),
	.w7(32'hbbaa14e8),
	.w8(32'hbbbaf34e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6edbc),
	.w1(32'h3b8fea37),
	.w2(32'h3ad606b9),
	.w3(32'hbc14cdc7),
	.w4(32'h3b2c5149),
	.w5(32'h3acff4ce),
	.w6(32'hbbeeaf44),
	.w7(32'hba427eea),
	.w8(32'hbaa69b9f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba680f0f),
	.w1(32'h3ba8b999),
	.w2(32'h3b267343),
	.w3(32'hbb4247eb),
	.w4(32'h3ac7410c),
	.w5(32'h3b85cde3),
	.w6(32'hba139cb6),
	.w7(32'h3bfe52c8),
	.w8(32'h3ba35d6f),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfab5d),
	.w1(32'h3b1dbaf0),
	.w2(32'h3b27cbfb),
	.w3(32'h3abbcae9),
	.w4(32'h3941506e),
	.w5(32'hbc8a50df),
	.w6(32'h3b1ebe98),
	.w7(32'h39f8303c),
	.w8(32'h3b7fb6d5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8950d),
	.w1(32'h3a1304d2),
	.w2(32'hbad44f93),
	.w3(32'hba0b0371),
	.w4(32'hbb05b05d),
	.w5(32'hbc44b2d7),
	.w6(32'h3bfbc5ed),
	.w7(32'h3a2b491a),
	.w8(32'hbba06074),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1bb03a),
	.w1(32'h3b7169ea),
	.w2(32'hbb7477c9),
	.w3(32'hbb82c1a7),
	.w4(32'h3bc72716),
	.w5(32'hba51c4b0),
	.w6(32'h399cafaf),
	.w7(32'hbb68a6dd),
	.w8(32'hbad17f3e),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb729ebc),
	.w1(32'h3b244208),
	.w2(32'h3a9a2504),
	.w3(32'h3a9e1f8c),
	.w4(32'hba3fe337),
	.w5(32'h3ba901f9),
	.w6(32'hb9959f45),
	.w7(32'h3a99d576),
	.w8(32'hbba19cb5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3b5a4),
	.w1(32'h3a7ce7a4),
	.w2(32'hbaba11e4),
	.w3(32'h3c8ab0cc),
	.w4(32'h3b5aca7f),
	.w5(32'h3ae05ca6),
	.w6(32'h3b822c8e),
	.w7(32'h3b0eba52),
	.w8(32'h3b6cb01a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb372f99),
	.w1(32'h3aebdb2c),
	.w2(32'hbb7775ef),
	.w3(32'hbab5c626),
	.w4(32'hbadfa017),
	.w5(32'h3c869119),
	.w6(32'h3b98bdc3),
	.w7(32'hbbff8b63),
	.w8(32'h3abe5139),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b6e71),
	.w1(32'hbbf26119),
	.w2(32'hba6dc9a8),
	.w3(32'hbac369dc),
	.w4(32'hbbd57faf),
	.w5(32'h3bc1076f),
	.w6(32'h3c357e03),
	.w7(32'hbc04216d),
	.w8(32'hbc5c548d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb440f71),
	.w1(32'h3b02cd67),
	.w2(32'h3c28cae2),
	.w3(32'hbb86aede),
	.w4(32'h3a303d87),
	.w5(32'h3c82ee12),
	.w6(32'hbb5c014b),
	.w7(32'hbb19d40f),
	.w8(32'h3ad6acd5),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b936b32),
	.w1(32'h3b3c034f),
	.w2(32'hbbcba11b),
	.w3(32'h3b1255dd),
	.w4(32'hbbb6a27b),
	.w5(32'h3c7a8cd8),
	.w6(32'h3bef5ed5),
	.w7(32'hbb6b4ee6),
	.w8(32'h39cba487),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77f3d3),
	.w1(32'h3bb83cb2),
	.w2(32'h3bc9c0c2),
	.w3(32'hbb75eb2e),
	.w4(32'h3bf734e0),
	.w5(32'hbb96e2dc),
	.w6(32'hbc3165f5),
	.w7(32'h3ab4f13b),
	.w8(32'h3b3c4da3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1814fb),
	.w1(32'h3bde5ba5),
	.w2(32'h3c4d5656),
	.w3(32'hbb1248c9),
	.w4(32'h3a7d81a5),
	.w5(32'h3d03d1a9),
	.w6(32'hbb8c6596),
	.w7(32'h3bd9df60),
	.w8(32'h3c57f7e2),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc2260),
	.w1(32'h3bf25186),
	.w2(32'h3c23cc3f),
	.w3(32'h3c74a81d),
	.w4(32'h3c8af484),
	.w5(32'h3ceb460a),
	.w6(32'h3b32925f),
	.w7(32'hb9a07929),
	.w8(32'h3c2129d5),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c345a7f),
	.w1(32'hbbb68f1a),
	.w2(32'hb9789be0),
	.w3(32'h3c2b6f33),
	.w4(32'hbbb66b7d),
	.w5(32'hbb8a5342),
	.w6(32'hbc01fa9b),
	.w7(32'hbc171d07),
	.w8(32'hbc999962),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc81ed2),
	.w1(32'hba2fcccd),
	.w2(32'hbb6910e6),
	.w3(32'hbc35ade5),
	.w4(32'hbaa5bac8),
	.w5(32'hbb280f2c),
	.w6(32'hbc3f847b),
	.w7(32'h3a3f545d),
	.w8(32'hbb014778),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afee503),
	.w1(32'hb9b301dc),
	.w2(32'hbc4f6aaa),
	.w3(32'h3ad18482),
	.w4(32'hbbf1fb53),
	.w5(32'h3bf473ad),
	.w6(32'hbbd87047),
	.w7(32'hbabecc8c),
	.w8(32'h3a72acd2),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba69e7a),
	.w1(32'h3b52f5b7),
	.w2(32'h3b7fb52e),
	.w3(32'h3b2b7f60),
	.w4(32'h3b6a9bf5),
	.w5(32'h3ba03e5b),
	.w6(32'h3a444c97),
	.w7(32'h3ba5c5a2),
	.w8(32'hbbc8ab6f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53b91e),
	.w1(32'hbb6a4a04),
	.w2(32'hbc02383e),
	.w3(32'h3b28dfdd),
	.w4(32'h3b54d39e),
	.w5(32'h3c5d2643),
	.w6(32'hbabfbd17),
	.w7(32'hbbc07b26),
	.w8(32'hbc270fa3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa27d3),
	.w1(32'h3bdb5430),
	.w2(32'hb967503b),
	.w3(32'h3a9c50d3),
	.w4(32'h3b441d15),
	.w5(32'hbc17ec4d),
	.w6(32'hbbdb9349),
	.w7(32'h3b65d97a),
	.w8(32'hbb3652ce),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb847a14),
	.w1(32'hba7cb1ea),
	.w2(32'hbbe31d68),
	.w3(32'hbb11c162),
	.w4(32'h3b9ffd88),
	.w5(32'hbb5b5491),
	.w6(32'hbb0912bf),
	.w7(32'hbc0f3ff5),
	.w8(32'hbb99b254),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b11ff),
	.w1(32'h3c07cd7e),
	.w2(32'hba81b064),
	.w3(32'hbb67c994),
	.w4(32'hb818b8fd),
	.w5(32'h3ad857e6),
	.w6(32'hbb47f327),
	.w7(32'hbba24a17),
	.w8(32'hbc21411e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97174c),
	.w1(32'h3a78ec94),
	.w2(32'h3baef25f),
	.w3(32'hbc2afe75),
	.w4(32'h3a5748b2),
	.w5(32'h3bbccf11),
	.w6(32'hbc2f5eed),
	.w7(32'h3b677d3b),
	.w8(32'h3b40db04),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f2979),
	.w1(32'hbc037614),
	.w2(32'hbb7304b4),
	.w3(32'hbb7ab31f),
	.w4(32'hbb9cb624),
	.w5(32'hbc0a6286),
	.w6(32'hbb04ab01),
	.w7(32'hbb882b39),
	.w8(32'hbbbf8be7),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e2e5),
	.w1(32'h3b7e72ba),
	.w2(32'h3c12b24d),
	.w3(32'hbbc894d6),
	.w4(32'hbb62e393),
	.w5(32'h3c6806da),
	.w6(32'hbb4b8a79),
	.w7(32'h3a5bad47),
	.w8(32'h3bbd72ba),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca7cbb),
	.w1(32'h3c0e3372),
	.w2(32'h3b471eef),
	.w3(32'h3aa8b9d1),
	.w4(32'h3be72017),
	.w5(32'h3c443b40),
	.w6(32'hbb33fa4f),
	.w7(32'h3aeaed3e),
	.w8(32'h3bee8d03),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389d3e68),
	.w1(32'hb8a38b1a),
	.w2(32'hbc0b0b14),
	.w3(32'hbbbdea97),
	.w4(32'hbb0eed3a),
	.w5(32'hbc612422),
	.w6(32'h3bb3fdb1),
	.w7(32'hbb7c9479),
	.w8(32'hbb7a0f54),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816ff4),
	.w1(32'h3ab4a509),
	.w2(32'hb93abf4e),
	.w3(32'hbb66015f),
	.w4(32'h3b10d904),
	.w5(32'h3b48ac83),
	.w6(32'h39c7d85c),
	.w7(32'h3ae022fd),
	.w8(32'hbb03e32a),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84ad39),
	.w1(32'hbb307453),
	.w2(32'h3b87bd5f),
	.w3(32'hbbea4d89),
	.w4(32'h3be96e6f),
	.w5(32'h3b02fe73),
	.w6(32'hbc07a006),
	.w7(32'hb9f231cf),
	.w8(32'h3b4ef37e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6817e5),
	.w1(32'hbb37a184),
	.w2(32'h3bf83d4e),
	.w3(32'hbb730ce4),
	.w4(32'h3b264921),
	.w5(32'h3c5286e4),
	.w6(32'h3b4f1344),
	.w7(32'hbaf56ca2),
	.w8(32'h3b74e46d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82638b),
	.w1(32'hbba836de),
	.w2(32'hba403f53),
	.w3(32'hbbf0b934),
	.w4(32'hbb84e37c),
	.w5(32'h3a93e284),
	.w6(32'hbb9e11f6),
	.w7(32'hb976113a),
	.w8(32'hbb7b84bc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa23aa0),
	.w1(32'hbb23d48d),
	.w2(32'hbb94730c),
	.w3(32'h3a87cd21),
	.w4(32'hba02d2eb),
	.w5(32'h3ab87979),
	.w6(32'h39e19add),
	.w7(32'h3addd539),
	.w8(32'h3b6f6b3a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17fd3b),
	.w1(32'hbc2274f7),
	.w2(32'hbb9d0e0a),
	.w3(32'hbb81089b),
	.w4(32'hbbde4327),
	.w5(32'h3b00b9a5),
	.w6(32'hbb66f0c8),
	.w7(32'hbb95daf0),
	.w8(32'h3b0054d8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44cc47),
	.w1(32'hb8bfc5fc),
	.w2(32'hbaed229f),
	.w3(32'h3a219517),
	.w4(32'hbadbbf3b),
	.w5(32'hbc3c5447),
	.w6(32'hbbfc6a99),
	.w7(32'hb9f57378),
	.w8(32'hbbc92f71),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55099f),
	.w1(32'hbb1f67ad),
	.w2(32'hba92d23e),
	.w3(32'hbba059c3),
	.w4(32'h3c001838),
	.w5(32'hbb1035c0),
	.w6(32'hbb073a04),
	.w7(32'h3b63c639),
	.w8(32'h3ac3314a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba50b6ef),
	.w1(32'hbb001d09),
	.w2(32'hbbbb4375),
	.w3(32'h3a8a5ab7),
	.w4(32'hbb5ae5b0),
	.w5(32'hbc168356),
	.w6(32'h3b5a5d7e),
	.w7(32'hbb7ab3ed),
	.w8(32'hbbb66019),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ab570),
	.w1(32'h3bc63b12),
	.w2(32'h3b419b7b),
	.w3(32'hba39bb17),
	.w4(32'h3b770482),
	.w5(32'h3bb1e8b7),
	.w6(32'h3ac42600),
	.w7(32'h3a8c8b19),
	.w8(32'h3b8308cf),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57cdab),
	.w1(32'h3c064d73),
	.w2(32'h3bd7d564),
	.w3(32'h3bdd2330),
	.w4(32'h3c2a4576),
	.w5(32'h3aaa1721),
	.w6(32'h3b715fb2),
	.w7(32'h3c0c20a7),
	.w8(32'h3bb722a4),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a27da5),
	.w1(32'hbb544794),
	.w2(32'h3bb6b32f),
	.w3(32'h39c38526),
	.w4(32'hbbf5bcd3),
	.w5(32'h3c5bc500),
	.w6(32'h3bacdbcb),
	.w7(32'hbb8cd35c),
	.w8(32'h3b05bcd2),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ff66c),
	.w1(32'h3ad65e15),
	.w2(32'hbc3f1845),
	.w3(32'hbbdc2327),
	.w4(32'hbaab4a7b),
	.w5(32'hbc702d2f),
	.w6(32'hbadee711),
	.w7(32'h3b0f46e1),
	.w8(32'hbbad2f61),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23b35a),
	.w1(32'h3b3ea10c),
	.w2(32'h3b775e1b),
	.w3(32'hbc436ada),
	.w4(32'h3bef0caa),
	.w5(32'h3c170af3),
	.w6(32'hbbe9cb93),
	.w7(32'h3bac61cb),
	.w8(32'hb9dab939),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda4d4c),
	.w1(32'h3bc9621b),
	.w2(32'h3a82fc16),
	.w3(32'h3bd8a7a4),
	.w4(32'h3b61f6f2),
	.w5(32'h3c3c3bf6),
	.w6(32'hbaf83cd2),
	.w7(32'hba088742),
	.w8(32'h3bd42db5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18dc67),
	.w1(32'hb9987aa1),
	.w2(32'h3a6cc7ef),
	.w3(32'h3ba1cefa),
	.w4(32'hbc12b60a),
	.w5(32'h3b4233b6),
	.w6(32'hba51899f),
	.w7(32'hbc5e0cec),
	.w8(32'hbb5acc72),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c35c1),
	.w1(32'h3b419931),
	.w2(32'h3abc43f6),
	.w3(32'hbbccce73),
	.w4(32'hbbb5e3ec),
	.w5(32'h3b6d953d),
	.w6(32'hbb5c5c08),
	.w7(32'hbb82819a),
	.w8(32'h3a25336a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1adb16),
	.w1(32'hbb839607),
	.w2(32'h3a910d5a),
	.w3(32'h3af31a06),
	.w4(32'hbb8f60fe),
	.w5(32'hbae4db35),
	.w6(32'h3b17b3a1),
	.w7(32'hbb6af681),
	.w8(32'hb98fd6cf),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f8c40),
	.w1(32'h3bc9098b),
	.w2(32'h3c0be3d3),
	.w3(32'hbb22c742),
	.w4(32'h3c21f57c),
	.w5(32'h3c826a63),
	.w6(32'h3b6bdb42),
	.w7(32'h3be34c1c),
	.w8(32'h3c3a407b),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac81df2),
	.w1(32'hbbb20881),
	.w2(32'h3abb1775),
	.w3(32'hb906a487),
	.w4(32'hbbc4e471),
	.w5(32'h3c4c97e8),
	.w6(32'h3b499919),
	.w7(32'hbba01542),
	.w8(32'h3acb4aa3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b12e),
	.w1(32'h3a9a2d49),
	.w2(32'h3c2ba403),
	.w3(32'h3b508ee2),
	.w4(32'h3aa54803),
	.w5(32'hbba740fc),
	.w6(32'h3b93a620),
	.w7(32'hbc09cf33),
	.w8(32'hbb249bf9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2af821),
	.w1(32'h3ba19242),
	.w2(32'h3b8668a3),
	.w3(32'h3c0d2d18),
	.w4(32'h3bf6decb),
	.w5(32'h3aa15905),
	.w6(32'h3a439dc5),
	.w7(32'hbba9e273),
	.w8(32'h3be39581),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3927ec),
	.w1(32'h3ac57c9b),
	.w2(32'h3b7ba8f5),
	.w3(32'h3ba94f1a),
	.w4(32'h3a997111),
	.w5(32'h3b2bc463),
	.w6(32'hbabb7068),
	.w7(32'hb892c892),
	.w8(32'h3b8300b0),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b9592),
	.w1(32'hba9818f1),
	.w2(32'hba34e369),
	.w3(32'h3b5b1c41),
	.w4(32'hbb8f9a75),
	.w5(32'hbb8833ad),
	.w6(32'h3b344aa4),
	.w7(32'h3b2353bb),
	.w8(32'h3c1c32b8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12625a),
	.w1(32'hbbc796c7),
	.w2(32'hbbdc8f8b),
	.w3(32'h3bf315fc),
	.w4(32'hbbf7212d),
	.w5(32'hbbc7ba79),
	.w6(32'h3bac3768),
	.w7(32'hbb82fbb9),
	.w8(32'hbb7ee9d3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1eeb7),
	.w1(32'h3b934e98),
	.w2(32'h39d9b822),
	.w3(32'hbc1163ca),
	.w4(32'h3afee3fa),
	.w5(32'hbb6bf089),
	.w6(32'hbb9cef3b),
	.w7(32'h3be7276e),
	.w8(32'h3b9a0765),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f25a1),
	.w1(32'hbb8e07b3),
	.w2(32'hbba0e944),
	.w3(32'h3b161db5),
	.w4(32'h3a9aaf0f),
	.w5(32'h3c048753),
	.w6(32'h3b8b8ab5),
	.w7(32'hbae4244d),
	.w8(32'h3b8ebb20),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9789a0),
	.w1(32'hbb4d0ea0),
	.w2(32'h3c2c8e3c),
	.w3(32'h394ecc31),
	.w4(32'h3ae2d161),
	.w5(32'h3c6260d3),
	.w6(32'h39a0790c),
	.w7(32'hbb842373),
	.w8(32'hbc53eee5),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b2729),
	.w1(32'h3a220f4f),
	.w2(32'h3959ebbf),
	.w3(32'hbb2d086b),
	.w4(32'hb9e5de18),
	.w5(32'hbb27f082),
	.w6(32'hbc2b860c),
	.w7(32'h3bcd8031),
	.w8(32'h3a4e2f54),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf40330),
	.w1(32'hbc5ce1cd),
	.w2(32'h3a7cad99),
	.w3(32'h3bbfff5a),
	.w4(32'hbcab8718),
	.w5(32'h3b97e180),
	.w6(32'h3ab96c2b),
	.w7(32'hbc30a3d9),
	.w8(32'h3b79a579),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae5de7),
	.w1(32'hbe20e4f1),
	.w2(32'hbf2f43bf),
	.w3(32'hb7dc117c),
	.w4(32'hbf527053),
	.w5(32'hbda28f06),
	.w6(32'hbad6c14f),
	.w7(32'hbeb234f6),
	.w8(32'hbe3d0cce),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbefc5c35),
	.w1(32'hbf226c72),
	.w2(32'hbf6e23e2),
	.w3(32'hbcaebb86),
	.w4(32'hbe8e01d9),
	.w5(32'hbec16356),
	.w6(32'hbe9a9890),
	.w7(32'hbe5433b3),
	.w8(32'hbefa527f),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbed41e86),
	.w1(32'hbf1a917d),
	.w2(32'hbe8e84a8),
	.w3(32'hbe4ae1e3),
	.w4(32'hbe1a2cbb),
	.w5(32'hbe9f9604),
	.w6(32'hbecd6e23),
	.w7(32'hbe61c1cc),
	.w8(32'hbd7f6e00),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe926e11),
	.w1(32'hbe925567),
	.w2(32'hbf1da255),
	.w3(32'hbe4c0e21),
	.w4(32'hbf086bd6),
	.w5(32'hbf1edfa5),
	.w6(32'hbf1a8632),
	.w7(32'hbf26af68),
	.w8(32'hbed8370c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe750c99),
	.w1(32'hbdae1fe6),
	.w2(32'hbdba2001),
	.w3(32'hbe6611d8),
	.w4(32'hbf30ab96),
	.w5(32'hbf12239b),
	.w6(32'hbe69c041),
	.w7(32'hbe7e56eb),
	.w8(32'hbe8b7054),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdb7606a),
	.w1(32'hbe26970c),
	.w2(32'hbda7caa5),
	.w3(32'hbdf59403),
	.w4(32'hbe29dc31),
	.w5(32'hbe7b6953),
	.w6(32'hbebca467),
	.w7(32'hbf066a9f),
	.w8(32'hbe494912),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e4fa2b5),
	.w1(32'hbf5b86ba),
	.w2(32'hbf023046),
	.w3(32'hbee3373d),
	.w4(32'hbf6a0eac),
	.w5(32'hbef1526b),
	.w6(32'hbe6daafe),
	.w7(32'h3d7b358c),
	.w8(32'hbf36370e),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0ae516),
	.w1(32'hbf197905),
	.w2(32'hbed551b6),
	.w3(32'hbed087ec),
	.w4(32'hbf997b7a),
	.w5(32'h3eecfd8f),
	.w6(32'hbdb23b38),
	.w7(32'hbf3913bd),
	.w8(32'hbef1a86c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbed6d06c),
	.w1(32'hbef67dba),
	.w2(32'hbf4282f0),
	.w3(32'h3da87d91),
	.w4(32'hbeb9f8d4),
	.w5(32'hbe79417e),
	.w6(32'hbf175ece),
	.w7(32'hbe43cf70),
	.w8(32'h3dd2998c),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe4ef6ed),
	.w1(32'hbdb27a77),
	.w2(32'hbee3329f),
	.w3(32'hbeca4267),
	.w4(32'hbf2aaea0),
	.w5(32'h3e89f259),
	.w6(32'hbec04fce),
	.w7(32'hbe9d57f9),
	.w8(32'h3db1fed0),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe919d46),
	.w1(32'hbed60881),
	.w2(32'hbd9aa1db),
	.w3(32'hbf24a774),
	.w4(32'h3bf08241),
	.w5(32'hbee5adf6),
	.w6(32'hbf0533c9),
	.w7(32'hbe7170fc),
	.w8(32'hbf243ea3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbec389f9),
	.w1(32'hbf099348),
	.w2(32'hbe60a215),
	.w3(32'hbfa53219),
	.w4(32'hbf19b5a9),
	.w5(32'hbe4ee80b),
	.w6(32'hbe91b65d),
	.w7(32'hbd1b5fcb),
	.w8(32'hbfafa0f1),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe8b8ed2),
	.w1(32'hbf251e60),
	.w2(32'hbe47712f),
	.w3(32'hbeb8df23),
	.w4(32'hbcca3d52),
	.w5(32'hbebbc8e0),
	.w6(32'hbeef8a90),
	.w7(32'hbea7d594),
	.w8(32'hbe2ee6aa),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ecc86c0),
	.w1(32'hbee9d7fe),
	.w2(32'hbe5d6de5),
	.w3(32'hbf7047a0),
	.w4(32'hbe49fccd),
	.w5(32'hbf227f6f),
	.w6(32'hbf387807),
	.w7(32'h3e24a355),
	.w8(32'hbec19af1),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbed8374f),
	.w1(32'hbf05aa2f),
	.w2(32'h3f905963),
	.w3(32'hbea23bcd),
	.w4(32'hbe7036b5),
	.w5(32'h3f52bf25),
	.w6(32'h3ad26077),
	.w7(32'h3f376dfd),
	.w8(32'h3f62552e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f27b2fc),
	.w1(32'h3f39a565),
	.w2(32'h3f52c0d9),
	.w3(32'h3f229257),
	.w4(32'h3f4f5134),
	.w5(32'h3f4310d4),
	.w6(32'h3f3b4acb),
	.w7(32'h3f87145f),
	.w8(32'h3f63271c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4ddb67),
	.w1(32'h3f193f79),
	.w2(32'h3f43be9a),
	.w3(32'h3f575df6),
	.w4(32'h3f49f9e3),
	.w5(32'h3f251c8c),
	.w6(32'h3f4926b3),
	.w7(32'h3f75f693),
	.w8(32'h3f8562ac),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f55c069),
	.w1(32'h3f46523f),
	.w2(32'h3f829dbc),
	.w3(32'h3f2452be),
	.w4(32'h3f86dcdd),
	.w5(32'h3f94a8d0),
	.w6(32'h3f5552cb),
	.w7(32'h3f4c296e),
	.w8(32'h3f7b1ad1),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f63b96d),
	.w1(32'h3f07e610),
	.w2(32'h3f796a88),
	.w3(32'h3f612672),
	.w4(32'h3f6eff11),
	.w5(32'h3f3eb5f3),
	.w6(32'h3f475a7f),
	.w7(32'h3f262912),
	.w8(32'h3f6e6e9c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f824b76),
	.w1(32'h3f6e09ab),
	.w2(32'h3f33d31c),
	.w3(32'h3f2d3e42),
	.w4(32'h3f551484),
	.w5(32'h3f5cd94f),
	.w6(32'h3f1865ca),
	.w7(32'h3f78a71d),
	.w8(32'h3f2ef61c),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f5cad61),
	.w1(32'h3f4fd597),
	.w2(32'h3fac72c3),
	.w3(32'h3f461177),
	.w4(32'h3f418917),
	.w5(32'h3f4d2e10),
	.w6(32'h3f224a5f),
	.w7(32'h3f8d870d),
	.w8(32'h3f6541f5),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f58535e),
	.w1(32'h3f807153),
	.w2(32'h3fa57483),
	.w3(32'h3f6a7c47),
	.w4(32'h3f3d7ea9),
	.w5(32'h3f7f0bf9),
	.w6(32'h3f450281),
	.w7(32'h3f6f85b2),
	.w8(32'h3f5e6325),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f67a77d),
	.w1(32'h3f5b1e79),
	.w2(32'h3f6549ba),
	.w3(32'h3f5b0942),
	.w4(32'h3f84fbe7),
	.w5(32'h3f2b98c5),
	.w6(32'h3f3fc215),
	.w7(32'h3f70e579),
	.w8(32'h3f951a0d),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f580010),
	.w1(32'h3f62e592),
	.w2(32'h3f884ffb),
	.w3(32'h3f5ebe5e),
	.w4(32'h3f2d854a),
	.w5(32'h3f51abba),
	.w6(32'h3f1fa0c5),
	.w7(32'h3f5febc1),
	.w8(32'h3f4e37c0),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4a7f00),
	.w1(32'h3f81ddda),
	.w2(32'h3f2c85ce),
	.w3(32'h3f4aa0af),
	.w4(32'h3f4f2aa1),
	.w5(32'h3f3ee0c3),
	.w6(32'h3f4c02cb),
	.w7(32'h3f849a49),
	.w8(32'h3f27af23),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f6b0168),
	.w1(32'h3f9c7fe0),
	.w2(32'h3f811f23),
	.w3(32'h3f7d9cb1),
	.w4(32'h3f38b152),
	.w5(32'h3f29c973),
	.w6(32'h3f64313d),
	.w7(32'h3f5d73a7),
	.w8(32'h3f2b0101),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f41a2a8),
	.w1(32'h3f7e31f6),
	.w2(32'h3f29eab5),
	.w3(32'h3fabb227),
	.w4(32'h3f6db7da),
	.w5(32'h3f378162),
	.w6(32'h3f3416ec),
	.w7(32'h3f8932f2),
	.w8(32'h3f415ff4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f544992),
	.w1(32'h3fa696f8),
	.w2(32'h3f427452),
	.w3(32'h3f45d2e8),
	.w4(32'h3f68115d),
	.w5(32'h3f35f98c),
	.w6(32'h3f2c467f),
	.w7(32'h3f6cb461),
	.w8(32'h3f420450),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f73a800),
	.w1(32'h3f5a1e16),
	.w2(32'h3f59f719),
	.w3(32'h3f4b423b),
	.w4(32'h3f37d07b),
	.w5(32'hbe0317c0),
	.w6(32'h3f5e433b),
	.w7(32'h3f5b2909),
	.w8(32'hbe5a7617),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5a6c5c),
	.w1(32'hbc828361),
	.w2(32'hbd50c3af),
	.w3(32'hbd6c2a7a),
	.w4(32'hbdb9300a),
	.w5(32'hbd49279e),
	.w6(32'hbd75bb87),
	.w7(32'h3c055fd2),
	.w8(32'hbe8998fe),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeac70d5),
	.w1(32'h3ee24b9b),
	.w2(32'hbe207bd1),
	.w3(32'h3e16eae4),
	.w4(32'hbe119581),
	.w5(32'hbe53c6fd),
	.w6(32'h3e1de482),
	.w7(32'h3b6f1b9b),
	.w8(32'hbda5ffb7),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd93671a),
	.w1(32'h3d190424),
	.w2(32'hbe6e16a1),
	.w3(32'h3eb1aa4a),
	.w4(32'hbdc645f6),
	.w5(32'hbe3bcda9),
	.w6(32'h3d7f0ab4),
	.w7(32'hbcd6d6ff),
	.w8(32'hbdc326a9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe570c23),
	.w1(32'hbd435ca7),
	.w2(32'hbee0c59b),
	.w3(32'hbd0334a3),
	.w4(32'hbe471bdf),
	.w5(32'h3dad0717),
	.w6(32'hbd01e906),
	.w7(32'hbe2abfd7),
	.w8(32'hbe5779d9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe0e604c),
	.w1(32'hbe4921e0),
	.w2(32'h3b926edc),
	.w3(32'hbd2073bd),
	.w4(32'hbd9fa110),
	.w5(32'h3da67d52),
	.w6(32'hbd4988ae),
	.w7(32'h3c7adffa),
	.w8(32'hbce3eb60),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e080c5e),
	.w1(32'h3c2535a4),
	.w2(32'hbe02b67b),
	.w3(32'hbe2f8095),
	.w4(32'hbcf5cf69),
	.w5(32'hbdd71d15),
	.w6(32'hbe940b9b),
	.w7(32'hbea36c50),
	.w8(32'hbe688f3a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe64e002),
	.w1(32'h3de4f4ea),
	.w2(32'hbd9f1275),
	.w3(32'h3df10482),
	.w4(32'h3db09233),
	.w5(32'hbe0ffaa5),
	.w6(32'h3d9ffbee),
	.w7(32'hbe221f43),
	.w8(32'h3d1ee433),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9715f2),
	.w1(32'hbea6c05e),
	.w2(32'hbdb0d57b),
	.w3(32'h3e26d03c),
	.w4(32'hbd0a313c),
	.w5(32'hbcc0d07a),
	.w6(32'hbedffd11),
	.w7(32'hbe27ca34),
	.w8(32'hbd8d0090),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbc9e17),
	.w1(32'hbe40bce7),
	.w2(32'h3e5f943b),
	.w3(32'hbeafc029),
	.w4(32'hbd7b8357),
	.w5(32'h3e478f1a),
	.w6(32'h3d6a0923),
	.w7(32'hbe90d6d6),
	.w8(32'hbe12a262),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57c53b),
	.w1(32'hbdaf78e4),
	.w2(32'hba69cbfb),
	.w3(32'h3e422fe5),
	.w4(32'h3d359143),
	.w5(32'h3d47ceed),
	.w6(32'h3d9f22dc),
	.w7(32'hbdf4afdf),
	.w8(32'hbdd739a1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe3911be),
	.w1(32'hbe55c954),
	.w2(32'hbd98f045),
	.w3(32'hbe496ffc),
	.w4(32'hbe867fea),
	.w5(32'hbcd7c87b),
	.w6(32'hbd173841),
	.w7(32'hbd83bd00),
	.w8(32'hbe92e06e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1f13b9),
	.w1(32'h3d37b218),
	.w2(32'hbe8d0f1d),
	.w3(32'hbe6f6393),
	.w4(32'hbe636923),
	.w5(32'hbda35894),
	.w6(32'h3e03602a),
	.w7(32'hbd96d43c),
	.w8(32'h3c948253),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e293997),
	.w1(32'hbe076194),
	.w2(32'h3e19a6ff),
	.w3(32'h3db3eefe),
	.w4(32'hbd22213f),
	.w5(32'hbe1153e3),
	.w6(32'h3e2f2024),
	.w7(32'hbe927c07),
	.w8(32'hbd258ca3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9e55f5),
	.w1(32'h3d87640e),
	.w2(32'h3c288aee),
	.w3(32'hbd427481),
	.w4(32'hbb709eaa),
	.w5(32'hbbf263a5),
	.w6(32'hbd5493ee),
	.w7(32'hbd777def),
	.w8(32'hbe69001d),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca859ea),
	.w1(32'h3c9e5d7f),
	.w2(32'h3c974207),
	.w3(32'h3cffcf6e),
	.w4(32'h3cb15598),
	.w5(32'h3cfda8bb),
	.w6(32'h3c9d759c),
	.w7(32'h3c80a9b3),
	.w8(32'h3ccf730b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd4a3bd),
	.w1(32'h3cac2b74),
	.w2(32'h3c903016),
	.w3(32'h3cd89e02),
	.w4(32'h3c9e074e),
	.w5(32'h3c77605c),
	.w6(32'h3d1cebde),
	.w7(32'h3cd78d54),
	.w8(32'h3cbff825),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc1edc3),
	.w1(32'h3d0bec76),
	.w2(32'h3ced39a0),
	.w3(32'h3cd62495),
	.w4(32'h3cd4c9b6),
	.w5(32'h3cc628dc),
	.w6(32'h3c873bd6),
	.w7(32'h3c98d0db),
	.w8(32'h3d02c1f9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb2353b),
	.w1(32'h3cda0bb6),
	.w2(32'h3cb3fe71),
	.w3(32'h3d0f53ea),
	.w4(32'h3c9bdcef),
	.w5(32'h3c1fafff),
	.w6(32'h3d5b6dba),
	.w7(32'h3cd5dadd),
	.w8(32'h3d66dc96),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc72bc2),
	.w1(32'h3d2e0e06),
	.w2(32'h3c71c0eb),
	.w3(32'h3cc7fe47),
	.w4(32'h3d09db7c),
	.w5(32'h3d1896d3),
	.w6(32'h3ccfaf1c),
	.w7(32'h3ca4bd3d),
	.w8(32'h3caf5112),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d5cc165),
	.w1(32'h3cf6d382),
	.w2(32'h3d19e45b),
	.w3(32'h3cccc173),
	.w4(32'h3ce1fc89),
	.w5(32'h3cae1152),
	.w6(32'h3cb5fd66),
	.w7(32'h3d0da8d9),
	.w8(32'h3cbc7c53),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccfde35),
	.w1(32'h3c9da1cf),
	.w2(32'h3d3d8ac3),
	.w3(32'h3d188116),
	.w4(32'h3cbf76ed),
	.w5(32'h3d66a357),
	.w6(32'h3d054ec2),
	.w7(32'h3ca7f69e),
	.w8(32'h3d2c4995),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd8b9f9),
	.w1(32'h3ca531e9),
	.w2(32'h3caf4945),
	.w3(32'h3d160f4c),
	.w4(32'h3d4601f7),
	.w5(32'h3d1af200),
	.w6(32'h3cde2804),
	.w7(32'h3cbe1561),
	.w8(32'h3d21152a),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce532a5),
	.w1(32'h3d05cc16),
	.w2(32'h3c8d4c9a),
	.w3(32'h3d072d4c),
	.w4(32'h3cde4e52),
	.w5(32'h3cf471fa),
	.w6(32'h3c7243b9),
	.w7(32'h3d42d586),
	.w8(32'h3c85ff3f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d225699),
	.w1(32'h3c9dfe09),
	.w2(32'h3d19f41e),
	.w3(32'h3d0d70dd),
	.w4(32'h3d53ddd0),
	.w5(32'h3cedfa34),
	.w6(32'h3cd86489),
	.w7(32'h3d2301ad),
	.w8(32'h3cb3dd76),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d352b52),
	.w1(32'h3cb471c1),
	.w2(32'h3d316802),
	.w3(32'h3c9fe720),
	.w4(32'h3c931e60),
	.w5(32'h3d15efc6),
	.w6(32'h3ca9a0a1),
	.w7(32'h3d04df98),
	.w8(32'h3cb3437f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd70f1a),
	.w1(32'h3c750b52),
	.w2(32'h3ca18c26),
	.w3(32'h3d12b398),
	.w4(32'h3cc25950),
	.w5(32'h3d1ee640),
	.w6(32'h3cd94d06),
	.w7(32'h3d0df771),
	.w8(32'h3ce938f4),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d057a47),
	.w1(32'h3ca9b7ff),
	.w2(32'h3d1d382a),
	.w3(32'h3cb9debb),
	.w4(32'h3d1c4310),
	.w5(32'h3d234a6f),
	.w6(32'h3c70f343),
	.w7(32'h3cb80afd),
	.w8(32'h3cbab7dd),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d00dc3b),
	.w1(32'h3cf611ef),
	.w2(32'h3cd7ee89),
	.w3(32'h3cda97c5),
	.w4(32'h3cbc5e04),
	.w5(32'h3cf4e455),
	.w6(32'h3d10e4be),
	.w7(32'h3cb779dc),
	.w8(32'h3cfde8b7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c966596),
	.w1(32'h3ca1e7e1),
	.w2(32'hbc0a2363),
	.w3(32'h3d26700b),
	.w4(32'hbce01d50),
	.w5(32'hbc55430e),
	.w6(32'hbc52f97c),
	.w7(32'hbba4dbfd),
	.w8(32'h3aab1571),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01a628),
	.w1(32'hbc2b1651),
	.w2(32'hbaa3dafa),
	.w3(32'h3bf6edc7),
	.w4(32'hbb809b3c),
	.w5(32'hb9de044b),
	.w6(32'hbb879a42),
	.w7(32'hbcb2512e),
	.w8(32'hbcae3867),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule