module layer_10_featuremap_402(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28ee2c),
	.w1(32'hb8940ace),
	.w2(32'h39acdaf6),
	.w3(32'hb8bf7972),
	.w4(32'h3c057655),
	.w5(32'h3c3bc9d7),
	.w6(32'h3b9a8526),
	.w7(32'hbba9f28a),
	.w8(32'hbab9477f),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0d823),
	.w1(32'h3ae80a0e),
	.w2(32'hba3316ce),
	.w3(32'h3b8f8330),
	.w4(32'hbae473ac),
	.w5(32'hb908a01a),
	.w6(32'hbbc598b1),
	.w7(32'hba4923b7),
	.w8(32'h3984e3aa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ea8b),
	.w1(32'h3b93fa00),
	.w2(32'hb9f09f61),
	.w3(32'hbbaff84a),
	.w4(32'hba9ad7b5),
	.w5(32'h3adb3be2),
	.w6(32'hbb13c657),
	.w7(32'h3ae8ab36),
	.w8(32'hbb6ddd91),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b77e2),
	.w1(32'h3bef172f),
	.w2(32'hbb16b10d),
	.w3(32'h3a9e0899),
	.w4(32'h3caf6b8f),
	.w5(32'hbb2360bc),
	.w6(32'hbb6adc8a),
	.w7(32'h3b8d2a3f),
	.w8(32'hbb1ff0dc),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96f17c),
	.w1(32'h3b27e6fe),
	.w2(32'hbae1430f),
	.w3(32'h3aa92622),
	.w4(32'h3b652005),
	.w5(32'hbb6b8765),
	.w6(32'h3b005c89),
	.w7(32'hb90b837d),
	.w8(32'hbb1ff82b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302b97),
	.w1(32'h3c2f962b),
	.w2(32'hba8e7d40),
	.w3(32'hb988a20f),
	.w4(32'hbaf729de),
	.w5(32'h3b808644),
	.w6(32'hba58015f),
	.w7(32'h3ada5930),
	.w8(32'h397bf521),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf291e5),
	.w1(32'h3adb4548),
	.w2(32'h37fa09f5),
	.w3(32'hbb81b006),
	.w4(32'h3bb9f6b4),
	.w5(32'h3b87dde8),
	.w6(32'hbab16718),
	.w7(32'h3b991941),
	.w8(32'h3909ba77),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b412243),
	.w1(32'hbb96d976),
	.w2(32'hbbceb9c6),
	.w3(32'h3c5a511e),
	.w4(32'hbafa302f),
	.w5(32'h3c28d319),
	.w6(32'h3bbc223c),
	.w7(32'hbaeef35b),
	.w8(32'hbb7cc991),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9b42f),
	.w1(32'h3b3b7cd0),
	.w2(32'h3bb223e3),
	.w3(32'h3b02e4d8),
	.w4(32'h3c08568b),
	.w5(32'h3c2557d3),
	.w6(32'hbb179e54),
	.w7(32'h3af3aeba),
	.w8(32'h3b909bf8),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab20bc),
	.w1(32'h3bb1e1f3),
	.w2(32'hba8d5635),
	.w3(32'h3c3fd5f6),
	.w4(32'h3b3e6cb7),
	.w5(32'hbb0671bf),
	.w6(32'h3b8393e6),
	.w7(32'hbb1462c7),
	.w8(32'h3b0c151f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fb79b),
	.w1(32'h3bba5c11),
	.w2(32'h3adc83e1),
	.w3(32'h3b7ff640),
	.w4(32'h3a378adb),
	.w5(32'hbbaecfa9),
	.w6(32'h3b4bf848),
	.w7(32'h3b8deb2b),
	.w8(32'h3a772a92),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff43ad),
	.w1(32'hbb5a5c0c),
	.w2(32'h39a8dbe9),
	.w3(32'hbbb5b9f0),
	.w4(32'hbc3a9da1),
	.w5(32'hbc5c358f),
	.w6(32'hb8af297e),
	.w7(32'hbba8dd96),
	.w8(32'hbb48ee15),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fdb53),
	.w1(32'hbaaffb09),
	.w2(32'hbbac6b74),
	.w3(32'hbc0625bd),
	.w4(32'hbc1b25ee),
	.w5(32'hbba7f824),
	.w6(32'hbac09cd5),
	.w7(32'hbbbb4ea0),
	.w8(32'h3b6ba94c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4429bc),
	.w1(32'hbb78c384),
	.w2(32'hbb656b93),
	.w3(32'hbc52da60),
	.w4(32'h3b15c2c6),
	.w5(32'hbb959c1f),
	.w6(32'hbc1e59b4),
	.w7(32'hba545036),
	.w8(32'hbbd914be),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925025f),
	.w1(32'hbbbbce8a),
	.w2(32'h3b02a5e9),
	.w3(32'h3b8209d4),
	.w4(32'hbc112aad),
	.w5(32'hbbb82ce9),
	.w6(32'h3b1fd564),
	.w7(32'hbb241959),
	.w8(32'hbad8b0bc),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac21b68),
	.w1(32'hbb994fc8),
	.w2(32'h3bdb70bb),
	.w3(32'hbbbc9179),
	.w4(32'hbba3526b),
	.w5(32'h3bb5b510),
	.w6(32'hbb096b2e),
	.w7(32'hbabaa73b),
	.w8(32'h3b908b71),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cfadb),
	.w1(32'hbb82c271),
	.w2(32'h3b6ef33d),
	.w3(32'hbbbeaea3),
	.w4(32'hbb6eabc1),
	.w5(32'hbba15159),
	.w6(32'h39377cd0),
	.w7(32'h3b84e39c),
	.w8(32'h3b3a0e52),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f27d0),
	.w1(32'h3920eb8f),
	.w2(32'hba3afd89),
	.w3(32'h3b07f244),
	.w4(32'h3ca29c87),
	.w5(32'h3c8938c2),
	.w6(32'h3a5b0fd7),
	.w7(32'h39c22679),
	.w8(32'hbb5ce7f1),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ba962),
	.w1(32'hbb8da374),
	.w2(32'hbb03a9c4),
	.w3(32'h3c3a2df3),
	.w4(32'hbbe749ed),
	.w5(32'hbc006bb8),
	.w6(32'hba4a24aa),
	.w7(32'hbbeb389d),
	.w8(32'hbb86b377),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16e780),
	.w1(32'h3a87c2ba),
	.w2(32'hbb7d7023),
	.w3(32'hbc51fa3b),
	.w4(32'h3bdd71d4),
	.w5(32'hbc1125ba),
	.w6(32'hbc0eec82),
	.w7(32'h3bb2679b),
	.w8(32'hbba6b53f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb628c60),
	.w1(32'hbb670d5c),
	.w2(32'hbb5c7930),
	.w3(32'hbc0d863e),
	.w4(32'hbc50f354),
	.w5(32'hbc213238),
	.w6(32'hbc1aa60f),
	.w7(32'hbad8e222),
	.w8(32'hbb8134a3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb371e4c),
	.w1(32'hbb8803d9),
	.w2(32'h3ba62b03),
	.w3(32'hbba4ffe7),
	.w4(32'hbbd64fa0),
	.w5(32'h3ae3a645),
	.w6(32'hbb1201ff),
	.w7(32'hbb8ab21e),
	.w8(32'h3b61b705),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79e37c),
	.w1(32'h3c2d71ad),
	.w2(32'h3c5fc447),
	.w3(32'h3bcf68fd),
	.w4(32'h3b947f87),
	.w5(32'hbb95ea3b),
	.w6(32'h3b8123ad),
	.w7(32'h39c4f9c1),
	.w8(32'hba55fcc8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eb253),
	.w1(32'h3c180bf5),
	.w2(32'hbc0b4f45),
	.w3(32'h3a27f88e),
	.w4(32'h3c51130b),
	.w5(32'hbb3719cf),
	.w6(32'hbb564cc5),
	.w7(32'h3b32ea4b),
	.w8(32'hbc201666),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba045a5a),
	.w1(32'h3b4bebfb),
	.w2(32'h3aa696f9),
	.w3(32'h3b60dafb),
	.w4(32'hbba204e8),
	.w5(32'hbc7635db),
	.w6(32'hbb73af32),
	.w7(32'hbbefe80b),
	.w8(32'hbbf612fa),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38270e77),
	.w1(32'hba3564ab),
	.w2(32'h3b4409de),
	.w3(32'h3c567673),
	.w4(32'h3a96ac66),
	.w5(32'h3ac54683),
	.w6(32'h3c08e1d8),
	.w7(32'h3b257ba1),
	.w8(32'h3aed7b8c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf76b48),
	.w1(32'hbbba37f6),
	.w2(32'hbba0cb11),
	.w3(32'h3ab252f1),
	.w4(32'hbbf04133),
	.w5(32'hbb8201eb),
	.w6(32'hb998a251),
	.w7(32'hbb546208),
	.w8(32'hbb270d0b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65629d),
	.w1(32'h3b21e944),
	.w2(32'h3b646136),
	.w3(32'hbc465187),
	.w4(32'h3b305442),
	.w5(32'h3bd72bce),
	.w6(32'hbc0cd7f5),
	.w7(32'hb5425840),
	.w8(32'h3ae3f19d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99cecb2),
	.w1(32'hbc046a39),
	.w2(32'hbb7f9366),
	.w3(32'hb9376f7c),
	.w4(32'hbbaf722f),
	.w5(32'hbbde07f5),
	.w6(32'hba75aea6),
	.w7(32'h3ba3f0bf),
	.w8(32'h3ba39aae),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26d60),
	.w1(32'hbc1f6ab8),
	.w2(32'hbbc26547),
	.w3(32'hbbcf32be),
	.w4(32'hbca93fa4),
	.w5(32'hbc8393d6),
	.w6(32'hbb1481d8),
	.w7(32'hbc2df9ae),
	.w8(32'hba97e04d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc99342),
	.w1(32'h3b839a15),
	.w2(32'h3c0ffa34),
	.w3(32'hbc8d4ef7),
	.w4(32'h3c2490a7),
	.w5(32'h3c38fdc6),
	.w6(32'hbbdef36c),
	.w7(32'h3bfe8c62),
	.w8(32'h3b89961e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09a5a5),
	.w1(32'h3ade1e5e),
	.w2(32'hbba34523),
	.w3(32'h3ba9d99f),
	.w4(32'hbb255257),
	.w5(32'hbb7f8928),
	.w6(32'h3a856a9d),
	.w7(32'hbabb508f),
	.w8(32'hbb8fc93b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66dab6),
	.w1(32'hbaa30a06),
	.w2(32'hbb8a96ac),
	.w3(32'hbbad7a6b),
	.w4(32'hbb1eaa53),
	.w5(32'hbb72bc8c),
	.w6(32'hbbdf939f),
	.w7(32'hbb71012e),
	.w8(32'hbbe61948),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3a246),
	.w1(32'hbb085f97),
	.w2(32'hba48509d),
	.w3(32'hbb4d435b),
	.w4(32'hba03cf34),
	.w5(32'h3b0ac047),
	.w6(32'hbba670a4),
	.w7(32'hbb2ebc3f),
	.w8(32'hbaf5faba),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6d8ee),
	.w1(32'hbaaca4ca),
	.w2(32'hbb233e67),
	.w3(32'h3b7618e6),
	.w4(32'h3beb0211),
	.w5(32'h3c1ea427),
	.w6(32'h3b8b0565),
	.w7(32'hb9a33bda),
	.w8(32'hbb8ddf99),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ee1fa),
	.w1(32'h3bc6a49e),
	.w2(32'h3c40b129),
	.w3(32'h3b61a334),
	.w4(32'h3c6043df),
	.w5(32'h3c78efce),
	.w6(32'hba1c56ec),
	.w7(32'h3bcdc0c8),
	.w8(32'h3c22de13),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f613b),
	.w1(32'h3bac4d59),
	.w2(32'hbb6e86f0),
	.w3(32'h3c93890a),
	.w4(32'h3bc15dee),
	.w5(32'hbc0d3d95),
	.w6(32'h3c84f8c7),
	.w7(32'h3b02ece1),
	.w8(32'hbbe43c49),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae5075),
	.w1(32'hbae89eb4),
	.w2(32'hbaffe510),
	.w3(32'hbc667ae6),
	.w4(32'hbbf4eb90),
	.w5(32'hbb85e8ec),
	.w6(32'hbc1ab1eb),
	.w7(32'hbb7185d6),
	.w8(32'hbac46da0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00249b),
	.w1(32'hbbb292e4),
	.w2(32'h3a039d32),
	.w3(32'hbc3fca9d),
	.w4(32'h3b73d502),
	.w5(32'h3c0c2008),
	.w6(32'hbb4ca1ae),
	.w7(32'hbb4bfd18),
	.w8(32'h39c52fcc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d9fc8),
	.w1(32'h3a9b2def),
	.w2(32'hba498f65),
	.w3(32'h3c864767),
	.w4(32'h3bec6fdb),
	.w5(32'h3bc5e45b),
	.w6(32'h3b1672fc),
	.w7(32'h3bd2d222),
	.w8(32'h3bbb0738),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8060d),
	.w1(32'h3ad96aa6),
	.w2(32'hbb0f060b),
	.w3(32'h3b57e135),
	.w4(32'h3c260dff),
	.w5(32'hbb89ce58),
	.w6(32'hba98aa47),
	.w7(32'h3b68543e),
	.w8(32'hbb227a54),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73c1cb),
	.w1(32'hbb49844e),
	.w2(32'h3b8bdb4a),
	.w3(32'h3adf89d3),
	.w4(32'hbbe669f6),
	.w5(32'h3bb5e636),
	.w6(32'h3ad277df),
	.w7(32'hba363351),
	.w8(32'h3b702bc0),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb152f9c),
	.w1(32'hbb2aa84c),
	.w2(32'hbbd68450),
	.w3(32'hbc0b0da1),
	.w4(32'hbb348c91),
	.w5(32'hbb1b4baa),
	.w6(32'hbb145c55),
	.w7(32'hbb8e74a8),
	.w8(32'h3ace6600),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b994b11),
	.w1(32'hbc49a95c),
	.w2(32'hbc77c747),
	.w3(32'h3c06ede8),
	.w4(32'h3b8b5651),
	.w5(32'hbb61aff3),
	.w6(32'h3b93bd07),
	.w7(32'hbc2f6413),
	.w8(32'hbc59f8aa),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc321b72),
	.w1(32'hbb29288e),
	.w2(32'hba82ca77),
	.w3(32'hba8e26af),
	.w4(32'hbbe04f0c),
	.w5(32'hbab1b159),
	.w6(32'hbc750700),
	.w7(32'hbb3d902e),
	.w8(32'hba382c67),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad74219),
	.w1(32'h3ae04e39),
	.w2(32'h3bee78b1),
	.w3(32'h37681a5d),
	.w4(32'hbb0a88b3),
	.w5(32'h3bdb789e),
	.w6(32'hbb2b8f94),
	.w7(32'h3a98eb61),
	.w8(32'h3ba220cf),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a19e),
	.w1(32'hbb4d0251),
	.w2(32'hbb8bf1a9),
	.w3(32'hbb4b5864),
	.w4(32'hbb49f974),
	.w5(32'hbb57aa6b),
	.w6(32'h3b83c0c3),
	.w7(32'h3b853d4a),
	.w8(32'h3b0e65a2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce584e),
	.w1(32'hbc064bc5),
	.w2(32'hbc1f480d),
	.w3(32'h3ba4842f),
	.w4(32'h3bab8317),
	.w5(32'hbbae1088),
	.w6(32'h38c958a9),
	.w7(32'hbbb3b5bb),
	.w8(32'hbc27d148),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23fc1a),
	.w1(32'hb9cffbb6),
	.w2(32'h3bad263c),
	.w3(32'hbbf5c029),
	.w4(32'hb9c049df),
	.w5(32'h3c026f68),
	.w6(32'hbbf824e3),
	.w7(32'h3baec6fd),
	.w8(32'h3c071316),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be53a1d),
	.w1(32'h3b9a39c9),
	.w2(32'h3c70a315),
	.w3(32'h3c7db394),
	.w4(32'hbb4f4391),
	.w5(32'h3ca33e6e),
	.w6(32'h3c702d93),
	.w7(32'hba9b072a),
	.w8(32'h3c4583b1),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f136d),
	.w1(32'h3aa1004e),
	.w2(32'h3acf274f),
	.w3(32'h3cb0ec7d),
	.w4(32'h3ab38ee2),
	.w5(32'hba76db03),
	.w6(32'h3c8366b2),
	.w7(32'h3ac6a2b9),
	.w8(32'h3a0dcc84),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6f61a),
	.w1(32'hbb6899ae),
	.w2(32'hbbfd8a2a),
	.w3(32'h3aa6fd88),
	.w4(32'h3a7dbaaa),
	.w5(32'hbbc6b859),
	.w6(32'h3aff91c5),
	.w7(32'hbbd1ee3b),
	.w8(32'hbc00a976),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cd4bd),
	.w1(32'h3b92cc82),
	.w2(32'h3ba57666),
	.w3(32'h3a40e596),
	.w4(32'hba89554c),
	.w5(32'h3c680fcc),
	.w6(32'hba25b57f),
	.w7(32'hba8516b0),
	.w8(32'h3bc1e170),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c04fb),
	.w1(32'h3bb1b23f),
	.w2(32'hba52889c),
	.w3(32'h3c59c54d),
	.w4(32'h3bc0b662),
	.w5(32'h3aecfc9b),
	.w6(32'h3c2c6a8e),
	.w7(32'h3a8de233),
	.w8(32'hbbcd1cb8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5ae2d),
	.w1(32'hbb6608ba),
	.w2(32'hb9c8b73d),
	.w3(32'hba6a82d9),
	.w4(32'hbc0f8a7e),
	.w5(32'hbb05c2a1),
	.w6(32'hb9a42110),
	.w7(32'h39b085ae),
	.w8(32'h3b169784),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4d56d),
	.w1(32'hbbc6b3b9),
	.w2(32'hbb1527dc),
	.w3(32'hba3a4837),
	.w4(32'hbbd6c1e3),
	.w5(32'h3acfe3fa),
	.w6(32'h3ada5d4b),
	.w7(32'hbc054d0a),
	.w8(32'hb990ecdf),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eac08),
	.w1(32'hbb3be6ea),
	.w2(32'hbbe55d5c),
	.w3(32'hba0c9fd5),
	.w4(32'hbbb3a997),
	.w5(32'hbc8c56fd),
	.w6(32'hbbb3e646),
	.w7(32'hbb87e2fe),
	.w8(32'hbbbc72bb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e7b8f),
	.w1(32'h3adc89fa),
	.w2(32'h3bcfa353),
	.w3(32'hbbd80a8e),
	.w4(32'hb851cd14),
	.w5(32'h3b63c38a),
	.w6(32'hbb44aaaf),
	.w7(32'hbab41f8c),
	.w8(32'h3b528603),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd2fff),
	.w1(32'hbbcf29c7),
	.w2(32'hbc22a05d),
	.w3(32'hbb9b9a6d),
	.w4(32'hbbb287c6),
	.w5(32'hbc27fc6d),
	.w6(32'hbb962cf7),
	.w7(32'hbc0e9052),
	.w8(32'hbc14b3fe),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44aea),
	.w1(32'h3b7274c2),
	.w2(32'h3adcd1dc),
	.w3(32'hbc018086),
	.w4(32'hbb6be18e),
	.w5(32'hbbab95b6),
	.w6(32'hbc247f40),
	.w7(32'hb9f02121),
	.w8(32'h3bef4c97),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b0680),
	.w1(32'hbb8f7a89),
	.w2(32'hbba23b47),
	.w3(32'hb9b8a73d),
	.w4(32'hbb403899),
	.w5(32'h39e4ba24),
	.w6(32'h3c13c19d),
	.w7(32'hba2e5c2e),
	.w8(32'h3b143e0c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d325e),
	.w1(32'hbb481c5e),
	.w2(32'hbb4d570f),
	.w3(32'h3bd11dc2),
	.w4(32'hbb0a64a7),
	.w5(32'hbb9211c6),
	.w6(32'h3c11a775),
	.w7(32'hbb57f3b3),
	.w8(32'hbb62bf7f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15203d),
	.w1(32'h3ba9e8b3),
	.w2(32'hbb9d9351),
	.w3(32'hbaac2389),
	.w4(32'h3c75a861),
	.w5(32'hbb81993d),
	.w6(32'hb93db817),
	.w7(32'h37583f1e),
	.w8(32'hbb64fc5a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1141d),
	.w1(32'hbac208c0),
	.w2(32'hbb078e22),
	.w3(32'h3c25d614),
	.w4(32'hbc11bafe),
	.w5(32'hbc1e6681),
	.w6(32'h3b768471),
	.w7(32'hbbc1ab2d),
	.w8(32'hbb86d05f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388498dc),
	.w1(32'hbba71ea9),
	.w2(32'hbbde234a),
	.w3(32'hbb9e80e4),
	.w4(32'hbaa6102a),
	.w5(32'hba88ac38),
	.w6(32'hbb604939),
	.w7(32'hbbb1fbf7),
	.w8(32'hbb9e70a0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab358d3),
	.w1(32'hba3ada2a),
	.w2(32'h3b888009),
	.w3(32'h3b825573),
	.w4(32'h3bedfb55),
	.w5(32'h3c5ce9c6),
	.w6(32'h38c46e45),
	.w7(32'h3b8eb093),
	.w8(32'h3a87abb6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb68237),
	.w1(32'h3ba5bfe1),
	.w2(32'h3b22f7d3),
	.w3(32'h3c3f2e82),
	.w4(32'h3b5a25fe),
	.w5(32'hb971d7f3),
	.w6(32'h3c17d2e2),
	.w7(32'h3bfc3f0d),
	.w8(32'h3a84fc07),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb337c39),
	.w1(32'hbbe329ef),
	.w2(32'hbbdaa2ac),
	.w3(32'hbb1d92dc),
	.w4(32'h3a3bce8a),
	.w5(32'h3c2f12b7),
	.w6(32'hbb1598e5),
	.w7(32'hbb6480ae),
	.w8(32'h3b6dd2fd),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf2a2a),
	.w1(32'hbb87c4cc),
	.w2(32'hbbe0c9ea),
	.w3(32'h3c43d8d9),
	.w4(32'h38896e41),
	.w5(32'hbbb70825),
	.w6(32'h3bbc6200),
	.w7(32'hbba37cf9),
	.w8(32'hbb749b9a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0702c),
	.w1(32'hbbeffdd2),
	.w2(32'h3c60faa5),
	.w3(32'hbb78edf6),
	.w4(32'hbb7461ef),
	.w5(32'h3c670a4a),
	.w6(32'hbc0fd02a),
	.w7(32'h3b1738f2),
	.w8(32'h3c1cfc66),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7f144),
	.w1(32'hbb299efc),
	.w2(32'hbc2e9884),
	.w3(32'h39c04674),
	.w4(32'h3aa4b0f1),
	.w5(32'hbc0ac8d9),
	.w6(32'hbbd49469),
	.w7(32'h3a346ce5),
	.w8(32'hbba2e7d2),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc102944),
	.w1(32'h39d1962b),
	.w2(32'hbbcbbac3),
	.w3(32'hbb8cb3d3),
	.w4(32'h3ba08058),
	.w5(32'hbb8a53ed),
	.w6(32'hbc04e365),
	.w7(32'hbb53d865),
	.w8(32'hbc29ed1b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e5e72),
	.w1(32'h3c2084cf),
	.w2(32'h3c3dc9c5),
	.w3(32'hbc4f7fea),
	.w4(32'h3c2fbb3d),
	.w5(32'h3cba7a28),
	.w6(32'hbc04894f),
	.w7(32'h3b896895),
	.w8(32'h3c40fb45),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfb75c3),
	.w1(32'hbb988a6a),
	.w2(32'h39afeb9e),
	.w3(32'hbb4443b4),
	.w4(32'h3a5fe8e6),
	.w5(32'hbbe264d3),
	.w6(32'hba433723),
	.w7(32'hb8b1039a),
	.w8(32'h3b41c876),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69e1a2),
	.w1(32'hbaed8f00),
	.w2(32'hbac2f491),
	.w3(32'h3b778b90),
	.w4(32'h3b9117e1),
	.w5(32'h3b9698fd),
	.w6(32'h3b665685),
	.w7(32'hbb78f1f6),
	.w8(32'hbbc36e84),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa3c8e),
	.w1(32'h3a242360),
	.w2(32'hbb738905),
	.w3(32'h3b246b62),
	.w4(32'hba51d60d),
	.w5(32'h399d8676),
	.w6(32'h3a8740b5),
	.w7(32'hba2b4ff4),
	.w8(32'h3b450a5f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fee05),
	.w1(32'h3bd7504a),
	.w2(32'hbbbfd8b5),
	.w3(32'h3b80016c),
	.w4(32'h3c000182),
	.w5(32'hbb868d7e),
	.w6(32'h3c1be28f),
	.w7(32'h3b18a18b),
	.w8(32'hbb1161d7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff016c),
	.w1(32'h3bbad012),
	.w2(32'hbc0838a4),
	.w3(32'hbc639d2b),
	.w4(32'h3bc8b33b),
	.w5(32'h3b1262b6),
	.w6(32'hbbb118a5),
	.w7(32'h3bf5e7c4),
	.w8(32'h3affce7e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00a90),
	.w1(32'hbbdb2eda),
	.w2(32'hbc281877),
	.w3(32'h3b38b47d),
	.w4(32'hbb0f4b9e),
	.w5(32'h3aaada21),
	.w6(32'h3b8bd72f),
	.w7(32'hba4a9857),
	.w8(32'hb83cf5cc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cdd06),
	.w1(32'h3b525da2),
	.w2(32'hbbb0398f),
	.w3(32'hbae7c335),
	.w4(32'h3c364efc),
	.w5(32'h3c7a9a22),
	.w6(32'h3b5d7cc4),
	.w7(32'h3b89f8c4),
	.w8(32'h3c5f882f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb31afd),
	.w1(32'h3c0ff3f0),
	.w2(32'h3b3d6190),
	.w3(32'hbc097bba),
	.w4(32'h3aa41714),
	.w5(32'hbc5cd995),
	.w6(32'hb7a4a748),
	.w7(32'h3a82706f),
	.w8(32'hbaa9e5fd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81caf9),
	.w1(32'h3b9b67b0),
	.w2(32'hba94c8cc),
	.w3(32'h39cafaff),
	.w4(32'hba5274cf),
	.w5(32'h3ad2a00c),
	.w6(32'h3ba7eee7),
	.w7(32'hbb6c2441),
	.w8(32'hbb3c4f2f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b1f78),
	.w1(32'h3b74c49d),
	.w2(32'hbb3b3807),
	.w3(32'h39996d32),
	.w4(32'hbb216a23),
	.w5(32'hbb97bf0e),
	.w6(32'h3b130d85),
	.w7(32'h3b18baab),
	.w8(32'h3abbdc00),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd46be7),
	.w1(32'h3b49864b),
	.w2(32'hbba0d32b),
	.w3(32'h3b834d7b),
	.w4(32'hbb1612b6),
	.w5(32'hbc15a3e4),
	.w6(32'h3bb8d278),
	.w7(32'hbb6c9c5a),
	.w8(32'hbc318338),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8a2da),
	.w1(32'h3a859ec4),
	.w2(32'h3a528796),
	.w3(32'hbc20cb8f),
	.w4(32'hbb27cc0e),
	.w5(32'h3b9bf3d3),
	.w6(32'hbc00f9c6),
	.w7(32'hbb0e96f5),
	.w8(32'h3b11b81b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1fda),
	.w1(32'hbc4b1f10),
	.w2(32'hbc37e6e8),
	.w3(32'hbc05a381),
	.w4(32'hbc028e72),
	.w5(32'hbbecaf75),
	.w6(32'hbb3ab91c),
	.w7(32'hbc143603),
	.w8(32'hbb843a19),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c1b2),
	.w1(32'h3b3cdce4),
	.w2(32'h3c287d06),
	.w3(32'hbc2f45d5),
	.w4(32'h3be0bb9d),
	.w5(32'h3c7559b8),
	.w6(32'hbbf4adf2),
	.w7(32'h3b15fae2),
	.w8(32'h3c27dc9f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0acdad),
	.w1(32'hbacdbb5f),
	.w2(32'hb991b6ba),
	.w3(32'h3c334843),
	.w4(32'h3ac17d7a),
	.w5(32'hb93a53cf),
	.w6(32'h3b175d88),
	.w7(32'hbbc2f110),
	.w8(32'hbb0cf28f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90b5564),
	.w1(32'hbb980406),
	.w2(32'hbc1abd21),
	.w3(32'h3bf07c4f),
	.w4(32'h3a69454d),
	.w5(32'hbc2da3a3),
	.w6(32'h3b8bb8bc),
	.w7(32'hbaa9cfd3),
	.w8(32'hbb90fc9e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc036c24),
	.w1(32'h3b293770),
	.w2(32'hbb240c0f),
	.w3(32'hbc77259c),
	.w4(32'hba34076f),
	.w5(32'h396cce72),
	.w6(32'hbc0e0b6c),
	.w7(32'h3a83dcab),
	.w8(32'hbb219c94),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b270d3e),
	.w1(32'hbb57cff4),
	.w2(32'h3c16a56f),
	.w3(32'h3af7dbd2),
	.w4(32'hbb9a65e9),
	.w5(32'h3c1f72db),
	.w6(32'h37f3a345),
	.w7(32'hbac0fbf6),
	.w8(32'h3bf447c2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b6aa0),
	.w1(32'h3aaa88bb),
	.w2(32'hbb43b79a),
	.w3(32'h3c29e165),
	.w4(32'h3c102158),
	.w5(32'h3ba576e0),
	.w6(32'h3bad6f0d),
	.w7(32'hba5a9a00),
	.w8(32'hbc416164),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc094c3a),
	.w1(32'hbb25df85),
	.w2(32'hbc2802a8),
	.w3(32'h3bd6bae1),
	.w4(32'hbc20b668),
	.w5(32'hba8ea33c),
	.w6(32'hbc485f99),
	.w7(32'hbc49a4a7),
	.w8(32'hbc294610),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391b8355),
	.w1(32'hbc44bb30),
	.w2(32'hbc1ddda1),
	.w3(32'h3b34b6f3),
	.w4(32'hbb7a08f3),
	.w5(32'hbc0750c0),
	.w6(32'h3b2defc1),
	.w7(32'hbb5f57e1),
	.w8(32'hbb44459a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1749),
	.w1(32'hbc65ad1d),
	.w2(32'hbc3b08b1),
	.w3(32'hbbcbf962),
	.w4(32'h3ad1c953),
	.w5(32'h3b82e9f4),
	.w6(32'hbc0db591),
	.w7(32'h3ae02559),
	.w8(32'hbb909490),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e188),
	.w1(32'h3afab9fa),
	.w2(32'h3ca6f547),
	.w3(32'hbc1c6506),
	.w4(32'hbb3b996b),
	.w5(32'h3bf0bd20),
	.w6(32'hbb2b9b3e),
	.w7(32'h3b7b1abf),
	.w8(32'h3c279998),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf7609),
	.w1(32'hba996068),
	.w2(32'hbb85a870),
	.w3(32'hbbd472c2),
	.w4(32'h3a9d342f),
	.w5(32'hbb63ed9d),
	.w6(32'h3a0c8f92),
	.w7(32'hbbe0071b),
	.w8(32'hbbf27290),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16d002),
	.w1(32'h3b3fbe76),
	.w2(32'h3b06d2f5),
	.w3(32'h3bc182dc),
	.w4(32'h386d8f67),
	.w5(32'h3b2370cf),
	.w6(32'h3bba77b9),
	.w7(32'h39876c24),
	.w8(32'hbaa3005c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba878c6),
	.w1(32'hbc324cdd),
	.w2(32'hbba3cbcd),
	.w3(32'hbbd8760a),
	.w4(32'hbc59e586),
	.w5(32'hba1f1ad5),
	.w6(32'hbb8599a7),
	.w7(32'hbc519237),
	.w8(32'h3b780fc5),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8b0b5),
	.w1(32'hb850dd50),
	.w2(32'h3a73a39a),
	.w3(32'h3ba105f6),
	.w4(32'hbbc8ac88),
	.w5(32'hbc383140),
	.w6(32'h3b412981),
	.w7(32'h3bbb51d6),
	.w8(32'hbb8ff105),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee29d3),
	.w1(32'hbb2e9bef),
	.w2(32'hbc0b2c03),
	.w3(32'hbbeb862f),
	.w4(32'h3b164e87),
	.w5(32'hbb946dbf),
	.w6(32'hbbd2bb18),
	.w7(32'hbaa199a1),
	.w8(32'hbb253483),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86335d),
	.w1(32'hba66138a),
	.w2(32'h3b7faaad),
	.w3(32'hbbf17a60),
	.w4(32'hba5182f0),
	.w5(32'h3c14e5cd),
	.w6(32'hbb03aa19),
	.w7(32'h3a96c669),
	.w8(32'h3a81dd14),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a64ce),
	.w1(32'h3a09d494),
	.w2(32'hbb944ba4),
	.w3(32'hbc0f4502),
	.w4(32'hbabffeb2),
	.w5(32'hbc2444a1),
	.w6(32'hbb68b686),
	.w7(32'hbb6a9c81),
	.w8(32'hbb8988af),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3383b),
	.w1(32'hba8062be),
	.w2(32'hbb3ea44a),
	.w3(32'h3b243a91),
	.w4(32'h395793ff),
	.w5(32'h3baffea2),
	.w6(32'hbac65b81),
	.w7(32'hbb82c772),
	.w8(32'hbae8ded8),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb331943),
	.w1(32'h3ba8934b),
	.w2(32'hbbaf68fb),
	.w3(32'hba0bd7bf),
	.w4(32'h3ca8781e),
	.w5(32'h3c1870b2),
	.w6(32'h3bba4ccb),
	.w7(32'h3c167588),
	.w8(32'h3b71ef94),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc48a0c),
	.w1(32'hbbadd198),
	.w2(32'hbb7f9966),
	.w3(32'h3ae689f5),
	.w4(32'hbb378083),
	.w5(32'hbb28b8de),
	.w6(32'h3b8ee694),
	.w7(32'hba41e4d2),
	.w8(32'hba95641d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f7af3),
	.w1(32'h3b0c39e5),
	.w2(32'hbb95ab35),
	.w3(32'hbacd4917),
	.w4(32'h3b6112c8),
	.w5(32'hbb4e8cf0),
	.w6(32'h3b5254be),
	.w7(32'h3b543fca),
	.w8(32'hbb071b37),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc82b49),
	.w1(32'h3a61e09e),
	.w2(32'h3bf1642d),
	.w3(32'h3b2701a6),
	.w4(32'hbbec360e),
	.w5(32'h3af5b8f5),
	.w6(32'hbacec55b),
	.w7(32'hbbb62870),
	.w8(32'h3b545362),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9bf0ac),
	.w1(32'hbb60343a),
	.w2(32'h3ad953f5),
	.w3(32'h3c9b2218),
	.w4(32'h3923c7f8),
	.w5(32'h3a379f6d),
	.w6(32'h3b5c8d9f),
	.w7(32'h3a590285),
	.w8(32'h3aa050cd),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7608a),
	.w1(32'h3c0ffc5a),
	.w2(32'h3c4b9b8d),
	.w3(32'hbc2c4f06),
	.w4(32'h3c4e82a0),
	.w5(32'h3cce81cc),
	.w6(32'hbb9945f0),
	.w7(32'h3b9c6395),
	.w8(32'h3c429cfc),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a600b),
	.w1(32'h3c2dfa7a),
	.w2(32'h3c13f59d),
	.w3(32'h3c78405d),
	.w4(32'h3b6cd766),
	.w5(32'h3c41ccc9),
	.w6(32'h3b5a3efb),
	.w7(32'h3a4afe6a),
	.w8(32'hb9e526f8),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b921dab),
	.w1(32'h3a313f94),
	.w2(32'hbb592d26),
	.w3(32'h3b635505),
	.w4(32'hbb80dab0),
	.w5(32'hbb23d750),
	.w6(32'hbbeb7e53),
	.w7(32'h3b4f3ca9),
	.w8(32'hb9b0f27b),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5139a3),
	.w1(32'hbb9bc42c),
	.w2(32'h3b0fa76e),
	.w3(32'h3c2217ba),
	.w4(32'hbb5358a9),
	.w5(32'hbc2ab15d),
	.w6(32'h3be86d29),
	.w7(32'hba9f5106),
	.w8(32'hbba5d0d7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f57d9),
	.w1(32'hba9c4818),
	.w2(32'h3ae73edb),
	.w3(32'h3c1d4c4c),
	.w4(32'h3bdf3e99),
	.w5(32'h3807ed66),
	.w6(32'h3c4e5ddc),
	.w7(32'h3ae0b7c5),
	.w8(32'h3ae9dc14),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb937a7a),
	.w1(32'h3ac3d378),
	.w2(32'hb88d9f78),
	.w3(32'hbc02c4fb),
	.w4(32'h3a97540f),
	.w5(32'hbbac2982),
	.w6(32'hb9771a87),
	.w7(32'h3b126de2),
	.w8(32'hba6b803b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb582fad),
	.w1(32'hbb844f8c),
	.w2(32'hbb9b5e2f),
	.w3(32'hbb54b05b),
	.w4(32'hbbe260c5),
	.w5(32'h3ac9a1c7),
	.w6(32'h398671cc),
	.w7(32'hbb735cd9),
	.w8(32'hb8b3df3b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad87cf),
	.w1(32'h3ba23cc3),
	.w2(32'h3c656bd0),
	.w3(32'hbb653c4c),
	.w4(32'h3be57659),
	.w5(32'h3cd2bbdb),
	.w6(32'hba7844fd),
	.w7(32'h3ba0a993),
	.w8(32'h3bbae22a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c2d45),
	.w1(32'h3aa47b4e),
	.w2(32'hba2f7a25),
	.w3(32'hbb750151),
	.w4(32'h3afa76aa),
	.w5(32'hbc185730),
	.w6(32'h3bef0b9d),
	.w7(32'h3bf62ac6),
	.w8(32'hbb2d097a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8408fe),
	.w1(32'h3ae33d7e),
	.w2(32'hbb6219d8),
	.w3(32'h3bf550be),
	.w4(32'h39e49342),
	.w5(32'h3b2fb54c),
	.w6(32'h3ae234e8),
	.w7(32'hbaf52603),
	.w8(32'hba0a8f01),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ffd71),
	.w1(32'hbc29f41d),
	.w2(32'h3c132fe6),
	.w3(32'hbb26d466),
	.w4(32'hbbba4f0f),
	.w5(32'h3bc37fc8),
	.w6(32'h3af9fead),
	.w7(32'hbb0b75f7),
	.w8(32'h3ac16a96),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa1c90),
	.w1(32'hba3fd805),
	.w2(32'hbb3a5edb),
	.w3(32'h3a298127),
	.w4(32'hbb2cedf1),
	.w5(32'hbb26c043),
	.w6(32'hbb8cb679),
	.w7(32'hbaaeadca),
	.w8(32'hbb1eb5d5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10ce53),
	.w1(32'hbc8696f8),
	.w2(32'hbc20db36),
	.w3(32'hbc578972),
	.w4(32'hbc24dd49),
	.w5(32'hbc5516cd),
	.w6(32'hbbaf3a04),
	.w7(32'hbc331f83),
	.w8(32'hbbb8abe4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773d07),
	.w1(32'hbba1ce80),
	.w2(32'hbb409e0a),
	.w3(32'hbc4634b7),
	.w4(32'h3b9df9fb),
	.w5(32'hbb169e13),
	.w6(32'hbc2c0603),
	.w7(32'h3aa0b97a),
	.w8(32'hb9b02a85),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1aff5),
	.w1(32'hbbd2602f),
	.w2(32'hbbd51da8),
	.w3(32'h3b90844b),
	.w4(32'hbbe8f42f),
	.w5(32'hbb9a6836),
	.w6(32'h3ad93048),
	.w7(32'hbb973b02),
	.w8(32'hbbb51f4e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a480),
	.w1(32'h3a14f923),
	.w2(32'hbbe90c6a),
	.w3(32'hb9cee43e),
	.w4(32'h3bda8c65),
	.w5(32'hbaceb6af),
	.w6(32'h39083cc3),
	.w7(32'h3aa6b2cb),
	.w8(32'hbb419a32),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad79436),
	.w1(32'h3b669488),
	.w2(32'hbbb302e6),
	.w3(32'hbc345ff6),
	.w4(32'h3c199fca),
	.w5(32'h3a8cfd18),
	.w6(32'hbb08ba6c),
	.w7(32'hba0ad383),
	.w8(32'hbb02ed9e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad54fc2),
	.w1(32'hbc52beb3),
	.w2(32'hbbeb991c),
	.w3(32'h39cbebf6),
	.w4(32'h3b5375e0),
	.w5(32'hbc290060),
	.w6(32'hbb5d02bc),
	.w7(32'h3bc4eade),
	.w8(32'h3bed6d62),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2456fb),
	.w1(32'hbc0d66ef),
	.w2(32'hbc44725e),
	.w3(32'hb982eee5),
	.w4(32'h39dfbfa7),
	.w5(32'hbbe8ef2a),
	.w6(32'hba7744d1),
	.w7(32'hbbc63d3d),
	.w8(32'hbbcf7776),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3e876),
	.w1(32'h3b8cc80c),
	.w2(32'h3c1fb671),
	.w3(32'hbbf800cf),
	.w4(32'h3c465157),
	.w5(32'h3b12ef4d),
	.w6(32'hbbeb81f1),
	.w7(32'h3c119ed5),
	.w8(32'h3c016354),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c102915),
	.w1(32'hbbf2b4c9),
	.w2(32'hba00be28),
	.w3(32'h3bee9189),
	.w4(32'hbaa850fd),
	.w5(32'h3ab54f95),
	.w6(32'h3b46fba2),
	.w7(32'h3b90c2a0),
	.w8(32'hba9d1fe6),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5579d),
	.w1(32'h3b750f85),
	.w2(32'hbb96f183),
	.w3(32'h3b9a374b),
	.w4(32'h3c0385be),
	.w5(32'h3c47c836),
	.w6(32'hba1b96c8),
	.w7(32'hbb96afd4),
	.w8(32'h3c15c2b6),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d1f88),
	.w1(32'hbc4d9608),
	.w2(32'h390f75cb),
	.w3(32'hbb800e75),
	.w4(32'hbb6e876c),
	.w5(32'h3bb9baac),
	.w6(32'hbb615456),
	.w7(32'hbb783319),
	.w8(32'h3be98639),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a345c1c),
	.w1(32'hb9952980),
	.w2(32'h3a8195c5),
	.w3(32'hbc0c3b4b),
	.w4(32'h3b25331a),
	.w5(32'h3a28478e),
	.w6(32'h3b7f61ae),
	.w7(32'h3bb0c62c),
	.w8(32'h3a4a6625),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e67ca),
	.w1(32'hbc2315b4),
	.w2(32'hbb5f89fd),
	.w3(32'hbbae7878),
	.w4(32'hbc2ec9c3),
	.w5(32'hbc04da80),
	.w6(32'hba8aa856),
	.w7(32'h3b8a0e2f),
	.w8(32'hbb567f17),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68274c),
	.w1(32'hbb9783f7),
	.w2(32'hbb869f6d),
	.w3(32'h3775f8a2),
	.w4(32'hbb20f199),
	.w5(32'hbc082e62),
	.w6(32'h3ae12a19),
	.w7(32'hbb307a7a),
	.w8(32'hbbafdb40),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc378986),
	.w1(32'hbb5c109f),
	.w2(32'hba30315d),
	.w3(32'hbc3642b8),
	.w4(32'hba817dae),
	.w5(32'hbb84b721),
	.w6(32'hbb8ae75c),
	.w7(32'hbb1cfb85),
	.w8(32'h3abc32f6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf91013),
	.w1(32'hbb8c427a),
	.w2(32'h3bd547c9),
	.w3(32'h3b896dfd),
	.w4(32'h3b9dfa2e),
	.w5(32'h3bc7a45b),
	.w6(32'hb9d27e5c),
	.w7(32'h3b10abf9),
	.w8(32'h3c075bc6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb826669),
	.w1(32'hbb5f3a5f),
	.w2(32'hb985d56c),
	.w3(32'hbc1b63c0),
	.w4(32'hbbb830a2),
	.w5(32'hbbf2c917),
	.w6(32'h3b25355e),
	.w7(32'h3ae040df),
	.w8(32'hbbaefab1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d8751),
	.w1(32'h3b6c1d6b),
	.w2(32'h38f972d6),
	.w3(32'hbbe603b2),
	.w4(32'h3bb631ea),
	.w5(32'h3c7916ef),
	.w6(32'h39973fde),
	.w7(32'h3bdc0f33),
	.w8(32'h3bc61567),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cc1c),
	.w1(32'hbae661b4),
	.w2(32'hbc225b96),
	.w3(32'h3b4190e7),
	.w4(32'h3a957e79),
	.w5(32'hbaca3468),
	.w6(32'h3c069070),
	.w7(32'hba51618e),
	.w8(32'hbb8a9820),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf86bd3),
	.w1(32'h3ae82cc2),
	.w2(32'hbc400271),
	.w3(32'hbbf51cfa),
	.w4(32'h3a0e5b92),
	.w5(32'hbbbd027f),
	.w6(32'hbb47b0b7),
	.w7(32'h3a9ab92f),
	.w8(32'hbbb843a6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7c051),
	.w1(32'hb9b0f345),
	.w2(32'h3afd67b0),
	.w3(32'hbb98cd43),
	.w4(32'h3b9ea1fb),
	.w5(32'h3c1ebc16),
	.w6(32'hbb346458),
	.w7(32'hb9c89810),
	.w8(32'h3bfd8407),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953fef0),
	.w1(32'h3b183aaa),
	.w2(32'hbabcba6c),
	.w3(32'hbb0543e7),
	.w4(32'h3bb84e2c),
	.w5(32'hb9dc3438),
	.w6(32'h3bad623e),
	.w7(32'hbb25afe6),
	.w8(32'hbad1076e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9163c),
	.w1(32'h3a609cb8),
	.w2(32'hbc2fcf80),
	.w3(32'h39e62682),
	.w4(32'h3b607b41),
	.w5(32'hbbfbe25b),
	.w6(32'hbaa05df6),
	.w7(32'hb9fab59e),
	.w8(32'hbb1f1e4b),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba5848),
	.w1(32'hbb1ebefc),
	.w2(32'hbbf1267d),
	.w3(32'h3b077fde),
	.w4(32'hbb299a52),
	.w5(32'hbb220b5c),
	.w6(32'hbb8029fb),
	.w7(32'hbbc6f75f),
	.w8(32'hbb566793),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ac87b),
	.w1(32'h3bc57cc3),
	.w2(32'h3ba01d75),
	.w3(32'hbc11ca1d),
	.w4(32'h3b99d757),
	.w5(32'h3a46a147),
	.w6(32'hbbbdb989),
	.w7(32'h3b7290b9),
	.w8(32'h3b4371c9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d15f7),
	.w1(32'hbb158ed9),
	.w2(32'hbbce60f9),
	.w3(32'hbb23f591),
	.w4(32'h3a0cc7fb),
	.w5(32'h38ac515e),
	.w6(32'hb787d273),
	.w7(32'h3bc6ca92),
	.w8(32'hba4c3c41),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b1e4f),
	.w1(32'h3c8c5fa1),
	.w2(32'h391bcd47),
	.w3(32'hbb7889b9),
	.w4(32'h3bed53e9),
	.w5(32'hbb1f59f5),
	.w6(32'h3a174b5e),
	.w7(32'h3baab05f),
	.w8(32'h3b1bb74e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bc323),
	.w1(32'hbb76db77),
	.w2(32'hbba9c0dc),
	.w3(32'hbbfe0a25),
	.w4(32'h3aa5e7bf),
	.w5(32'hbb5288d6),
	.w6(32'hbb74d44f),
	.w7(32'h3b5a06e7),
	.w8(32'hbb9cdaf4),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade81ff),
	.w1(32'h3bcdb4a8),
	.w2(32'hbb912543),
	.w3(32'hbabdd752),
	.w4(32'h3b0fd499),
	.w5(32'hbbdc9b63),
	.w6(32'hbb0a5c56),
	.w7(32'h3ba9b177),
	.w8(32'hbbfbc3ee),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c5ab6),
	.w1(32'hbc2056ae),
	.w2(32'hbc0af4f2),
	.w3(32'hbb56b005),
	.w4(32'hbc024072),
	.w5(32'hbbf5dea6),
	.w6(32'h3ba14418),
	.w7(32'hbbbbe782),
	.w8(32'hbbc538be),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b151c),
	.w1(32'h3bc1b2a2),
	.w2(32'hbb535e2a),
	.w3(32'hbc18cee2),
	.w4(32'hbbb441d7),
	.w5(32'hbc826706),
	.w6(32'h3b1b9fad),
	.w7(32'h3b530c18),
	.w8(32'hbb484fa5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6d32c9),
	.w1(32'h3a178b26),
	.w2(32'h3caa6021),
	.w3(32'hbc57c3ff),
	.w4(32'h3b27b67d),
	.w5(32'h3c765a7d),
	.w6(32'hbbbc34b2),
	.w7(32'h3c0b20ae),
	.w8(32'h3cb9b764),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82c40b),
	.w1(32'hbc0c7e51),
	.w2(32'hbbf6ce89),
	.w3(32'h3a867845),
	.w4(32'hbc7f5c86),
	.w5(32'hbc8cc5ce),
	.w6(32'hba927b89),
	.w7(32'hbba83a80),
	.w8(32'hbb20c65e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26950d),
	.w1(32'hbac1f2a9),
	.w2(32'hbb8642aa),
	.w3(32'hb965ec15),
	.w4(32'hb9e83312),
	.w5(32'hbc21373e),
	.w6(32'h3aeffb06),
	.w7(32'hbc0f027c),
	.w8(32'hbc210e7d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb139a52),
	.w1(32'hbc0eb647),
	.w2(32'h3b1c777c),
	.w3(32'h3bb3896b),
	.w4(32'hbb12837e),
	.w5(32'hbb06f1f4),
	.w6(32'hbb187a3d),
	.w7(32'hbb91153c),
	.w8(32'h3aa00928),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd56948),
	.w1(32'hbc75c1e9),
	.w2(32'hbc5c738a),
	.w3(32'hbac36219),
	.w4(32'hbc77f4ba),
	.w5(32'hbcb9a85a),
	.w6(32'hbad555d2),
	.w7(32'hbcbcb1b2),
	.w8(32'hbcbf5bbb),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8dd1f1),
	.w1(32'h39ab92d5),
	.w2(32'hbb9aad7e),
	.w3(32'hbc6d84e2),
	.w4(32'hbb9ac14c),
	.w5(32'hbb7e3f4d),
	.w6(32'hbc87cc69),
	.w7(32'hbadc7f52),
	.w8(32'hbbbc6104),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b783761),
	.w1(32'hbc1a5e93),
	.w2(32'hbc030da6),
	.w3(32'h3b408b61),
	.w4(32'hbba622e9),
	.w5(32'hbbcc3a43),
	.w6(32'hba6b0082),
	.w7(32'hbb5fe812),
	.w8(32'hbba676ce),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63adfe),
	.w1(32'hbb677726),
	.w2(32'h3ab9eda1),
	.w3(32'hbbe336a6),
	.w4(32'h3ae4447f),
	.w5(32'h3ae7bcd8),
	.w6(32'hba3724ab),
	.w7(32'h3998fb57),
	.w8(32'hba2984da),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a998bc2),
	.w1(32'h3b3bdfe1),
	.w2(32'h3bd94571),
	.w3(32'h3b8781bd),
	.w4(32'h3b09208b),
	.w5(32'h3ac3751e),
	.w6(32'h3b29e17a),
	.w7(32'h3c0eebad),
	.w8(32'h3be28b63),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269c7a),
	.w1(32'hbb99a7ba),
	.w2(32'hbb9a8c94),
	.w3(32'h38c9bc8c),
	.w4(32'hbb76bb0c),
	.w5(32'hba3c86d1),
	.w6(32'h3b84c7ee),
	.w7(32'hba0c94ca),
	.w8(32'h39537c7c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb185cf),
	.w1(32'h38ceca0c),
	.w2(32'hbb1ed7db),
	.w3(32'hbab6b130),
	.w4(32'hbaae6481),
	.w5(32'hbc16fce8),
	.w6(32'h3b38b59b),
	.w7(32'h3aa3c230),
	.w8(32'hbb161e03),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcfac99),
	.w1(32'h39f37026),
	.w2(32'hbaed6119),
	.w3(32'hba6b817a),
	.w4(32'hbb341816),
	.w5(32'hb9907383),
	.w6(32'hbb17f6c6),
	.w7(32'hba4ebb3b),
	.w8(32'h3a609591),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dbfff),
	.w1(32'hbc03b904),
	.w2(32'hb9582203),
	.w3(32'hbbdc6d85),
	.w4(32'hba5cdb90),
	.w5(32'h3c7d4410),
	.w6(32'h3b2a2432),
	.w7(32'h3b7323f2),
	.w8(32'h3ba3a604),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b63ce),
	.w1(32'hbae230c4),
	.w2(32'hbb99746f),
	.w3(32'h3aca5437),
	.w4(32'hbbce23dd),
	.w5(32'h3baf0787),
	.w6(32'h3babd6ad),
	.w7(32'hba9ac469),
	.w8(32'hbbbf87af),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd07f89),
	.w1(32'h3b30accc),
	.w2(32'h3c8689c9),
	.w3(32'hbad97a5e),
	.w4(32'h3b1236d0),
	.w5(32'h3bc6f269),
	.w6(32'hba36dc83),
	.w7(32'h3aed6a64),
	.w8(32'h3c099118),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c494b18),
	.w1(32'h3a06c194),
	.w2(32'h3bfb1bbd),
	.w3(32'h3c84dd02),
	.w4(32'h3b83626e),
	.w5(32'h3b9430d9),
	.w6(32'h3c6006b8),
	.w7(32'hbb210abc),
	.w8(32'h3b91a2ef),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bc001),
	.w1(32'h3b5dafb4),
	.w2(32'hbc0287a0),
	.w3(32'h3c573e9b),
	.w4(32'h3c1c63e9),
	.w5(32'hbbda9857),
	.w6(32'h3c27cbb4),
	.w7(32'h3baeb42c),
	.w8(32'h3b12a0ba),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59ad7c),
	.w1(32'hbb3175b3),
	.w2(32'hbaa530a3),
	.w3(32'h3b86715a),
	.w4(32'hba3c16e2),
	.w5(32'h3adf137f),
	.w6(32'h3aa679b1),
	.w7(32'h3accf7e0),
	.w8(32'hbb37de08),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac4e70),
	.w1(32'hba5e308c),
	.w2(32'hbb8b669f),
	.w3(32'hbb1c1af2),
	.w4(32'hba79cb30),
	.w5(32'h3bc72a4d),
	.w6(32'hbb926ef3),
	.w7(32'h3a864ac8),
	.w8(32'h3b4a9afb),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a6ea1),
	.w1(32'h3b38ef4a),
	.w2(32'h3c8abba6),
	.w3(32'hbc21ee13),
	.w4(32'h3b7ef5bc),
	.w5(32'h3b9cc67f),
	.w6(32'hbbc5e4d6),
	.w7(32'h3c11d8f4),
	.w8(32'h3c2b1a21),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c283d06),
	.w1(32'hb9ced16c),
	.w2(32'h3b8ea204),
	.w3(32'h3c354532),
	.w4(32'h3ab05158),
	.w5(32'h3a15b090),
	.w6(32'h3c29dc63),
	.w7(32'h3b48f165),
	.w8(32'h3c18c5cc),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd58af),
	.w1(32'hbb8724f8),
	.w2(32'hbc1d973a),
	.w3(32'hbb3172ed),
	.w4(32'hba3ba323),
	.w5(32'hbc3de0d0),
	.w6(32'hbb0f8009),
	.w7(32'hbb55c3f1),
	.w8(32'hbc3a9bad),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d1201),
	.w1(32'h3c386a4c),
	.w2(32'h3c02f12c),
	.w3(32'h3bf26459),
	.w4(32'h3c357ef0),
	.w5(32'h3beca866),
	.w6(32'h3a0b88a4),
	.w7(32'hbb8b7e80),
	.w8(32'hbc0d03ee),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3c663),
	.w1(32'hbb25a024),
	.w2(32'h3bd86f71),
	.w3(32'h3ca0c521),
	.w4(32'hbabb71fe),
	.w5(32'h3a7bdef4),
	.w6(32'hbbd57ef0),
	.w7(32'hbb6023aa),
	.w8(32'hbb68f0fb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ceb7),
	.w1(32'h3bd9ef2d),
	.w2(32'h3b447df6),
	.w3(32'hbb289523),
	.w4(32'h3ba2c9f6),
	.w5(32'hba773110),
	.w6(32'hbbd92f06),
	.w7(32'h38346de3),
	.w8(32'hbb2cf4ea),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862488c),
	.w1(32'h3a7f06be),
	.w2(32'h3bb3a393),
	.w3(32'hbbb11f24),
	.w4(32'h392ee415),
	.w5(32'hbbba6375),
	.w6(32'hbae2ede5),
	.w7(32'h3b3c8967),
	.w8(32'h3b6fa140),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a202c1a),
	.w1(32'h3b51463e),
	.w2(32'hbaf2ddaa),
	.w3(32'hbaf25550),
	.w4(32'h3c7e2ae0),
	.w5(32'hbbcce7c8),
	.w6(32'hbace2335),
	.w7(32'h3c5c1d38),
	.w8(32'hb82edc1e),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0a70b),
	.w1(32'hbb93285f),
	.w2(32'h3a2f09f2),
	.w3(32'hbb680992),
	.w4(32'hbb7b26ec),
	.w5(32'h3b524ab3),
	.w6(32'hbb9010e6),
	.w7(32'h3bbbf7b1),
	.w8(32'h3b7fac33),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b4ff),
	.w1(32'hbbcc5c36),
	.w2(32'hbba6f684),
	.w3(32'hbbd102b6),
	.w4(32'hbb58b6cf),
	.w5(32'hbc0ef15c),
	.w6(32'h3b1563cc),
	.w7(32'hbbba4bc0),
	.w8(32'hbabe3519),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16219c),
	.w1(32'hbb93a1c0),
	.w2(32'hbb67cd19),
	.w3(32'h3b8d939d),
	.w4(32'hbbcef3df),
	.w5(32'hba1436b2),
	.w6(32'h3b97343c),
	.w7(32'hbc079d3b),
	.w8(32'hbac5e887),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa2080),
	.w1(32'h3b392efa),
	.w2(32'h3b8177e9),
	.w3(32'hbaf89ba4),
	.w4(32'h3c0198cf),
	.w5(32'h3cae9075),
	.w6(32'hbbeab3ce),
	.w7(32'hbb9392ba),
	.w8(32'h3c737667),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb81c30),
	.w1(32'hbb3409df),
	.w2(32'h3b7499c0),
	.w3(32'hb84199fd),
	.w4(32'hbb23349a),
	.w5(32'h3c0a4627),
	.w6(32'h3ace76b1),
	.w7(32'h3b7e1306),
	.w8(32'h3b860861),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc289da2),
	.w1(32'hbae3ec6d),
	.w2(32'hbb834a3a),
	.w3(32'hbc3d206c),
	.w4(32'hbb3f53e3),
	.w5(32'hba692931),
	.w6(32'hbbdaecae),
	.w7(32'hbb677d38),
	.w8(32'hbb92bc39),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b803bab),
	.w1(32'h3b89d512),
	.w2(32'hbb95e923),
	.w3(32'h38df7f3c),
	.w4(32'hbb8394d0),
	.w5(32'hbc247215),
	.w6(32'h3b146989),
	.w7(32'h3c0b0744),
	.w8(32'hbc5fdd16),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3ae08),
	.w1(32'hbc137c6a),
	.w2(32'hbc1ce781),
	.w3(32'h3bee3d0a),
	.w4(32'hbc21eda8),
	.w5(32'h3af8b06a),
	.w6(32'h3ae6bff8),
	.w7(32'hbc00436e),
	.w8(32'hbb1910fc),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1f37c),
	.w1(32'h3bddab6a),
	.w2(32'h3ca2fa6a),
	.w3(32'h3b75225e),
	.w4(32'h3c2a86bb),
	.w5(32'h3ca7518f),
	.w6(32'h3b863f07),
	.w7(32'h3b4385da),
	.w8(32'h3bbea797),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae86d06),
	.w1(32'h3b49bd1b),
	.w2(32'h3c7670ea),
	.w3(32'h3cb8d5ca),
	.w4(32'hbc0dcd7d),
	.w5(32'h3b952f05),
	.w6(32'h3c1be76d),
	.w7(32'hbc06ab54),
	.w8(32'h3ba89365),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d079),
	.w1(32'hbbd94668),
	.w2(32'h3bfcab61),
	.w3(32'h3be9c64b),
	.w4(32'hbb6d55b6),
	.w5(32'h3bab8b3e),
	.w6(32'hbb050cfb),
	.w7(32'hbb766527),
	.w8(32'h3b8dae9b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fd256f),
	.w1(32'h3952b96e),
	.w2(32'h3bd1d13d),
	.w3(32'hba2eb642),
	.w4(32'hba05e425),
	.w5(32'h3b21a8ae),
	.w6(32'hbb122d4e),
	.w7(32'h38112f9e),
	.w8(32'h3b9945b4),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd5b53),
	.w1(32'hbbd6013f),
	.w2(32'hbbd10e0f),
	.w3(32'hbc3e6e8c),
	.w4(32'hbae4d8f2),
	.w5(32'h3ac75091),
	.w6(32'hbc3ca318),
	.w7(32'h3b037aad),
	.w8(32'h3b682427),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce43cc),
	.w1(32'h3c3fa2fd),
	.w2(32'h3b27486a),
	.w3(32'hbb55b189),
	.w4(32'h3bb99609),
	.w5(32'hbb9234a0),
	.w6(32'h3b922428),
	.w7(32'h3b56fe78),
	.w8(32'hbb0428db),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42fa6d),
	.w1(32'h3b047379),
	.w2(32'hba86619b),
	.w3(32'h3ba74b1a),
	.w4(32'hba86ffa0),
	.w5(32'hb9c10825),
	.w6(32'h3bf3e206),
	.w7(32'hbb713c1d),
	.w8(32'hbad9b377),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1adaea),
	.w1(32'hbc411f62),
	.w2(32'hbb43228a),
	.w3(32'hbc4a7385),
	.w4(32'hbc379839),
	.w5(32'hbc5af939),
	.w6(32'hbc09281a),
	.w7(32'hba6c75f0),
	.w8(32'hbb12767f),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a96cd),
	.w1(32'h3b1bd8a6),
	.w2(32'h3b89685c),
	.w3(32'h3a51a92d),
	.w4(32'h3a8fd307),
	.w5(32'hbbf7c3b3),
	.w6(32'h3b3b4c58),
	.w7(32'hbbc020cf),
	.w8(32'hbb3c3b4f),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83e056),
	.w1(32'hbab3bc47),
	.w2(32'h3c89f8d4),
	.w3(32'hbb07ba20),
	.w4(32'h3c27a027),
	.w5(32'h3c2ebe47),
	.w6(32'hbbcdf2f1),
	.w7(32'h3b57e51a),
	.w8(32'h3c18ba67),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afd80),
	.w1(32'hbb288616),
	.w2(32'hba97e231),
	.w3(32'hbbb9c36c),
	.w4(32'hba2ca53d),
	.w5(32'h3916da83),
	.w6(32'hbc1a5a87),
	.w7(32'h3beeaddd),
	.w8(32'h3b5ec78a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ad450),
	.w1(32'h3b6b9de5),
	.w2(32'h3b3920c9),
	.w3(32'h3b86adde),
	.w4(32'hb8a3ab9c),
	.w5(32'hbb4ddb93),
	.w6(32'h39986388),
	.w7(32'hbb9624fa),
	.w8(32'hbb997f65),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1f1c6),
	.w1(32'h3a4e8de7),
	.w2(32'h3993ffa9),
	.w3(32'hbb2e619f),
	.w4(32'h3b3119b9),
	.w5(32'h3ba8a32e),
	.w6(32'hb8108877),
	.w7(32'hbb4a9525),
	.w8(32'hbb0ccc55),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50b72),
	.w1(32'hbb25d562),
	.w2(32'hbae44416),
	.w3(32'h3c139e9a),
	.w4(32'hbb851009),
	.w5(32'hbba1115e),
	.w6(32'h380bd404),
	.w7(32'hba14546e),
	.w8(32'h399d9e27),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf6830),
	.w1(32'hbb226f57),
	.w2(32'hbae6f790),
	.w3(32'hb98d06ad),
	.w4(32'hb9965521),
	.w5(32'h3b33aed2),
	.w6(32'h3adf6ab1),
	.w7(32'hbad9a017),
	.w8(32'hba7711ac),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04c987),
	.w1(32'hbb5a216a),
	.w2(32'hbb4a469a),
	.w3(32'hbaf65dc9),
	.w4(32'hbb8a0088),
	.w5(32'h3b9fe840),
	.w6(32'hbb499bbb),
	.w7(32'hbbbd4fe7),
	.w8(32'h3b2a01e2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a535436),
	.w1(32'hbc023918),
	.w2(32'hbba54a3a),
	.w3(32'hbbd4d429),
	.w4(32'hbbba987e),
	.w5(32'hb96174da),
	.w6(32'hbbe49e5a),
	.w7(32'hbb8a21f2),
	.w8(32'hbb28b947),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3100e3),
	.w1(32'h39d537d6),
	.w2(32'h3acf3b02),
	.w3(32'hbb7bb14e),
	.w4(32'h3b915998),
	.w5(32'h3a354d65),
	.w6(32'hbb0fc392),
	.w7(32'h3b121a53),
	.w8(32'h3b45c606),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24d64b),
	.w1(32'hba944da1),
	.w2(32'hbb4896dd),
	.w3(32'h3ba9f32e),
	.w4(32'hbb93da9d),
	.w5(32'hbb4c5ffe),
	.w6(32'h3ba4708d),
	.w7(32'hbbac6a44),
	.w8(32'h3b9d0ae1),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86c345),
	.w1(32'h3aad58da),
	.w2(32'h3b604ffb),
	.w3(32'h3b0f625f),
	.w4(32'hba092d4d),
	.w5(32'h39f7d015),
	.w6(32'h3be25048),
	.w7(32'hbb94c0b3),
	.w8(32'hba67eedf),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e8069),
	.w1(32'hb9f53d34),
	.w2(32'hba6c224a),
	.w3(32'h3a8e5965),
	.w4(32'h3bd82f58),
	.w5(32'hba5a6fd7),
	.w6(32'h3b49e117),
	.w7(32'h3b9f0eb3),
	.w8(32'h3afa47c2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacf7da),
	.w1(32'h3aa17c5f),
	.w2(32'h3b669620),
	.w3(32'hbb5725ea),
	.w4(32'h39c7da57),
	.w5(32'h3a8ece7c),
	.w6(32'hbaadc228),
	.w7(32'h3b94eaaa),
	.w8(32'h3bdafe0d),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fe0e4),
	.w1(32'h3b9d4b09),
	.w2(32'h3b70920d),
	.w3(32'h3ba62e22),
	.w4(32'h3b3c98b2),
	.w5(32'h3b3730ff),
	.w6(32'h3bb8e70e),
	.w7(32'h39422fc1),
	.w8(32'h3b1eb062),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39effa3d),
	.w1(32'hba71275a),
	.w2(32'hba4b2b35),
	.w3(32'h3992903c),
	.w4(32'hba23e1fa),
	.w5(32'hbb5dcf6d),
	.w6(32'h3b826912),
	.w7(32'hbb45ddc7),
	.w8(32'hbb23dd0f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba5a56),
	.w1(32'h3bf6ab60),
	.w2(32'h3c55ef7a),
	.w3(32'hbb4ea378),
	.w4(32'hbb75e1b2),
	.w5(32'h3b9e3b59),
	.w6(32'hbb401952),
	.w7(32'hbbecdd86),
	.w8(32'hbb0ad8c6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a872f),
	.w1(32'h3bd10d16),
	.w2(32'h39f01f72),
	.w3(32'h3bf9160f),
	.w4(32'h3b4f8dc3),
	.w5(32'h3bb7da32),
	.w6(32'h3b43a9bc),
	.w7(32'hb983aa8b),
	.w8(32'h3b5a7762),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a406653),
	.w1(32'h39e07049),
	.w2(32'h3b73194e),
	.w3(32'hb84a950e),
	.w4(32'hbaaacf7d),
	.w5(32'hbc00e3fc),
	.w6(32'h3b8f3da9),
	.w7(32'hba3f62d5),
	.w8(32'h3a6edb9b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89dffa),
	.w1(32'hbb9c81f9),
	.w2(32'hba99af16),
	.w3(32'hbbe1c727),
	.w4(32'hbc0ee753),
	.w5(32'hbc0b30af),
	.w6(32'hba8ea766),
	.w7(32'hbb7f4ce2),
	.w8(32'hbbb0f0c4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87e2df),
	.w1(32'hba2abae5),
	.w2(32'hba833313),
	.w3(32'h3af46c63),
	.w4(32'hbb394d7b),
	.w5(32'h3ae8e96f),
	.w6(32'hb91c5b1f),
	.w7(32'hba3f86d2),
	.w8(32'h39170a73),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7448bf),
	.w1(32'hbb304214),
	.w2(32'h3b5e7684),
	.w3(32'hb7ec800d),
	.w4(32'h3ab3e95e),
	.w5(32'h3b8b4726),
	.w6(32'hbae0e2c4),
	.w7(32'hba25a252),
	.w8(32'hb84471db),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe8fb4),
	.w1(32'h3aad8822),
	.w2(32'hb8bfed63),
	.w3(32'hba05320f),
	.w4(32'h3c4f326b),
	.w5(32'hbb076caf),
	.w6(32'hbaa0799f),
	.w7(32'h3c2c4818),
	.w8(32'h3b0e96f8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b315683),
	.w1(32'h3bb96110),
	.w2(32'h3b947dd1),
	.w3(32'hb8a6af36),
	.w4(32'h3ae554a0),
	.w5(32'hbc041139),
	.w6(32'hba9b47bc),
	.w7(32'hbabcc625),
	.w8(32'hbbf76562),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86d4f3),
	.w1(32'h3af62208),
	.w2(32'h3bb5145a),
	.w3(32'hba9f4b4a),
	.w4(32'hb986c107),
	.w5(32'hb9e83002),
	.w6(32'hbb68de21),
	.w7(32'hba5dd082),
	.w8(32'h3af79e94),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c55450),
	.w1(32'hbba5c0a0),
	.w2(32'hbb25ba42),
	.w3(32'hbb850c87),
	.w4(32'hbc1935d7),
	.w5(32'hbbd7724d),
	.w6(32'h3b28a04d),
	.w7(32'hbc09f466),
	.w8(32'hbbc78b00),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e644),
	.w1(32'hbb66693f),
	.w2(32'h39ed54aa),
	.w3(32'hba96d4b9),
	.w4(32'hbb11456d),
	.w5(32'hbb8c9ca9),
	.w6(32'hb9859c17),
	.w7(32'h3b60d16b),
	.w8(32'h3bc5aba7),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae3a1f),
	.w1(32'h3b36d107),
	.w2(32'h3ba95fa4),
	.w3(32'hb87136a7),
	.w4(32'hbad1a2e5),
	.w5(32'hbadfaa19),
	.w6(32'h3a95afdf),
	.w7(32'hbb0b0e80),
	.w8(32'h3ae0c7c9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beacbfd),
	.w1(32'hbbacfaa9),
	.w2(32'hbb23b848),
	.w3(32'hba9f45d7),
	.w4(32'hbbb8aff0),
	.w5(32'hbb02f174),
	.w6(32'hba4fe321),
	.w7(32'hbb8942b8),
	.w8(32'hbbacf9bf),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8575b9),
	.w1(32'h3a251cdf),
	.w2(32'hb99b199d),
	.w3(32'h3ac0a219),
	.w4(32'h3a1942a9),
	.w5(32'h3b0b1017),
	.w6(32'hbbf805ac),
	.w7(32'h3a220831),
	.w8(32'h3a9a1098),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba9c36),
	.w1(32'h3ba88036),
	.w2(32'h3b7865f4),
	.w3(32'h3a700980),
	.w4(32'h3c7c0ce0),
	.w5(32'h3b9a7c8d),
	.w6(32'h3b1e1f7c),
	.w7(32'h3bfabdf4),
	.w8(32'h3c016799),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acac187),
	.w1(32'hbb39b7ef),
	.w2(32'h3a797577),
	.w3(32'h3b90b887),
	.w4(32'h3bcce9d7),
	.w5(32'h3b00f886),
	.w6(32'h3ba0ad46),
	.w7(32'h3c5b6e88),
	.w8(32'hbac69596),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98c692),
	.w1(32'h3bd18762),
	.w2(32'h3afe49b4),
	.w3(32'h3c0c75e4),
	.w4(32'h3c6a7d0c),
	.w5(32'h3c05dad7),
	.w6(32'h3bcc8272),
	.w7(32'h3c03cbf9),
	.w8(32'h3ccfb411),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5c285),
	.w1(32'hbad2a2f9),
	.w2(32'hba7c0463),
	.w3(32'hbb5a8c70),
	.w4(32'hbb4f42e6),
	.w5(32'hba9e89fd),
	.w6(32'h3c284113),
	.w7(32'hbac02a0d),
	.w8(32'hbb28041b),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07a317),
	.w1(32'hbb92a126),
	.w2(32'hbae8470b),
	.w3(32'hbb3d519c),
	.w4(32'hba92b597),
	.w5(32'hba3ea999),
	.w6(32'hbba13cd6),
	.w7(32'hbb504484),
	.w8(32'hbb5e92d6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba29d2e),
	.w1(32'hbb03ce56),
	.w2(32'hba7fc71b),
	.w3(32'hbb211176),
	.w4(32'h3baa975e),
	.w5(32'hbafa3acd),
	.w6(32'hba0328d8),
	.w7(32'h3a34a502),
	.w8(32'hbb7a196f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f8e6),
	.w1(32'h3b09f468),
	.w2(32'h3bb342d5),
	.w3(32'h3b18b154),
	.w4(32'h3a410fa7),
	.w5(32'h3bdf55a1),
	.w6(32'h3ab3fe4a),
	.w7(32'h3a3b3b64),
	.w8(32'h3bc3b47b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1eadf1),
	.w1(32'hba0848ce),
	.w2(32'h3bc5f55c),
	.w3(32'h3a051375),
	.w4(32'hba915e69),
	.w5(32'hbad989f4),
	.w6(32'h3c098ed8),
	.w7(32'hbb0494b2),
	.w8(32'hbb2b555a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77ab0),
	.w1(32'h3a62dbff),
	.w2(32'h3b2dd166),
	.w3(32'hbb53be58),
	.w4(32'hba3421e2),
	.w5(32'hbae35b26),
	.w6(32'hbb2b20b9),
	.w7(32'h38b474d3),
	.w8(32'hb9ba8c05),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15f03b),
	.w1(32'h3b064370),
	.w2(32'hb8e2ec7d),
	.w3(32'hbaeee76c),
	.w4(32'h3a60eeb7),
	.w5(32'hbb3cd7c8),
	.w6(32'hbad86aa6),
	.w7(32'hba2f2ead),
	.w8(32'hba765c86),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb347b8c),
	.w1(32'hbb4387df),
	.w2(32'hbba53748),
	.w3(32'hbb605b49),
	.w4(32'hbb7536b4),
	.w5(32'hbb230449),
	.w6(32'hbabac22b),
	.w7(32'hbb748093),
	.w8(32'hbb07a3be),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80e38a),
	.w1(32'hbb3d5c20),
	.w2(32'hbb15e216),
	.w3(32'hbb3a52c2),
	.w4(32'hbae28da6),
	.w5(32'h3a810612),
	.w6(32'hbb863d86),
	.w7(32'h3b4ad4e7),
	.w8(32'h3bc16e53),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81a101),
	.w1(32'hbb11870d),
	.w2(32'hbb7c898f),
	.w3(32'h3a93d3bd),
	.w4(32'hbb457c06),
	.w5(32'h3a49182b),
	.w6(32'h3b9c2a99),
	.w7(32'hbb888c4d),
	.w8(32'hbb958a1f),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbaf21),
	.w1(32'h3b29fe9b),
	.w2(32'hb98740d7),
	.w3(32'h3abcbb24),
	.w4(32'hbb8b5a04),
	.w5(32'hbb31770e),
	.w6(32'hbb00043d),
	.w7(32'hbb00c438),
	.w8(32'hb986496c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa07821),
	.w1(32'hba7094d4),
	.w2(32'h3b2cfa9f),
	.w3(32'h3b0ac9df),
	.w4(32'h3b7f5eb7),
	.w5(32'hb9a29184),
	.w6(32'h3bac61a5),
	.w7(32'h3b5cca98),
	.w8(32'h3acdd9cb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77cab4),
	.w1(32'hbab01d5a),
	.w2(32'hbaa3728c),
	.w3(32'h3b900001),
	.w4(32'h398c4563),
	.w5(32'h3b2f9c22),
	.w6(32'h3a298962),
	.w7(32'h3b786294),
	.w8(32'h3b9ea274),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fbc837),
	.w1(32'hbbfe7350),
	.w2(32'hbb8d1ff7),
	.w3(32'h39bc2e41),
	.w4(32'h3a8ae432),
	.w5(32'h3ae12a18),
	.w6(32'h3b9bfa72),
	.w7(32'hbb4c43f6),
	.w8(32'hbaf4fa47),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12c2b),
	.w1(32'hba749ed3),
	.w2(32'hbb87fe29),
	.w3(32'hbb432312),
	.w4(32'hbad017dd),
	.w5(32'hbb902076),
	.w6(32'hbb78bc83),
	.w7(32'hbb2fec40),
	.w8(32'hb96dfc3c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074b6e),
	.w1(32'hb8a699d9),
	.w2(32'h39ae2390),
	.w3(32'h3b7dedc4),
	.w4(32'hbb83373c),
	.w5(32'hbb82c294),
	.w6(32'h3bb189a3),
	.w7(32'hbb906064),
	.w8(32'hbb1f10ce),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af74351),
	.w1(32'h3aa92362),
	.w2(32'hbb35d2e8),
	.w3(32'hbb09120e),
	.w4(32'hba859f00),
	.w5(32'h3ac81838),
	.w6(32'hbaf78e27),
	.w7(32'hbb13e953),
	.w8(32'hbb527315),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae342b2),
	.w1(32'hbb1e9000),
	.w2(32'hbb5e724a),
	.w3(32'h3ba65cea),
	.w4(32'h3a8e3cbc),
	.w5(32'hbb99e748),
	.w6(32'h39b6942e),
	.w7(32'hb90cffa7),
	.w8(32'hbad153d7),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba17f36c),
	.w1(32'hbb8e0135),
	.w2(32'hbb189a4a),
	.w3(32'h3a156591),
	.w4(32'hbb6c41d7),
	.w5(32'hbb14dffd),
	.w6(32'h39faa6a3),
	.w7(32'hbb77bebf),
	.w8(32'hbbdf7a03),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925db03),
	.w1(32'hbb898ced),
	.w2(32'hbb8486f3),
	.w3(32'hba973b05),
	.w4(32'hbb444877),
	.w5(32'hbb4c3dc8),
	.w6(32'hbb916c19),
	.w7(32'hb9ea2d16),
	.w8(32'hbb3373ea),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007719),
	.w1(32'h399db103),
	.w2(32'h3b963867),
	.w3(32'hbaac98f3),
	.w4(32'hba0e3717),
	.w5(32'h3b27202c),
	.w6(32'hbb3609c5),
	.w7(32'hba51812d),
	.w8(32'h3a2d790f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fd0b4),
	.w1(32'hbb970165),
	.w2(32'hbb259f73),
	.w3(32'h3aa4984d),
	.w4(32'hbb19b9df),
	.w5(32'hbb5f0295),
	.w6(32'h3af49070),
	.w7(32'h3ba70ffd),
	.w8(32'h3b5a56bf),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb476993),
	.w1(32'hb9c54d62),
	.w2(32'h3b136042),
	.w3(32'h3a6f6a90),
	.w4(32'hbb25a017),
	.w5(32'hba30b797),
	.w6(32'h3bbdaec5),
	.w7(32'hbb68cdf1),
	.w8(32'hba01296d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397cd3e6),
	.w1(32'hbb84118b),
	.w2(32'h3911a480),
	.w3(32'hb915bbea),
	.w4(32'hbb57b8ce),
	.w5(32'hbadd7d9c),
	.w6(32'h39613913),
	.w7(32'h3950ab5a),
	.w8(32'h3b024f13),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988c660),
	.w1(32'hba09d65a),
	.w2(32'h3a94225c),
	.w3(32'h3b062405),
	.w4(32'h3a996340),
	.w5(32'h3c102d22),
	.w6(32'hb8d0ed68),
	.w7(32'hbb9ede21),
	.w8(32'h3a2b188d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b817d77),
	.w1(32'hb955c277),
	.w2(32'h3b5d6e10),
	.w3(32'h3be552c5),
	.w4(32'h3bfaf0c5),
	.w5(32'h3b834703),
	.w6(32'h3b623dd7),
	.w7(32'hbac56aaf),
	.w8(32'hba51413f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20773f),
	.w1(32'hbad47107),
	.w2(32'hbb995200),
	.w3(32'hbab96fd2),
	.w4(32'h3b1c3187),
	.w5(32'hbb8687dc),
	.w6(32'hbaeea5d9),
	.w7(32'h3b02f97e),
	.w8(32'h3974a517),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc306d65),
	.w1(32'hbb4d6f0c),
	.w2(32'hbb24a98a),
	.w3(32'hbc62be83),
	.w4(32'hbbc08234),
	.w5(32'hbb9815d0),
	.w6(32'hbb8038cd),
	.w7(32'hbbbb262a),
	.w8(32'hbbc753aa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule