module layer_8_featuremap_73(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8780a),
	.w1(32'hbc06b163),
	.w2(32'h3b2ee97d),
	.w3(32'hbba2eb67),
	.w4(32'hbbd5dbba),
	.w5(32'h3a63e4d8),
	.w6(32'hbb38e3d9),
	.w7(32'hbb0a3941),
	.w8(32'hbb8623bb),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30bec6),
	.w1(32'hba943c17),
	.w2(32'hba986baf),
	.w3(32'hbada9653),
	.w4(32'hb90701e7),
	.w5(32'h39829ddd),
	.w6(32'hba1e235f),
	.w7(32'h389cd733),
	.w8(32'hb9d5cae3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a831393),
	.w1(32'h3a529864),
	.w2(32'hb89c5162),
	.w3(32'h3aa2dfc3),
	.w4(32'h3b4aba69),
	.w5(32'h3b1ee7e3),
	.w6(32'hb9a3f3a6),
	.w7(32'h3adc7306),
	.w8(32'hbc0203a9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29a300),
	.w1(32'h3cbf71e6),
	.w2(32'hbb45ae7c),
	.w3(32'hbc079bd2),
	.w4(32'hbbb17be2),
	.w5(32'hbbd87840),
	.w6(32'hbbea207f),
	.w7(32'hbbe3375a),
	.w8(32'h3a8efe7a),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a5f86),
	.w1(32'hbbf6d192),
	.w2(32'h39073f2c),
	.w3(32'hbb287974),
	.w4(32'hbb2cd5cc),
	.w5(32'hbb01e855),
	.w6(32'hbb38ebae),
	.w7(32'hbb38e0e7),
	.w8(32'h3bdde2b3),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844a12),
	.w1(32'h3b32a8b5),
	.w2(32'h3c3ba4e2),
	.w3(32'h3c6b7dc9),
	.w4(32'h3b86b954),
	.w5(32'h3c3720d2),
	.w6(32'h3bc43187),
	.w7(32'h3c9491eb),
	.w8(32'h3ba69568),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d8699),
	.w1(32'hbbbf2976),
	.w2(32'hba1442b9),
	.w3(32'hbbb2dc2b),
	.w4(32'hbba7bb70),
	.w5(32'h3afda5b4),
	.w6(32'hbb034070),
	.w7(32'hbb3e4c86),
	.w8(32'h3b104e63),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb6dfa),
	.w1(32'hbba485be),
	.w2(32'h3ab6bbe2),
	.w3(32'hbb48b4fe),
	.w4(32'hbb5bc90d),
	.w5(32'hbbb3d6ad),
	.w6(32'hbb2c4e3c),
	.w7(32'hbba88e83),
	.w8(32'hba9dacab),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5cf7f5),
	.w1(32'hbba901b2),
	.w2(32'hbba1627a),
	.w3(32'hbb1a766f),
	.w4(32'hbb74f557),
	.w5(32'hbb1345bd),
	.w6(32'hb9b8e911),
	.w7(32'hbb1c2091),
	.w8(32'hbb88e504),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50f868),
	.w1(32'h3d7f6e53),
	.w2(32'h3ba080d3),
	.w3(32'hbc32336d),
	.w4(32'hbb8cb58c),
	.w5(32'h3b8ea729),
	.w6(32'hbbd25397),
	.w7(32'h3b9aeb91),
	.w8(32'h3a088a56),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a189a),
	.w1(32'h3b4c882f),
	.w2(32'hba8703f0),
	.w3(32'hbae2d807),
	.w4(32'hbb0d698b),
	.w5(32'hba1f137d),
	.w6(32'hbb25380e),
	.w7(32'hbb95ab2d),
	.w8(32'hbba3b27f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9992deb),
	.w1(32'hbb2db76e),
	.w2(32'hbadcd6f8),
	.w3(32'hbae4eb34),
	.w4(32'hbb5a0e11),
	.w5(32'hbaf15b90),
	.w6(32'h39bf7280),
	.w7(32'h3905458c),
	.w8(32'h3b227989),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b269704),
	.w1(32'hba88608f),
	.w2(32'h3a00f0a3),
	.w3(32'hbba09af1),
	.w4(32'hb89e0b3e),
	.w5(32'hba02c82e),
	.w6(32'hba8b3a00),
	.w7(32'hbb39898b),
	.w8(32'h3c460662),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad43fb8),
	.w1(32'hba7335d7),
	.w2(32'h3c0e94eb),
	.w3(32'h3c7be92e),
	.w4(32'h3a8a8af8),
	.w5(32'h3c257e8b),
	.w6(32'h3bac32aa),
	.w7(32'h3c8479d6),
	.w8(32'h3b3cceb7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0270c2),
	.w1(32'h39d0687d),
	.w2(32'h3be24dbf),
	.w3(32'h3b67de00),
	.w4(32'h37b42c18),
	.w5(32'h3bb671be),
	.w6(32'h398290d7),
	.w7(32'h3be3928f),
	.w8(32'h3adb89c5),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1c33),
	.w1(32'hbbcf4172),
	.w2(32'h3888374c),
	.w3(32'hbb824d0f),
	.w4(32'hbc0fc9c9),
	.w5(32'hbaca2127),
	.w6(32'hbbde4d13),
	.w7(32'hbb14f407),
	.w8(32'hbb7d98c7),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995f45),
	.w1(32'h3cae8ff5),
	.w2(32'hbc58cfc0),
	.w3(32'hbc1a0dbf),
	.w4(32'h3c3d4b7a),
	.w5(32'hbb6d0387),
	.w6(32'h3b6c7a66),
	.w7(32'h3b343894),
	.w8(32'hb9fac731),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3eb6b),
	.w1(32'h39dc1b87),
	.w2(32'h3b809402),
	.w3(32'hbad25612),
	.w4(32'h3997acda),
	.w5(32'h3aae836d),
	.w6(32'h3ae33f01),
	.w7(32'hbb688995),
	.w8(32'h3b799848),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0260c4),
	.w1(32'hbcc6c14f),
	.w2(32'hbc5d6443),
	.w3(32'hb9e13ff5),
	.w4(32'hbc6e2295),
	.w5(32'hbc7dfc60),
	.w6(32'hbb598dca),
	.w7(32'hbc8f52d6),
	.w8(32'hbd1661ad),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f60b6),
	.w1(32'h3d4adc9f),
	.w2(32'hbb0193ab),
	.w3(32'h3b102ef2),
	.w4(32'h3c51d0ae),
	.w5(32'hbcdb32bf),
	.w6(32'h3c271156),
	.w7(32'h3ac9a2f3),
	.w8(32'hbbf342bf),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926a0fb),
	.w1(32'h3b5579d2),
	.w2(32'h3bf5aed7),
	.w3(32'hbacf9f3e),
	.w4(32'h3c0053bb),
	.w5(32'h3c30ae7a),
	.w6(32'h3b6db71d),
	.w7(32'h3bc79ba7),
	.w8(32'h3b943342),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0da33e),
	.w1(32'hbbbb6710),
	.w2(32'h3b89db2d),
	.w3(32'hbadedd41),
	.w4(32'h3a130733),
	.w5(32'h3ad5d1df),
	.w6(32'hbaace22d),
	.w7(32'h3a460772),
	.w8(32'h3ca32c3d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0f60d),
	.w1(32'h3b04df27),
	.w2(32'hbc119de1),
	.w3(32'h3cca1150),
	.w4(32'h3bf2ce61),
	.w5(32'hb919059f),
	.w6(32'h3c9b93cf),
	.w7(32'hbb42adc6),
	.w8(32'hbc151383),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfb184),
	.w1(32'hbc0011df),
	.w2(32'h3bd2c4f2),
	.w3(32'h3ad5bb5b),
	.w4(32'hbb29c4b3),
	.w5(32'h3bc134a4),
	.w6(32'hbb365fa8),
	.w7(32'h399d7cd7),
	.w8(32'hba04e023),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7c4c5),
	.w1(32'hbca4b4ad),
	.w2(32'hbc32ab20),
	.w3(32'hbc2939a8),
	.w4(32'hbbc96d89),
	.w5(32'h3a8aad06),
	.w6(32'hbc5455ff),
	.w7(32'hbc1c8f77),
	.w8(32'h3c9723fe),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c850f09),
	.w1(32'h3b245492),
	.w2(32'hbbb68b86),
	.w3(32'h3c8f6f20),
	.w4(32'h3bccb23b),
	.w5(32'h3b4ca249),
	.w6(32'h3c277160),
	.w7(32'hbb827c92),
	.w8(32'h3c14682f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72c91f),
	.w1(32'h3b62a101),
	.w2(32'hbb0d000e),
	.w3(32'h3c7b923f),
	.w4(32'h3c0a63dd),
	.w5(32'h3bf301ce),
	.w6(32'h3c1168b2),
	.w7(32'hb9404ac2),
	.w8(32'h3b4989a1),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63751b),
	.w1(32'hbcc68f25),
	.w2(32'h3b9585f0),
	.w3(32'hbc41159f),
	.w4(32'h3ba6f258),
	.w5(32'hbc134cdc),
	.w6(32'h3c5982c1),
	.w7(32'h3b99f149),
	.w8(32'hbc4799c4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcadd6e7),
	.w1(32'h3d3cca92),
	.w2(32'h3cd3a316),
	.w3(32'h3b5e7485),
	.w4(32'h3c912456),
	.w5(32'h3bbea4b2),
	.w6(32'h3d1a3ec6),
	.w7(32'hbb40039d),
	.w8(32'hbb215956),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93fdcac),
	.w1(32'h3a71d94b),
	.w2(32'h3aa0793d),
	.w3(32'hbaebea1c),
	.w4(32'hb9f9a3cf),
	.w5(32'hb92d66d4),
	.w6(32'hbaddbf79),
	.w7(32'hb9200881),
	.w8(32'hbb9f7f7b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d4545),
	.w1(32'h3d3e9223),
	.w2(32'h3c46df5b),
	.w3(32'hbb1af3e8),
	.w4(32'h3c31ffd5),
	.w5(32'hbc874d2c),
	.w6(32'hbc06f87b),
	.w7(32'h3c05c20f),
	.w8(32'hba9a4cfb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6170b1),
	.w1(32'hbca8b5f7),
	.w2(32'h3c709817),
	.w3(32'hbc54c1be),
	.w4(32'hb926d2e4),
	.w5(32'h3ca78511),
	.w6(32'hbc05aa1a),
	.w7(32'hbb52f227),
	.w8(32'hba2ec145),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb296d),
	.w1(32'h3c18bd0d),
	.w2(32'hbb8e2add),
	.w3(32'h3bb6952f),
	.w4(32'h3c91c831),
	.w5(32'h3c7f8ca9),
	.w6(32'h39a4d8bc),
	.w7(32'hbb75f646),
	.w8(32'hbbe5905f),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07b7e5),
	.w1(32'h3d1aa052),
	.w2(32'h3c58c1d6),
	.w3(32'hb906f2d0),
	.w4(32'h3b815d37),
	.w5(32'h3b5dcd56),
	.w6(32'h3ce4a119),
	.w7(32'h3c87fe11),
	.w8(32'h3c301598),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f07a2),
	.w1(32'hb9790f03),
	.w2(32'h3beef7dc),
	.w3(32'h3c6a29c9),
	.w4(32'h3b3ba8a5),
	.w5(32'h3c28bc04),
	.w6(32'h3bb07c70),
	.w7(32'h3c8daf55),
	.w8(32'h3b697b7b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b558bd),
	.w1(32'hbc89f617),
	.w2(32'hbb19a123),
	.w3(32'hbb9305a6),
	.w4(32'hbbde245e),
	.w5(32'hba9ed589),
	.w6(32'h39f55133),
	.w7(32'hbbe22abc),
	.w8(32'hbb9577c3),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a904c0c),
	.w1(32'h3b2ddc41),
	.w2(32'hbc4e368b),
	.w3(32'hbc21a734),
	.w4(32'h3908f7fc),
	.w5(32'hbc188f78),
	.w6(32'hbb9e271e),
	.w7(32'hbc9501c2),
	.w8(32'h3a5713ff),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12daac),
	.w1(32'h3ae313c1),
	.w2(32'h3b554f8a),
	.w3(32'hba389585),
	.w4(32'h39431f34),
	.w5(32'h3af63097),
	.w6(32'h398aa413),
	.w7(32'h39c23469),
	.w8(32'h3b657f8e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba4b23c),
	.w1(32'h3b6ac34d),
	.w2(32'h3c737286),
	.w3(32'h3b95a043),
	.w4(32'h3b80fbc3),
	.w5(32'h3c4a680a),
	.w6(32'h3b93959e),
	.w7(32'h3c2bec12),
	.w8(32'hbad1c8e0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf07395),
	.w1(32'hbc703c50),
	.w2(32'hbb1acbad),
	.w3(32'hbc1a0e5d),
	.w4(32'hbba43660),
	.w5(32'hba2a8eb0),
	.w6(32'hbbe0efd9),
	.w7(32'hbbe72b99),
	.w8(32'h3bddac72),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ebd3e),
	.w1(32'h380848c3),
	.w2(32'hbbc0bc97),
	.w3(32'h3c2150ce),
	.w4(32'hb9c2cda3),
	.w5(32'hbb4c53c7),
	.w6(32'h3c043bbb),
	.w7(32'hbb0285ca),
	.w8(32'hbb16853f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba019f27),
	.w1(32'hb88cc100),
	.w2(32'h3a42d921),
	.w3(32'hb8e4aab9),
	.w4(32'hb902fc15),
	.w5(32'hba322cb3),
	.w6(32'h3a51bcf6),
	.w7(32'h398aaa85),
	.w8(32'hba23d2ea),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf47ad),
	.w1(32'hba504c95),
	.w2(32'hba5f701d),
	.w3(32'hba038aaf),
	.w4(32'hb97cfe21),
	.w5(32'hba7a4521),
	.w6(32'hba8e7f29),
	.w7(32'hb9e901b2),
	.w8(32'h3a5980f7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8df4f6),
	.w1(32'hbadb18dc),
	.w2(32'hba802a9e),
	.w3(32'hbabdf604),
	.w4(32'hbb1e3711),
	.w5(32'hbb502d0b),
	.w6(32'h38e10d80),
	.w7(32'hbb01cf41),
	.w8(32'hbb06e2ae),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3992dedc),
	.w1(32'hbaad07de),
	.w2(32'hbafee0b5),
	.w3(32'h3ace13b0),
	.w4(32'hba8a2af5),
	.w5(32'hbba58181),
	.w6(32'h3b17d809),
	.w7(32'hbab4383e),
	.w8(32'hbba91761),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84543e),
	.w1(32'hbb4e9d2f),
	.w2(32'hba9c7a32),
	.w3(32'hba536cc6),
	.w4(32'hbb13903a),
	.w5(32'hbb16c265),
	.w6(32'hb9889320),
	.w7(32'hba80653b),
	.w8(32'hba0c73e9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8024f),
	.w1(32'hbb94a7ef),
	.w2(32'hbb7f1d80),
	.w3(32'hbabd147c),
	.w4(32'hbb2cd586),
	.w5(32'hbb2577c7),
	.w6(32'h3a120fec),
	.w7(32'h39b10b20),
	.w8(32'h3a79b75d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fb46a3),
	.w1(32'hbb20dfa6),
	.w2(32'hbb0b13e4),
	.w3(32'h3adb4a73),
	.w4(32'hba0fc9f3),
	.w5(32'hbb33df16),
	.w6(32'h3b5ad629),
	.w7(32'h38b1aecf),
	.w8(32'hbbdaa50b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9540f),
	.w1(32'hbad08743),
	.w2(32'hbae8ff25),
	.w3(32'hba398ee0),
	.w4(32'hba8fa08a),
	.w5(32'hbabe8f9b),
	.w6(32'hba773a8a),
	.w7(32'hba864dd5),
	.w8(32'hb920533e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d6f7b),
	.w1(32'h3b302dbc),
	.w2(32'h3a5173e2),
	.w3(32'h3b07a819),
	.w4(32'h3a833314),
	.w5(32'hbae296dd),
	.w6(32'h3acbb129),
	.w7(32'h3ab5fee8),
	.w8(32'hbb044d18),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafae5f),
	.w1(32'h3ba8cf60),
	.w2(32'h3b0ce8f8),
	.w3(32'h3b6158e6),
	.w4(32'h3b960625),
	.w5(32'h3b3ff7be),
	.w6(32'h3b680f76),
	.w7(32'h3b839a35),
	.w8(32'h3b2c0495),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5279ee),
	.w1(32'hbb6dfb60),
	.w2(32'h3a2e2121),
	.w3(32'hbabffdf9),
	.w4(32'hbbb8a5f6),
	.w5(32'hbbc48499),
	.w6(32'h3b1e74e4),
	.w7(32'hbbba7539),
	.w8(32'hbbbd0792),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964ccca),
	.w1(32'hbb3dd838),
	.w2(32'hbb76864d),
	.w3(32'hba1a34b7),
	.w4(32'hbb614430),
	.w5(32'hbb1e72a3),
	.w6(32'hba896681),
	.w7(32'hbb102f9f),
	.w8(32'hbbc4a010),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392472aa),
	.w1(32'h3a948ecb),
	.w2(32'hbb2a5f45),
	.w3(32'h399d2d33),
	.w4(32'hb930711a),
	.w5(32'hbb427405),
	.w6(32'h3a0f2f28),
	.w7(32'hba99023a),
	.w8(32'h3ad02203),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a800d34),
	.w1(32'hbb7e22e6),
	.w2(32'hbb2fc42c),
	.w3(32'hb94f6100),
	.w4(32'hba9d052c),
	.w5(32'hba92f8e4),
	.w6(32'hbafac258),
	.w7(32'hbacb0697),
	.w8(32'hb9e24ff0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389c9dee),
	.w1(32'hbbb2f599),
	.w2(32'hbbff0036),
	.w3(32'hb7385a75),
	.w4(32'hbb137c93),
	.w5(32'hbbf4696a),
	.w6(32'h3b80c621),
	.w7(32'hbacd9e31),
	.w8(32'hbbd47684),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d0c02),
	.w1(32'hb9bbaa52),
	.w2(32'h3b129f78),
	.w3(32'h3a62395c),
	.w4(32'h3abb3a69),
	.w5(32'h3b02c1f0),
	.w6(32'h3ac694de),
	.w7(32'h3b06cdf4),
	.w8(32'hba1bb489),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c9f3a),
	.w1(32'hb8a76dcd),
	.w2(32'hb983af5e),
	.w3(32'hb9af1b82),
	.w4(32'hbb5bc488),
	.w5(32'hbb7ab6ef),
	.w6(32'hba62ad6d),
	.w7(32'hb9df967a),
	.w8(32'hbaf3648c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb933a680),
	.w1(32'hbac57e40),
	.w2(32'h37a5d542),
	.w3(32'hb9d663ee),
	.w4(32'hbabeb06e),
	.w5(32'hbb0d2ddb),
	.w6(32'h3a95b9f6),
	.w7(32'hb89bb64b),
	.w8(32'hbb09b114),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac5504a),
	.w1(32'h3a4c9456),
	.w2(32'hba33a21d),
	.w3(32'h3b100ed0),
	.w4(32'hb907a807),
	.w5(32'h39026346),
	.w6(32'h3ac96715),
	.w7(32'h38fd2a1a),
	.w8(32'h390c35dd),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb282c60),
	.w1(32'hbb7f3f6a),
	.w2(32'hb9d056ae),
	.w3(32'h3ab3edb4),
	.w4(32'h3ad71382),
	.w5(32'hb99fa0ad),
	.w6(32'hbb32d5e1),
	.w7(32'hbb6cdf07),
	.w8(32'h39788444),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d115a6),
	.w1(32'hbad90c7e),
	.w2(32'hbaad6ea1),
	.w3(32'hb9d2b46d),
	.w4(32'hba9db6df),
	.w5(32'hba953031),
	.w6(32'h3a189047),
	.w7(32'hb86e8551),
	.w8(32'h3a5c5112),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7adc35),
	.w1(32'hba306045),
	.w2(32'hbb7167fa),
	.w3(32'h3afc76ab),
	.w4(32'hbaab8399),
	.w5(32'hbbaefb0a),
	.w6(32'h3b183e18),
	.w7(32'hbab1396c),
	.w8(32'hbb872dfb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e56e0),
	.w1(32'h3af20294),
	.w2(32'hbb715699),
	.w3(32'h3b5d0293),
	.w4(32'h3a97af64),
	.w5(32'h39cf0772),
	.w6(32'hbb0a81da),
	.w7(32'h3afb894a),
	.w8(32'h3948b775),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdf5b0),
	.w1(32'hba91d936),
	.w2(32'hba38f41f),
	.w3(32'hbab74635),
	.w4(32'hbb102067),
	.w5(32'hbaa485c9),
	.w6(32'hba6c7af8),
	.w7(32'hbb0dc7de),
	.w8(32'hba6f5a3d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafd365),
	.w1(32'hba918c4d),
	.w2(32'hbac6dd21),
	.w3(32'hba29a181),
	.w4(32'hb9f3f8fa),
	.w5(32'hbad4678b),
	.w6(32'h39e68a9d),
	.w7(32'hb993de99),
	.w8(32'hbadb7530),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a928d6f),
	.w1(32'h3a9487e0),
	.w2(32'hbaa0eab9),
	.w3(32'h3ab22a2b),
	.w4(32'h3ad49ec6),
	.w5(32'hba21f0f3),
	.w6(32'h3a9f6d43),
	.w7(32'h3aa46816),
	.w8(32'hbb24f574),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fa9f9),
	.w1(32'hbb17b805),
	.w2(32'hbb7f434b),
	.w3(32'hb9e72a36),
	.w4(32'hbaddd1b3),
	.w5(32'hbb800c27),
	.w6(32'h3a8d6fca),
	.w7(32'hb9d77374),
	.w8(32'h372e3a23),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f091d),
	.w1(32'h39b89b52),
	.w2(32'h3a05e761),
	.w3(32'h39601a96),
	.w4(32'h398a42c9),
	.w5(32'h39a781b4),
	.w6(32'h395dbcb5),
	.w7(32'h39b2fa49),
	.w8(32'h3a0d40d1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d7275),
	.w1(32'hbbbc883c),
	.w2(32'hbb7a1403),
	.w3(32'hbaf5c537),
	.w4(32'hbac33fd3),
	.w5(32'hbb9a4eac),
	.w6(32'h3b5f07ad),
	.w7(32'hbab47a9c),
	.w8(32'hbbb3dbf2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75d5e6),
	.w1(32'h3a89d3b5),
	.w2(32'h3a7632f7),
	.w3(32'h392d8567),
	.w4(32'h39feb4de),
	.w5(32'h3a1f84ec),
	.w6(32'h3a4b2899),
	.w7(32'h3a0a6cbd),
	.w8(32'h3a7d9380),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a8253),
	.w1(32'hbb213b5e),
	.w2(32'hbb125834),
	.w3(32'hbaa8086b),
	.w4(32'hbae7841d),
	.w5(32'hbac8d084),
	.w6(32'hbaee2a7f),
	.w7(32'hbb18acdf),
	.w8(32'hbb52489a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ffb43),
	.w1(32'h3a544d3c),
	.w2(32'h3a534051),
	.w3(32'hb84b9d3a),
	.w4(32'h388c1575),
	.w5(32'h39da28c7),
	.w6(32'h39f9a4a0),
	.w7(32'h37624eb8),
	.w8(32'hbb739af4),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb314f),
	.w1(32'h3b0334b5),
	.w2(32'hbb7e15c2),
	.w3(32'h3b08f923),
	.w4(32'h3a74ed10),
	.w5(32'hbb5a9eba),
	.w6(32'hbb31f2d3),
	.w7(32'hbb277a47),
	.w8(32'hbaa72c2a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393aff81),
	.w1(32'hb8cdd163),
	.w2(32'hb96674cb),
	.w3(32'hb97958bc),
	.w4(32'hb9c2617e),
	.w5(32'hb98869d9),
	.w6(32'hb9197c6b),
	.w7(32'h38c75968),
	.w8(32'h3a10ad7f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae55da),
	.w1(32'hba79bc9d),
	.w2(32'hb9e07add),
	.w3(32'hbb19468c),
	.w4(32'hbaebf613),
	.w5(32'hbac63590),
	.w6(32'h39979bb6),
	.w7(32'hba1fbad1),
	.w8(32'hbb1d8daf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b2ce9),
	.w1(32'h39b83b77),
	.w2(32'h3981c564),
	.w3(32'hb959d017),
	.w4(32'hb8e50f76),
	.w5(32'hb8af56c7),
	.w6(32'h39ada70a),
	.w7(32'h39536fa9),
	.w8(32'h3a18ab9c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cca4b4),
	.w1(32'hbae198d7),
	.w2(32'hb98e0cbc),
	.w3(32'h3932bc3f),
	.w4(32'hbaf9ae28),
	.w5(32'hbb64805a),
	.w6(32'h3b06ba9e),
	.w7(32'hba8d6870),
	.w8(32'hbba6547f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ea239),
	.w1(32'h39e2f441),
	.w2(32'hb9ea9683),
	.w3(32'h395bb337),
	.w4(32'hb9e0e4b0),
	.w5(32'hbb4d5543),
	.w6(32'h3ab3b1d4),
	.w7(32'h3a3ae5a9),
	.w8(32'h3a1b1b77),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994774a),
	.w1(32'h38307d13),
	.w2(32'h38c04e48),
	.w3(32'hb8b4f236),
	.w4(32'h398dd64e),
	.w5(32'h398b2077),
	.w6(32'h3929dd93),
	.w7(32'h39d68603),
	.w8(32'hbad3a27e),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ee7a7),
	.w1(32'hbaa5a2f6),
	.w2(32'hbb8eca58),
	.w3(32'h3a901c39),
	.w4(32'h3a128357),
	.w5(32'hbb17a400),
	.w6(32'hb9d90551),
	.w7(32'hba8e8918),
	.w8(32'h381b03c1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0b66),
	.w1(32'hbb0c3252),
	.w2(32'hba73ea60),
	.w3(32'hbabedad8),
	.w4(32'hbb0f7631),
	.w5(32'hbaeb6f4d),
	.w6(32'hba485390),
	.w7(32'hba6f44ef),
	.w8(32'hbac38e46),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8dcf17),
	.w1(32'hbb918179),
	.w2(32'hbb511970),
	.w3(32'hbae402fc),
	.w4(32'hbbad53ce),
	.w5(32'hbbcace56),
	.w6(32'h39299f62),
	.w7(32'hbb402ef5),
	.w8(32'hbbe36614),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a4c55),
	.w1(32'hba8a576c),
	.w2(32'hbbebfb40),
	.w3(32'hbaba80b3),
	.w4(32'hbba225a5),
	.w5(32'hbbcbaa64),
	.w6(32'hba712a2e),
	.w7(32'hbb4cd732),
	.w8(32'h39b0f955),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dfb37),
	.w1(32'hbbae7e86),
	.w2(32'hbbe4c715),
	.w3(32'hbb2ea107),
	.w4(32'hbc0c32bd),
	.w5(32'hbc55209f),
	.w6(32'hba6c7c3a),
	.w7(32'hbbf863e4),
	.w8(32'hbc19b664),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c83a),
	.w1(32'hbae31e68),
	.w2(32'hba89df30),
	.w3(32'hbaccd6c0),
	.w4(32'hbb7a88cd),
	.w5(32'hbb52deb2),
	.w6(32'h3a7e78b6),
	.w7(32'hbb790bb8),
	.w8(32'hbbcc7207),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa64a6e),
	.w1(32'hbac8b63a),
	.w2(32'hba43e32b),
	.w3(32'hba9650f9),
	.w4(32'hbabd1081),
	.w5(32'hba1e4a56),
	.w6(32'hba9eea21),
	.w7(32'hba947ac0),
	.w8(32'h39ec4385),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88d8a3e),
	.w1(32'hba4099d3),
	.w2(32'h3a084501),
	.w3(32'hb970f89e),
	.w4(32'hba1b1ebb),
	.w5(32'h39419ffc),
	.w6(32'hb9a6bce8),
	.w7(32'h39eafe52),
	.w8(32'hb9131af7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3f51f),
	.w1(32'h3a19f0e2),
	.w2(32'hb9998a7e),
	.w3(32'h3a980c58),
	.w4(32'h37d56c1b),
	.w5(32'h38191f9d),
	.w6(32'h39aa7c67),
	.w7(32'h39d97755),
	.w8(32'hbaab1daf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9654db),
	.w1(32'hba673ca9),
	.w2(32'hb9a92118),
	.w3(32'hba91f139),
	.w4(32'hbac221f5),
	.w5(32'hb9c32c2a),
	.w6(32'h394a3b0f),
	.w7(32'hba71db95),
	.w8(32'hbb204177),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a3fc55),
	.w1(32'hba694bee),
	.w2(32'hba947eb8),
	.w3(32'hba52f2bf),
	.w4(32'hbace2449),
	.w5(32'hba9598a3),
	.w6(32'h395b92e0),
	.w7(32'h3a05ddab),
	.w8(32'hba410137),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8680b6a),
	.w1(32'h38fb61dc),
	.w2(32'hb8623c5a),
	.w3(32'hb8dc0fd9),
	.w4(32'h39517233),
	.w5(32'h3981c5f2),
	.w6(32'h38cff021),
	.w7(32'hba18cd09),
	.w8(32'h3982df69),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96a06e),
	.w1(32'hbaaebf76),
	.w2(32'h3a3aa51b),
	.w3(32'hba5b46c3),
	.w4(32'h3a6d3252),
	.w5(32'h3a68935c),
	.w6(32'hb8df075c),
	.w7(32'h3b0de0eb),
	.w8(32'hb8a2b2d3),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bbaa61),
	.w1(32'hb98c7809),
	.w2(32'hbabbb27e),
	.w3(32'hb92186e7),
	.w4(32'hbaab8252),
	.w5(32'hbb2af3d6),
	.w6(32'hb60f0b6f),
	.w7(32'hbac07f53),
	.w8(32'hbaf01ab4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0895d),
	.w1(32'hbb6f6d93),
	.w2(32'hbb830df4),
	.w3(32'h3acbfcf7),
	.w4(32'hba3ea1e5),
	.w5(32'hbb29029b),
	.w6(32'h3b12dbbd),
	.w7(32'h3b2042a7),
	.w8(32'h381c0be8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c007d),
	.w1(32'hbaa0f988),
	.w2(32'hba2e52ce),
	.w3(32'hbabfbee8),
	.w4(32'hbb2c1f8a),
	.w5(32'hbb2d89fb),
	.w6(32'h37ca927d),
	.w7(32'hbb196ccf),
	.w8(32'hb965340a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e54ea),
	.w1(32'hbb603427),
	.w2(32'hbbe80e14),
	.w3(32'hbb11e9e1),
	.w4(32'hbbd8694f),
	.w5(32'hbc287db1),
	.w6(32'h3b49da09),
	.w7(32'hbb162e20),
	.w8(32'hbc0e7545),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c24b20),
	.w1(32'hbb213362),
	.w2(32'hbb20248f),
	.w3(32'hbada9197),
	.w4(32'hbb4e5217),
	.w5(32'hbb05ba2b),
	.w6(32'h39aeb059),
	.w7(32'h3a7fe80e),
	.w8(32'h3a0f35b0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e64bd),
	.w1(32'h3ab3a39c),
	.w2(32'h3b03beb8),
	.w3(32'h393ec7fc),
	.w4(32'h3a14b368),
	.w5(32'h3a1619df),
	.w6(32'h3a972f64),
	.w7(32'h3ae00a42),
	.w8(32'h3959e2c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f205fc),
	.w1(32'hba1edbfe),
	.w2(32'h39d9773f),
	.w3(32'hba3681d8),
	.w4(32'hb9e3a956),
	.w5(32'h39375e57),
	.w6(32'hb89f6498),
	.w7(32'h39c9baae),
	.w8(32'hb9e46ac8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf8805),
	.w1(32'hbacb3528),
	.w2(32'hbad5b4c7),
	.w3(32'hb9864ad1),
	.w4(32'hbac13654),
	.w5(32'hbaa99c32),
	.w6(32'hba362147),
	.w7(32'hba61a336),
	.w8(32'hb93f4d63),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c6419d),
	.w1(32'hb918cec9),
	.w2(32'hba28dec5),
	.w3(32'hb901b53c),
	.w4(32'hb9feae6e),
	.w5(32'hba6fafb6),
	.w6(32'hb880c1d0),
	.w7(32'hba50c0a0),
	.w8(32'hba4f8cc3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fe1ff),
	.w1(32'h3a2d2699),
	.w2(32'h3ab32360),
	.w3(32'hba2071cc),
	.w4(32'hb9893e53),
	.w5(32'hba03f971),
	.w6(32'h3a31995a),
	.w7(32'h3a679042),
	.w8(32'hb76adc36),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf46b6b),
	.w1(32'hbaf30c7b),
	.w2(32'hbafd7d3f),
	.w3(32'hbb08f5d9),
	.w4(32'hbab0a04a),
	.w5(32'hba476427),
	.w6(32'hbafb9e3e),
	.w7(32'hbb2c760d),
	.w8(32'hbb0bf5b9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba002f98),
	.w1(32'hb9235065),
	.w2(32'hb8f62b58),
	.w3(32'hb9f0b88c),
	.w4(32'h3999ff2b),
	.w5(32'h39cb9795),
	.w6(32'hba16288e),
	.w7(32'h3978b979),
	.w8(32'hb9a43ba3),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a52d6),
	.w1(32'hbb845a52),
	.w2(32'hbb54a61e),
	.w3(32'hbb4e57e2),
	.w4(32'hbb6c1810),
	.w5(32'hbba921a1),
	.w6(32'hbb37a592),
	.w7(32'hbb8aaa2c),
	.w8(32'hbb49062a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb188b82),
	.w1(32'hb9a6a296),
	.w2(32'hb9d0f1fb),
	.w3(32'hba566d7e),
	.w4(32'hbae80880),
	.w5(32'hbb9c12bc),
	.w6(32'h3b64e7dc),
	.w7(32'h3a6ffa22),
	.w8(32'hbbbf017e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabac53f),
	.w1(32'hba066db3),
	.w2(32'hba0f9bae),
	.w3(32'hbaade6f6),
	.w4(32'hba29f8c5),
	.w5(32'hba78790f),
	.w6(32'hbaca05c7),
	.w7(32'hba039f32),
	.w8(32'hba9ca1be),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a828c),
	.w1(32'h3a81a2ca),
	.w2(32'h3acc7a23),
	.w3(32'h3a99532b),
	.w4(32'h3af6bedb),
	.w5(32'h3b08ef0d),
	.w6(32'hb9e1dd72),
	.w7(32'h3a57754d),
	.w8(32'h39cc0b30),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bbb23),
	.w1(32'h3ab34ccd),
	.w2(32'hbae5124d),
	.w3(32'h3b00fe8a),
	.w4(32'h3a889af1),
	.w5(32'hba64ef3b),
	.w6(32'h3a815c00),
	.w7(32'hba95686d),
	.w8(32'hbbdb3e48),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05eb73),
	.w1(32'h3b73f34d),
	.w2(32'hbb1b00be),
	.w3(32'hbb9893f3),
	.w4(32'hbb3f5ff4),
	.w5(32'hba28167b),
	.w6(32'h38c56e01),
	.w7(32'h3aa2b77b),
	.w8(32'h3ab7cfa6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ff627),
	.w1(32'hbb53263f),
	.w2(32'hbb250d40),
	.w3(32'hbb0465a3),
	.w4(32'hba92374c),
	.w5(32'hba3a1c38),
	.w6(32'hbad01e72),
	.w7(32'hba90af8a),
	.w8(32'h3a67a745),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059c74),
	.w1(32'h3b28332b),
	.w2(32'h3b06c2a6),
	.w3(32'h3a852839),
	.w4(32'h3b258efa),
	.w5(32'h3aaf9faf),
	.w6(32'h3af4a0e5),
	.w7(32'h3af3371d),
	.w8(32'h3b12346f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d71c4),
	.w1(32'hb8b044f1),
	.w2(32'h39fb3859),
	.w3(32'h399e1ca1),
	.w4(32'h3a53b921),
	.w5(32'h3ab853de),
	.w6(32'hba12423d),
	.w7(32'h39c37395),
	.w8(32'hb9b8161b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ada90d),
	.w1(32'h396024fc),
	.w2(32'hb83be0f0),
	.w3(32'h3a6a6627),
	.w4(32'hb9e155f0),
	.w5(32'hba6f294c),
	.w6(32'h3938a24f),
	.w7(32'hb98c9994),
	.w8(32'hbae472a7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a5e9d0),
	.w1(32'hb9b52061),
	.w2(32'hb9c9f595),
	.w3(32'h38ef764c),
	.w4(32'hb94945e8),
	.w5(32'hba701a13),
	.w6(32'hba04a182),
	.w7(32'h393a4b7f),
	.w8(32'hbb155289),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47ed8a),
	.w1(32'hbb17368c),
	.w2(32'hbb2c24a0),
	.w3(32'hbb8b2e39),
	.w4(32'hbb7670a5),
	.w5(32'hbb1f7e3e),
	.w6(32'h3acd6c18),
	.w7(32'hbae42ebf),
	.w8(32'h3b570701),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e3263),
	.w1(32'h3b28b2ed),
	.w2(32'h3a957c64),
	.w3(32'h3b3daf77),
	.w4(32'h39af24ff),
	.w5(32'hbb348bbf),
	.w6(32'h3b79bb0c),
	.w7(32'h3a972112),
	.w8(32'hbb3c6054),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92cdf46),
	.w1(32'hba3c75eb),
	.w2(32'hbab822a6),
	.w3(32'hba80b702),
	.w4(32'hb8662873),
	.w5(32'hb807aff7),
	.w6(32'hb844a535),
	.w7(32'h3b536f83),
	.w8(32'hba6ac7f8),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4ff20),
	.w1(32'hbac7dd64),
	.w2(32'hb88d79e9),
	.w3(32'hb9a35ce0),
	.w4(32'hbb02cacf),
	.w5(32'h3a971f76),
	.w6(32'hba082df1),
	.w7(32'hb9d328b2),
	.w8(32'hba5348fe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a844f47),
	.w1(32'h3ad54708),
	.w2(32'hbb08ac69),
	.w3(32'h39ebbf92),
	.w4(32'hbb009289),
	.w5(32'hbb0f2ef2),
	.w6(32'h3b5d25fd),
	.w7(32'h398dda41),
	.w8(32'h3b2a766d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5181bd),
	.w1(32'hb8e4cb76),
	.w2(32'h3afda841),
	.w3(32'h3a909270),
	.w4(32'h3b2bee7e),
	.w5(32'h3aa70704),
	.w6(32'h3b44891c),
	.w7(32'h3a01a76b),
	.w8(32'hbaca016b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49bcf4),
	.w1(32'hb86236ee),
	.w2(32'h38c49760),
	.w3(32'hb962a357),
	.w4(32'h3a3e1f07),
	.w5(32'h3a31fc3e),
	.w6(32'h3a475bba),
	.w7(32'h3a02d5c5),
	.w8(32'hbae41122),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395760b8),
	.w1(32'h3b3ea788),
	.w2(32'hba412f6d),
	.w3(32'hba5bcbdc),
	.w4(32'h3a307a0f),
	.w5(32'hbaec86a5),
	.w6(32'h39902c72),
	.w7(32'hba43050a),
	.w8(32'h3ac1714b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ab1fa),
	.w1(32'h3c7a3685),
	.w2(32'h3be9a36c),
	.w3(32'h3bb7871a),
	.w4(32'h3b348973),
	.w5(32'hba664870),
	.w6(32'h3b314649),
	.w7(32'h3bb72ca7),
	.w8(32'hb9a8df1a),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98eea04),
	.w1(32'hb9cca6b2),
	.w2(32'hba860b31),
	.w3(32'hb9b0e526),
	.w4(32'h3b0ba77b),
	.w5(32'h3a37ff77),
	.w6(32'h39ce94cf),
	.w7(32'hba54bac9),
	.w8(32'hba13a946),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47207),
	.w1(32'h3ac8fc3b),
	.w2(32'h3aba1d0d),
	.w3(32'h3b3e1d29),
	.w4(32'h3af8fa23),
	.w5(32'h3a3f0502),
	.w6(32'h3a4a77cf),
	.w7(32'h3abff711),
	.w8(32'h3996b2b9),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb56fdd0),
	.w1(32'hbbd81854),
	.w2(32'hbb874436),
	.w3(32'hbb9d75da),
	.w4(32'hbb84e0f9),
	.w5(32'hbba53b16),
	.w6(32'h3b8fb9ad),
	.w7(32'h38e04eb6),
	.w8(32'hbab88ecd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule