module layer_10_featuremap_215(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828443f),
	.w1(32'h394fcc9f),
	.w2(32'h3a36d74c),
	.w3(32'h380383b7),
	.w4(32'h397d6169),
	.w5(32'h39e53436),
	.w6(32'h396b706c),
	.w7(32'h39736ec7),
	.w8(32'h39430329),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a5e59),
	.w1(32'h39ed3fd7),
	.w2(32'h3a900447),
	.w3(32'h38376b83),
	.w4(32'h3a7e26c0),
	.w5(32'h3ad4ec6e),
	.w6(32'h39540391),
	.w7(32'h3aed6ea4),
	.w8(32'h3b307dc6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e579b),
	.w1(32'hb9855e9f),
	.w2(32'hb91f5234),
	.w3(32'hb8854c6c),
	.w4(32'h380db7a5),
	.w5(32'hb8df9bc3),
	.w6(32'hb803cb4f),
	.w7(32'hb959bb4d),
	.w8(32'hb9375699),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894bf9f),
	.w1(32'hba869bfd),
	.w2(32'hba8727cb),
	.w3(32'h3a24877c),
	.w4(32'hba017610),
	.w5(32'hb95a4b80),
	.w6(32'hbb07e8cf),
	.w7(32'hbad3d03a),
	.w8(32'h381293a0),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97621ae),
	.w1(32'h3a068154),
	.w2(32'h39a13b4b),
	.w3(32'h38b65084),
	.w4(32'h39c432f2),
	.w5(32'h393d114c),
	.w6(32'h39eb1b6e),
	.w7(32'h39def3d7),
	.w8(32'h39b5fcc0),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d139cc),
	.w1(32'h396a05fd),
	.w2(32'h37468cf9),
	.w3(32'h39c997aa),
	.w4(32'h3983bc01),
	.w5(32'h391a2d0a),
	.w6(32'h396ef711),
	.w7(32'h38df3651),
	.w8(32'h3907cd6f),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e47e34),
	.w1(32'hbb605506),
	.w2(32'h3af3b2f4),
	.w3(32'hbaac019c),
	.w4(32'hbb1521ef),
	.w5(32'h3b3abd2a),
	.w6(32'hbb066ef8),
	.w7(32'hbad4d1e3),
	.w8(32'h3b1d0760),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50204d),
	.w1(32'hbabe77fa),
	.w2(32'hb9911255),
	.w3(32'h3b5f8666),
	.w4(32'hbadddbeb),
	.w5(32'h38dd1f39),
	.w6(32'hbba71199),
	.w7(32'hb857e054),
	.w8(32'hbb86c052),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d0689),
	.w1(32'hb9addfbd),
	.w2(32'h38b43814),
	.w3(32'hb9ea5aed),
	.w4(32'hb99a0827),
	.w5(32'hb911e0c2),
	.w6(32'h38ac7925),
	.w7(32'h37f0ec7c),
	.w8(32'hb7902d25),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98f2940),
	.w1(32'h3a1e5043),
	.w2(32'h3b969fff),
	.w3(32'h3ac65497),
	.w4(32'h3a5ee3e4),
	.w5(32'h3b0b6cc1),
	.w6(32'hba803812),
	.w7(32'hbaa5838f),
	.w8(32'h3b5bd082),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30a86b),
	.w1(32'hb9a95842),
	.w2(32'hba41f7b4),
	.w3(32'hb9dd4006),
	.w4(32'hb9a6817e),
	.w5(32'hba302e29),
	.w6(32'hb9c89fe2),
	.w7(32'hb9e011d1),
	.w8(32'hba457f1d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90a952),
	.w1(32'hbbbd7df8),
	.w2(32'h3a8c4d62),
	.w3(32'h3a4e1175),
	.w4(32'hbb8100f5),
	.w5(32'h3b33b3ca),
	.w6(32'hbb69b448),
	.w7(32'hbba9a2a9),
	.w8(32'h3b158a00),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6739b8),
	.w1(32'hba802f7e),
	.w2(32'h3b1ae079),
	.w3(32'hba344563),
	.w4(32'hbb0fac6b),
	.w5(32'hb806068b),
	.w6(32'hbb4a7841),
	.w7(32'hbb63c85c),
	.w8(32'hb7b66838),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab80a56),
	.w1(32'hb833a628),
	.w2(32'h3a2cc687),
	.w3(32'h35f2ef88),
	.w4(32'h3aebbc76),
	.w5(32'h3aaa38cf),
	.w6(32'hb9b595fb),
	.w7(32'h3ad7491d),
	.w8(32'h3a56ffbe),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9981e6c),
	.w1(32'h3a8fa3c2),
	.w2(32'h3b240810),
	.w3(32'hba6571b3),
	.w4(32'hb945ed35),
	.w5(32'h3ad7baaa),
	.w6(32'h39288295),
	.w7(32'h3ae83fda),
	.w8(32'h3b5808f6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa315de),
	.w1(32'h3b20401f),
	.w2(32'h3bb4b235),
	.w3(32'h3a593cf4),
	.w4(32'h3aea5cbe),
	.w5(32'h3b0bfe8c),
	.w6(32'h3a8f7176),
	.w7(32'h3b1e03cc),
	.w8(32'h3b48dc4b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397b1da2),
	.w1(32'h39cf4d11),
	.w2(32'hb630ab3e),
	.w3(32'h39b6c7dc),
	.w4(32'h39d4d16e),
	.w5(32'hb9c43a4b),
	.w6(32'h39bd2628),
	.w7(32'h39ecda61),
	.w8(32'hb82664cf),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e8529),
	.w1(32'hbad9824a),
	.w2(32'h3b7a4fe9),
	.w3(32'hbb3d58ae),
	.w4(32'hbb993c9a),
	.w5(32'h3b454471),
	.w6(32'hbbf2d809),
	.w7(32'hbb8f7c80),
	.w8(32'hbb27b90d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7e55b),
	.w1(32'hbb0240a5),
	.w2(32'h3ac76c66),
	.w3(32'hbac02444),
	.w4(32'hbb129a96),
	.w5(32'h39d191e6),
	.w6(32'hbb5ba1e3),
	.w7(32'hbb5fd1a5),
	.w8(32'hbad4c6b9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b2eb1b),
	.w1(32'hb8efd577),
	.w2(32'hb70d3c3c),
	.w3(32'hb9357ccf),
	.w4(32'hb8fee613),
	.w5(32'hb956cd0a),
	.w6(32'hb890920c),
	.w7(32'hb8f28a15),
	.w8(32'hb9012df5),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c03ea),
	.w1(32'hb7c6b140),
	.w2(32'hb8165cb5),
	.w3(32'hb8b7dcda),
	.w4(32'hb8568122),
	.w5(32'h381e4d57),
	.w6(32'hb90dec89),
	.w7(32'hb95838eb),
	.w8(32'hb9062993),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c6a4c),
	.w1(32'hb9e09161),
	.w2(32'h3997388c),
	.w3(32'hb9b0fe84),
	.w4(32'hb96547cb),
	.w5(32'h3a3a2984),
	.w6(32'h39c70ce3),
	.w7(32'h37c13977),
	.w8(32'h39978c48),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47840f),
	.w1(32'hbb3fb919),
	.w2(32'h3bf61192),
	.w3(32'hbaaced60),
	.w4(32'hbbccdd6e),
	.w5(32'h3bb3f48e),
	.w6(32'hbbee85ca),
	.w7(32'hbbd53c2b),
	.w8(32'h3bbd55fd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c548c7),
	.w1(32'h387c3be1),
	.w2(32'h3b3b1b20),
	.w3(32'h3a4d27e1),
	.w4(32'hbade7d4a),
	.w5(32'hba9de8e0),
	.w6(32'hbae6ed50),
	.w7(32'hbb090b1d),
	.w8(32'h3a584e69),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa9137a),
	.w1(32'hbabe4986),
	.w2(32'h39d19153),
	.w3(32'h3a6c661e),
	.w4(32'hba91ee6e),
	.w5(32'hba51e09b),
	.w6(32'h3af76532),
	.w7(32'h3aacee57),
	.w8(32'h3b432d74),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ae6829),
	.w1(32'hb8b30fe7),
	.w2(32'h37a6d74a),
	.w3(32'h38859413),
	.w4(32'h383393f7),
	.w5(32'h39485960),
	.w6(32'h39c49f52),
	.w7(32'h39cec3f4),
	.w8(32'h39c91266),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91b6312),
	.w1(32'hb940c6c0),
	.w2(32'hb94b0f1b),
	.w3(32'hb91bbb3a),
	.w4(32'hb9252895),
	.w5(32'hb9750466),
	.w6(32'hb91b96a0),
	.w7(32'hb9611463),
	.w8(32'hb981ea3a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b723092),
	.w1(32'hbab190d0),
	.w2(32'h39ec48a6),
	.w3(32'h3baaac89),
	.w4(32'h3a5ff85a),
	.w5(32'h3a89095f),
	.w6(32'h3c0fcd51),
	.w7(32'h3b1a441f),
	.w8(32'h3b360d14),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d319a),
	.w1(32'hbb03934f),
	.w2(32'hbb0c3541),
	.w3(32'hb98063b3),
	.w4(32'hba9d6593),
	.w5(32'hba97972c),
	.w6(32'h39b7b038),
	.w7(32'hba857552),
	.w8(32'hba5bd605),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8fb70),
	.w1(32'h3a4a47e8),
	.w2(32'h3b410468),
	.w3(32'h3b8b5ca6),
	.w4(32'h3aeb1639),
	.w5(32'h3b38c176),
	.w6(32'h3ba77f8f),
	.w7(32'h3b632a13),
	.w8(32'h3b920fb2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390efb64),
	.w1(32'hb810faa2),
	.w2(32'h366bfd46),
	.w3(32'h38b459d7),
	.w4(32'h35ba3282),
	.w5(32'hb5fe6699),
	.w6(32'hb78bfc2c),
	.w7(32'hb8aeb6b8),
	.w8(32'hb7952a03),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37dbad32),
	.w1(32'h378d2e3a),
	.w2(32'h37de2224),
	.w3(32'h3756a798),
	.w4(32'h37c1a4a6),
	.w5(32'hb81d4a2a),
	.w6(32'h389cf165),
	.w7(32'h380948a0),
	.w8(32'hb7e2fc02),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dc7d94),
	.w1(32'h39add06d),
	.w2(32'h3b1624dc),
	.w3(32'h390e6d35),
	.w4(32'h3a0888c0),
	.w5(32'h3ac24c7d),
	.w6(32'hba2e0a21),
	.w7(32'hb968b462),
	.w8(32'h3ac9d708),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22e50e),
	.w1(32'h39cb62d5),
	.w2(32'h3a0aeaa5),
	.w3(32'h39dc5a33),
	.w4(32'h38bff544),
	.w5(32'h3a4e0c73),
	.w6(32'h3a725d71),
	.w7(32'h3a9f0c0d),
	.w8(32'h3ad6cde7),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad3923),
	.w1(32'hb9632f83),
	.w2(32'h390b69e0),
	.w3(32'hb9fce35e),
	.w4(32'hb7a4adc3),
	.w5(32'h37e1578a),
	.w6(32'h3877da45),
	.w7(32'hb8be0354),
	.w8(32'h3a475aa8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885f259),
	.w1(32'hbad5f056),
	.w2(32'h3a1315d8),
	.w3(32'hba0780f6),
	.w4(32'hba8d4de1),
	.w5(32'h38ce8d3a),
	.w6(32'hbb17c9ca),
	.w7(32'hbb10abb9),
	.w8(32'hba754a99),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c99bc),
	.w1(32'hbc2c7dd8),
	.w2(32'h3b528bef),
	.w3(32'h3ba02ee2),
	.w4(32'hbbb99484),
	.w5(32'h3b42b459),
	.w6(32'hbadbb428),
	.w7(32'hbba81750),
	.w8(32'h3b56b478),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3758cb),
	.w1(32'hbb2368ca),
	.w2(32'hbafffbb1),
	.w3(32'h3ae16664),
	.w4(32'hb9b49a74),
	.w5(32'h39fe2ad1),
	.w6(32'h3bb2fd8f),
	.w7(32'h3b15f3d7),
	.w8(32'h3bb20736),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8e08a),
	.w1(32'hbab98558),
	.w2(32'hba1c461b),
	.w3(32'h3b8b2c53),
	.w4(32'h3b0acbb1),
	.w5(32'h3b1a0a2a),
	.w6(32'h3bb38f6a),
	.w7(32'h3b7a1a22),
	.w8(32'h3babf758),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72590a4),
	.w1(32'hba4b4a13),
	.w2(32'hba16c257),
	.w3(32'h3822e7cb),
	.w4(32'hb9e4dbd7),
	.w5(32'hb995578f),
	.w6(32'h3a0a5286),
	.w7(32'h39914929),
	.w8(32'h3a243217),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bacad1),
	.w1(32'h39383645),
	.w2(32'h397a1c9e),
	.w3(32'hb9740125),
	.w4(32'h392d19f5),
	.w5(32'h39343464),
	.w6(32'hb9042943),
	.w7(32'h382a2567),
	.w8(32'hb8897143),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392511b4),
	.w1(32'h38c36102),
	.w2(32'hb9547546),
	.w3(32'h392ae59e),
	.w4(32'hb86a1742),
	.w5(32'hb9a6ce4d),
	.w6(32'hb9222e67),
	.w7(32'hb91683ed),
	.w8(32'hb78c9570),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a999e1),
	.w1(32'hba270ae5),
	.w2(32'hb8cce13d),
	.w3(32'hb972437f),
	.w4(32'hba4a9ddf),
	.w5(32'hb8a92fb3),
	.w6(32'hb9419c25),
	.w7(32'hba5eccf5),
	.w8(32'h38dd2906),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377fb03e),
	.w1(32'h3b3e20d1),
	.w2(32'h3baca9bf),
	.w3(32'h3b1bbaaf),
	.w4(32'h3aaa3777),
	.w5(32'h3b3913f4),
	.w6(32'h3b706982),
	.w7(32'h3afda57f),
	.w8(32'h3b1260ff),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe1b7d),
	.w1(32'h39ecf176),
	.w2(32'h3b133b83),
	.w3(32'h3aa70003),
	.w4(32'hb82fcef8),
	.w5(32'h3a8832b1),
	.w6(32'h3ac06b93),
	.w7(32'hb95a59a8),
	.w8(32'h3b1b25c7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb60f5),
	.w1(32'h3a011ae5),
	.w2(32'h3b76d6b5),
	.w3(32'h3ad4f1a4),
	.w4(32'hbabb2a4d),
	.w5(32'h3a7d0810),
	.w6(32'hb90f1ec8),
	.w7(32'hba8f5f6b),
	.w8(32'h3b34e689),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39257fa2),
	.w1(32'h3aa84f82),
	.w2(32'h3b8eca49),
	.w3(32'h3a08125c),
	.w4(32'h363f6d95),
	.w5(32'h3ae93782),
	.w6(32'hb9874876),
	.w7(32'hb98cd2ce),
	.w8(32'h3b0d5d0b),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58d87e),
	.w1(32'hbbddd7fb),
	.w2(32'h3a650b1d),
	.w3(32'hbb62624d),
	.w4(32'hbbdd1311),
	.w5(32'h3897992b),
	.w6(32'hbc54621a),
	.w7(32'hbc479c69),
	.w8(32'hbbcf9c04),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901c8a2),
	.w1(32'h38a5baad),
	.w2(32'h39394347),
	.w3(32'hb7ee5cf8),
	.w4(32'hb8dc5a45),
	.w5(32'hb88263e3),
	.w6(32'hb7cff46d),
	.w7(32'hb8664650),
	.w8(32'hb82a6166),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938fd9c),
	.w1(32'h39bc64cd),
	.w2(32'h3a0bc9ae),
	.w3(32'hb97f15b0),
	.w4(32'hb9926337),
	.w5(32'h390bd297),
	.w6(32'hb95ea752),
	.w7(32'hb918e134),
	.w8(32'hb8a467fa),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382a87c6),
	.w1(32'h3922f5ce),
	.w2(32'hb8a3d812),
	.w3(32'h3893d602),
	.w4(32'h3980a3c5),
	.w5(32'h37b19a05),
	.w6(32'h3917446d),
	.w7(32'hb82fe540),
	.w8(32'hb81ba81d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f02e69),
	.w1(32'h3af8ea2e),
	.w2(32'h3b54f27e),
	.w3(32'h3989af4d),
	.w4(32'h38f23c09),
	.w5(32'h3a890ddb),
	.w6(32'h3a6fcf44),
	.w7(32'h3ae43ad0),
	.w8(32'h3abbe99c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5eda97),
	.w1(32'h3a595e28),
	.w2(32'h3a5a8744),
	.w3(32'h3a11e859),
	.w4(32'hb91f1951),
	.w5(32'h39f25641),
	.w6(32'h39ce8ab3),
	.w7(32'h390d6651),
	.w8(32'hb74770f8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3849decd),
	.w1(32'hbb1d3ecc),
	.w2(32'h3b30ecab),
	.w3(32'h3a99f027),
	.w4(32'hba978cf7),
	.w5(32'h3b1c6b7b),
	.w6(32'hbbdf25d1),
	.w7(32'hbbe8726f),
	.w8(32'hbb5c7aac),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a011cea),
	.w1(32'hba24ee47),
	.w2(32'hb8be1d3b),
	.w3(32'h39d7d413),
	.w4(32'hba0002e0),
	.w5(32'h3927ba54),
	.w6(32'h3a1fde59),
	.w7(32'hb97d02f5),
	.w8(32'hba484c3b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb69f6),
	.w1(32'hb941fb35),
	.w2(32'h3997aad4),
	.w3(32'hb82d330a),
	.w4(32'h38b5521f),
	.w5(32'h393a11d7),
	.w6(32'hb9962a24),
	.w7(32'hb86d8983),
	.w8(32'h37975817),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390837c6),
	.w1(32'hb9b181c5),
	.w2(32'hb9d2fd2b),
	.w3(32'h399060a4),
	.w4(32'hb9131be1),
	.w5(32'hb957661a),
	.w6(32'hb998195a),
	.w7(32'hb9529b18),
	.w8(32'hb8dc9225),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00b8bd),
	.w1(32'h3a166a4a),
	.w2(32'h39ada8d6),
	.w3(32'hb9c839c7),
	.w4(32'h3a0c93a9),
	.w5(32'hb879d2be),
	.w6(32'h3996d7d4),
	.w7(32'h3a23ff11),
	.w8(32'h3a3cc7f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d5df4),
	.w1(32'hb9d7d57d),
	.w2(32'hb8ecbef9),
	.w3(32'h3986a006),
	.w4(32'hb9238ce6),
	.w5(32'h395db6a5),
	.w6(32'h39ae4ae7),
	.w7(32'hb8054bbc),
	.w8(32'h396c1a93),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e5a42f),
	.w1(32'h388be14e),
	.w2(32'h38f5639f),
	.w3(32'h393a0c1c),
	.w4(32'h38971077),
	.w5(32'h384e0b1e),
	.w6(32'h39982bf7),
	.w7(32'h39946164),
	.w8(32'h391bed0b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94bc30),
	.w1(32'hb9aa2a61),
	.w2(32'h3b092339),
	.w3(32'hb9e1fc1b),
	.w4(32'hba3c2686),
	.w5(32'h3a1090ae),
	.w6(32'hbb43ccea),
	.w7(32'hbb0b5757),
	.w8(32'hb9c3e810),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c01c20),
	.w1(32'h3accdcfd),
	.w2(32'h3ac41522),
	.w3(32'h3a7f59c8),
	.w4(32'hba20e610),
	.w5(32'hb93f89d9),
	.w6(32'h3b0055b1),
	.w7(32'hb8d77e05),
	.w8(32'hba4cb1f5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb840e837),
	.w1(32'h39970a7f),
	.w2(32'h3a0d8413),
	.w3(32'hb868a0d1),
	.w4(32'hb8d24f3e),
	.w5(32'h37b0d220),
	.w6(32'h39e25ec3),
	.w7(32'h39862132),
	.w8(32'h394df235),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4b211),
	.w1(32'h3956cf35),
	.w2(32'h3831e095),
	.w3(32'h38419cc6),
	.w4(32'h39e11794),
	.w5(32'h396c78d4),
	.w6(32'h396e5932),
	.w7(32'h391bb868),
	.w8(32'h39853061),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2f0ed),
	.w1(32'hb9265408),
	.w2(32'hb91d1914),
	.w3(32'h3915812f),
	.w4(32'hb824f279),
	.w5(32'hb8bc47b6),
	.w6(32'hb8b2bb09),
	.w7(32'h37294d16),
	.w8(32'h379e526e),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82fc347),
	.w1(32'h39dfaa7d),
	.w2(32'h39863777),
	.w3(32'hb9270edd),
	.w4(32'hb7dca4b3),
	.w5(32'hb98f5f50),
	.w6(32'h3940f868),
	.w7(32'h39d4a9ab),
	.w8(32'h398a380b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f6cb1),
	.w1(32'hba3bb46f),
	.w2(32'h3ba510eb),
	.w3(32'hba8afe9c),
	.w4(32'h3ab33a12),
	.w5(32'h3b12ff4e),
	.w6(32'hbb93a8cf),
	.w7(32'hba97cf2c),
	.w8(32'h3b5212b0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8c8ae),
	.w1(32'h3a21e025),
	.w2(32'h3b70b142),
	.w3(32'hba584506),
	.w4(32'hbab72887),
	.w5(32'h3aec451e),
	.w6(32'hbb338666),
	.w7(32'h38cab283),
	.w8(32'h3b3f184e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a838fed),
	.w1(32'h3b0ff6ee),
	.w2(32'h3b8c5a69),
	.w3(32'h399d3d29),
	.w4(32'hba3f8c33),
	.w5(32'h3b49aa79),
	.w6(32'hba43bc0b),
	.w7(32'hb91d9db7),
	.w8(32'h3afba43f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74908e),
	.w1(32'hbb058aad),
	.w2(32'hba8bd0ad),
	.w3(32'h3b359249),
	.w4(32'hbae95148),
	.w5(32'hbac3512c),
	.w6(32'h3b844cdd),
	.w7(32'h3b21ed0e),
	.w8(32'h3bbc146f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84a49b7),
	.w1(32'hb81a3c8e),
	.w2(32'hb7875fab),
	.w3(32'h37b53dfe),
	.w4(32'h38a8d6a0),
	.w5(32'h37d7e9d6),
	.w6(32'hb881a0a5),
	.w7(32'hb9020edf),
	.w8(32'hb8e74443),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8677e1c),
	.w1(32'h38a4e95e),
	.w2(32'h3845da22),
	.w3(32'hb8cbdc63),
	.w4(32'hb83ef72d),
	.w5(32'hb8ca70b5),
	.w6(32'hb771a5a8),
	.w7(32'hb63a9220),
	.w8(32'hb8ad7a9a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c79bde),
	.w1(32'h39321965),
	.w2(32'h3905cfb7),
	.w3(32'hb60352c3),
	.w4(32'h3822ad7e),
	.w5(32'hb7d22c6d),
	.w6(32'h37a9cf07),
	.w7(32'h38aa8493),
	.w8(32'hb8f38517),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3038cb),
	.w1(32'hba1e7528),
	.w2(32'h3a04f76f),
	.w3(32'hb9b6ee83),
	.w4(32'hba81e85a),
	.w5(32'h3910ecd7),
	.w6(32'hba39c53a),
	.w7(32'hba7d02f6),
	.w8(32'hba0aa0df),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810114c),
	.w1(32'hb8ff642f),
	.w2(32'hb94b0db1),
	.w3(32'hb89b0b2c),
	.w4(32'hb7908d22),
	.w5(32'hb95a1795),
	.w6(32'h3699a7df),
	.w7(32'hb8aaf9b2),
	.w8(32'hb94536b5),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71d99b4),
	.w1(32'hbabff3a0),
	.w2(32'h39fc901f),
	.w3(32'h3a9dc768),
	.w4(32'hbaea2ced),
	.w5(32'h3a5d9c64),
	.w6(32'hbb973877),
	.w7(32'hbbaa8d7b),
	.w8(32'hbb1a7481),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d5433),
	.w1(32'hbb2bd7c8),
	.w2(32'h3b18998c),
	.w3(32'hba08345e),
	.w4(32'hbaf9212d),
	.w5(32'h3ae1e53a),
	.w6(32'hbba016cb),
	.w7(32'hbbaa2ae2),
	.w8(32'hbaaca960),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3af56d),
	.w1(32'hb993dcb7),
	.w2(32'h3a34d91a),
	.w3(32'h39b35fd9),
	.w4(32'hb9e8e97f),
	.w5(32'hb9891353),
	.w6(32'h3aa285a9),
	.w7(32'hba291719),
	.w8(32'h3a0c771d),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab9dc6),
	.w1(32'h386770e0),
	.w2(32'h3aa7e9e2),
	.w3(32'h3a28bb3a),
	.w4(32'h3a35a470),
	.w5(32'h3abd9cf6),
	.w6(32'h3a0347c1),
	.w7(32'h3a09022b),
	.w8(32'h3a99ad6c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ecde1),
	.w1(32'hbb1258ac),
	.w2(32'h3b0673e4),
	.w3(32'hba85b49f),
	.w4(32'hbaeee6a2),
	.w5(32'h39281d64),
	.w6(32'hbabe0cc5),
	.w7(32'hba99069a),
	.w8(32'h3b03c7d9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f82a3a),
	.w1(32'h3a3772cf),
	.w2(32'h3a80a807),
	.w3(32'h3a0744b1),
	.w4(32'h395dbc51),
	.w5(32'h39e49b94),
	.w6(32'h3a83eb56),
	.w7(32'h394736da),
	.w8(32'h3a80341a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39985c57),
	.w1(32'hbaa0462e),
	.w2(32'h3a6af664),
	.w3(32'hba0432bc),
	.w4(32'hbac7b25a),
	.w5(32'h39d920dc),
	.w6(32'hbb126174),
	.w7(32'hbb713bab),
	.w8(32'hbafa4fbb),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb967ac83),
	.w1(32'hb90ca42c),
	.w2(32'hb939ec52),
	.w3(32'hb9adba83),
	.w4(32'h32d81288),
	.w5(32'hb922aa12),
	.w6(32'hb8bdfefe),
	.w7(32'hb92066df),
	.w8(32'hb9255651),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb901be0d),
	.w1(32'h37cf885b),
	.w2(32'h383a1699),
	.w3(32'hb89adc9c),
	.w4(32'h3796f78d),
	.w5(32'hb72ef286),
	.w6(32'h3905acb9),
	.w7(32'hb848bc31),
	.w8(32'hb8cbd116),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38761daf),
	.w1(32'hb91a52c2),
	.w2(32'hb7f434da),
	.w3(32'hb8c0a00e),
	.w4(32'hb8fa7a76),
	.w5(32'hb9061b29),
	.w6(32'h3a48301e),
	.w7(32'h34efd21d),
	.w8(32'h390abf26),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391dcf9c),
	.w1(32'hb9751739),
	.w2(32'hb90b7bbe),
	.w3(32'h38488386),
	.w4(32'h39207206),
	.w5(32'h398a5632),
	.w6(32'h39368305),
	.w7(32'h38c9d24e),
	.w8(32'h3984f39d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1da59),
	.w1(32'hb9a7d01d),
	.w2(32'hb7c7f49d),
	.w3(32'h3afa4bbf),
	.w4(32'h39b34d8f),
	.w5(32'h39e7a694),
	.w6(32'h3b326bcf),
	.w7(32'h3afaf478),
	.w8(32'h3b1a9af3),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb897ef9c),
	.w1(32'hba3087e9),
	.w2(32'hb8c20fac),
	.w3(32'hb9adbc6e),
	.w4(32'hba147e5c),
	.w5(32'h38c2b1d6),
	.w6(32'h3960a87b),
	.w7(32'hb9a8d22e),
	.w8(32'h397720d5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82d2cc),
	.w1(32'h39321a5b),
	.w2(32'h3a0cc88d),
	.w3(32'h398a2359),
	.w4(32'hb95feb9c),
	.w5(32'h392887a4),
	.w6(32'h39639af9),
	.w7(32'h3a1384e0),
	.w8(32'h3a97ac83),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38458621),
	.w1(32'h3801bc56),
	.w2(32'h3b953a06),
	.w3(32'h3aba49de),
	.w4(32'h39237d43),
	.w5(32'h3b8cea38),
	.w6(32'hbb60c77a),
	.w7(32'hbb71640b),
	.w8(32'h3a13a1f4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad5d13),
	.w1(32'hbae2de0d),
	.w2(32'hbaa9e608),
	.w3(32'h3a8dc978),
	.w4(32'hbae3254a),
	.w5(32'h37d0c88e),
	.w6(32'h3adf9131),
	.w7(32'hbaea2648),
	.w8(32'h3901608d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaac57),
	.w1(32'hbb964672),
	.w2(32'h3b7b1262),
	.w3(32'h3ae188b4),
	.w4(32'hba8e553b),
	.w5(32'h3b6859cf),
	.w6(32'hbba0c0dc),
	.w7(32'hba28d15f),
	.w8(32'h3bdf10ad),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a276b),
	.w1(32'hba0a477c),
	.w2(32'hba9d1a7a),
	.w3(32'h39ca9f37),
	.w4(32'h39fa7c8d),
	.w5(32'h388714a7),
	.w6(32'h3a4023a5),
	.w7(32'h3a3b6248),
	.w8(32'h3add0c24),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd0412),
	.w1(32'h3a8b5c74),
	.w2(32'h3baa7eee),
	.w3(32'h3a77593f),
	.w4(32'h3acc7450),
	.w5(32'h3b868fe0),
	.w6(32'hbabc2e7c),
	.w7(32'h3a179092),
	.w8(32'h3b5ace29),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6cd0a),
	.w1(32'h38bb66f1),
	.w2(32'h3a98077d),
	.w3(32'hb981c9f6),
	.w4(32'h394c0140),
	.w5(32'h3a10e708),
	.w6(32'h3a61fc02),
	.w7(32'h3a44298a),
	.w8(32'h3b434072),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb6dbe),
	.w1(32'h3a832c65),
	.w2(32'h3a6ca42b),
	.w3(32'h3a032abb),
	.w4(32'h3a05f638),
	.w5(32'h3afe7a2c),
	.w6(32'h3b5e02d9),
	.w7(32'h3b151917),
	.w8(32'h3b61765b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f7fa3),
	.w1(32'h38ed1b72),
	.w2(32'h3a016724),
	.w3(32'h3a136b3c),
	.w4(32'hb856aa7b),
	.w5(32'h388e0b00),
	.w6(32'h3999c8ae),
	.w7(32'h3991bb78),
	.w8(32'h3a364ee1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f982d),
	.w1(32'hb8b25890),
	.w2(32'h3bb8d4e9),
	.w3(32'hba0463e3),
	.w4(32'hbad816fa),
	.w5(32'h3b49dd80),
	.w6(32'hbb3a0713),
	.w7(32'hbb15bf9d),
	.w8(32'h3ae27917),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9eab7),
	.w1(32'hba278713),
	.w2(32'h3bb293e8),
	.w3(32'h396412ca),
	.w4(32'hbac2c2fe),
	.w5(32'h3a67ccac),
	.w6(32'hbbaf1c55),
	.w7(32'hbb5d050c),
	.w8(32'h3b1a4685),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac848ef),
	.w1(32'hbb73daeb),
	.w2(32'h3b3cfa3b),
	.w3(32'h3b1b43d9),
	.w4(32'hba44db89),
	.w5(32'h3b036951),
	.w6(32'hbbc9806e),
	.w7(32'hbbda8aae),
	.w8(32'hba860dfb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49eec1),
	.w1(32'hba89a3bf),
	.w2(32'h3a23d1e4),
	.w3(32'h3aff30d5),
	.w4(32'hba8593b3),
	.w5(32'hb910d3d2),
	.w6(32'h3bc7fca3),
	.w7(32'h3b0da8b9),
	.w8(32'h3bb2ee0b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe7702),
	.w1(32'h3abe6e50),
	.w2(32'h3b392058),
	.w3(32'h3a9e89b1),
	.w4(32'hba4bb3b6),
	.w5(32'hba6f153a),
	.w6(32'h39b6b514),
	.w7(32'h3a8204e9),
	.w8(32'h3b3eece3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39085717),
	.w1(32'hbb9f3492),
	.w2(32'h3b486d7c),
	.w3(32'h3b21130c),
	.w4(32'hbb5e0c38),
	.w5(32'h3a87bf17),
	.w6(32'hbc0406c5),
	.w7(32'hbbc8b311),
	.w8(32'hba02461d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a266dfe),
	.w1(32'h3a64e462),
	.w2(32'h3a269100),
	.w3(32'h3a417b61),
	.w4(32'h394f843f),
	.w5(32'hb90bbe22),
	.w6(32'h3a7d57e8),
	.w7(32'h3a26f2f2),
	.w8(32'h39949c46),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c8413),
	.w1(32'hbb635539),
	.w2(32'h3b187297),
	.w3(32'h3afe2c97),
	.w4(32'hbbea7b2e),
	.w5(32'h3aa27bba),
	.w6(32'hbc22d247),
	.w7(32'hbc66896c),
	.w8(32'hb96ff76b),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3688a4),
	.w1(32'hba9b6a4c),
	.w2(32'hba39cd3f),
	.w3(32'h3b11077b),
	.w4(32'h3a8f210b),
	.w5(32'hb95c43bb),
	.w6(32'hbac9ee1c),
	.w7(32'hba19da7c),
	.w8(32'h3a81fc9f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c67f2),
	.w1(32'hb93d1fd6),
	.w2(32'hb9a6a783),
	.w3(32'hb9176c2f),
	.w4(32'h387af02a),
	.w5(32'hb94c88c8),
	.w6(32'h39de92c0),
	.w7(32'h357f29fc),
	.w8(32'hb964fa7d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac153ff),
	.w1(32'h39a7cfd2),
	.w2(32'h3a699e20),
	.w3(32'hbab1d05a),
	.w4(32'hb9d3831e),
	.w5(32'h39ff0073),
	.w6(32'h392c4c3a),
	.w7(32'h393db72e),
	.w8(32'h3a388001),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f1b3ab),
	.w1(32'hba326fb4),
	.w2(32'h3b1a424c),
	.w3(32'hba1b22f8),
	.w4(32'hbaa747a4),
	.w5(32'h3a8a10af),
	.w6(32'hbacd4747),
	.w7(32'hbac80c52),
	.w8(32'h3a982062),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae491d5),
	.w1(32'h3a03f74c),
	.w2(32'h3a6fc56c),
	.w3(32'h3aa7a478),
	.w4(32'h38b7cd90),
	.w5(32'h38e7e7a0),
	.w6(32'h3a507a76),
	.w7(32'h39c08707),
	.w8(32'h3aae4bc2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a41c8),
	.w1(32'h3aba4429),
	.w2(32'h3b1280f6),
	.w3(32'h3aba315d),
	.w4(32'h3a9da237),
	.w5(32'h3b18d09b),
	.w6(32'h3acd963d),
	.w7(32'h3af41ee3),
	.w8(32'h3b64904a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f70d5),
	.w1(32'h3a68d0d9),
	.w2(32'h3b18193d),
	.w3(32'h3a4f0fb9),
	.w4(32'h399732eb),
	.w5(32'h3b0c64fe),
	.w6(32'h3ae4edfa),
	.w7(32'h3aa266a3),
	.w8(32'h3afea8ca),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07d35d),
	.w1(32'hbb82e68f),
	.w2(32'hbacbd192),
	.w3(32'hbb0290fe),
	.w4(32'hbb599188),
	.w5(32'hbaba9c22),
	.w6(32'hbb958c50),
	.w7(32'hbb805146),
	.w8(32'hbb06a2a9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb252019),
	.w1(32'h3a580e74),
	.w2(32'h3b7d44a6),
	.w3(32'hb80bb91c),
	.w4(32'h3a7e35a2),
	.w5(32'h3af85be1),
	.w6(32'h3a88cd34),
	.w7(32'h3a9bc9b3),
	.w8(32'h3b06451e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39251262),
	.w1(32'hb993f5c4),
	.w2(32'h3a2b059c),
	.w3(32'h394036d8),
	.w4(32'hba673109),
	.w5(32'h39051855),
	.w6(32'hba02c241),
	.w7(32'hba20aa3d),
	.w8(32'h3a32a386),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915d769),
	.w1(32'h378317bd),
	.w2(32'hb80d54e6),
	.w3(32'hb84863dc),
	.w4(32'hb9015e99),
	.w5(32'hb934df44),
	.w6(32'hb7a3721a),
	.w7(32'hb800f2ce),
	.w8(32'hb913a0b3),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9977a89),
	.w1(32'hb7d5564e),
	.w2(32'h3979adc0),
	.w3(32'hb93196c8),
	.w4(32'hb87cfe57),
	.w5(32'h392ffe87),
	.w6(32'h385455ec),
	.w7(32'h392e117e),
	.w8(32'h3997f91e),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a69e81),
	.w1(32'h381deee0),
	.w2(32'hb7e96cde),
	.w3(32'h380da63e),
	.w4(32'hb814755a),
	.w5(32'hb8d4f19b),
	.w6(32'h38c859a1),
	.w7(32'hb80924de),
	.w8(32'hb8a85a7b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abb472),
	.w1(32'hb9dc25d3),
	.w2(32'hb9a59c5f),
	.w3(32'hb918b88e),
	.w4(32'hb945809b),
	.w5(32'hb9796d78),
	.w6(32'hb90570e8),
	.w7(32'hb94f4cd6),
	.w8(32'hb8b8c21c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84f195),
	.w1(32'h3a98f28c),
	.w2(32'h3aee2fb2),
	.w3(32'h3a66ae79),
	.w4(32'h3947e632),
	.w5(32'h384be694),
	.w6(32'h3a069baa),
	.w7(32'h399c4bb2),
	.w8(32'h3a906e55),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fa02e2),
	.w1(32'h398cbd55),
	.w2(32'hb92649f5),
	.w3(32'hb702660b),
	.w4(32'h39a8335d),
	.w5(32'hb8b70706),
	.w6(32'h3a53aaeb),
	.w7(32'h39944b52),
	.w8(32'hb819a6ed),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd59d4),
	.w1(32'hbb0559d3),
	.w2(32'h3959dfa9),
	.w3(32'hba26fe1f),
	.w4(32'hbb0a6dc1),
	.w5(32'hba886ee1),
	.w6(32'hbb4f2be8),
	.w7(32'hbb3247c2),
	.w8(32'hbac2dcb7),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c5cc5),
	.w1(32'h3a90bea0),
	.w2(32'h3b4680b8),
	.w3(32'hba3ecec5),
	.w4(32'h3ac538c5),
	.w5(32'h3b8a9699),
	.w6(32'h3aa15d2f),
	.w7(32'h3b66b641),
	.w8(32'h3bc70976),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf1295),
	.w1(32'h3a68b498),
	.w2(32'h3a26792b),
	.w3(32'hb8c95914),
	.w4(32'h3a1221d2),
	.w5(32'h39c135bd),
	.w6(32'h3a50d78c),
	.w7(32'h3a2781dc),
	.w8(32'h3a52bed2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1ae75),
	.w1(32'h39ab712d),
	.w2(32'h38630749),
	.w3(32'h398ecc67),
	.w4(32'h39c6fa04),
	.w5(32'h3944addd),
	.w6(32'h3a0e89d9),
	.w7(32'h39ac7397),
	.w8(32'h396f674f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f84f9),
	.w1(32'hb8ac5fde),
	.w2(32'hb86bf7bc),
	.w3(32'hb935831d),
	.w4(32'hb8efcdcd),
	.w5(32'hb911f9c3),
	.w6(32'hb88c71c1),
	.w7(32'hb9386b19),
	.w8(32'hb90dc576),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89b19b3),
	.w1(32'hb9b2f9c1),
	.w2(32'hb9c63fbe),
	.w3(32'h3798f4b1),
	.w4(32'hb90301dd),
	.w5(32'hb9572ec1),
	.w6(32'h396bc4ee),
	.w7(32'h38fac54b),
	.w8(32'h3948e4b3),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb607764),
	.w1(32'hbb0fec92),
	.w2(32'h3bb4c9c4),
	.w3(32'hbace5b3b),
	.w4(32'hbaf43d04),
	.w5(32'h3b7ed770),
	.w6(32'hbc3153cf),
	.w7(32'hbb74a1d0),
	.w8(32'h3aaf3304),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd94f9),
	.w1(32'h3a059e66),
	.w2(32'h3b5a982c),
	.w3(32'h3a49381a),
	.w4(32'h3a320da1),
	.w5(32'h3ad4e815),
	.w6(32'hba81ae5d),
	.w7(32'hb807f029),
	.w8(32'h3af3e8d0),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba263458),
	.w1(32'hb9cb07e4),
	.w2(32'h3a0276c4),
	.w3(32'hb9b8ca36),
	.w4(32'hb938ac21),
	.w5(32'h3990c9a1),
	.w6(32'hbaa9c2bb),
	.w7(32'hba7bba90),
	.w8(32'h3858309a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0478d1),
	.w1(32'hb922842c),
	.w2(32'h3a17a963),
	.w3(32'hba13d9b2),
	.w4(32'hba462e22),
	.w5(32'h39563754),
	.w6(32'hba4cf930),
	.w7(32'h382ec465),
	.w8(32'h39e3e686),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f4bf2),
	.w1(32'h39d36abc),
	.w2(32'h399dc10e),
	.w3(32'h39af3af4),
	.w4(32'hb8373f0d),
	.w5(32'h398ddccd),
	.w6(32'h3999327e),
	.w7(32'hb97116a4),
	.w8(32'h3999d3f7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7885b3e),
	.w1(32'h391db695),
	.w2(32'h3a9c623b),
	.w3(32'h39f832b9),
	.w4(32'h3989fea4),
	.w5(32'h3a7baa98),
	.w6(32'h3967698c),
	.w7(32'hb84df5be),
	.w8(32'h3a25a169),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70ee02),
	.w1(32'h3af39d96),
	.w2(32'h3a852d41),
	.w3(32'h3ab2de42),
	.w4(32'h3ad5b73d),
	.w5(32'h3a9b769c),
	.w6(32'h3acbd3af),
	.w7(32'h3a889238),
	.w8(32'h3ad5df28),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa26dd8),
	.w1(32'hbb1e143e),
	.w2(32'h3b26b70f),
	.w3(32'hba5ff4f9),
	.w4(32'hbb513bf7),
	.w5(32'h3b4c0bb5),
	.w6(32'hbc0a9072),
	.w7(32'hbbc32f70),
	.w8(32'hbb1ff15a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a279414),
	.w1(32'hb9b2c7db),
	.w2(32'h39ba0f94),
	.w3(32'h39934409),
	.w4(32'hb98ad36f),
	.w5(32'h3a7b8781),
	.w6(32'h3a796700),
	.w7(32'h3a1c104c),
	.w8(32'h3b120907),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad52747),
	.w1(32'h39e776a2),
	.w2(32'h3b611ee3),
	.w3(32'hba965afc),
	.w4(32'hb8e419e6),
	.w5(32'h3afd13f7),
	.w6(32'hbaf8269b),
	.w7(32'hb9c2a68d),
	.w8(32'h3b44335f),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3eb9d6),
	.w1(32'hbb58d58b),
	.w2(32'h3aa3fb28),
	.w3(32'hbadbae0f),
	.w4(32'hbb9fbc0b),
	.w5(32'h3b3c39ee),
	.w6(32'hbc331e93),
	.w7(32'hbc1d40be),
	.w8(32'hbb790bdb),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ceca28),
	.w1(32'hbabe3132),
	.w2(32'hb9700a78),
	.w3(32'hb90525f2),
	.w4(32'hbaaa29ae),
	.w5(32'hba4332b5),
	.w6(32'hba633718),
	.w7(32'hba571077),
	.w8(32'h39fba598),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93ee4dd),
	.w1(32'h391854bb),
	.w2(32'h3b5cc177),
	.w3(32'h3a26df55),
	.w4(32'h3a12706c),
	.w5(32'h3b175e7d),
	.w6(32'hba89c342),
	.w7(32'hb9a861ed),
	.w8(32'h3b254ac1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db1300),
	.w1(32'h38bd5ef3),
	.w2(32'h3a01d99d),
	.w3(32'hb8a8a3a7),
	.w4(32'hb8e352cb),
	.w5(32'h390f9c7e),
	.w6(32'h393a5dae),
	.w7(32'hb8d27922),
	.w8(32'h3994a44e),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad79ba5),
	.w1(32'hba665928),
	.w2(32'h3a8a0647),
	.w3(32'h3b520a1c),
	.w4(32'h3943c343),
	.w5(32'h3b39f2e4),
	.w6(32'h3bb5a63c),
	.w7(32'h3b482ce6),
	.w8(32'h3b853331),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e5991d),
	.w1(32'hb8a611b8),
	.w2(32'h3a11fa90),
	.w3(32'h3957f951),
	.w4(32'hb992a03d),
	.w5(32'h3a160123),
	.w6(32'hba2645eb),
	.w7(32'hb9d827d6),
	.w8(32'h39451352),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82e7e23),
	.w1(32'hb864487e),
	.w2(32'hb7e36367),
	.w3(32'hb8ef47fb),
	.w4(32'hb8bb4c71),
	.w5(32'hb7f342d9),
	.w6(32'hb8a20110),
	.w7(32'hb711b0a3),
	.w8(32'h378fcaab),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb821e84b),
	.w1(32'hb7b6287c),
	.w2(32'hb8dbf775),
	.w3(32'hb858cb4e),
	.w4(32'hb884aff8),
	.w5(32'hb8bbca89),
	.w6(32'hb8800298),
	.w7(32'hb90f34ab),
	.w8(32'hb9114e5a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952163d),
	.w1(32'hba82dd60),
	.w2(32'hba3ede84),
	.w3(32'h3a07805c),
	.w4(32'hba216d1c),
	.w5(32'hba69d200),
	.w6(32'hba6f0cae),
	.w7(32'h3927a178),
	.w8(32'h3a1e35ca),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58abd2),
	.w1(32'hbafb13e0),
	.w2(32'hb8be26a4),
	.w3(32'hb5acab9c),
	.w4(32'hbb105e90),
	.w5(32'h39174820),
	.w6(32'hb9bbb66e),
	.w7(32'hbb0cde38),
	.w8(32'h3a0a30e9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb007c),
	.w1(32'hba5b4ba9),
	.w2(32'h3a9f9404),
	.w3(32'hba00de52),
	.w4(32'hba39d850),
	.w5(32'h3a073d3d),
	.w6(32'hba6e4fff),
	.w7(32'hbabfbdd9),
	.w8(32'h39a5df97),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb718ee0a),
	.w1(32'h388589ab),
	.w2(32'h36cf92c5),
	.w3(32'hb78d8004),
	.w4(32'h3843ef6c),
	.w5(32'hb6d60dd5),
	.w6(32'h38769595),
	.w7(32'h3726a7ca),
	.w8(32'hb76e52dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c53dd5),
	.w1(32'h399e2337),
	.w2(32'h3b6ea71d),
	.w3(32'h3ab4dcfc),
	.w4(32'h3a67ef96),
	.w5(32'h3b13434b),
	.w6(32'hb709d875),
	.w7(32'h37e3b1ff),
	.w8(32'h3b121e78),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc9308),
	.w1(32'hb87340b2),
	.w2(32'h3a830dc3),
	.w3(32'h3a249f30),
	.w4(32'h3819d8d4),
	.w5(32'h3996925d),
	.w6(32'h3800ec66),
	.w7(32'h38a65942),
	.w8(32'h3ad5837e),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96bce9),
	.w1(32'hbbaacf77),
	.w2(32'h3b0d0ef9),
	.w3(32'hbb37e8aa),
	.w4(32'hbb866a4f),
	.w5(32'hba4414d5),
	.w6(32'hbc069be4),
	.w7(32'hbbce0414),
	.w8(32'hbb92bd9f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34469b),
	.w1(32'h398b8c27),
	.w2(32'h3b2f1158),
	.w3(32'h3b324dd3),
	.w4(32'h39d23535),
	.w5(32'h3a95ba30),
	.w6(32'h3ba19d44),
	.w7(32'h3b176532),
	.w8(32'h3b08c10e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b31dd9),
	.w1(32'h3a228dc6),
	.w2(32'h3a7299d1),
	.w3(32'h3a0001b5),
	.w4(32'h3a8d3440),
	.w5(32'h3acb1fca),
	.w6(32'h3a1da134),
	.w7(32'h3aa77742),
	.w8(32'h3b016e23),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a671b51),
	.w1(32'h3a0a7497),
	.w2(32'hb8e2ca4e),
	.w3(32'h3a0a8f43),
	.w4(32'h38b91233),
	.w5(32'hb9179e92),
	.w6(32'h3a85d7bb),
	.w7(32'h3a1d8d50),
	.w8(32'h39076aa5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94654d9),
	.w1(32'hba8cb086),
	.w2(32'h39a49389),
	.w3(32'hb91708fc),
	.w4(32'hbaefb47b),
	.w5(32'hba1d98a1),
	.w6(32'hb9f1f464),
	.w7(32'hbad11485),
	.w8(32'hba077f67),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ba007),
	.w1(32'hb9ada571),
	.w2(32'h39a1f038),
	.w3(32'h397604b3),
	.w4(32'h3a0106b7),
	.w5(32'h39d41a54),
	.w6(32'h3b002362),
	.w7(32'h3a3d1872),
	.w8(32'h3a95f17b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388460c2),
	.w1(32'hba0d49d0),
	.w2(32'hba3797ce),
	.w3(32'hb762f77b),
	.w4(32'hb98ca6d4),
	.w5(32'hb81cb545),
	.w6(32'h3a681289),
	.w7(32'h39810e1f),
	.w8(32'h3a667a5e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986f62b),
	.w1(32'hba4574c7),
	.w2(32'h3a01b5dd),
	.w3(32'hb921abcd),
	.w4(32'hba0a2a5d),
	.w5(32'h39cb581a),
	.w6(32'hbacd3f7a),
	.w7(32'hbacbd131),
	.w8(32'hb9c238a5),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9861d3f),
	.w1(32'hb7e28cf4),
	.w2(32'hb8c30a10),
	.w3(32'hb944dd74),
	.w4(32'h38a9c451),
	.w5(32'h394eb6b5),
	.w6(32'hb9280189),
	.w7(32'h38a70fd6),
	.w8(32'h398aea47),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b72154),
	.w1(32'h398a2c89),
	.w2(32'h3b5c16aa),
	.w3(32'h3a0e6fc0),
	.w4(32'h38c7e513),
	.w5(32'h3b2f50d5),
	.w6(32'hbb3c6e90),
	.w7(32'hbb1dd63b),
	.w8(32'h3a86bcea),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bdc434),
	.w1(32'hba2e2a46),
	.w2(32'h38f30815),
	.w3(32'hb991f97d),
	.w4(32'hb99fa64b),
	.w5(32'h3968ea1c),
	.w6(32'hba1f3dec),
	.w7(32'hba2b9886),
	.w8(32'h39d2364c),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3538e),
	.w1(32'h38814689),
	.w2(32'h387f7bf7),
	.w3(32'h39fe8d55),
	.w4(32'hb894e709),
	.w5(32'hba26f98d),
	.w6(32'h3972c018),
	.w7(32'hba010350),
	.w8(32'hb9bd60f8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85cbd08),
	.w1(32'hb98cb0d5),
	.w2(32'hba297d17),
	.w3(32'h3952dd5c),
	.w4(32'hb7ff0405),
	.w5(32'hba13f608),
	.w6(32'h3997b202),
	.w7(32'h372f1e3b),
	.w8(32'hb9dc69a8),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabfa1dc),
	.w1(32'hba1e6ceb),
	.w2(32'h3a8e3a02),
	.w3(32'hb96425a0),
	.w4(32'h3a8667f4),
	.w5(32'h3affa3b7),
	.w6(32'hba04ed79),
	.w7(32'hb92a6f61),
	.w8(32'h3ae232a1),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d10e91),
	.w1(32'h37f4c982),
	.w2(32'hb8679ca2),
	.w3(32'h3886e858),
	.w4(32'hb6f509d2),
	.w5(32'hb8ad871f),
	.w6(32'hb49a694a),
	.w7(32'hb8ab9e1b),
	.w8(32'hb909c0e3),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88aeeeb),
	.w1(32'hb928ee18),
	.w2(32'hb98bfe06),
	.w3(32'hb8b8a635),
	.w4(32'hb91e87b9),
	.w5(32'hb9600bdc),
	.w6(32'hb932c50b),
	.w7(32'hb8a797c4),
	.w8(32'hb8ba175a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f39213),
	.w1(32'hba5bac12),
	.w2(32'hb913d2b5),
	.w3(32'hba701c63),
	.w4(32'hba80e3e5),
	.w5(32'hb9e56160),
	.w6(32'h37e81906),
	.w7(32'hb9afc0e3),
	.w8(32'h3a52141b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a286b7e),
	.w1(32'h39dbaefe),
	.w2(32'h3ba14f9c),
	.w3(32'hbad17744),
	.w4(32'hbafc2213),
	.w5(32'h3afed281),
	.w6(32'hbb963f34),
	.w7(32'hbb85f823),
	.w8(32'h3abd0bb1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71db825),
	.w1(32'hba915f8a),
	.w2(32'hba62cdac),
	.w3(32'h39999cd8),
	.w4(32'hba03e108),
	.w5(32'hb8e96e13),
	.w6(32'h39d99cca),
	.w7(32'hb9a57bdc),
	.w8(32'hb79d943f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39515b6c),
	.w1(32'hb9fbe9bf),
	.w2(32'hb99a5cb7),
	.w3(32'hba7575c1),
	.w4(32'hbaa1d324),
	.w5(32'hb9b25868),
	.w6(32'h38d4bd9b),
	.w7(32'h39698f64),
	.w8(32'h3aea0129),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb616c3d4),
	.w1(32'hb92e4e33),
	.w2(32'h394a123e),
	.w3(32'h39c76b79),
	.w4(32'h39cd039b),
	.w5(32'h39312ba2),
	.w6(32'h3ab3c2d0),
	.w7(32'h39e60134),
	.w8(32'h3a1e7849),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d90fda),
	.w1(32'h3ad09234),
	.w2(32'h3b2b0c6b),
	.w3(32'h3ac850d8),
	.w4(32'hb9761c1a),
	.w5(32'h38f2dcd4),
	.w6(32'h3b0bc79f),
	.w7(32'h39b158f5),
	.w8(32'h39a23f43),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4026d),
	.w1(32'h39d9e518),
	.w2(32'h3b0c3393),
	.w3(32'h39811ae7),
	.w4(32'h3a52d402),
	.w5(32'h3ae3c571),
	.w6(32'hba58b05d),
	.w7(32'hb975acea),
	.w8(32'h3a94e9ab),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ca085),
	.w1(32'h3aedfa38),
	.w2(32'h3b93196c),
	.w3(32'h3abcfce1),
	.w4(32'h3aa379f3),
	.w5(32'h3b68d3b3),
	.w6(32'hba4cf820),
	.w7(32'hb9fddeac),
	.w8(32'h3aedf1e4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae142e),
	.w1(32'h3a117b86),
	.w2(32'hb8384387),
	.w3(32'h39d304f6),
	.w4(32'h3a0949dd),
	.w5(32'hb6c1b2b2),
	.w6(32'h39fc0bb7),
	.w7(32'h39bbed24),
	.w8(32'hb821cd7c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39ba07),
	.w1(32'h39c62e75),
	.w2(32'h3b223564),
	.w3(32'hb9cfd4ca),
	.w4(32'h39d2fbcc),
	.w5(32'h3adcc989),
	.w6(32'hba845767),
	.w7(32'hba7eb788),
	.w8(32'h39b8d476),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782061a),
	.w1(32'h37f0bcac),
	.w2(32'hb7909bbe),
	.w3(32'hb76193d4),
	.w4(32'h37117884),
	.w5(32'hb7d0eb5d),
	.w6(32'hb56465a1),
	.w7(32'h37027576),
	.w8(32'hb779ba9d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82ef704),
	.w1(32'h39945201),
	.w2(32'h3a3270c9),
	.w3(32'h3845ee1f),
	.w4(32'h38b418ba),
	.w5(32'h393e3be7),
	.w6(32'h38b2e082),
	.w7(32'h380cec0c),
	.w8(32'h3a161cab),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91374fe),
	.w1(32'hb9594bed),
	.w2(32'h396120f8),
	.w3(32'hb7f038de),
	.w4(32'hb9c43818),
	.w5(32'h3959341d),
	.w6(32'h39100da0),
	.w7(32'h39f1f024),
	.w8(32'h3a1c8f56),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fb02d),
	.w1(32'h3a02ff49),
	.w2(32'h3b393c59),
	.w3(32'h3899ac79),
	.w4(32'h3a23d3e9),
	.w5(32'h3a6aaa52),
	.w6(32'hb80924c6),
	.w7(32'h3a5b1f0a),
	.w8(32'h3af13517),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64d1f68),
	.w1(32'h37a840b7),
	.w2(32'hb868f7d7),
	.w3(32'h378ccbc3),
	.w4(32'h37a7b029),
	.w5(32'hb810eb7f),
	.w6(32'h37bed89a),
	.w7(32'hb821052c),
	.w8(32'hb7e21efd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3861d05e),
	.w1(32'h38d2541f),
	.w2(32'h38e37500),
	.w3(32'h38759a52),
	.w4(32'h388a6118),
	.w5(32'h38990cd5),
	.w6(32'h383e15db),
	.w7(32'h3850b9b1),
	.w8(32'h38d2dbf4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55622f),
	.w1(32'hba570302),
	.w2(32'h3a270889),
	.w3(32'hb9f7780e),
	.w4(32'hbb0d3416),
	.w5(32'hbac8642b),
	.w6(32'hbb11769a),
	.w7(32'hbacff6be),
	.w8(32'hba1d5ff8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a992464),
	.w1(32'h3a2f11e8),
	.w2(32'h3b833de5),
	.w3(32'h3a8f4b35),
	.w4(32'h3a2b0aa4),
	.w5(32'h3b1eb760),
	.w6(32'hbb0eb335),
	.w7(32'h398e8881),
	.w8(32'h3b277229),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84e93e),
	.w1(32'hbb87c50d),
	.w2(32'hbaeecd76),
	.w3(32'h3b2485ee),
	.w4(32'hbad51eff),
	.w5(32'hbad64acc),
	.w6(32'hbb5b23c9),
	.w7(32'hbb6a5b0f),
	.w8(32'hba482b6d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0f255),
	.w1(32'hb9bd4c96),
	.w2(32'hb9e86633),
	.w3(32'h38be79fd),
	.w4(32'hb93dae96),
	.w5(32'hb97b2a5b),
	.w6(32'h39563165),
	.w7(32'hb78c8c33),
	.w8(32'hb9adf38c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c9cfc),
	.w1(32'h3a9b37f0),
	.w2(32'h3bcda7e7),
	.w3(32'hbab6bfee),
	.w4(32'hbb0a824a),
	.w5(32'hb9e8748c),
	.w6(32'hbc15d4f0),
	.w7(32'hbbf2f114),
	.w8(32'hbae7f4c9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cdb2b),
	.w1(32'hb76ea547),
	.w2(32'h3a8f5759),
	.w3(32'h39548bbb),
	.w4(32'h3815fa95),
	.w5(32'h39763f3c),
	.w6(32'h3a85252f),
	.w7(32'hba1de4fc),
	.w8(32'h3b4ccbdd),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba849529),
	.w1(32'hbae5b505),
	.w2(32'h39868c9e),
	.w3(32'hba68e75a),
	.w4(32'hba906edb),
	.w5(32'hb80ec2d1),
	.w6(32'hbae603d8),
	.w7(32'hbac66f1c),
	.w8(32'h39c3fa95),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c6b246),
	.w1(32'h36510f12),
	.w2(32'h38e207f7),
	.w3(32'h3751b0f6),
	.w4(32'h37f0df03),
	.w5(32'h38b91371),
	.w6(32'h363b175c),
	.w7(32'h38f81a09),
	.w8(32'hb5a48fc6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de243c),
	.w1(32'h38d8f47a),
	.w2(32'h390df4eb),
	.w3(32'hb6d5e684),
	.w4(32'hb79fafff),
	.w5(32'h38a8bc65),
	.w6(32'h37826815),
	.w7(32'h38b03edb),
	.w8(32'h3955b398),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385756fd),
	.w1(32'hb7b4923a),
	.w2(32'hb824a687),
	.w3(32'h382c18dc),
	.w4(32'hb7c6946e),
	.w5(32'hb8005d81),
	.w6(32'hb784bcfa),
	.w7(32'hb6be8ce3),
	.w8(32'hb756fbce),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7257378),
	.w1(32'hbb181132),
	.w2(32'h39f32391),
	.w3(32'hba367984),
	.w4(32'hbb073345),
	.w5(32'h3a13c779),
	.w6(32'hbb2cddcd),
	.w7(32'hbb147537),
	.w8(32'h3a3b9bca),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bf7de),
	.w1(32'hb98b0d8d),
	.w2(32'h3a06613d),
	.w3(32'hb9374647),
	.w4(32'hba97cd09),
	.w5(32'h3921f162),
	.w6(32'hba047a42),
	.w7(32'hba8c6d2b),
	.w8(32'h392c980e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a4c73),
	.w1(32'h3927fc42),
	.w2(32'h39d2502a),
	.w3(32'h3a93e8d4),
	.w4(32'hb6df3a00),
	.w5(32'hb9ae800a),
	.w6(32'h3b0dc5f8),
	.w7(32'h3a04ff9f),
	.w8(32'h3a840a68),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39868bd6),
	.w1(32'hb94424b5),
	.w2(32'h36ec6df3),
	.w3(32'h390b124b),
	.w4(32'hb987bdf4),
	.w5(32'hb8199de1),
	.w6(32'h391cec3a),
	.w7(32'hb8a6436f),
	.w8(32'h396f5b03),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada75b1),
	.w1(32'hbb0e6f61),
	.w2(32'h3b0f8654),
	.w3(32'hbae4c003),
	.w4(32'hbb309178),
	.w5(32'h39941f3a),
	.w6(32'hbb651e81),
	.w7(32'hbb8342f5),
	.w8(32'h39f6d2a8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ab629),
	.w1(32'hba2f4191),
	.w2(32'hb958bd83),
	.w3(32'h3aca404f),
	.w4(32'h39c5859b),
	.w5(32'hb96e3adf),
	.w6(32'hb90bdfb4),
	.w7(32'hb86c79aa),
	.w8(32'hb9c56587),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3796b7b6),
	.w1(32'h37c72637),
	.w2(32'hb7fa8745),
	.w3(32'h37d65fd8),
	.w4(32'h37081529),
	.w5(32'hb81e8d34),
	.w6(32'h36fa6ecb),
	.w7(32'hb79c6b71),
	.w8(32'hb831800c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917185f),
	.w1(32'hba32cd01),
	.w2(32'h3a5eca6d),
	.w3(32'h39fdf1d4),
	.w4(32'hba878c86),
	.w5(32'h3a1b5f42),
	.w6(32'hbb19c936),
	.w7(32'hbb343002),
	.w8(32'hba852500),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb391c72b),
	.w1(32'h387ad3e9),
	.w2(32'hb7e94922),
	.w3(32'hb8072890),
	.w4(32'h37bc29d8),
	.w5(32'hb85da5be),
	.w6(32'hb60a1d6a),
	.w7(32'h35e3bf7e),
	.w8(32'hb84c93ee),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9825dd),
	.w1(32'hb84eb9ee),
	.w2(32'h3b3f8821),
	.w3(32'hba3a74fd),
	.w4(32'h38e5cafb),
	.w5(32'h3b3d45ed),
	.w6(32'hbaba0c9c),
	.w7(32'hb9017938),
	.w8(32'h3aff4f12),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1dd05),
	.w1(32'h398d09eb),
	.w2(32'h3ad6389a),
	.w3(32'h395bbca1),
	.w4(32'h39814c72),
	.w5(32'h3aa9f969),
	.w6(32'h3b0833d0),
	.w7(32'h3b1b5d0a),
	.w8(32'h3b7ea7b5),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e77cca),
	.w1(32'hba8b7fb2),
	.w2(32'h39259ad6),
	.w3(32'h39abf8c2),
	.w4(32'hba526015),
	.w5(32'h38cfcc68),
	.w6(32'h39bc7b4b),
	.w7(32'hba0e7b36),
	.w8(32'h3aa7d0aa),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24e367),
	.w1(32'hba6b3f06),
	.w2(32'hb9e79a93),
	.w3(32'hba21829d),
	.w4(32'hba3941d4),
	.w5(32'hb97a27aa),
	.w6(32'hb9cac9fc),
	.w7(32'hba06ebda),
	.w8(32'hb9527aa8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65abe2),
	.w1(32'hba69e46c),
	.w2(32'hb97e9bf8),
	.w3(32'h3aa1b3a8),
	.w4(32'hb9213ab5),
	.w5(32'h392b39dd),
	.w6(32'h3ae96e06),
	.w7(32'h399075c5),
	.w8(32'h3a4fbd01),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890eaf8),
	.w1(32'h39f24ebd),
	.w2(32'h3b334c03),
	.w3(32'h3a24bc8c),
	.w4(32'h3a567a16),
	.w5(32'h3a874aaa),
	.w6(32'hb90510f4),
	.w7(32'hb8704979),
	.w8(32'h3ad1f359),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89e4c84),
	.w1(32'h3a298362),
	.w2(32'h3b1111d6),
	.w3(32'h39786dae),
	.w4(32'h39b81184),
	.w5(32'h3a1faf59),
	.w6(32'hba53d356),
	.w7(32'hbab4a01d),
	.w8(32'h39e3ad01),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82c641d),
	.w1(32'hb833e7a3),
	.w2(32'hb7e29f89),
	.w3(32'hb845d9a4),
	.w4(32'hb881b40b),
	.w5(32'hb7d051a8),
	.w6(32'hb8ad7f87),
	.w7(32'hb8050dfc),
	.w8(32'h36e0aeef),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80fa0be),
	.w1(32'hb829172f),
	.w2(32'h375ec207),
	.w3(32'h3753b4c4),
	.w4(32'h38747fd3),
	.w5(32'h38c56225),
	.w6(32'hb6999864),
	.w7(32'hb8085ae1),
	.w8(32'hb7f6deea),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb788f1ad),
	.w1(32'hbad15595),
	.w2(32'h3aeb6021),
	.w3(32'hbac70dcb),
	.w4(32'hbacc88b4),
	.w5(32'h3b22c240),
	.w6(32'hbb0aa562),
	.w7(32'hba3d8a20),
	.w8(32'h3b6c10b6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d52e8),
	.w1(32'h3aa6f1ab),
	.w2(32'h3b89b8f3),
	.w3(32'hba314590),
	.w4(32'hbaad4235),
	.w5(32'h3adc27e1),
	.w6(32'hbb3c9f9c),
	.w7(32'hba60d6f8),
	.w8(32'h3b0c820a),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a8e02),
	.w1(32'hba732145),
	.w2(32'h3afff7b2),
	.w3(32'h39b24937),
	.w4(32'hbadbd615),
	.w5(32'hba1286ba),
	.w6(32'hbad108f2),
	.w7(32'hbabea4d4),
	.w8(32'h39f791e3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac72e63),
	.w1(32'hbb8681c9),
	.w2(32'h3b55dd48),
	.w3(32'hbaa7e351),
	.w4(32'hbb59f6af),
	.w5(32'h3adbd1bf),
	.w6(32'hbbbaadd5),
	.w7(32'hbb393711),
	.w8(32'h3ae9f1b8),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92e927a),
	.w1(32'h393e6171),
	.w2(32'h38f2dac1),
	.w3(32'hb974416d),
	.w4(32'h3910cee4),
	.w5(32'h38c4cee6),
	.w6(32'hb93d67e6),
	.w7(32'h394392ce),
	.w8(32'h395480c6),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cdc29),
	.w1(32'h39eeadd2),
	.w2(32'h3a5b6cd4),
	.w3(32'hb98b9fe0),
	.w4(32'h3a183168),
	.w5(32'h3a830600),
	.w6(32'hb92bf4c4),
	.w7(32'h3a3b2c68),
	.w8(32'h3a41a3c3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8345fb),
	.w1(32'hbc149fdc),
	.w2(32'h39fa732a),
	.w3(32'h3b167219),
	.w4(32'hbbb109fb),
	.w5(32'h3b731c86),
	.w6(32'hba4e3e51),
	.w7(32'hbbdb574f),
	.w8(32'h3b295206),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa37dd),
	.w1(32'hbb013f01),
	.w2(32'h3b12a638),
	.w3(32'hbac1278b),
	.w4(32'hbb80ec76),
	.w5(32'hba84f87a),
	.w6(32'hbbeb22d6),
	.w7(32'hbbcd9424),
	.w8(32'hbb3dd8ed),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2181cb),
	.w1(32'hbb5e1a01),
	.w2(32'hb88f740f),
	.w3(32'h3964a46d),
	.w4(32'hbae292f1),
	.w5(32'h375ab080),
	.w6(32'hbc09ff2b),
	.w7(32'hbbd8ffc8),
	.w8(32'hbb5bb60c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a898a4a),
	.w1(32'hb9e9f63a),
	.w2(32'hba62d8eb),
	.w3(32'h3a8f44f0),
	.w4(32'h390d3970),
	.w5(32'h38a6f908),
	.w6(32'h3aef2993),
	.w7(32'h3a8ce01c),
	.w8(32'h3adb25a9),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae139c),
	.w1(32'h3aae5932),
	.w2(32'h3ab71aa4),
	.w3(32'h394e76c7),
	.w4(32'h3a653f26),
	.w5(32'h3a7e84ac),
	.w6(32'h3b0dfaa1),
	.w7(32'h3ad7e11d),
	.w8(32'h3b5f8b27),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d1966),
	.w1(32'hb74c05ca),
	.w2(32'hb81b274f),
	.w3(32'h374531be),
	.w4(32'hb6a81bdb),
	.w5(32'hb7b6e5fb),
	.w6(32'hb66cc68d),
	.w7(32'hb7a63614),
	.w8(32'hb7a8159b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8004782),
	.w1(32'hb86f9738),
	.w2(32'hb8b33fca),
	.w3(32'hb79735c2),
	.w4(32'hb847fe71),
	.w5(32'hb867d30a),
	.w6(32'hb81f2f69),
	.w7(32'hb863e7ff),
	.w8(32'hb86f1d20),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12ad7c),
	.w1(32'hb9e5a23f),
	.w2(32'hb9085929),
	.w3(32'h3a0317d5),
	.w4(32'h39bd350d),
	.w5(32'h39a5ada2),
	.w6(32'hb9846cde),
	.w7(32'hba124457),
	.w8(32'h395ea9f4),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76f7d2d),
	.w1(32'h381dd2d1),
	.w2(32'h38021a58),
	.w3(32'h360ad730),
	.w4(32'h382aaeae),
	.w5(32'h3773c407),
	.w6(32'hb6d1916f),
	.w7(32'h372dbbe1),
	.w8(32'hb778fa78),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba661d8a),
	.w1(32'hbaecfc97),
	.w2(32'h39c2d92f),
	.w3(32'hb9a95ad3),
	.w4(32'hb9c9c7dc),
	.w5(32'h3a683b74),
	.w6(32'hbaab8540),
	.w7(32'hb9e8f039),
	.w8(32'h3a615932),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd99bb),
	.w1(32'h3993bf23),
	.w2(32'h3baec316),
	.w3(32'hbb0674ee),
	.w4(32'hba931c99),
	.w5(32'h3b868d60),
	.w6(32'hbb942598),
	.w7(32'hba92d39d),
	.w8(32'h3b0eeb33),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f3c4b),
	.w1(32'hb8a012d0),
	.w2(32'h3aa574c0),
	.w3(32'h39b5e470),
	.w4(32'hb9bb381a),
	.w5(32'h3a85a237),
	.w6(32'hba514a50),
	.w7(32'hba0bdef6),
	.w8(32'h3a927421),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e3d26b),
	.w1(32'hb7370729),
	.w2(32'hb8e068e4),
	.w3(32'hb6bbf13f),
	.w4(32'hb83fca23),
	.w5(32'hb8b62af8),
	.w6(32'h38035ea6),
	.w7(32'hb8410b91),
	.w8(32'hb88ef7fa),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa92441),
	.w1(32'hbbb32985),
	.w2(32'h3aba9ed4),
	.w3(32'hbae6cecc),
	.w4(32'hbb922968),
	.w5(32'h3b0abd60),
	.w6(32'hbc3d04fd),
	.w7(32'hbc1c330d),
	.w8(32'hbb8d4640),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b02cf5),
	.w1(32'h39cb490a),
	.w2(32'h3b0e65ba),
	.w3(32'hb9a7c92a),
	.w4(32'h38ce5855),
	.w5(32'h3aa9f99d),
	.w6(32'hbae8a101),
	.w7(32'hba6b2c5b),
	.w8(32'h3a5309c8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f5ad30),
	.w1(32'h38cb2261),
	.w2(32'hb8214422),
	.w3(32'h3951964c),
	.w4(32'h392ee2eb),
	.w5(32'h38944b25),
	.w6(32'h394f7e1d),
	.w7(32'h39056dbf),
	.w8(32'h39136c88),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae893),
	.w1(32'hbae0b682),
	.w2(32'h3a6e18f8),
	.w3(32'hbad7883a),
	.w4(32'hbae3c656),
	.w5(32'h3954da59),
	.w6(32'hbb59c0b4),
	.w7(32'hbb73363b),
	.w8(32'hba83bd94),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390eb99b),
	.w1(32'h38ffadcf),
	.w2(32'h3878555f),
	.w3(32'h380f00f2),
	.w4(32'h3880103c),
	.w5(32'h37f279e7),
	.w6(32'h38d6d0a7),
	.w7(32'h38c9b6a3),
	.w8(32'h38a9a097),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cb0df8),
	.w1(32'h388fd3d1),
	.w2(32'h388001cb),
	.w3(32'hb9342c45),
	.w4(32'h38767cbd),
	.w5(32'h3944dc8a),
	.w6(32'hb807b828),
	.w7(32'h38f1b59d),
	.w8(32'h39904fd9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78606d6),
	.w1(32'h37f1ff9b),
	.w2(32'hb844962f),
	.w3(32'h36256874),
	.w4(32'h3774d0b5),
	.w5(32'hb7e0fe90),
	.w6(32'h380901ff),
	.w7(32'hb777de34),
	.w8(32'hb7b6aaf9),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cd8094),
	.w1(32'hb80b6877),
	.w2(32'h36ed34ef),
	.w3(32'h371030a1),
	.w4(32'h33bd2ead),
	.w5(32'h376d3903),
	.w6(32'hb800f60b),
	.w7(32'h380d48b8),
	.w8(32'h373f7c52),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d479fe),
	.w1(32'hba8ab155),
	.w2(32'hba94ef4e),
	.w3(32'h3a8017b9),
	.w4(32'hba03c0cc),
	.w5(32'hba5e7a91),
	.w6(32'h399626c9),
	.w7(32'hba33ef84),
	.w8(32'hb9e8c353),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7acb77),
	.w1(32'h3aa4df76),
	.w2(32'h3bc82d2f),
	.w3(32'h3b01c727),
	.w4(32'h3a8fcc72),
	.w5(32'h3b3a63e9),
	.w6(32'h3a52e171),
	.w7(32'h3a070f85),
	.w8(32'h3b7e71ca),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acda86),
	.w1(32'h36b43516),
	.w2(32'h3b450baf),
	.w3(32'hb8687d60),
	.w4(32'hba1afbed),
	.w5(32'h3af29b4f),
	.w6(32'hbb24f3a0),
	.w7(32'hbb324937),
	.w8(32'hb8d4d029),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba828854),
	.w1(32'hba1af308),
	.w2(32'h3b474871),
	.w3(32'h38a19b19),
	.w4(32'hb99179f5),
	.w5(32'h3abf2ccd),
	.w6(32'hbb12bc58),
	.w7(32'hbb275073),
	.w8(32'h39b39f41),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63e65f3),
	.w1(32'hb8d52b6a),
	.w2(32'hb90cc86c),
	.w3(32'h3891b00f),
	.w4(32'hb7c95b02),
	.w5(32'hb8a33f85),
	.w6(32'h39171f1f),
	.w7(32'h385bd5a3),
	.w8(32'hb8a6c0c4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bf19f6),
	.w1(32'h398161eb),
	.w2(32'h38a140b8),
	.w3(32'h37a8832d),
	.w4(32'h39a7a9f8),
	.w5(32'h397e9202),
	.w6(32'h38960e08),
	.w7(32'h39a6b2ca),
	.w8(32'h395fd83e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3606ecf4),
	.w1(32'h377a532f),
	.w2(32'hb7b4e3f9),
	.w3(32'h370d4286),
	.w4(32'h34e0ba91),
	.w5(32'hb78d63f3),
	.w6(32'h36f63962),
	.w7(32'hb70b0783),
	.w8(32'hb6f96775),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79ec4c5),
	.w1(32'h378cdbd5),
	.w2(32'hb7b0bbcb),
	.w3(32'hb7051152),
	.w4(32'h37eb8460),
	.w5(32'hb782a738),
	.w6(32'h37e3ad4c),
	.w7(32'h37973ca2),
	.w8(32'hb7052152),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c4340),
	.w1(32'h3a49dae7),
	.w2(32'h3b34014d),
	.w3(32'h37e20f2d),
	.w4(32'h3a53fefc),
	.w5(32'h3b08d087),
	.w6(32'hbaee7d2d),
	.w7(32'hba3b8ba9),
	.w8(32'hb95e8367),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85786d0),
	.w1(32'h394c17d1),
	.w2(32'h38f3e56e),
	.w3(32'hb90dcc81),
	.w4(32'h37e44855),
	.w5(32'h37b2d0b7),
	.w6(32'h376a876e),
	.w7(32'h382613c8),
	.w8(32'h38682bb3),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944f737),
	.w1(32'hba2a3366),
	.w2(32'hba158258),
	.w3(32'hb7ba6d77),
	.w4(32'hb9ca9bb2),
	.w5(32'hb9e1143e),
	.w6(32'h39e1430c),
	.w7(32'hb8a4d265),
	.w8(32'hb928fe79),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37eab5a6),
	.w1(32'h3a90b8fa),
	.w2(32'hb88b309d),
	.w3(32'h3a851950),
	.w4(32'h3a2b27a7),
	.w5(32'h399a9845),
	.w6(32'h3a42fab0),
	.w7(32'h3a18c221),
	.w8(32'hb98f6bee),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3724d634),
	.w1(32'h3771094c),
	.w2(32'hb6227731),
	.w3(32'h36bd9199),
	.w4(32'hb79d70d6),
	.w5(32'hb77c8e06),
	.w6(32'hb69d24a5),
	.w7(32'hb81c6599),
	.w8(32'hb81b92e0),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5a2365),
	.w1(32'hba0462cd),
	.w2(32'h3a32a15b),
	.w3(32'hba28d1b2),
	.w4(32'hba6795ca),
	.w5(32'h39261e87),
	.w6(32'hbaf2fb49),
	.w7(32'hbab41e77),
	.w8(32'hb9e626c1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3859c5ec),
	.w1(32'h397f9535),
	.w2(32'h392e8e36),
	.w3(32'h3987205c),
	.w4(32'h39cc8f9a),
	.w5(32'h39a1ef98),
	.w6(32'h39bd5ffb),
	.w7(32'h3a01eb74),
	.w8(32'h39baf001),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80b1b7),
	.w1(32'h3a64be7f),
	.w2(32'h3bac535c),
	.w3(32'hb72f1470),
	.w4(32'h39939af0),
	.w5(32'h3b095a71),
	.w6(32'h3a800fef),
	.w7(32'hba195f57),
	.w8(32'h3ad14d1d),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c8c3c9),
	.w1(32'hb8cb009e),
	.w2(32'hb8288bbe),
	.w3(32'hb77835fd),
	.w4(32'hb8225afa),
	.w5(32'hb7d22786),
	.w6(32'hb7d271a4),
	.w7(32'hb86bb85b),
	.w8(32'hb84977c7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb888d01d),
	.w1(32'hbb7f6efe),
	.w2(32'hbac0fcef),
	.w3(32'hbac72280),
	.w4(32'hbbac0105),
	.w5(32'hbb433bb4),
	.w6(32'hbb108b52),
	.w7(32'hbb467418),
	.w8(32'hbaf51f7a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule