module layer_10_featuremap_72(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d732),
	.w1(32'hba49f5a2),
	.w2(32'h3a20e4b9),
	.w3(32'h3aab0d9f),
	.w4(32'hbb0172d8),
	.w5(32'h3a333ae4),
	.w6(32'h3b8ca3e9),
	.w7(32'hba418db0),
	.w8(32'h3bff0cc0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc0614),
	.w1(32'hbb677807),
	.w2(32'hbae1caa7),
	.w3(32'hbba22450),
	.w4(32'hba82ec68),
	.w5(32'h396b2052),
	.w6(32'hba4528ad),
	.w7(32'h3b22292b),
	.w8(32'h3b063424),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becefa0),
	.w1(32'h3ab77ce4),
	.w2(32'h3ad42faa),
	.w3(32'h3c143130),
	.w4(32'h3af597b8),
	.w5(32'h3af9b451),
	.w6(32'h3becf43a),
	.w7(32'h3b05c4a9),
	.w8(32'hba7efb4a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70856c),
	.w1(32'h3ba480c5),
	.w2(32'h3ba9ebe4),
	.w3(32'h3a54e580),
	.w4(32'h3bc318e5),
	.w5(32'h3b8eb012),
	.w6(32'hbb424a9c),
	.w7(32'h3b394255),
	.w8(32'h37389d28),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ea2c4),
	.w1(32'hba0c57fb),
	.w2(32'h3b877c58),
	.w3(32'hbaa2b8bd),
	.w4(32'hbaa46066),
	.w5(32'h3b4ada8d),
	.w6(32'hbbd58502),
	.w7(32'hbbf37c22),
	.w8(32'hba19511f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208ac4),
	.w1(32'h3ac87481),
	.w2(32'h3ad99190),
	.w3(32'hbba3dd8c),
	.w4(32'h39c85986),
	.w5(32'hbbb98d77),
	.w6(32'hbb77a9cb),
	.w7(32'hba4dc7c2),
	.w8(32'h3a19a116),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9969a7),
	.w1(32'h3b99d86b),
	.w2(32'hbb4d28c4),
	.w3(32'h3b94b3ab),
	.w4(32'hbc0d4b7a),
	.w5(32'hbbba0aec),
	.w6(32'h390504b9),
	.w7(32'hbb3cce52),
	.w8(32'hbb8ff2f3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc939f74),
	.w1(32'hbbf13939),
	.w2(32'hbc891851),
	.w3(32'hbc577c01),
	.w4(32'hbbca6a9c),
	.w5(32'hbc241850),
	.w6(32'hbc9338f8),
	.w7(32'hbca7bdfc),
	.w8(32'hbcafdd69),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba327973),
	.w1(32'hbb0d14eb),
	.w2(32'hbb73d3b1),
	.w3(32'hb94f7006),
	.w4(32'hbb80054b),
	.w5(32'h3aa05011),
	.w6(32'h39575df8),
	.w7(32'hbb0d3eba),
	.w8(32'hba5786bd),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c4e4d),
	.w1(32'hbb9f0376),
	.w2(32'hbca5e2e2),
	.w3(32'h3c4bda7e),
	.w4(32'h3c482aa1),
	.w5(32'hb9879d42),
	.w6(32'h3c1ed671),
	.w7(32'h3c6094c2),
	.w8(32'hbb6392c9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd74f73),
	.w1(32'h3b77eec3),
	.w2(32'h3b40b16b),
	.w3(32'h3c709c7a),
	.w4(32'h3c32cd30),
	.w5(32'h3a193703),
	.w6(32'h3c0eab5d),
	.w7(32'h3bc6c7a9),
	.w8(32'h3a854118),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc34a4d),
	.w1(32'h3c888728),
	.w2(32'hbcfdee4e),
	.w3(32'h3ca8ea27),
	.w4(32'h3c3b8880),
	.w5(32'hbd0179ab),
	.w6(32'h3c092633),
	.w7(32'h3c5589d3),
	.w8(32'hbcb63ade),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5e778),
	.w1(32'hbcba26cc),
	.w2(32'hbcc2a76f),
	.w3(32'hbc4f366f),
	.w4(32'hbc920dd6),
	.w5(32'hbc8c966c),
	.w6(32'hbc49871a),
	.w7(32'hbc493bf8),
	.w8(32'hbc309d6b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb927c01),
	.w1(32'hbc4e8700),
	.w2(32'hbae3b0f5),
	.w3(32'hbc26507c),
	.w4(32'hbc6a08ea),
	.w5(32'hbbbca026),
	.w6(32'hbb781142),
	.w7(32'hbc46060f),
	.w8(32'hbb8547b6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3dea5),
	.w1(32'h3b811f69),
	.w2(32'h3b261c41),
	.w3(32'hbae7ab5b),
	.w4(32'h3b30e5bd),
	.w5(32'h3b42b5b6),
	.w6(32'h3b248c9d),
	.w7(32'h3bdb3df5),
	.w8(32'h3bd4db27),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80f1d7),
	.w1(32'hbc8327d3),
	.w2(32'hbcd8e788),
	.w3(32'h3b85f46a),
	.w4(32'hbb518676),
	.w5(32'hbc5b452b),
	.w6(32'hb98d137c),
	.w7(32'hbb889c95),
	.w8(32'hbc6fc914),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f84a6),
	.w1(32'h3b14209d),
	.w2(32'h3ac3a1ed),
	.w3(32'h3c2fb143),
	.w4(32'h3bfe627d),
	.w5(32'h3ae9face),
	.w6(32'h3bee80bf),
	.w7(32'h3bb0a544),
	.w8(32'h3b7967e3),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c053718),
	.w1(32'hbbc3cda1),
	.w2(32'hbcaf8595),
	.w3(32'h3bab6de1),
	.w4(32'h3b3efc48),
	.w5(32'hbc7f252b),
	.w6(32'hbbcc428d),
	.w7(32'h3a95dd6a),
	.w8(32'hbc8989cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d8919d),
	.w1(32'hbc2886a1),
	.w2(32'hbb83540b),
	.w3(32'h3b25975c),
	.w4(32'hbae5f21a),
	.w5(32'hbaed0ab6),
	.w6(32'hbb7b4e5c),
	.w7(32'hbb301b79),
	.w8(32'h3b093909),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babddbe),
	.w1(32'h3b9eac68),
	.w2(32'hbb09422d),
	.w3(32'hba561b30),
	.w4(32'h3b6a9d28),
	.w5(32'hbb1210fb),
	.w6(32'h3afd4fd7),
	.w7(32'h3b325529),
	.w8(32'hbb4a4b95),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa77e6),
	.w1(32'hbaedd529),
	.w2(32'h3acea5ef),
	.w3(32'h39be0543),
	.w4(32'hbb258aa0),
	.w5(32'hbaf261de),
	.w6(32'hb73216f6),
	.w7(32'hbb36e7a1),
	.w8(32'h390f7c1a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb223acf),
	.w1(32'hbabb14e6),
	.w2(32'h3b667a80),
	.w3(32'h378f7c8c),
	.w4(32'h3b6af192),
	.w5(32'h3b9a317b),
	.w6(32'h3a4912a1),
	.w7(32'h3b8b89f5),
	.w8(32'h3bda2df3),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b238389),
	.w1(32'hbb31fabb),
	.w2(32'hbd1a180b),
	.w3(32'h3b28e833),
	.w4(32'h3c55cc19),
	.w5(32'hbc2d5699),
	.w6(32'h3b9bb29f),
	.w7(32'h3c9e619f),
	.w8(32'hbccd2670),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb134c1),
	.w1(32'hbbdcf8c9),
	.w2(32'hbc6986df),
	.w3(32'h3beb2e7e),
	.w4(32'h3bd979ad),
	.w5(32'hbb9c546e),
	.w6(32'h3b9daacd),
	.w7(32'h3baa9d5f),
	.w8(32'hbb1564c2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e1387),
	.w1(32'hbb91864b),
	.w2(32'hbba6f760),
	.w3(32'hbc74efe7),
	.w4(32'hbbed7f84),
	.w5(32'hbb0b7576),
	.w6(32'hbbe9d0d4),
	.w7(32'hbb1dea3b),
	.w8(32'h3b9e88e4),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a5564),
	.w1(32'h3b0a9175),
	.w2(32'hbac9a07f),
	.w3(32'hbbc50b75),
	.w4(32'hbaee858e),
	.w5(32'hb9fef2fc),
	.w6(32'hbb48f5d4),
	.w7(32'hbae31256),
	.w8(32'h3b197365),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bdc50),
	.w1(32'h3a67bb97),
	.w2(32'h3a89f6e2),
	.w3(32'hbb591f67),
	.w4(32'hba23f664),
	.w5(32'h3b9b6140),
	.w6(32'hb9f2c814),
	.w7(32'hb9e48f8a),
	.w8(32'h3a5d3eb4),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820fba),
	.w1(32'hbb9b1a7c),
	.w2(32'h3bbce212),
	.w3(32'h3bb8f0aa),
	.w4(32'hba0ef793),
	.w5(32'h3c064136),
	.w6(32'h3c9a6b53),
	.w7(32'h3b35645a),
	.w8(32'h3cb9cf23),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8c2f4),
	.w1(32'h3c526a41),
	.w2(32'hbc7004cf),
	.w3(32'h3c0ae671),
	.w4(32'h3c2158a1),
	.w5(32'hbc695992),
	.w6(32'h3b3045c2),
	.w7(32'h3bbdeb39),
	.w8(32'h3b0a5a90),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0da4ca),
	.w1(32'hbbc4238f),
	.w2(32'h3c11dc04),
	.w3(32'hbc620f42),
	.w4(32'hbcc5086b),
	.w5(32'h3c5ed348),
	.w6(32'h3cbe9852),
	.w7(32'h3bb6d8e5),
	.w8(32'h3c94be17),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9bb16),
	.w1(32'h3b66cbe7),
	.w2(32'h3b68ee2a),
	.w3(32'h3c644144),
	.w4(32'h3c25bfab),
	.w5(32'h3c5bad92),
	.w6(32'h3c305116),
	.w7(32'h3c2697e4),
	.w8(32'hbb299ecb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc9b83d),
	.w1(32'hbb8f9567),
	.w2(32'hbad2e405),
	.w3(32'h3c2bd9dc),
	.w4(32'hbbbf8a8b),
	.w5(32'hbbda91da),
	.w6(32'h3b8563e6),
	.w7(32'h3b3942a9),
	.w8(32'h3a9540d1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a5ad),
	.w1(32'h3a71ad2a),
	.w2(32'hbbfda776),
	.w3(32'h3b883eac),
	.w4(32'hba3deeae),
	.w5(32'hbba5b4fd),
	.w6(32'hb9df12a5),
	.w7(32'h3bcf098c),
	.w8(32'hbaedecb9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb091),
	.w1(32'hbb2fb582),
	.w2(32'hbb2d4c61),
	.w3(32'hbc1f0425),
	.w4(32'hbbab71ad),
	.w5(32'h3c4e69c6),
	.w6(32'hbb18885a),
	.w7(32'hbabdb0b2),
	.w8(32'h3b7ab8db),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac830),
	.w1(32'h3c390245),
	.w2(32'hbc19d3bb),
	.w3(32'h3cc2e75d),
	.w4(32'h3b77a02a),
	.w5(32'hbc89c442),
	.w6(32'hbc051687),
	.w7(32'hbc932c40),
	.w8(32'hbc189c86),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5403bb0),
	.w1(32'hbb09abf4),
	.w2(32'hbb84d980),
	.w3(32'hbc1c2d1c),
	.w4(32'hbc48e283),
	.w5(32'hbb0135ec),
	.w6(32'hbc5c1837),
	.w7(32'hbc87a254),
	.w8(32'hbc973603),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c636bfb),
	.w1(32'h3bbb409a),
	.w2(32'hbd2ac092),
	.w3(32'h3bddce69),
	.w4(32'h3c257d70),
	.w5(32'hbc812c24),
	.w6(32'hbccdbf57),
	.w7(32'h3c121881),
	.w8(32'hbc672205),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca82ccb),
	.w1(32'h3c5d38b0),
	.w2(32'hbc528158),
	.w3(32'h3c066eed),
	.w4(32'h3ce942ab),
	.w5(32'h3ad6adf3),
	.w6(32'h3cb03726),
	.w7(32'h3d12bffc),
	.w8(32'h3c97bbf0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b5ee7),
	.w1(32'hbc3dae64),
	.w2(32'hbc196ef2),
	.w3(32'h3b0be8ba),
	.w4(32'hbcaf6db2),
	.w5(32'hbbdee997),
	.w6(32'h3c40ece2),
	.w7(32'h3c274077),
	.w8(32'h3c939e25),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc291417),
	.w1(32'h3b37eb78),
	.w2(32'hbbb60b4e),
	.w3(32'hbcd87a23),
	.w4(32'hbb95b942),
	.w5(32'hbb9b7f02),
	.w6(32'hbb621e9c),
	.w7(32'h3bac82bb),
	.w8(32'h3c093e77),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4453f7),
	.w1(32'hbaaedcb6),
	.w2(32'hbbfb5db2),
	.w3(32'hbc73cb03),
	.w4(32'hbc138fe4),
	.w5(32'hbc6e18d9),
	.w6(32'hbbd2b21f),
	.w7(32'hbaf1648f),
	.w8(32'hbbd191f4),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43e9d4),
	.w1(32'hbbfe8b12),
	.w2(32'h3b89c0d0),
	.w3(32'hbca6383b),
	.w4(32'hbc01438a),
	.w5(32'h3c7f39ba),
	.w6(32'hbc448833),
	.w7(32'hbb72445e),
	.w8(32'h3c1a4ad9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4fe87),
	.w1(32'h390ebf9a),
	.w2(32'hbb146e5d),
	.w3(32'h3ce1526d),
	.w4(32'h3c8b5e2f),
	.w5(32'hbbaa25a3),
	.w6(32'h3ccdd3ff),
	.w7(32'h3c976098),
	.w8(32'hb8a4e362),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b870c62),
	.w1(32'hbba26bf4),
	.w2(32'hbcac9074),
	.w3(32'h3bf15733),
	.w4(32'h3c237be5),
	.w5(32'hbc1cb95a),
	.w6(32'hbb30a4bc),
	.w7(32'h38d47196),
	.w8(32'hbc1c7870),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf867f2),
	.w1(32'h3af6bda4),
	.w2(32'hbcea5d18),
	.w3(32'h3bae6e74),
	.w4(32'h3b918541),
	.w5(32'hbd1e5517),
	.w6(32'h3ca72fcf),
	.w7(32'h3ca88e97),
	.w8(32'hbc35098e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7a168),
	.w1(32'hbc707e12),
	.w2(32'h3ba83b63),
	.w3(32'hbcef7142),
	.w4(32'hbb26e863),
	.w5(32'h3c301dd7),
	.w6(32'hb9f2a8b6),
	.w7(32'h3c66961e),
	.w8(32'hbaf501ec),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2daed8),
	.w1(32'hb958cd6e),
	.w2(32'hbc61997e),
	.w3(32'h3caed89f),
	.w4(32'h3c6a7950),
	.w5(32'hbb288cc3),
	.w6(32'h3bde0ba6),
	.w7(32'h3c7d34e3),
	.w8(32'hbbd573dc),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7747e),
	.w1(32'hbc925f61),
	.w2(32'hbc9fd40b),
	.w3(32'h3b6683f0),
	.w4(32'hbc2d711a),
	.w5(32'hbc0dd889),
	.w6(32'hbc407acc),
	.w7(32'hbc06873d),
	.w8(32'hbc0f9726),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9a3b1),
	.w1(32'h3c0c6ebb),
	.w2(32'hbb2e3155),
	.w3(32'h3bcc305f),
	.w4(32'h3bfe56b9),
	.w5(32'h3c4833f8),
	.w6(32'h3b90a671),
	.w7(32'h3bb5ad94),
	.w8(32'h3bc6e337),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc7798),
	.w1(32'hb7e5b31b),
	.w2(32'h3bdf006f),
	.w3(32'h3c8df151),
	.w4(32'h3bb8f8be),
	.w5(32'h3ba486ef),
	.w6(32'h3b7e1c83),
	.w7(32'h3b60ec83),
	.w8(32'h3aa93ea7),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08d397),
	.w1(32'hbc1f6867),
	.w2(32'h3c9cd53b),
	.w3(32'hbcb5a6af),
	.w4(32'hbd01fb5b),
	.w5(32'h3c014163),
	.w6(32'hbd0cc08a),
	.w7(32'hbcd0c2ab),
	.w8(32'hbbecfe88),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8078d),
	.w1(32'hbbc7c249),
	.w2(32'hbc09fb15),
	.w3(32'hbc40ab64),
	.w4(32'h3c504c02),
	.w5(32'hbcb08019),
	.w6(32'hbb6dc93e),
	.w7(32'h3c504b7b),
	.w8(32'hbc9c2408),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdd8b),
	.w1(32'hbc96ab2a),
	.w2(32'hbb946ab0),
	.w3(32'hbd512904),
	.w4(32'hbd4685aa),
	.w5(32'h3b5c2e9f),
	.w6(32'hbd43c10e),
	.w7(32'hbcf471b0),
	.w8(32'hba0dc6f2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b3f53),
	.w1(32'hbc30c6ca),
	.w2(32'hbcb8d07c),
	.w3(32'h3c8b0e2c),
	.w4(32'h3b642e7b),
	.w5(32'hbc03bd46),
	.w6(32'hb87805ba),
	.w7(32'h3b0532e4),
	.w8(32'hbc1104d7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb773e91),
	.w1(32'hbc2596e9),
	.w2(32'hbbb785c4),
	.w3(32'h3b0b1d44),
	.w4(32'h3b41af46),
	.w5(32'h3b825236),
	.w6(32'h3ba41906),
	.w7(32'h3a167d96),
	.w8(32'hba8e6d3d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16dc6e),
	.w1(32'h3c0735bd),
	.w2(32'hbbaada03),
	.w3(32'h3bb1f1e1),
	.w4(32'hbb0b51c5),
	.w5(32'h3b48c01c),
	.w6(32'h3be4ec53),
	.w7(32'h3c26e983),
	.w8(32'h3bec7735),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87fbd18),
	.w1(32'h3aa58159),
	.w2(32'h3bc26e6f),
	.w3(32'h3b8675ab),
	.w4(32'hbadefef8),
	.w5(32'hba4b1c4a),
	.w6(32'h3c51d49a),
	.w7(32'h3bd81732),
	.w8(32'hbaba2c88),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b52fb89),
	.w1(32'hbb891f59),
	.w2(32'hbb293c39),
	.w3(32'hbb6b7178),
	.w4(32'hbb8478e7),
	.w5(32'hbbc4b480),
	.w6(32'h3a72e2f2),
	.w7(32'h3a65c113),
	.w8(32'h3b9ae22e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb823ef3),
	.w1(32'h3be8cb74),
	.w2(32'h3b21602b),
	.w3(32'hbbf19812),
	.w4(32'h3bc956ce),
	.w5(32'hbc145420),
	.w6(32'h3bc44804),
	.w7(32'h3c93cc50),
	.w8(32'hba8187b3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28c52),
	.w1(32'hbb879d20),
	.w2(32'h39f98895),
	.w3(32'hbc8c1049),
	.w4(32'hbc319ee4),
	.w5(32'h3b14c781),
	.w6(32'hbbfc8040),
	.w7(32'hbbef8ea1),
	.w8(32'hba0f9269),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad53ce9),
	.w1(32'h3a6bb8af),
	.w2(32'hbc22f37b),
	.w3(32'h3b877ed7),
	.w4(32'h3bc2fe5e),
	.w5(32'h3ae61d70),
	.w6(32'h3b335bfa),
	.w7(32'h3bbbe421),
	.w8(32'hbba6fc77),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed699),
	.w1(32'hbb8a48d1),
	.w2(32'hbd12968b),
	.w3(32'h3c47c0fd),
	.w4(32'h3bdfda4c),
	.w5(32'hbc8f39ea),
	.w6(32'h3b66a654),
	.w7(32'h3ba951fb),
	.w8(32'h3aa2dd85),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4cc519),
	.w1(32'hbba6b956),
	.w2(32'h3c09ddb1),
	.w3(32'h3c4bed05),
	.w4(32'h3c0594f4),
	.w5(32'h3c32f102),
	.w6(32'h3c938c3f),
	.w7(32'hba496e3c),
	.w8(32'h3bf5396e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30c61b),
	.w1(32'h3b1e8230),
	.w2(32'h39166d06),
	.w3(32'h3cc449ee),
	.w4(32'h3c3cab9c),
	.w5(32'hbc3967a2),
	.w6(32'h3c1c9d6e),
	.w7(32'h3a63324b),
	.w8(32'hbc7c4a4d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc327981),
	.w1(32'hbc522a13),
	.w2(32'hbbc22f7b),
	.w3(32'hbcfd6d68),
	.w4(32'hbc73404f),
	.w5(32'hbc1c95d2),
	.w6(32'hbcf518c4),
	.w7(32'hbcbce4c5),
	.w8(32'hbc0f5e5a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8eecab),
	.w1(32'hbba413b2),
	.w2(32'h3bfa0824),
	.w3(32'hbc0badca),
	.w4(32'hbba08c27),
	.w5(32'h3c18b9da),
	.w6(32'hbc45182d),
	.w7(32'hbc133397),
	.w8(32'h3c09963f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd6c2fc),
	.w1(32'hbc9453a4),
	.w2(32'hbd1e1371),
	.w3(32'h3cd9fcc6),
	.w4(32'h3c28e774),
	.w5(32'hbcb76173),
	.w6(32'h3caca129),
	.w7(32'h3c2aabf4),
	.w8(32'hbc73b91b),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1d252),
	.w1(32'hbb6c412c),
	.w2(32'hbd0ffaad),
	.w3(32'hbcee0ead),
	.w4(32'hbcadc984),
	.w5(32'hbd6e1ce5),
	.w6(32'hbc97e286),
	.w7(32'hbccfc313),
	.w8(32'hbd885c49),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd10b352),
	.w1(32'hbd0b1b4c),
	.w2(32'hbc679150),
	.w3(32'hbd7d76dc),
	.w4(32'hbd44932c),
	.w5(32'hbb42d638),
	.w6(32'hbd3c7d0d),
	.w7(32'hbd22f60c),
	.w8(32'hbb60c4df),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c49d3),
	.w1(32'h3c66695e),
	.w2(32'hbbe49e03),
	.w3(32'h3b8c6d72),
	.w4(32'h3cb1abc0),
	.w5(32'h3c615b2d),
	.w6(32'h3c4d113f),
	.w7(32'h3cc58b02),
	.w8(32'h3c0b87c9),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e05ef),
	.w1(32'h3c7b0f97),
	.w2(32'hbbaaf2de),
	.w3(32'h3c1e26ad),
	.w4(32'h3c132484),
	.w5(32'hbb22f053),
	.w6(32'h3b1f9c29),
	.w7(32'h3c209ca7),
	.w8(32'hbb57de4c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4b0519),
	.w1(32'hbbe134ee),
	.w2(32'h3c7019b7),
	.w3(32'hbc006146),
	.w4(32'hbbc44f8c),
	.w5(32'h3c674a4a),
	.w6(32'hbb9d0e7f),
	.w7(32'hbb149649),
	.w8(32'h3a6dd5a0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbeb710),
	.w1(32'h3c83aa9d),
	.w2(32'hba983880),
	.w3(32'h3ceb998e),
	.w4(32'h3ca32e6f),
	.w5(32'h3b9d34ef),
	.w6(32'h3c647e19),
	.w7(32'h3c687837),
	.w8(32'h3bb65a18),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcea77),
	.w1(32'h3b1b69e3),
	.w2(32'h3ba97a89),
	.w3(32'h3ca53095),
	.w4(32'h3cb8d467),
	.w5(32'h3bbb7fb3),
	.w6(32'h3c482f71),
	.w7(32'h3caa45a8),
	.w8(32'h3c0dca10),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8dafb),
	.w1(32'h3b956fd1),
	.w2(32'hbc9fc74b),
	.w3(32'h3beb3235),
	.w4(32'h3beda55e),
	.w5(32'hbcc9bf41),
	.w6(32'h3bc9c073),
	.w7(32'h3bbfa1c4),
	.w8(32'hbc8765dc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbf6a04),
	.w1(32'hbca8378f),
	.w2(32'hbc20435b),
	.w3(32'hbd0d285d),
	.w4(32'hbca74a3c),
	.w5(32'hbbd0a0d5),
	.w6(32'hbcf6d829),
	.w7(32'hbc06a5ef),
	.w8(32'hbcd12490),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c953c06),
	.w1(32'h3c653e5f),
	.w2(32'h3a858af8),
	.w3(32'hbc618d49),
	.w4(32'hbc70424c),
	.w5(32'hbaa3b8da),
	.w6(32'hbd3ccbac),
	.w7(32'hbcec9162),
	.w8(32'hbc0ce242),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9aa9d2),
	.w1(32'hbbe49ced),
	.w2(32'hbcaba451),
	.w3(32'hbc670e4e),
	.w4(32'hbc9f6df4),
	.w5(32'hbcad2d5d),
	.w6(32'hbc8270e3),
	.w7(32'hbc657749),
	.w8(32'hbba36dbd),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8b94),
	.w1(32'hbc0ca9ab),
	.w2(32'hbc1c57ac),
	.w3(32'h3b173221),
	.w4(32'h3aa60eca),
	.w5(32'hbb774aa3),
	.w6(32'h3b3974c4),
	.w7(32'h3bfca2f2),
	.w8(32'hbbf384be),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ee5cb),
	.w1(32'h3a024b28),
	.w2(32'hba622ba3),
	.w3(32'h3beb479c),
	.w4(32'h3bde8525),
	.w5(32'hbba6ea18),
	.w6(32'h3be081a2),
	.w7(32'h3bd1c7a4),
	.w8(32'hbbf553dd),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f9d46),
	.w1(32'h3baf21a3),
	.w2(32'hbbef64ce),
	.w3(32'h3bf3cf01),
	.w4(32'hba1590bf),
	.w5(32'hbba3795e),
	.w6(32'hbaaf0c74),
	.w7(32'hbbabd442),
	.w8(32'hbbc4650e),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b034aff),
	.w1(32'hbc4e3341),
	.w2(32'h3b2d5168),
	.w3(32'h3b998d1d),
	.w4(32'hbb1c8bbc),
	.w5(32'h3c07623e),
	.w6(32'hb88ec5d6),
	.w7(32'hbafc0d45),
	.w8(32'hb815cdfa),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c377582),
	.w1(32'h3aac38de),
	.w2(32'hbbb2b5f6),
	.w3(32'h3c4f8a1f),
	.w4(32'h3bd030b1),
	.w5(32'hbc1a9587),
	.w6(32'h3afcc149),
	.w7(32'h3b3e655d),
	.w8(32'hbbd8b035),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4862a3),
	.w1(32'hbbbe5645),
	.w2(32'h3c6b5c06),
	.w3(32'hbc078fc6),
	.w4(32'hbc38cab1),
	.w5(32'h3c3f4926),
	.w6(32'hbc59f7bd),
	.w7(32'hbb86ced3),
	.w8(32'h3bdda65a),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c955281),
	.w1(32'h3c626da5),
	.w2(32'h3c6d02e0),
	.w3(32'h3cc81f4b),
	.w4(32'h3c987691),
	.w5(32'h3b94dd7c),
	.w6(32'h3c97be57),
	.w7(32'h3c7eb2f2),
	.w8(32'hbc970139),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00a1f3),
	.w1(32'hbb2a283c),
	.w2(32'hb92950be),
	.w3(32'hbc067075),
	.w4(32'hbb783ffd),
	.w5(32'hba311df2),
	.w6(32'hbcaf4844),
	.w7(32'h3c4d3c0e),
	.w8(32'h38ec2292),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2023cf),
	.w1(32'hbb497d1c),
	.w2(32'hbc1de15d),
	.w3(32'hbc44f259),
	.w4(32'h3adad16d),
	.w5(32'hbbb7532b),
	.w6(32'hbc1cabe1),
	.w7(32'hb99582bb),
	.w8(32'h392076fb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ea557),
	.w1(32'hba947347),
	.w2(32'h3bfce8f0),
	.w3(32'hbbf3513a),
	.w4(32'hbbbf62ad),
	.w5(32'hbaf61afc),
	.w6(32'hbb8d33aa),
	.w7(32'h3a1cf622),
	.w8(32'hbbc4f924),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf81ad),
	.w1(32'hbc2036de),
	.w2(32'hbb5eda62),
	.w3(32'hbd0c18d7),
	.w4(32'hbcfe2c22),
	.w5(32'h3b8f8adc),
	.w6(32'hbd148d9f),
	.w7(32'hbcbbd513),
	.w8(32'h38129be4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb034f23),
	.w1(32'hbbe0a727),
	.w2(32'hbc4c500b),
	.w3(32'h3b29dc17),
	.w4(32'h3aeb1abc),
	.w5(32'hbc69ed1e),
	.w6(32'hbc15685c),
	.w7(32'h3b6a4d81),
	.w8(32'hbc3b53a7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018b0d),
	.w1(32'h3b26d1a5),
	.w2(32'h3b0d4f5b),
	.w3(32'hbc5d0218),
	.w4(32'h3b21dc4d),
	.w5(32'h3c1ed5c8),
	.w6(32'h39969349),
	.w7(32'h3c63cac5),
	.w8(32'h3ce51d79),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeac8a),
	.w1(32'h3a50266a),
	.w2(32'hbcefbdee),
	.w3(32'h3ced6480),
	.w4(32'h3c64afdf),
	.w5(32'hbc853f96),
	.w6(32'h3c99dea8),
	.w7(32'h3b6c0aa1),
	.w8(32'hbc4a021b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfab098),
	.w1(32'h3c2558de),
	.w2(32'h3c0fb2ac),
	.w3(32'hbadeaa94),
	.w4(32'h3c818648),
	.w5(32'h3c0b705a),
	.w6(32'h38fd1468),
	.w7(32'h3ca7fbe5),
	.w8(32'h3c213970),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ec575),
	.w1(32'hbc028c6e),
	.w2(32'hbd364ae6),
	.w3(32'h3b744a78),
	.w4(32'hbb794a49),
	.w5(32'hbd5c69bc),
	.w6(32'hbb9126dd),
	.w7(32'hbb5d4631),
	.w8(32'hbd4ffdab),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd053859),
	.w1(32'hbd086dc8),
	.w2(32'hbc7fc193),
	.w3(32'hbd8b43bf),
	.w4(32'hbd6f9cb7),
	.w5(32'hbab7b009),
	.w6(32'hbd5ab137),
	.w7(32'hbd33be94),
	.w8(32'h3c07213f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7499bb),
	.w1(32'h3c1db48e),
	.w2(32'h3b60bbd1),
	.w3(32'h3ad03124),
	.w4(32'h3b9eba97),
	.w5(32'h3b8204a0),
	.w6(32'h3b124c56),
	.w7(32'h3bdb1615),
	.w8(32'h3cbd9340),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ebd89),
	.w1(32'hbb55fbc1),
	.w2(32'hb93489d9),
	.w3(32'hbc5100cc),
	.w4(32'hbbb5b643),
	.w5(32'h3afc9a97),
	.w6(32'h3b037de0),
	.w7(32'h3c1248ad),
	.w8(32'h3bb51bd8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42d44b),
	.w1(32'hbb9d945a),
	.w2(32'h3c02e51a),
	.w3(32'h3b157bca),
	.w4(32'h3bedca7a),
	.w5(32'h3ce5e081),
	.w6(32'h3c4ffc08),
	.w7(32'h3889a80d),
	.w8(32'hba5ea6e5),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d4bf5cf),
	.w1(32'h3c9ed813),
	.w2(32'hbc4121f7),
	.w3(32'h3d629708),
	.w4(32'h3c9e6ff8),
	.w5(32'hbbd618d0),
	.w6(32'h3cdff67e),
	.w7(32'h3bdfa6ee),
	.w8(32'hbba73edb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda85af),
	.w1(32'h3c34df0b),
	.w2(32'hbbd23128),
	.w3(32'hbcc927dd),
	.w4(32'hbc0ab3b2),
	.w5(32'hbc4b4680),
	.w6(32'hbcb8f9ba),
	.w7(32'h3c245165),
	.w8(32'hbc9bc3dd),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990b25b),
	.w1(32'h3cde862d),
	.w2(32'h3c6f3100),
	.w3(32'h3a9c989a),
	.w4(32'h3d1ff12f),
	.w5(32'h3cca33e7),
	.w6(32'h3c9ad0fb),
	.w7(32'h3d4c59ce),
	.w8(32'h3d2d83c7),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9003),
	.w1(32'h3a297094),
	.w2(32'hbac9d016),
	.w3(32'hbb2b859e),
	.w4(32'h3bfd1663),
	.w5(32'h3b13a0f9),
	.w6(32'hba86b9e0),
	.w7(32'h3be52b8c),
	.w8(32'h3a7c33b8),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95cc56),
	.w1(32'h3c2e23b0),
	.w2(32'hbbaf7818),
	.w3(32'h3cd83572),
	.w4(32'h3c8c69be),
	.w5(32'hbc01f3d1),
	.w6(32'hba9d9964),
	.w7(32'h3c967d2c),
	.w8(32'hbc2955a0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9260c),
	.w1(32'hbab082b2),
	.w2(32'h3c8e1ad0),
	.w3(32'h3bdbc9cf),
	.w4(32'hba0c3fa1),
	.w5(32'h3c30c73d),
	.w6(32'hbc049130),
	.w7(32'hbb4ad417),
	.w8(32'hbc218302),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb5c9a),
	.w1(32'hbbe69e20),
	.w2(32'hbc4bc25a),
	.w3(32'hbb7ce396),
	.w4(32'h3b3f29d7),
	.w5(32'hbb8efd69),
	.w6(32'hbd1b019c),
	.w7(32'hbaac6955),
	.w8(32'hbccdd57d),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c700269),
	.w1(32'h3c554e6e),
	.w2(32'hbbe88397),
	.w3(32'h3c8c91af),
	.w4(32'h3bd07536),
	.w5(32'h383a3a9a),
	.w6(32'h3b5d5ae2),
	.w7(32'h3c4663a5),
	.w8(32'hbba6f1d2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be614df),
	.w1(32'h3a639d57),
	.w2(32'hbc224c94),
	.w3(32'h3bc96ca5),
	.w4(32'h3b1accbe),
	.w5(32'hbc14f3ef),
	.w6(32'h39325653),
	.w7(32'h3b9c8a2c),
	.w8(32'h3b42d738),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b3b71),
	.w1(32'hbc2c0029),
	.w2(32'h3be08417),
	.w3(32'hbc80c795),
	.w4(32'hbb8bf029),
	.w5(32'h3c66810b),
	.w6(32'hbb941c4f),
	.w7(32'hbb87b005),
	.w8(32'h3bd27cf0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c433332),
	.w1(32'hbaf9a4e1),
	.w2(32'hbc3e9ab8),
	.w3(32'h3cbd2fc3),
	.w4(32'h3c504ee5),
	.w5(32'h3bb06c7b),
	.w6(32'h3cce9747),
	.w7(32'h3c8467f4),
	.w8(32'hbba46347),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ebf9b),
	.w1(32'hba907ed8),
	.w2(32'hbbcf6b03),
	.w3(32'h3c7c5ed6),
	.w4(32'h3c161003),
	.w5(32'h3bed1298),
	.w6(32'h3bc2dd36),
	.w7(32'h3b019d16),
	.w8(32'h3c76d3fb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3082b7),
	.w1(32'h3b3d417f),
	.w2(32'h3c89a414),
	.w3(32'h3bed64f7),
	.w4(32'h3c44e05d),
	.w5(32'h3cd67b60),
	.w6(32'h3c738769),
	.w7(32'h3cc079a9),
	.w8(32'h3baabdc3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83ebe9),
	.w1(32'hbb9f1f71),
	.w2(32'hbabda6c6),
	.w3(32'h3c9ff20a),
	.w4(32'h3b9019fd),
	.w5(32'h3c5348f1),
	.w6(32'h39920d63),
	.w7(32'hbb998a18),
	.w8(32'h3b230730),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb74aea),
	.w1(32'h3cbd8a0b),
	.w2(32'hbbdb614e),
	.w3(32'h3c9de25c),
	.w4(32'h3c07d370),
	.w5(32'hbbdc7f64),
	.w6(32'hbc7887cb),
	.w7(32'hbc7f614a),
	.w8(32'hbbddc72c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc946350),
	.w1(32'hbcebbe6f),
	.w2(32'hbcbb8f77),
	.w3(32'hbb273817),
	.w4(32'hbc653280),
	.w5(32'hbc3725d7),
	.w6(32'h3c10ce89),
	.w7(32'h3ba376b3),
	.w8(32'hbc261f93),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac0f77),
	.w1(32'h3b9f7aaa),
	.w2(32'hbba80844),
	.w3(32'h3c30ef0c),
	.w4(32'h3ad13eec),
	.w5(32'h3a9fde73),
	.w6(32'h3c0e53a5),
	.w7(32'hbbd042a1),
	.w8(32'h3b1a58ed),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b1c2),
	.w1(32'hb971d7cb),
	.w2(32'hbbac4f68),
	.w3(32'hbbb28d94),
	.w4(32'hbac9e490),
	.w5(32'hb9ec5a72),
	.w6(32'hbbbeba93),
	.w7(32'hbbc9c315),
	.w8(32'h3bcef46a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2344),
	.w1(32'h3b907615),
	.w2(32'h3b8eeb23),
	.w3(32'h3be78a2f),
	.w4(32'h3ba5674d),
	.w5(32'hba3a1af2),
	.w6(32'h3b5772b7),
	.w7(32'h3b368578),
	.w8(32'h3b6b62b1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf9cfe),
	.w1(32'h3b391bba),
	.w2(32'h3c60452c),
	.w3(32'hba8ed380),
	.w4(32'hbab205ba),
	.w5(32'h3ca14384),
	.w6(32'h3bc5bb09),
	.w7(32'h3b9e529f),
	.w8(32'h3c050cde),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca69f30),
	.w1(32'hbb91e820),
	.w2(32'h3c3a117d),
	.w3(32'h3c052591),
	.w4(32'hbab347f2),
	.w5(32'h3c2cf941),
	.w6(32'h3ace22a4),
	.w7(32'hbbe52ec7),
	.w8(32'h3c41a7a5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf0b66),
	.w1(32'h3bc3dcb9),
	.w2(32'hbc736f0e),
	.w3(32'h3cb4326c),
	.w4(32'h3c803386),
	.w5(32'hbbab08d2),
	.w6(32'h3ba96c02),
	.w7(32'h3c466614),
	.w8(32'h3b6c7815),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45b0af),
	.w1(32'h3a796f0c),
	.w2(32'hbb71ab2b),
	.w3(32'hba24362e),
	.w4(32'h3c1cbebe),
	.w5(32'hba5dd704),
	.w6(32'h3c4b7ac9),
	.w7(32'h3bd41580),
	.w8(32'h3b69c6c4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4f4df),
	.w1(32'hbafd77d6),
	.w2(32'hbbb75043),
	.w3(32'h3bd72b8e),
	.w4(32'h3be79726),
	.w5(32'h3adddc5c),
	.w6(32'h3bb45c39),
	.w7(32'h3bb12b8c),
	.w8(32'h3aae2321),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc349956),
	.w1(32'hbb489efe),
	.w2(32'h3b9933a6),
	.w3(32'hbc0eea1e),
	.w4(32'hbc461bb7),
	.w5(32'h3b7e92c3),
	.w6(32'hba71d41e),
	.w7(32'hba1baa64),
	.w8(32'h3c2ebdda),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a1c5d),
	.w1(32'h3c8f3334),
	.w2(32'hb9d83c82),
	.w3(32'h3b9caa9f),
	.w4(32'h3c05feb3),
	.w5(32'h3b5d1e44),
	.w6(32'h3b5f7671),
	.w7(32'hbaf30a02),
	.w8(32'h3be6b545),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1dfbb),
	.w1(32'h3bbfd861),
	.w2(32'h3ce2822a),
	.w3(32'h3c5c9bf8),
	.w4(32'h3c05d34a),
	.w5(32'h3ca13ccc),
	.w6(32'h3c4e269b),
	.w7(32'h3c34739d),
	.w8(32'hbc2a260c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccb16fd),
	.w1(32'h3b32f797),
	.w2(32'h3c872334),
	.w3(32'h3c143d08),
	.w4(32'h396190b0),
	.w5(32'h3c31209e),
	.w6(32'hbc53636a),
	.w7(32'hbc379a60),
	.w8(32'hb9f04279),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86894e),
	.w1(32'h3aee25b4),
	.w2(32'h3c6c8f15),
	.w3(32'hbb3a777e),
	.w4(32'hbc0af250),
	.w5(32'h3c3c2a90),
	.w6(32'hbc464db5),
	.w7(32'hbcb4d0ad),
	.w8(32'hbb7af938),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d409610),
	.w1(32'h3cbc1c03),
	.w2(32'hbc940953),
	.w3(32'h3c3fc771),
	.w4(32'hbc510899),
	.w5(32'hbd152e82),
	.w6(32'hbc7794e3),
	.w7(32'hbc1907bb),
	.w8(32'hbd044ec8),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b1bb7),
	.w1(32'hbcae3944),
	.w2(32'hbcc1dcec),
	.w3(32'hbc47b0c7),
	.w4(32'hbc26711a),
	.w5(32'hbc7c34f1),
	.w6(32'hbaced610),
	.w7(32'h3a883bdc),
	.w8(32'hbccd5d33),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ced75),
	.w1(32'hba00d0cd),
	.w2(32'hbc856614),
	.w3(32'hba65e8cd),
	.w4(32'h3c4b76eb),
	.w5(32'hbbc8ed79),
	.w6(32'hbc7a8907),
	.w7(32'h3c4df691),
	.w8(32'h3bb38670),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc964b7f),
	.w1(32'hbc4c2cfe),
	.w2(32'h3b094994),
	.w3(32'h3c568fbc),
	.w4(32'h3c404756),
	.w5(32'h3c83a848),
	.w6(32'h3c544a56),
	.w7(32'h3bdf8d53),
	.w8(32'h3c463028),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befb811),
	.w1(32'h3ba0ee0c),
	.w2(32'h3c8a938e),
	.w3(32'h3cb052de),
	.w4(32'h3c8576df),
	.w5(32'h39798f92),
	.w6(32'h3d077e4a),
	.w7(32'h3cdd5f33),
	.w8(32'hbb8226c8),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbcf6c),
	.w1(32'hbbdeb2d9),
	.w2(32'hba19c0ea),
	.w3(32'hbb936067),
	.w4(32'h39f8fa37),
	.w5(32'hbbf4c76a),
	.w6(32'hbbf9b0aa),
	.w7(32'h3bc4791f),
	.w8(32'hbc206d1f),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bb85c),
	.w1(32'hbc605310),
	.w2(32'hbc164f3a),
	.w3(32'hbaf787d9),
	.w4(32'hbc830f1a),
	.w5(32'hbbfd4da0),
	.w6(32'h3b338dff),
	.w7(32'h3b9ec3cb),
	.w8(32'hbb2ccaf1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50295c),
	.w1(32'hbc116c90),
	.w2(32'hbc63f0d4),
	.w3(32'h3c1fda17),
	.w4(32'h3ba4259d),
	.w5(32'hba0e7575),
	.w6(32'h3b26e29c),
	.w7(32'h39b05d14),
	.w8(32'hbba61695),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38642e60),
	.w1(32'h3ba97cc8),
	.w2(32'hbba6cb49),
	.w3(32'h3ae46a83),
	.w4(32'hbb3c7c82),
	.w5(32'h3b2b2577),
	.w6(32'hbbb79f1f),
	.w7(32'hbba0396c),
	.w8(32'h3ab33a13),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a760662),
	.w1(32'hbb934d86),
	.w2(32'hbd0047f4),
	.w3(32'hba0fad86),
	.w4(32'h3bdb7aff),
	.w5(32'hbd1cb13b),
	.w6(32'h3af0dc12),
	.w7(32'h3a1583ae),
	.w8(32'hbcd20647),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcff059a),
	.w1(32'hbcbb1dc9),
	.w2(32'hbbc7949f),
	.w3(32'hbd40f78d),
	.w4(32'hbd086b05),
	.w5(32'hbb141cbe),
	.w6(32'hbcfe4f1c),
	.w7(32'hbcedba6f),
	.w8(32'hbbc3126b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5af8),
	.w1(32'hb91f618d),
	.w2(32'h3b9abf91),
	.w3(32'hbc37dcb3),
	.w4(32'hbb938f0d),
	.w5(32'h3c82f3ba),
	.w6(32'hbc369d6d),
	.w7(32'hbb0ae068),
	.w8(32'h3c98fbef),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cc2c8),
	.w1(32'h3b10939e),
	.w2(32'hbc81b403),
	.w3(32'h3d0809dd),
	.w4(32'h3cafb5f5),
	.w5(32'hbc1d8983),
	.w6(32'h3d26ee05),
	.w7(32'h3d11cab3),
	.w8(32'hbb0e856a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb862658),
	.w1(32'h3be4836b),
	.w2(32'hbbcc94f7),
	.w3(32'hb951e83f),
	.w4(32'h3be7c78e),
	.w5(32'h3a43f7c2),
	.w6(32'h3bc49d9e),
	.w7(32'h3bfb350c),
	.w8(32'h3c05ce1c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0301b8),
	.w1(32'hbb98e93e),
	.w2(32'h3cd77dca),
	.w3(32'hbc425414),
	.w4(32'hbbb6ce66),
	.w5(32'h3c68bf3d),
	.w6(32'h3c2bcafd),
	.w7(32'h3c174c6d),
	.w8(32'h3c7c8036),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0efcc4),
	.w1(32'hba2a7eaa),
	.w2(32'h3ac41335),
	.w3(32'hbb84f4ed),
	.w4(32'hbb9dc57f),
	.w5(32'h3b29f6a4),
	.w6(32'hbbec96a4),
	.w7(32'h3c1ec94f),
	.w8(32'h3bef32e8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa9a044),
	.w1(32'hba7bd046),
	.w2(32'h3b4101c2),
	.w3(32'hbbdfb98b),
	.w4(32'h3a919781),
	.w5(32'h3af20911),
	.w6(32'h3b55b2a5),
	.w7(32'h3b51a748),
	.w8(32'hbaf4c680),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c1227),
	.w1(32'hbaf75614),
	.w2(32'h3b0fe76d),
	.w3(32'h3b31168e),
	.w4(32'h39f918a7),
	.w5(32'h3beba84b),
	.w6(32'h3a715be6),
	.w7(32'h3ae6f509),
	.w8(32'h3ae8a8dc),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58cfef),
	.w1(32'h3b2299cb),
	.w2(32'hbabc3b71),
	.w3(32'h3c6cf4c6),
	.w4(32'h3c45dfd6),
	.w5(32'h3bbe0300),
	.w6(32'h3a80e6fb),
	.w7(32'h3aaaf8d5),
	.w8(32'h3c8cc885),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1086bb),
	.w1(32'h3b1a5de2),
	.w2(32'hbc5104a5),
	.w3(32'h3c22c0cf),
	.w4(32'h3c8b9039),
	.w5(32'hbbb84a9e),
	.w6(32'h3c1ce434),
	.w7(32'h3ca8393c),
	.w8(32'h3bda2cd4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccf0bbc),
	.w1(32'hbca0eeeb),
	.w2(32'hbbc40fca),
	.w3(32'hbbee9718),
	.w4(32'hbc50033d),
	.w5(32'hbbb042b3),
	.w6(32'h3bebf015),
	.w7(32'hbb9ab515),
	.w8(32'hbba1f56d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caf432),
	.w1(32'hbad005ea),
	.w2(32'hbc1700a2),
	.w3(32'h3baa53b6),
	.w4(32'h3b1339cf),
	.w5(32'h3b0b735d),
	.w6(32'h3b5578e4),
	.w7(32'h3c2c8440),
	.w8(32'h388e0f28),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb0948),
	.w1(32'hbc452cd2),
	.w2(32'hbc85e8ed),
	.w3(32'hb8362ae1),
	.w4(32'hbadd0817),
	.w5(32'hbc14dcfd),
	.w6(32'h3c2bfb74),
	.w7(32'h3ba41541),
	.w8(32'h39cae651),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93d68),
	.w1(32'h3af505f0),
	.w2(32'hbbcef0e4),
	.w3(32'h3b763487),
	.w4(32'h3b3791f3),
	.w5(32'hb8aed377),
	.w6(32'h3ba8b2bc),
	.w7(32'h3c70f830),
	.w8(32'h3a3be436),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b548c65),
	.w1(32'hbbaecc68),
	.w2(32'hbc8d8652),
	.w3(32'h3c3ffe38),
	.w4(32'h3b002e65),
	.w5(32'hbc3a9e38),
	.w6(32'h3c2735c0),
	.w7(32'h3c149b3a),
	.w8(32'hbc22a55a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ca10),
	.w1(32'hbc889e05),
	.w2(32'hbc0ccb8f),
	.w3(32'hbb27f77c),
	.w4(32'hbc32a468),
	.w5(32'h3b3e3210),
	.w6(32'hbbfc9f43),
	.w7(32'hbacb1392),
	.w8(32'hbb3095ed),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd605ef),
	.w1(32'h3a038411),
	.w2(32'hbb6b3bf0),
	.w3(32'h3c32a40f),
	.w4(32'h3b813d7f),
	.w5(32'hbbfb882a),
	.w6(32'hbb559edd),
	.w7(32'h398a53f9),
	.w8(32'hbcd9dcbc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1dd5ff),
	.w1(32'hbba6f741),
	.w2(32'h3b8bac5e),
	.w3(32'hbce48311),
	.w4(32'hbcd775bd),
	.w5(32'h3b5ea511),
	.w6(32'hbd12fa42),
	.w7(32'hbce90fa7),
	.w8(32'h3b569ff0),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f62a1),
	.w1(32'h3adb1c5c),
	.w2(32'hbd3cc9b7),
	.w3(32'h3c6045a9),
	.w4(32'h3af7836e),
	.w5(32'hbd22dae7),
	.w6(32'h3ca30796),
	.w7(32'h3b8f542e),
	.w8(32'hbce1a1ef),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87b67a),
	.w1(32'h3befe6b9),
	.w2(32'h3a0a2dfd),
	.w3(32'hbbbaa2fb),
	.w4(32'h3cb6b018),
	.w5(32'h3c8c593d),
	.w6(32'h3c28a93d),
	.w7(32'h3cf72263),
	.w8(32'h3cc8c713),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80a064),
	.w1(32'hbc78930e),
	.w2(32'hbb49286d),
	.w3(32'h3b76c9fa),
	.w4(32'hbb55f7ee),
	.w5(32'hbb51ca25),
	.w6(32'h3cb07643),
	.w7(32'h3cb3f52c),
	.w8(32'h3bb76a32),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c227e7e),
	.w1(32'h3b544c7d),
	.w2(32'hbc56c8d5),
	.w3(32'h3c09b4c3),
	.w4(32'h3b17fa1c),
	.w5(32'hbaea294c),
	.w6(32'h3c2630c6),
	.w7(32'h3c07d416),
	.w8(32'hbbc83d8a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1dd0e6),
	.w1(32'hbc2e1ed7),
	.w2(32'h3c0532b2),
	.w3(32'hbb0293bb),
	.w4(32'h3a42ef70),
	.w5(32'h3c33a782),
	.w6(32'hba65be0f),
	.w7(32'hbbcba769),
	.w8(32'h3c822001),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ba946),
	.w1(32'h39e1b9a3),
	.w2(32'hbbb51061),
	.w3(32'h3c46e7d7),
	.w4(32'h3c0ac3bb),
	.w5(32'h3a1e2357),
	.w6(32'h3bf3206b),
	.w7(32'h3c01f959),
	.w8(32'h3bb293b5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14fbc7),
	.w1(32'h3c563b25),
	.w2(32'hbadfd33f),
	.w3(32'h3b97ec08),
	.w4(32'h3c217c3b),
	.w5(32'h3c6deeb8),
	.w6(32'h3c2d78b5),
	.w7(32'h3c7d121e),
	.w8(32'h3c0f663e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca94574),
	.w1(32'h3c188042),
	.w2(32'hbc496de4),
	.w3(32'h3c6e539f),
	.w4(32'hbb8f0f03),
	.w5(32'hbc64bac6),
	.w6(32'hbb203383),
	.w7(32'hbc7c7ad9),
	.w8(32'hbc417170),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdafb27),
	.w1(32'hbadf0004),
	.w2(32'hbc745393),
	.w3(32'hbc160f95),
	.w4(32'hb973762d),
	.w5(32'hbcb68c74),
	.w6(32'hbbb0e471),
	.w7(32'h3ae3fddc),
	.w8(32'hbcd3666a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d641a),
	.w1(32'h3be6755e),
	.w2(32'hbd6e6303),
	.w3(32'h3a510fac),
	.w4(32'h3a640487),
	.w5(32'hbd63b90e),
	.w6(32'hbc99922f),
	.w7(32'hbc471ca0),
	.w8(32'hbd4e48fd),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bb951),
	.w1(32'h3c5fc542),
	.w2(32'hbc05e9fe),
	.w3(32'h3c4ae049),
	.w4(32'h3c61260a),
	.w5(32'hbc22c6e9),
	.w6(32'h3caf76ab),
	.w7(32'h3c9cfa91),
	.w8(32'hbcb68e79),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925a52),
	.w1(32'hbb402a5e),
	.w2(32'hbc52e7cf),
	.w3(32'h3b59a7c3),
	.w4(32'h3c24127c),
	.w5(32'hbc33eefe),
	.w6(32'hbaf1914f),
	.w7(32'h3c343e3f),
	.w8(32'hbc38077b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a2e5),
	.w1(32'h3a4916a5),
	.w2(32'h3c51d774),
	.w3(32'h3ca4170e),
	.w4(32'h3c795113),
	.w5(32'h3ca02628),
	.w6(32'h3c1bc8d2),
	.w7(32'h3c62f3d7),
	.w8(32'h3ce2e5d1),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d310f90),
	.w1(32'h3cff3c4d),
	.w2(32'hbc90087a),
	.w3(32'h3d25a430),
	.w4(32'h3d072231),
	.w5(32'hbbcd2e38),
	.w6(32'h3d23486a),
	.w7(32'h3d126a62),
	.w8(32'hbc5d03dd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88e5a3),
	.w1(32'h3c55ef84),
	.w2(32'h3aac9665),
	.w3(32'h3cf73631),
	.w4(32'h3ce3d1d4),
	.w5(32'h3c39d63d),
	.w6(32'h3c1bf177),
	.w7(32'h3c8b4295),
	.w8(32'hba7b1f37),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fc524),
	.w1(32'h3bb47687),
	.w2(32'hbccd4f40),
	.w3(32'h3c5bc26f),
	.w4(32'h3c432354),
	.w5(32'hbc953b36),
	.w6(32'h3c90f0c3),
	.w7(32'h3c138dce),
	.w8(32'hbc8965dc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b987efe),
	.w1(32'h390dae5a),
	.w2(32'hbcf10202),
	.w3(32'h3c558a5e),
	.w4(32'h3bdee940),
	.w5(32'hbcd843f3),
	.w6(32'h3c5b4a61),
	.w7(32'h3b63b0ea),
	.w8(32'hbcad4367),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbea006),
	.w1(32'hbc571ee6),
	.w2(32'hbd0e4694),
	.w3(32'h39e064ec),
	.w4(32'h3c725084),
	.w5(32'hbc9eb5cd),
	.w6(32'h3c1dd3bf),
	.w7(32'h3c5ff4ed),
	.w8(32'h3c8eb22c),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695e91),
	.w1(32'h3c777c5a),
	.w2(32'hbc59311d),
	.w3(32'h3caf9fb0),
	.w4(32'h3cc45220),
	.w5(32'hbb215d1f),
	.w6(32'h3cba2f10),
	.w7(32'h3c3c0c5a),
	.w8(32'hbb4b7b0c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c975b7c),
	.w1(32'hbb5f92ce),
	.w2(32'hbc39ecb8),
	.w3(32'h3c9ebe2a),
	.w4(32'h3c070ece),
	.w5(32'hbbfd9ef6),
	.w6(32'h3b4b3b9e),
	.w7(32'h3ae4429a),
	.w8(32'hbc65dc9a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c968937),
	.w1(32'h3c82d150),
	.w2(32'hbc99dae9),
	.w3(32'h3c67a7e0),
	.w4(32'h3c693279),
	.w5(32'hbc8b941f),
	.w6(32'h3bc55c56),
	.w7(32'h3c246672),
	.w8(32'hbc8a3659),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f0b4),
	.w1(32'hb986a7ab),
	.w2(32'hbc7756f5),
	.w3(32'hbb77a2e0),
	.w4(32'h3ba4a622),
	.w5(32'hbc00688a),
	.w6(32'hb93a40bd),
	.w7(32'h3baba564),
	.w8(32'hbb972df6),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3c9ac),
	.w1(32'hbb7d4643),
	.w2(32'h3c28d422),
	.w3(32'hbc6280da),
	.w4(32'hbb9b6e5d),
	.w5(32'h3c4eefcf),
	.w6(32'hbc622b3f),
	.w7(32'hbbbdd15a),
	.w8(32'h3b2ba407),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b701c),
	.w1(32'hbb0a9cba),
	.w2(32'hbc8dca98),
	.w3(32'h3b1d2325),
	.w4(32'h3c3603b5),
	.w5(32'hbc920776),
	.w6(32'h3c1050ae),
	.w7(32'h3c290cb0),
	.w8(32'hbc085119),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef7229),
	.w1(32'hba61114d),
	.w2(32'h3c1715d7),
	.w3(32'h3c34cb35),
	.w4(32'h3c3fad64),
	.w5(32'h3c626786),
	.w6(32'h3c9d1c26),
	.w7(32'h3be346b1),
	.w8(32'h3b9aac2f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0e6b2),
	.w1(32'hbc0a37d9),
	.w2(32'hbca6eac1),
	.w3(32'h3b910d9e),
	.w4(32'h3b7f914f),
	.w5(32'hbb82200f),
	.w6(32'h3bf142f1),
	.w7(32'h3b8f6900),
	.w8(32'h3b230c14),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c83c),
	.w1(32'h3a1fc626),
	.w2(32'h3bf5b4d4),
	.w3(32'h3c17acbe),
	.w4(32'h3b44145b),
	.w5(32'h3bf24ba3),
	.w6(32'h3bd5dbc6),
	.w7(32'h3ad1c87e),
	.w8(32'hbbcd0ce4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6825),
	.w1(32'h3a501745),
	.w2(32'h3c32ac7a),
	.w3(32'h3b310ae0),
	.w4(32'hbb672af6),
	.w5(32'h3c11ed53),
	.w6(32'hbc4570c0),
	.w7(32'hbba3d1db),
	.w8(32'h3bb4bab3),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e21c6),
	.w1(32'h3bab4861),
	.w2(32'h3be432bf),
	.w3(32'h3bd3537a),
	.w4(32'h3c209778),
	.w5(32'h3c141b14),
	.w6(32'hbb878b8a),
	.w7(32'h3b17602c),
	.w8(32'h3c313a13),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c826412),
	.w1(32'hbcacd087),
	.w2(32'hbd242c1b),
	.w3(32'h3cb2ae09),
	.w4(32'hbc1b8a49),
	.w5(32'hbce03f08),
	.w6(32'h3c2c7aa7),
	.w7(32'hbadddad4),
	.w8(32'hbcfecd7e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94715b),
	.w1(32'h3c82f9c0),
	.w2(32'hbaef6663),
	.w3(32'h3bfee239),
	.w4(32'h3c24a4fb),
	.w5(32'h3be4a6f1),
	.w6(32'hbbbf9f4b),
	.w7(32'h3c3e968c),
	.w8(32'hbbbf53f3),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c965d02),
	.w1(32'h3bb0b10c),
	.w2(32'hbbac3bf7),
	.w3(32'h3c9abe39),
	.w4(32'h3bf5e9c8),
	.w5(32'hbc0d062a),
	.w6(32'h3c8e5f8c),
	.w7(32'h3bcb316a),
	.w8(32'hbc8a98e2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0eed32),
	.w1(32'h3cac50ad),
	.w2(32'hbd54b1ac),
	.w3(32'h3cc73e67),
	.w4(32'h3cb9cea6),
	.w5(32'hbd2147e2),
	.w6(32'h3ba230bb),
	.w7(32'h3c5ff306),
	.w8(32'hbcf98661),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc020ebe),
	.w1(32'hbb63cf90),
	.w2(32'hbcc4e16c),
	.w3(32'h3ca2c9e2),
	.w4(32'h3c89ba41),
	.w5(32'hb940a98a),
	.w6(32'h3cb2638c),
	.w7(32'h3cdecbbe),
	.w8(32'h3c075121),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b4c66),
	.w1(32'h3b83c67f),
	.w2(32'hbcc96a9a),
	.w3(32'h3c3d0388),
	.w4(32'h3ac85e53),
	.w5(32'hbd038240),
	.w6(32'h3ac83a9a),
	.w7(32'hbbe62fe4),
	.w8(32'hbcfb00d4),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95b1c2),
	.w1(32'hbca70828),
	.w2(32'h3b619b4d),
	.w3(32'hbd14d8e7),
	.w4(32'hbcc1cd02),
	.w5(32'h3bfdaab7),
	.w6(32'hbcbec9f4),
	.w7(32'hbc5a3fff),
	.w8(32'h3b0e342f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f13261),
	.w1(32'hbb384632),
	.w2(32'h3c328ab8),
	.w3(32'h3c145ee1),
	.w4(32'h3bb8f8b0),
	.w5(32'h3b66cc6f),
	.w6(32'h39c33c2e),
	.w7(32'hbb1b555d),
	.w8(32'h3c2ad923),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f078),
	.w1(32'h3c1ccf70),
	.w2(32'hba9eb9fe),
	.w3(32'h3cbf81b7),
	.w4(32'h3c915583),
	.w5(32'h39c7c03a),
	.w6(32'h3cb51d5d),
	.w7(32'h3c5a4799),
	.w8(32'h3b9fbf56),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c808e21),
	.w1(32'h3c2c551c),
	.w2(32'hbcf9ccb4),
	.w3(32'h3c3f567e),
	.w4(32'h3a2a5d14),
	.w5(32'hbcb86319),
	.w6(32'h3b764cc8),
	.w7(32'hbb74834c),
	.w8(32'hbcaf6ded),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11b454),
	.w1(32'h3b11a1b1),
	.w2(32'hbc08215b),
	.w3(32'h3c6e39c9),
	.w4(32'h3c101a47),
	.w5(32'hbb0f6d91),
	.w6(32'h3c87f1ab),
	.w7(32'h3bb2946e),
	.w8(32'h3a8c1984),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7332d),
	.w1(32'h3a9415b0),
	.w2(32'hbca8a01a),
	.w3(32'h3b07ed9b),
	.w4(32'hb8b34aa4),
	.w5(32'hbcd77159),
	.w6(32'h3bed1225),
	.w7(32'h3b5297fc),
	.w8(32'hbcd4b75e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb1b1bb),
	.w1(32'hbcb513fd),
	.w2(32'h3bb8f10c),
	.w3(32'hbd057089),
	.w4(32'hbce591f5),
	.w5(32'h3c3a9655),
	.w6(32'hbcc874c2),
	.w7(32'hbc8e82db),
	.w8(32'h3c5a54bb),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd62a4c),
	.w1(32'hba04e2de),
	.w2(32'hbd52ee11),
	.w3(32'h3d098e9d),
	.w4(32'h3c655b66),
	.w5(32'hbd37cdee),
	.w6(32'h3d0b792b),
	.w7(32'h3c980181),
	.w8(32'hbd192109),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b8258),
	.w1(32'h3c76a105),
	.w2(32'hbb8322b4),
	.w3(32'h3c3bcfb0),
	.w4(32'h3ce8ac0b),
	.w5(32'h3beebfe7),
	.w6(32'h3bc2767f),
	.w7(32'h3cc03eb8),
	.w8(32'h3a9f77dd),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf06587),
	.w1(32'h3bae5049),
	.w2(32'hbca1fcf5),
	.w3(32'h3b7b33bd),
	.w4(32'h3b72636c),
	.w5(32'hbc86298a),
	.w6(32'hba9b0484),
	.w7(32'h3ab82933),
	.w8(32'hbc27002c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de2ab),
	.w1(32'hbc2e0941),
	.w2(32'hbcb2a7ae),
	.w3(32'hbbd40000),
	.w4(32'hbc5608cd),
	.w5(32'hbcb1eab9),
	.w6(32'hbba0d436),
	.w7(32'hbbe42814),
	.w8(32'hbc852d15),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1de453),
	.w1(32'hbc094ce8),
	.w2(32'h3c0b2a05),
	.w3(32'hbc0bd7ed),
	.w4(32'hbc93def8),
	.w5(32'h3b3a83ec),
	.w6(32'hbbe39ee6),
	.w7(32'hbc43c21d),
	.w8(32'h3b4f91ec),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a43d6),
	.w1(32'h3b94d588),
	.w2(32'hbd1f8999),
	.w3(32'h3ce2f55c),
	.w4(32'h3b215322),
	.w5(32'hbce2e4d2),
	.w6(32'h3ce3b08a),
	.w7(32'h3b992429),
	.w8(32'hbd01dda6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce54966),
	.w1(32'hbc3e983c),
	.w2(32'hba985170),
	.w3(32'hbcbd594c),
	.w4(32'hbbb785dc),
	.w5(32'h3c038459),
	.w6(32'hbc439423),
	.w7(32'hbbbcb6f6),
	.w8(32'h3c3486f4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c4e32),
	.w1(32'h3bfc2c7d),
	.w2(32'h3b477b9c),
	.w3(32'h3be04996),
	.w4(32'h3c072081),
	.w5(32'h3abf6226),
	.w6(32'h3c22bc2b),
	.w7(32'h3ca33d8c),
	.w8(32'hbaafc2ce),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0780b),
	.w1(32'hbb0af2e0),
	.w2(32'hbb420340),
	.w3(32'h3bce9f56),
	.w4(32'h3c0d8676),
	.w5(32'h3b149ede),
	.w6(32'h3b962508),
	.w7(32'h3bb0b8aa),
	.w8(32'hbc2e7998),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83bb5e),
	.w1(32'hbbb45da2),
	.w2(32'h39066134),
	.w3(32'h3cecdb05),
	.w4(32'hb8c0ab02),
	.w5(32'h39741d70),
	.w6(32'h3cd29009),
	.w7(32'h3c3629b5),
	.w8(32'h3bfbc48c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbb7d3),
	.w1(32'hbb9ebbbb),
	.w2(32'hbc3e5604),
	.w3(32'h3c987094),
	.w4(32'hbb9bfd3e),
	.w5(32'hbc2f0507),
	.w6(32'h3cbe549b),
	.w7(32'hbaff28dc),
	.w8(32'hbc34e2a1),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388deded),
	.w1(32'hbca8b231),
	.w2(32'hbc876676),
	.w3(32'h3c4a0888),
	.w4(32'hbc58de03),
	.w5(32'hbbaa38fc),
	.w6(32'h3c4503ca),
	.w7(32'hbc8cc97c),
	.w8(32'hbb65edc4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d13a0eb),
	.w1(32'h3b208820),
	.w2(32'hbb275280),
	.w3(32'h3d19ace4),
	.w4(32'h3ad9d449),
	.w5(32'hbc2d07c8),
	.w6(32'h3d188859),
	.w7(32'h3b1530ac),
	.w8(32'hbc8a8aa5),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfdde8a),
	.w1(32'h3a989c3b),
	.w2(32'h3ad8db91),
	.w3(32'hbc4b175d),
	.w4(32'h3a6d2d93),
	.w5(32'hbbaa4cf4),
	.w6(32'hbc9ead2c),
	.w7(32'hbc134a9a),
	.w8(32'hbc455de4),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbe68a1),
	.w1(32'h3caaa71c),
	.w2(32'hbc220fc6),
	.w3(32'h3c9bd71b),
	.w4(32'h3c8f8bb3),
	.w5(32'hbaeef5a5),
	.w6(32'h3b3a797c),
	.w7(32'hbbea54a9),
	.w8(32'hbc457562),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94d1d9),
	.w1(32'h3c301b34),
	.w2(32'hbc11d640),
	.w3(32'h3c66c6a0),
	.w4(32'h3c9f71a0),
	.w5(32'hbc40aea2),
	.w6(32'h3c8f2cc8),
	.w7(32'h3c852d0b),
	.w8(32'hbc1766f1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7216cd),
	.w1(32'h3bb568f4),
	.w2(32'hbc27f14e),
	.w3(32'h3b975031),
	.w4(32'h3c1a6f3e),
	.w5(32'hbb59e58f),
	.w6(32'h3c64d26b),
	.w7(32'hb9b3d426),
	.w8(32'hbb3acd42),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2dbe5),
	.w1(32'hbc695ce0),
	.w2(32'hbb4873f6),
	.w3(32'h3cc364ba),
	.w4(32'hbba3bf63),
	.w5(32'hbb3fb8b3),
	.w6(32'h3cd259d4),
	.w7(32'hbc060c41),
	.w8(32'h3bf51699),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf08222),
	.w1(32'h3c2b1c58),
	.w2(32'h3c83bae9),
	.w3(32'h3b5da2ee),
	.w4(32'h3bf76fc9),
	.w5(32'h3c8300ed),
	.w6(32'h3b29ee70),
	.w7(32'h3c21c17c),
	.w8(32'h3c8bbca1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55ec06),
	.w1(32'h3b98661e),
	.w2(32'hbc92ee3d),
	.w3(32'h3c2ad9bf),
	.w4(32'h3c25981b),
	.w5(32'hbc215473),
	.w6(32'h3c816f2d),
	.w7(32'h3c2c6b15),
	.w8(32'hbc6a1585),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d012579),
	.w1(32'h3d1ff257),
	.w2(32'hbd08b173),
	.w3(32'h3caa8065),
	.w4(32'h3c910f4f),
	.w5(32'hbd02b7d9),
	.w6(32'hbbf7838c),
	.w7(32'h3c884675),
	.w8(32'hbd328af2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbbe363),
	.w1(32'h3c5cdc1e),
	.w2(32'hbd824391),
	.w3(32'h3cea814e),
	.w4(32'h3ca08a31),
	.w5(32'hbd5378a4),
	.w6(32'h392593aa),
	.w7(32'hbb5b4aad),
	.w8(32'hbd5ebf0f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfd090),
	.w1(32'hbc859358),
	.w2(32'hbcd81a4f),
	.w3(32'h3c997837),
	.w4(32'hbb7cd992),
	.w5(32'hbcb6521c),
	.w6(32'hbc0f3e9b),
	.w7(32'hbb95438c),
	.w8(32'hbc6a0508),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8420c5),
	.w1(32'hbacbe424),
	.w2(32'hbc502771),
	.w3(32'hbc41abbd),
	.w4(32'h3b18c71c),
	.w5(32'hbc0ef5c9),
	.w6(32'hba87c1c6),
	.w7(32'h3c3f3146),
	.w8(32'hbb2d216d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffa8f4),
	.w1(32'hbb028869),
	.w2(32'hbc8cabc1),
	.w3(32'hb8e40775),
	.w4(32'h3919b483),
	.w5(32'hbcc1698b),
	.w6(32'h3bfcef64),
	.w7(32'h3c400c17),
	.w8(32'hbc856aec),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81d747),
	.w1(32'hbcb516f8),
	.w2(32'hbbf416c2),
	.w3(32'hbd0e1e87),
	.w4(32'hbcef6b44),
	.w5(32'hbc6e79f3),
	.w6(32'hbcc2df9f),
	.w7(32'hbc5f95c4),
	.w8(32'hbae92b29),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd26aaa),
	.w1(32'h3b851716),
	.w2(32'hb8862a19),
	.w3(32'hbc33b63e),
	.w4(32'hbba5713b),
	.w5(32'h3c2ce46d),
	.w6(32'hbc418a5d),
	.w7(32'hbb7036ba),
	.w8(32'h3b64b760),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c557016),
	.w1(32'h3bd10584),
	.w2(32'h3c367445),
	.w3(32'h3c302ca4),
	.w4(32'h3c3207fe),
	.w5(32'h3c9c15ec),
	.w6(32'h3c01babc),
	.w7(32'h3b871f2c),
	.w8(32'h3c06f951),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf47c4f),
	.w1(32'h3c634c5c),
	.w2(32'h3b2215d5),
	.w3(32'h3d0023bc),
	.w4(32'h3caa66d4),
	.w5(32'h3b99b413),
	.w6(32'h3cbfd012),
	.w7(32'h3b5dbb19),
	.w8(32'hbc1f490f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0e01d),
	.w1(32'hbae1c6a2),
	.w2(32'hbcd05068),
	.w3(32'h3c55faea),
	.w4(32'hbb96e709),
	.w5(32'hbcb51ed2),
	.w6(32'h3c0eb39f),
	.w7(32'hb97a053d),
	.w8(32'hbcb24259),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a22db),
	.w1(32'h3ad2fd9b),
	.w2(32'hbc65618c),
	.w3(32'h3ba4f764),
	.w4(32'h3a19ba89),
	.w5(32'hbcb0a785),
	.w6(32'h3bb12d80),
	.w7(32'h3be84e99),
	.w8(32'hbcb6e1ff),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0079f),
	.w1(32'hbbb99265),
	.w2(32'hbbf89e42),
	.w3(32'hbba296b0),
	.w4(32'hbc255b37),
	.w5(32'hbcaf5e0b),
	.w6(32'hbbb97dc9),
	.w7(32'h399623ed),
	.w8(32'hbc71f87f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1070ee),
	.w1(32'hbaae11da),
	.w2(32'hb9c16e78),
	.w3(32'hbc3540de),
	.w4(32'hbc01bf36),
	.w5(32'h3b0b2077),
	.w6(32'hbc18164e),
	.w7(32'hbb964a7f),
	.w8(32'h3b202da4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb59961),
	.w1(32'h3b95a5e5),
	.w2(32'hbc0a590d),
	.w3(32'h3cc48b1f),
	.w4(32'h3b12b779),
	.w5(32'hbc0bae8d),
	.w6(32'h3c4a852e),
	.w7(32'h3c3fd5e5),
	.w8(32'hbc5af652),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01c9d5),
	.w1(32'h3aab9e77),
	.w2(32'hbc1b2847),
	.w3(32'h3c0e6e82),
	.w4(32'h3b22afa4),
	.w5(32'hbc1c30a7),
	.w6(32'hbbb66a27),
	.w7(32'hbb08c2fa),
	.w8(32'hbc3e42a8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad73bdb),
	.w1(32'h3b14550e),
	.w2(32'h3c245ac3),
	.w3(32'h3b643ea0),
	.w4(32'h3b414f01),
	.w5(32'h3b6b2b1e),
	.w6(32'h3b4787a8),
	.w7(32'h3b922524),
	.w8(32'h3ba0f351),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7fcb),
	.w1(32'h3bbb9cb8),
	.w2(32'h3b0b2539),
	.w3(32'hbaeed99c),
	.w4(32'h3b11e2ae),
	.w5(32'h3a9f76d3),
	.w6(32'hbc2dcd10),
	.w7(32'h3bef778a),
	.w8(32'h3b40f009),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab6091),
	.w1(32'h3bed0400),
	.w2(32'h3c0d465a),
	.w3(32'h3b308239),
	.w4(32'h3b551267),
	.w5(32'h3c787aa7),
	.w6(32'h3b091721),
	.w7(32'h3b890597),
	.w8(32'h3c8237bc),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66bdd1),
	.w1(32'h3a87409b),
	.w2(32'h3ae86632),
	.w3(32'hbbadff2a),
	.w4(32'hbb1f19ec),
	.w5(32'h3c150fcd),
	.w6(32'h3aa7e6a0),
	.w7(32'hba49518d),
	.w8(32'h3c09b5b6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6de93f),
	.w1(32'hbb6931aa),
	.w2(32'hbbd38108),
	.w3(32'h3be8d125),
	.w4(32'h3bfaf43e),
	.w5(32'hbb41962a),
	.w6(32'h386aa4c8),
	.w7(32'hbadf342e),
	.w8(32'hbb33b372),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5fd92),
	.w1(32'h3b4b2507),
	.w2(32'h3bb817ca),
	.w3(32'h3b9aab29),
	.w4(32'hbb48b1fc),
	.w5(32'h3c3e7b22),
	.w6(32'hb846c0b5),
	.w7(32'hbb942374),
	.w8(32'h3b72c49b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85894d),
	.w1(32'h3c73a348),
	.w2(32'hbc399f6b),
	.w3(32'h3cae6f3a),
	.w4(32'h3cb0e8c6),
	.w5(32'hbc2306a4),
	.w6(32'h3c9979c5),
	.w7(32'h3c6f764d),
	.w8(32'hba9aca14),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbae95),
	.w1(32'hbcbe6afc),
	.w2(32'hbcac23d5),
	.w3(32'h3c542735),
	.w4(32'hbc5bc39f),
	.w5(32'h3b4ac15a),
	.w6(32'h3befa4b6),
	.w7(32'hbbf00bf3),
	.w8(32'hbaaf502c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d063017),
	.w1(32'h3c91a82e),
	.w2(32'hbbebc371),
	.w3(32'h3d2c887f),
	.w4(32'h3c8eb983),
	.w5(32'h3b396957),
	.w6(32'h3cd1e900),
	.w7(32'h3c333010),
	.w8(32'h3c0c155f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c91c1),
	.w1(32'hbc2f429c),
	.w2(32'hbca2acb4),
	.w3(32'h3ca41fc8),
	.w4(32'h3c0f7cd6),
	.w5(32'hbc2d9e67),
	.w6(32'h3c832be8),
	.w7(32'h3b9ef63e),
	.w8(32'hbb86a5dc),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c44e1b3),
	.w1(32'h3c2c1ba8),
	.w2(32'hbc117244),
	.w3(32'h3bce464f),
	.w4(32'h3c435f4e),
	.w5(32'hbbbee369),
	.w6(32'hbc2a978d),
	.w7(32'hbb8c92a4),
	.w8(32'hba7369f2),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3affaa),
	.w1(32'h3b20fa96),
	.w2(32'hbd498574),
	.w3(32'hbaa40e6f),
	.w4(32'hb91174fa),
	.w5(32'hbcfa260c),
	.w6(32'h3bbaf261),
	.w7(32'h3bf3ad91),
	.w8(32'hbc8dad75),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7ea7e3),
	.w1(32'hba501809),
	.w2(32'h3ae6bbaf),
	.w3(32'h3bc7e9b8),
	.w4(32'h3c5e79f8),
	.w5(32'h3c06000a),
	.w6(32'h3c87f590),
	.w7(32'h3ca5eca8),
	.w8(32'hba82bd81),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdaae0a),
	.w1(32'h3b6fa1a6),
	.w2(32'hbb4d8ab1),
	.w3(32'h3c51c755),
	.w4(32'h3bba1eb8),
	.w5(32'h3b7adf96),
	.w6(32'h3ba949ae),
	.w7(32'h39428d50),
	.w8(32'hbbc072b2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabba94f),
	.w1(32'hbbb1dbd0),
	.w2(32'hbd02abff),
	.w3(32'hbae6197e),
	.w4(32'hb94bbfea),
	.w5(32'hbcf60d6a),
	.w6(32'hbbab931e),
	.w7(32'hbbba11ee),
	.w8(32'hbcb593ca),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b96c),
	.w1(32'hbbacca96),
	.w2(32'hbc3ea729),
	.w3(32'hbcab51ff),
	.w4(32'hbc24f3ed),
	.w5(32'hbc899db4),
	.w6(32'hbbec2399),
	.w7(32'hbbccf75f),
	.w8(32'hbc2ccfef),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc407ee1),
	.w1(32'hbaa4e6b5),
	.w2(32'h3be0cece),
	.w3(32'hbca7fd85),
	.w4(32'hbc1c8413),
	.w5(32'h3b9f0cdd),
	.w6(32'hbc3e16f3),
	.w7(32'hbc319cae),
	.w8(32'h3bebb248),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa51d57),
	.w1(32'h3b8bb624),
	.w2(32'hbc4c7046),
	.w3(32'hbb63870f),
	.w4(32'h3aa9d065),
	.w5(32'hbc374a54),
	.w6(32'hba81b271),
	.w7(32'h3b5fc6b3),
	.w8(32'hbc2af8cc),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0c786),
	.w1(32'hbbd9a337),
	.w2(32'h3ac3437d),
	.w3(32'hbc0dd795),
	.w4(32'hbbe71350),
	.w5(32'hbaae984d),
	.w6(32'hbbab894b),
	.w7(32'hbb9abd53),
	.w8(32'hbc1049d1),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24f6d5),
	.w1(32'h3bded5da),
	.w2(32'h3ad50b71),
	.w3(32'h3ce3595d),
	.w4(32'h3b7deaf6),
	.w5(32'h3b3c1f8f),
	.w6(32'h3bc92dce),
	.w7(32'h3b6aa110),
	.w8(32'h3a4e8b3a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaa269),
	.w1(32'hbb448acc),
	.w2(32'h3a6da52e),
	.w3(32'h3c1b3cc1),
	.w4(32'hbb26e7ec),
	.w5(32'hbba7e2e7),
	.w6(32'h3bff79b5),
	.w7(32'hbb22866e),
	.w8(32'hbbb5e5e9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c405a8f),
	.w1(32'hbc50a613),
	.w2(32'hbd1b5522),
	.w3(32'h3caabde8),
	.w4(32'h3bbb63d8),
	.w5(32'hbcf16bb3),
	.w6(32'h3b64a9ef),
	.w7(32'hbbfc94b8),
	.w8(32'hbca46c03),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb79c43),
	.w1(32'h3b5290bd),
	.w2(32'hbc949965),
	.w3(32'h3c0bbb57),
	.w4(32'hba340b47),
	.w5(32'hbc5e4c46),
	.w6(32'h3b5a9345),
	.w7(32'h3aec5fc9),
	.w8(32'hbc669bc7),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76ac14),
	.w1(32'h3c33793f),
	.w2(32'hb87e8af2),
	.w3(32'h3b936899),
	.w4(32'h3c006fdd),
	.w5(32'h3bc44e7e),
	.w6(32'hbc6a0645),
	.w7(32'hb99d98c5),
	.w8(32'hbba2e987),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule