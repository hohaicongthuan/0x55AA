module layer_8_featuremap_54(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ba4eb),
	.w1(32'h3b9cc47d),
	.w2(32'h3b06171d),
	.w3(32'h3b8aec51),
	.w4(32'h3b8626a5),
	.w5(32'hb94227fb),
	.w6(32'h3b8cff37),
	.w7(32'hba859f22),
	.w8(32'hbb72fa93),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba445880),
	.w1(32'hba24a1d4),
	.w2(32'hba8c100b),
	.w3(32'hba6c1841),
	.w4(32'hba2f71ff),
	.w5(32'hbaa22a6e),
	.w6(32'hb89925e2),
	.w7(32'hb8f555ba),
	.w8(32'hb982a2c5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a389523),
	.w1(32'h3a818de8),
	.w2(32'h39e2c880),
	.w3(32'h39dd106a),
	.w4(32'h3a9c1254),
	.w5(32'h3a2193c7),
	.w6(32'h3a82245b),
	.w7(32'h39f5b837),
	.w8(32'hbafef9c2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa909a5),
	.w1(32'hb7b22bde),
	.w2(32'hba5cac4c),
	.w3(32'hb96569ec),
	.w4(32'hba11cc3b),
	.w5(32'hbae1ccb4),
	.w6(32'hbbb6e9f0),
	.w7(32'hbb937515),
	.w8(32'hbb00c984),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4d19f),
	.w1(32'h3b2d3dc2),
	.w2(32'h3ae45998),
	.w3(32'hbad9d536),
	.w4(32'h3b0758c8),
	.w5(32'h3aa4da9c),
	.w6(32'hb8c42d44),
	.w7(32'h3a805634),
	.w8(32'h3b1acbd7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa413dd),
	.w1(32'h3b285f0a),
	.w2(32'h3b995e0a),
	.w3(32'h3b6a0f7f),
	.w4(32'h3b50a395),
	.w5(32'h3bf4ff19),
	.w6(32'h3b4a364e),
	.w7(32'h3ba90b3d),
	.w8(32'h39e5dab0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7c0200),
	.w1(32'h3b33fea9),
	.w2(32'h3adf5c1b),
	.w3(32'h3999434e),
	.w4(32'h3acc85cf),
	.w5(32'h3a6d5c29),
	.w6(32'h3a0a34c1),
	.w7(32'hb8c9a838),
	.w8(32'hbb0d4b8d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba990e66),
	.w1(32'h3a814858),
	.w2(32'hba944a53),
	.w3(32'hb827a56c),
	.w4(32'h3a86c310),
	.w5(32'hbb35a746),
	.w6(32'h3a453964),
	.w7(32'hba68b5ca),
	.w8(32'hbb28c32e),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22c038),
	.w1(32'h3aff7c7d),
	.w2(32'h3a359654),
	.w3(32'hba4b9c85),
	.w4(32'h3b13276c),
	.w5(32'h3a371d54),
	.w6(32'h39fe3eec),
	.w7(32'h39d8820b),
	.w8(32'hb906a90b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b09d),
	.w1(32'h396381ab),
	.w2(32'hbb1423a6),
	.w3(32'h3b400bc6),
	.w4(32'hb9b1e5df),
	.w5(32'hbb7e92bc),
	.w6(32'hba9b116e),
	.w7(32'hbb8b622b),
	.w8(32'hbb706df4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba945d88),
	.w1(32'h392a8da8),
	.w2(32'h398851cc),
	.w3(32'hb9d435cb),
	.w4(32'h3a6ee002),
	.w5(32'hb99ee49b),
	.w6(32'hb9adba00),
	.w7(32'hbb6401cd),
	.w8(32'hbb89a8f3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2932),
	.w1(32'h3af8887f),
	.w2(32'hb981f441),
	.w3(32'h3ad70b0b),
	.w4(32'h3b0945d2),
	.w5(32'hbacd8610),
	.w6(32'h3af788a3),
	.w7(32'hbad61870),
	.w8(32'hbb4ba1d2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9014c7e),
	.w1(32'h3ad1a85c),
	.w2(32'h39156bb9),
	.w3(32'hba69f58a),
	.w4(32'h3a49a9b1),
	.w5(32'hb9e6b35f),
	.w6(32'hb966806d),
	.w7(32'hba19b067),
	.w8(32'h3b078e6e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b020060),
	.w1(32'h3b8f2365),
	.w2(32'h3bca610d),
	.w3(32'h3b812dbd),
	.w4(32'h3ba2e150),
	.w5(32'h3be1d485),
	.w6(32'h3b553da3),
	.w7(32'h3bb59f95),
	.w8(32'h3a541c1f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a925540),
	.w1(32'h3b4a9b70),
	.w2(32'h3b46fffa),
	.w3(32'h3ad80b1a),
	.w4(32'h3b356057),
	.w5(32'h3b26f5de),
	.w6(32'h3b072295),
	.w7(32'h3b127385),
	.w8(32'hb998fbec),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a1e18),
	.w1(32'h3ac0b396),
	.w2(32'hb995ee73),
	.w3(32'hb9716455),
	.w4(32'h3a3d730a),
	.w5(32'hba71fccd),
	.w6(32'h3a17d858),
	.w7(32'hba1c4268),
	.w8(32'hbae31878),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab8772b),
	.w1(32'hbb5cb933),
	.w2(32'hbb630f19),
	.w3(32'hba21d064),
	.w4(32'hba063158),
	.w5(32'h3af77eef),
	.w6(32'hbb4fc37e),
	.w7(32'hbb8070cd),
	.w8(32'hbb87c12d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab48514),
	.w1(32'h3ac77a13),
	.w2(32'hba875d84),
	.w3(32'h3a4c31d4),
	.w4(32'h3ad16e22),
	.w5(32'hba75061f),
	.w6(32'h3afeea28),
	.w7(32'hb965a88d),
	.w8(32'hbb2cf893),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e7e47),
	.w1(32'hba9b20c9),
	.w2(32'hbb26408b),
	.w3(32'h3bea6e66),
	.w4(32'h3b34bfb4),
	.w5(32'hbbece3ab),
	.w6(32'h3b7afca5),
	.w7(32'hbc2c9b1b),
	.w8(32'hbc5de84b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac975f7),
	.w1(32'h38b58859),
	.w2(32'hbb2123a1),
	.w3(32'h3b246ecf),
	.w4(32'hbacaf8d2),
	.w5(32'hbb22c239),
	.w6(32'h3ad684c3),
	.w7(32'hb947cc93),
	.w8(32'hbb463d82),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3101),
	.w1(32'hbb9649bd),
	.w2(32'hbb3582d3),
	.w3(32'hbbad72ec),
	.w4(32'hbb546f6f),
	.w5(32'hbafc7c75),
	.w6(32'hb801a1fe),
	.w7(32'hbb7192ee),
	.w8(32'hbb832397),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c55f6b),
	.w1(32'h3ae5dfe5),
	.w2(32'h3a57e1b4),
	.w3(32'hba81bdb2),
	.w4(32'h3abec3da),
	.w5(32'h3a449db1),
	.w6(32'h3a824ade),
	.w7(32'h3a7d6166),
	.w8(32'h3b151dea),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8850b0),
	.w1(32'hbb6037e6),
	.w2(32'hbb33c6b6),
	.w3(32'h3c17cfb9),
	.w4(32'h3a91f062),
	.w5(32'hbaec4a30),
	.w6(32'h3bc43f34),
	.w7(32'hbac48780),
	.w8(32'hbb56f40a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c7eda),
	.w1(32'h3b940021),
	.w2(32'h3a9feeff),
	.w3(32'h398f51dc),
	.w4(32'h3b131a4e),
	.w5(32'h3a536b2f),
	.w6(32'h3af87ee6),
	.w7(32'h3a976151),
	.w8(32'h39faab1c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba126888),
	.w1(32'h3a3ec569),
	.w2(32'hb8f18520),
	.w3(32'hbabb0580),
	.w4(32'h3a205993),
	.w5(32'hb822fa66),
	.w6(32'hba1c3d22),
	.w7(32'hba30a384),
	.w8(32'h3a4be3fb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82cb31),
	.w1(32'hbb8839f4),
	.w2(32'hbb5fb9ee),
	.w3(32'h3b27f6ee),
	.w4(32'hbb2a84b8),
	.w5(32'hbb0e55d4),
	.w6(32'hba534b4a),
	.w7(32'hbb207563),
	.w8(32'hbaaf2dc4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07327d),
	.w1(32'hbb664a19),
	.w2(32'hbafdad60),
	.w3(32'h396dc389),
	.w4(32'hbb1bce99),
	.w5(32'h389a743d),
	.w6(32'hbb03db8d),
	.w7(32'hb98c332e),
	.w8(32'hbb3fcdab),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2176eb),
	.w1(32'hbcc38029),
	.w2(32'hbcbfc147),
	.w3(32'h3bc949d8),
	.w4(32'h3a33ccb2),
	.w5(32'hbc8d7f4d),
	.w6(32'h3c2acf73),
	.w7(32'hbc812df7),
	.w8(32'hbd43dc02),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba827598),
	.w1(32'h3b7c39fa),
	.w2(32'hbb089fd1),
	.w3(32'hb9f4ea9e),
	.w4(32'h3b231977),
	.w5(32'hbb12dc48),
	.w6(32'h3aaa2ae0),
	.w7(32'hbb1461a2),
	.w8(32'hbb3c9051),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be35eb),
	.w1(32'h39309c2e),
	.w2(32'h3875302a),
	.w3(32'hba1ebdb9),
	.w4(32'hb91f3ea2),
	.w5(32'hb9b7ba80),
	.w6(32'hb9abd084),
	.w7(32'hba103c1d),
	.w8(32'hbb114ba0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b33a7),
	.w1(32'h3b602408),
	.w2(32'h3a85b427),
	.w3(32'hb8283cbb),
	.w4(32'h391ee99b),
	.w5(32'hba545491),
	.w6(32'hb69974aa),
	.w7(32'hbb2ca136),
	.w8(32'hbb7b0890),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d1ba5),
	.w1(32'hbb37f2f9),
	.w2(32'hbb793adc),
	.w3(32'hbb9a2ca4),
	.w4(32'hbb7236cf),
	.w5(32'hbb81a6b8),
	.w6(32'hbb1d6a02),
	.w7(32'hbbb6ce72),
	.w8(32'hbb1f9d0e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa93a18),
	.w1(32'h3b81c7b7),
	.w2(32'h3b11ff0a),
	.w3(32'hba289a7f),
	.w4(32'hb9c2740f),
	.w5(32'hbad46165),
	.w6(32'hba39a8e2),
	.w7(32'hbb16bbac),
	.w8(32'hba33e36a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96204f),
	.w1(32'h3a01460e),
	.w2(32'hb93dec2b),
	.w3(32'h39d935da),
	.w4(32'hba9dece3),
	.w5(32'hbb05d013),
	.w6(32'hba324f5e),
	.w7(32'h3a0d6501),
	.w8(32'h3ad596fa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae22ebf),
	.w1(32'h3b85dd77),
	.w2(32'h3bc4417e),
	.w3(32'h3b5ed747),
	.w4(32'h3bafc452),
	.w5(32'h3c06c169),
	.w6(32'h3b26c124),
	.w7(32'h3be0b96e),
	.w8(32'h3a466243),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3925f741),
	.w1(32'h3aaa538f),
	.w2(32'hbaf95438),
	.w3(32'h3838e910),
	.w4(32'h398dc4a4),
	.w5(32'hbb8d6d52),
	.w6(32'h3b28f901),
	.w7(32'hbb65e720),
	.w8(32'hbbb8c316),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ff067),
	.w1(32'hba149d18),
	.w2(32'hbaade48c),
	.w3(32'hbaf9e6f5),
	.w4(32'hba9db887),
	.w5(32'hbb0628f5),
	.w6(32'hbaa8f89b),
	.w7(32'hbaee8a4d),
	.w8(32'hba1f08f4),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a718908),
	.w1(32'h3b0d46ec),
	.w2(32'h3ac02651),
	.w3(32'h3a3c579b),
	.w4(32'h3afa3bec),
	.w5(32'h3a9a9950),
	.w6(32'h3a77ec7c),
	.w7(32'h3a2c964f),
	.w8(32'h3aa7933d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae11594),
	.w1(32'h3bbcd2bd),
	.w2(32'h3ba659e6),
	.w3(32'h3b2573a6),
	.w4(32'h3b9b53a6),
	.w5(32'h3b6e4d1e),
	.w6(32'h3b71c5f2),
	.w7(32'h3b5bf485),
	.w8(32'hbb0859b0),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa772c1),
	.w1(32'hba5e11b7),
	.w2(32'hbaf5f813),
	.w3(32'hbb0afd73),
	.w4(32'hbaf1c6d5),
	.w5(32'hbb3578f3),
	.w6(32'hbab49dcb),
	.w7(32'hbb1f3850),
	.w8(32'h3996b806),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b169402),
	.w1(32'hbaaafa78),
	.w2(32'hbb5ed92e),
	.w3(32'h3b82fd56),
	.w4(32'hbaabe88f),
	.w5(32'hbabca284),
	.w6(32'h389ed908),
	.w7(32'hbbcf3dc9),
	.w8(32'hbb4ffe60),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ceefb),
	.w1(32'hbb00296b),
	.w2(32'h38223a1e),
	.w3(32'hbb0bc1c3),
	.w4(32'hbb3b2d9f),
	.w5(32'hbb197d95),
	.w6(32'hbaeb00ec),
	.w7(32'hba1c3f94),
	.w8(32'hbb49ba63),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9ef05),
	.w1(32'hbb0ac7e4),
	.w2(32'h3b8ffcc9),
	.w3(32'hbba3596c),
	.w4(32'hb9591d1b),
	.w5(32'h3ad77fad),
	.w6(32'hbaf79d34),
	.w7(32'h3c18d771),
	.w8(32'h39cb89c8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3cd79),
	.w1(32'hb8112e3e),
	.w2(32'hb88481af),
	.w3(32'h3b54f3cb),
	.w4(32'h3aa237b4),
	.w5(32'hb9e5f360),
	.w6(32'h3aff9090),
	.w7(32'hbb0c6092),
	.w8(32'h3b8392c1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6d96),
	.w1(32'h3c038276),
	.w2(32'h3c15e647),
	.w3(32'h3c24077b),
	.w4(32'h3bef39cd),
	.w5(32'h3b9be07d),
	.w6(32'h3c28f157),
	.w7(32'h3b734c8b),
	.w8(32'hbc2bb90d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897fff),
	.w1(32'hba3f5992),
	.w2(32'hbb37a70a),
	.w3(32'hbbb560b3),
	.w4(32'hba93b1c8),
	.w5(32'hbb995a29),
	.w6(32'hbbdb0f0d),
	.w7(32'hbc0d44f0),
	.w8(32'hbc27f0a6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818f20),
	.w1(32'h3b79d3a3),
	.w2(32'h3b9aa6d4),
	.w3(32'h3a128266),
	.w4(32'h3b9b1bbc),
	.w5(32'h3b530d37),
	.w6(32'hbbc1c997),
	.w7(32'hbab1dc5a),
	.w8(32'h393dc8ae),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d8212),
	.w1(32'h3b27ecf0),
	.w2(32'hbb7a7cab),
	.w3(32'h3ae80ccb),
	.w4(32'h3ac65e55),
	.w5(32'hbbbd56ea),
	.w6(32'h3bfe5bca),
	.w7(32'hbbf89c9e),
	.w8(32'hbbb39c43),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb543ce),
	.w1(32'hbc33f78d),
	.w2(32'hbc29d3bd),
	.w3(32'hbb66732d),
	.w4(32'hbc1091a7),
	.w5(32'hbbf04d5e),
	.w6(32'hbbe1d04c),
	.w7(32'hbb97c059),
	.w8(32'h3ae39fbb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe6b1e),
	.w1(32'h3c0fe0bd),
	.w2(32'h3ba3b217),
	.w3(32'h3bcd2ece),
	.w4(32'h3be6b4dc),
	.w5(32'h3b1d6130),
	.w6(32'h3b792872),
	.w7(32'h3aa40117),
	.w8(32'hbb0541ae),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82c3a89),
	.w1(32'h3ab792d2),
	.w2(32'h3b55999c),
	.w3(32'hbab7b003),
	.w4(32'h3aa4f55a),
	.w5(32'h3bb18f78),
	.w6(32'hba417807),
	.w7(32'h3abde68b),
	.w8(32'h3b05180a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a814793),
	.w1(32'h3a21858c),
	.w2(32'h3b850610),
	.w3(32'h3bc1c4da),
	.w4(32'h39b3ec3e),
	.w5(32'hbb20d501),
	.w6(32'h3bcad405),
	.w7(32'hbb900f25),
	.w8(32'hbb41550d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b275a02),
	.w1(32'hbbca1591),
	.w2(32'hbc1d91f2),
	.w3(32'h3af560db),
	.w4(32'hbc02117d),
	.w5(32'hbb55e9a9),
	.w6(32'hbb36098e),
	.w7(32'hbbb766a6),
	.w8(32'hbb773e90),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2e59d),
	.w1(32'h3af120ae),
	.w2(32'h37061b60),
	.w3(32'h39d75080),
	.w4(32'h396f0998),
	.w5(32'hbba56111),
	.w6(32'h3ac52b05),
	.w7(32'hbad82c92),
	.w8(32'hba670218),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6113a0),
	.w1(32'h3bee2e27),
	.w2(32'h3b62e19a),
	.w3(32'hbb8ae4d9),
	.w4(32'h3bacfc7c),
	.w5(32'hba282aff),
	.w6(32'h3bc9f432),
	.w7(32'h3bae3b4c),
	.w8(32'hb9e11f97),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b6255),
	.w1(32'hbb958034),
	.w2(32'hbbb8dce9),
	.w3(32'h3a0159f1),
	.w4(32'h3a207a2c),
	.w5(32'hbb7ff903),
	.w6(32'h3b2159d9),
	.w7(32'hbc3180e5),
	.w8(32'hbc0a7671),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c74f04),
	.w1(32'h3ae4af8c),
	.w2(32'h3b7be49a),
	.w3(32'h3816b24c),
	.w4(32'h3a378210),
	.w5(32'h3b48e857),
	.w6(32'h3b7731e0),
	.w7(32'h3b446187),
	.w8(32'h3ad78931),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8eb20),
	.w1(32'hba71baa4),
	.w2(32'hba94c0de),
	.w3(32'h3b912356),
	.w4(32'hbb78c798),
	.w5(32'hbc2c4831),
	.w6(32'h3c1a1e4d),
	.w7(32'h3b8c8d96),
	.w8(32'h3badd6b3),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf15e9),
	.w1(32'hbb3da61e),
	.w2(32'hbab655a6),
	.w3(32'h3b4d973a),
	.w4(32'hbacac374),
	.w5(32'hba300292),
	.w6(32'h3bbecb7f),
	.w7(32'h3b5a394b),
	.w8(32'h3beee0ac),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beacf2a),
	.w1(32'h3b28c072),
	.w2(32'h3c23db92),
	.w3(32'h3c1f3987),
	.w4(32'h3c040d1a),
	.w5(32'h3c15c55b),
	.w6(32'h3b80e86b),
	.w7(32'h3c552e2a),
	.w8(32'hbafdb1b9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9ad0),
	.w1(32'hbbe76cf0),
	.w2(32'h3a74d559),
	.w3(32'hbc181949),
	.w4(32'h3ad038fd),
	.w5(32'h3bee1b17),
	.w6(32'hbbe4c8e8),
	.w7(32'hbb79a1fa),
	.w8(32'h3a054e45),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae63897),
	.w1(32'h3bae99eb),
	.w2(32'h39b20751),
	.w3(32'hbbc055e8),
	.w4(32'hbb9bda62),
	.w5(32'hbb9ef345),
	.w6(32'h3b6e0bf5),
	.w7(32'hbb6614a6),
	.w8(32'h3bfec0f4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c183cbf),
	.w1(32'h3c19baaf),
	.w2(32'h3c012e85),
	.w3(32'h3c22f410),
	.w4(32'h3c19c740),
	.w5(32'h3baf8eea),
	.w6(32'h3c081249),
	.w7(32'h3b351502),
	.w8(32'hbb9b4da9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62b391),
	.w1(32'hbc21ffab),
	.w2(32'hbc048551),
	.w3(32'h3b67d0cd),
	.w4(32'hbbbcff8d),
	.w5(32'hbbce8ac2),
	.w6(32'h3b84d646),
	.w7(32'h3bff010f),
	.w8(32'hb9bdd094),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b9582),
	.w1(32'h3b7cb3c7),
	.w2(32'h3b5ac5f7),
	.w3(32'hb9ee5fba),
	.w4(32'h3b1ccb87),
	.w5(32'h3aa01c51),
	.w6(32'h3afb273c),
	.w7(32'h3a84abf2),
	.w8(32'hbaf89de2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2e05d),
	.w1(32'hbb87f449),
	.w2(32'hbb1c3d53),
	.w3(32'hb98b5262),
	.w4(32'hbb1c0f9e),
	.w5(32'hbb29ba20),
	.w6(32'hbab429ae),
	.w7(32'hbb1f8290),
	.w8(32'hbb16e6ce),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed349c),
	.w1(32'hbaa7af87),
	.w2(32'hb95daf8c),
	.w3(32'hba45326f),
	.w4(32'h38c77f99),
	.w5(32'h3ace395d),
	.w6(32'h386c7526),
	.w7(32'h3a0f8943),
	.w8(32'h3a6d3f13),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7fcd96),
	.w1(32'h3ba342eb),
	.w2(32'h3b358384),
	.w3(32'h39fb25cb),
	.w4(32'h38da2186),
	.w5(32'hba8f9ebf),
	.w6(32'hbab05e85),
	.w7(32'hbb8b6d5b),
	.w8(32'h3a098342),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa95ee),
	.w1(32'h3bda3c9d),
	.w2(32'h3bc56e00),
	.w3(32'h3b7024d0),
	.w4(32'h3ba508c8),
	.w5(32'h3b869ce2),
	.w6(32'h3bac982e),
	.w7(32'h3b7d15e7),
	.w8(32'h3c8f49e7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ee993),
	.w1(32'h3be04d70),
	.w2(32'h3c24ae13),
	.w3(32'h3c820971),
	.w4(32'h3c5a4081),
	.w5(32'h3c469206),
	.w6(32'h3cc30b97),
	.w7(32'h3c188fcd),
	.w8(32'hbc0885ed),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83b296),
	.w1(32'hba709118),
	.w2(32'h3ab9aa17),
	.w3(32'hbac33024),
	.w4(32'hba806046),
	.w5(32'h39b2ff17),
	.w6(32'hba8ef173),
	.w7(32'h3a299431),
	.w8(32'h3acfa5aa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c25e6),
	.w1(32'h3bae3c3a),
	.w2(32'h3b9a5582),
	.w3(32'h3b490de5),
	.w4(32'h3b795251),
	.w5(32'h3b4bdba5),
	.w6(32'h3b9a00b6),
	.w7(32'h3aed0676),
	.w8(32'hbba4834b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaeb77),
	.w1(32'hbbc0f1b9),
	.w2(32'hb9ecd7a1),
	.w3(32'hbb954fe7),
	.w4(32'hbb90d2e4),
	.w5(32'hba4ee48d),
	.w6(32'hbb99f551),
	.w7(32'hbab04f22),
	.w8(32'hbbc6b5fb),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be01bf0),
	.w1(32'hbacd0124),
	.w2(32'hbb8aed87),
	.w3(32'h3bcd68ab),
	.w4(32'hba9af0b6),
	.w5(32'hbb001e8b),
	.w6(32'hbc00fe4a),
	.w7(32'hbc0fbb93),
	.w8(32'hbb5ec489),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7351b),
	.w1(32'h3ade991d),
	.w2(32'h3bb4d6d9),
	.w3(32'hbb3e2a1a),
	.w4(32'h3a93e9bb),
	.w5(32'h3b887a14),
	.w6(32'hb9e99771),
	.w7(32'h3b326ddc),
	.w8(32'hba8b0e24),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7264e),
	.w1(32'hba17aaea),
	.w2(32'h3965eccb),
	.w3(32'hba21b04c),
	.w4(32'hb9a8b821),
	.w5(32'hb893e1c3),
	.w6(32'hba004b5f),
	.w7(32'hba44f531),
	.w8(32'hbb6eb254),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5aba8),
	.w1(32'hbab745b5),
	.w2(32'h3ad90b93),
	.w3(32'hbb67dbf6),
	.w4(32'hbb2a9b66),
	.w5(32'hb8db3680),
	.w6(32'hbaf7aeaf),
	.w7(32'h3a113f24),
	.w8(32'h3caa8357),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c672a16),
	.w1(32'h3c11c2c6),
	.w2(32'h3c1b990e),
	.w3(32'h3c68dcbb),
	.w4(32'h3c181578),
	.w5(32'h3bf4ee0c),
	.w6(32'h3caf4827),
	.w7(32'h3c2ea143),
	.w8(32'h3ba75450),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01148e),
	.w1(32'h3bde9aa3),
	.w2(32'h3bb81df4),
	.w3(32'h3bea00b5),
	.w4(32'h3b83a5b6),
	.w5(32'h3a75165d),
	.w6(32'h3c2cd955),
	.w7(32'h3b963ad8),
	.w8(32'hba6c8be0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38982e),
	.w1(32'h3a0a2a04),
	.w2(32'h3a54bfa2),
	.w3(32'h3adf4791),
	.w4(32'h3b06a9b2),
	.w5(32'h398bbce2),
	.w6(32'h3a894a6b),
	.w7(32'hb9910f2b),
	.w8(32'hbb899171),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea3edc),
	.w1(32'hbc62289f),
	.w2(32'hbc3a8cc2),
	.w3(32'hba0e4d8c),
	.w4(32'hbb3a8b09),
	.w5(32'h3b2ec2d9),
	.w6(32'hbc1b7d71),
	.w7(32'hbba6d3fe),
	.w8(32'hbb015896),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd1a34),
	.w1(32'h3a55c5ed),
	.w2(32'h3ba01830),
	.w3(32'hbb213672),
	.w4(32'hbad415ca),
	.w5(32'h3aee7351),
	.w6(32'h3b6344f0),
	.w7(32'h3b2f723f),
	.w8(32'h3ac35607),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ea701),
	.w1(32'h3b934972),
	.w2(32'h3a2ee2e1),
	.w3(32'h3b76c6c3),
	.w4(32'h3b3242c0),
	.w5(32'hbb457143),
	.w6(32'h3b4624f1),
	.w7(32'hbbdf2f16),
	.w8(32'h3b07545a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06ca3f),
	.w1(32'hbc8d95f0),
	.w2(32'hbb85597b),
	.w3(32'h3b325925),
	.w4(32'hbb89c6a0),
	.w5(32'hbb9b4d81),
	.w6(32'hbc286ba7),
	.w7(32'hbc14fabd),
	.w8(32'h3b6a36a6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b005cca),
	.w1(32'hbaa4107d),
	.w2(32'hbaf83a64),
	.w3(32'h3bb2f4ff),
	.w4(32'h3987767e),
	.w5(32'hbb815c47),
	.w6(32'h3b6f7952),
	.w7(32'hbbad8ff7),
	.w8(32'h3ac59597),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1767ec),
	.w1(32'h3c3d2ae0),
	.w2(32'h3c59e191),
	.w3(32'h3c163786),
	.w4(32'h3c1029e6),
	.w5(32'h3c1c6de4),
	.w6(32'h3c17d4b1),
	.w7(32'h3bfe04f3),
	.w8(32'hbb0125cb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefbdcd),
	.w1(32'hbc597e0d),
	.w2(32'hbc503ffa),
	.w3(32'hbb9ab231),
	.w4(32'hbc314d9f),
	.w5(32'hbc17ad15),
	.w6(32'hbc120eff),
	.w7(32'hbba16b1f),
	.w8(32'hbb4cbb18),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41c64a),
	.w1(32'h3b73c5ba),
	.w2(32'h3b341e17),
	.w3(32'h39f6461e),
	.w4(32'h3b706d5f),
	.w5(32'h3abada4f),
	.w6(32'h3aa03d94),
	.w7(32'h39e3b7da),
	.w8(32'h3b576e2e),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b173bbc),
	.w1(32'h3a495dab),
	.w2(32'h3b3f58a5),
	.w3(32'h3ba94fd5),
	.w4(32'h3ba4790b),
	.w5(32'h3bcc10e2),
	.w6(32'h3b026f72),
	.w7(32'h3bad0296),
	.w8(32'hbafc4090),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe05213),
	.w1(32'hbc48ced4),
	.w2(32'hbc42495b),
	.w3(32'hbb9ad494),
	.w4(32'hbc1d91ef),
	.w5(32'hbc070af4),
	.w6(32'hbc0e1957),
	.w7(32'hbb9ab98c),
	.w8(32'hbad38e73),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb23be),
	.w1(32'hbc3a99d5),
	.w2(32'hbc24bdd6),
	.w3(32'hbb7bad20),
	.w4(32'hbc144a2a),
	.w5(32'hbbf41021),
	.w6(32'hbbeb340f),
	.w7(32'hbb857417),
	.w8(32'hba8f908b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa703d5),
	.w1(32'hb9578a40),
	.w2(32'h3a88a660),
	.w3(32'hb9ffe8d7),
	.w4(32'h3a3ec30d),
	.w5(32'h3a942a6a),
	.w6(32'hba3774d8),
	.w7(32'h3ab8db56),
	.w8(32'h3b70d3ee),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c123c77),
	.w1(32'h3c023195),
	.w2(32'h3ba61095),
	.w3(32'h3b903dbb),
	.w4(32'h3c062b18),
	.w5(32'h3bbd43e4),
	.w6(32'h3bf02173),
	.w7(32'h3b18fdd4),
	.w8(32'h3933ff5c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b8c6f),
	.w1(32'hb946beef),
	.w2(32'h398ab35a),
	.w3(32'h39edbc98),
	.w4(32'hba356067),
	.w5(32'hb9f44967),
	.w6(32'h3a24ebfb),
	.w7(32'hba9b1c0a),
	.w8(32'h3a409816),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb489dc9),
	.w1(32'hbbd91896),
	.w2(32'hbc080140),
	.w3(32'hbb10f045),
	.w4(32'hbbe4d374),
	.w5(32'hbbd73579),
	.w6(32'h3be28faf),
	.w7(32'hb882f9f5),
	.w8(32'hba95ebc8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c952a),
	.w1(32'hbb1031a8),
	.w2(32'hbb24fbb9),
	.w3(32'h3b77ed4b),
	.w4(32'h3a94dac1),
	.w5(32'hbab79ca4),
	.w6(32'h39da0b13),
	.w7(32'hbb191c30),
	.w8(32'hbc3dda91),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c7a96),
	.w1(32'h3c1fcfce),
	.w2(32'h3b47dd04),
	.w3(32'hbb88edd7),
	.w4(32'hbbca4f46),
	.w5(32'hbc0164ec),
	.w6(32'h3aab6cd9),
	.w7(32'hbb97f4f5),
	.w8(32'h3ac40dbf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabe63d),
	.w1(32'hba9a1524),
	.w2(32'h3a82320f),
	.w3(32'h3b95e34e),
	.w4(32'h3b647a2e),
	.w5(32'h3aadd1e0),
	.w6(32'h3b07fb1b),
	.w7(32'h3b9aa444),
	.w8(32'h3c95526a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e3ed3),
	.w1(32'h3c20123e),
	.w2(32'h3c2abce3),
	.w3(32'h3c30d1b7),
	.w4(32'h3bffbe5b),
	.w5(32'h3bf5e3b7),
	.w6(32'h3c887399),
	.w7(32'h3c6332ad),
	.w8(32'hbb5b06c2),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c065a),
	.w1(32'h3a4524c8),
	.w2(32'h3abd4060),
	.w3(32'hbb21a6dd),
	.w4(32'h3987cf13),
	.w5(32'hba9126db),
	.w6(32'hb99b0de2),
	.w7(32'hba8dd5f3),
	.w8(32'h3a194c41),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9909c26),
	.w1(32'hba18b8aa),
	.w2(32'h3b249c4b),
	.w3(32'hb90a148d),
	.w4(32'h3b063bbc),
	.w5(32'h3b0fbf39),
	.w6(32'hba86a12e),
	.w7(32'h3b2d0272),
	.w8(32'hba257184),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba292b5d),
	.w1(32'h39a907ca),
	.w2(32'h3b20fdd3),
	.w3(32'hba887953),
	.w4(32'h3a41d770),
	.w5(32'h3b12ad68),
	.w6(32'h3982a8ad),
	.w7(32'h3acd2234),
	.w8(32'h3c687235),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c506ede),
	.w1(32'h3c9dbfdc),
	.w2(32'h3c83d2ef),
	.w3(32'h3c2a1097),
	.w4(32'h3c3fb91a),
	.w5(32'h3c13577d),
	.w6(32'h3ca119bf),
	.w7(32'h3c4a5932),
	.w8(32'hbae1bff4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95d5d6b),
	.w1(32'hb96c32ca),
	.w2(32'h3b27f0d0),
	.w3(32'h3847cea3),
	.w4(32'h3a4d40ce),
	.w5(32'h3b5643e0),
	.w6(32'h3aec6373),
	.w7(32'h3b64da0b),
	.w8(32'h39a084aa),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57389b),
	.w1(32'hbbaa1ed0),
	.w2(32'hbb9942ed),
	.w3(32'hbb016c7b),
	.w4(32'hbb69a3c8),
	.w5(32'hbb26ad8b),
	.w6(32'hbb6ba571),
	.w7(32'hbabefbe8),
	.w8(32'h3a399f7a),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb1655),
	.w1(32'hba453d18),
	.w2(32'hb9b57e8f),
	.w3(32'h3b54a512),
	.w4(32'h3ae3d464),
	.w5(32'hb98d5901),
	.w6(32'h3b79790b),
	.w7(32'hba28b38d),
	.w8(32'hbb2606ba),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91817bd),
	.w1(32'hba92494e),
	.w2(32'h3a9fc855),
	.w3(32'h3a235861),
	.w4(32'hba4de95c),
	.w5(32'h3ad5ed44),
	.w6(32'h3a6ed9a8),
	.w7(32'h3abbc19f),
	.w8(32'hba073a78),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87e53ce),
	.w1(32'h3a0b1888),
	.w2(32'h3a5f7f10),
	.w3(32'h3a206613),
	.w4(32'h3ab998bc),
	.w5(32'h3ab7f31f),
	.w6(32'h3a29e619),
	.w7(32'h3aa30a02),
	.w8(32'h3a2dd400),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920bc01),
	.w1(32'h398b2e96),
	.w2(32'h3a30ad21),
	.w3(32'h3990583b),
	.w4(32'h39eabe7b),
	.w5(32'h3a166f63),
	.w6(32'h3974fc29),
	.w7(32'h3a67c792),
	.w8(32'hb9e7dede),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948357),
	.w1(32'hba6afa43),
	.w2(32'hba8cedfd),
	.w3(32'hba88aad3),
	.w4(32'hb9be87a7),
	.w5(32'hb972fa39),
	.w6(32'hba9af025),
	.w7(32'hbab6dddc),
	.w8(32'hb826ec3c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38be48cc),
	.w1(32'h3aac2a5f),
	.w2(32'hbb149b5e),
	.w3(32'hb7584b72),
	.w4(32'h3a8cfa5b),
	.w5(32'h3a839d24),
	.w6(32'hb95f3eac),
	.w7(32'hbaec1ea4),
	.w8(32'hbb59fced),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dd70e),
	.w1(32'hbba344c3),
	.w2(32'hbb4eff0c),
	.w3(32'hbb1204fe),
	.w4(32'hbb81a04e),
	.w5(32'hbb5841a5),
	.w6(32'hbb409724),
	.w7(32'hbb4f891a),
	.w8(32'hba7da724),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b4cfd),
	.w1(32'hbaf39ccc),
	.w2(32'hb9fcb271),
	.w3(32'hb993c2ba),
	.w4(32'hb9e93e33),
	.w5(32'h3a7fed2f),
	.w6(32'hba42142c),
	.w7(32'h3a08ff10),
	.w8(32'h3a637c90),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c1dad3),
	.w1(32'h39fb62ed),
	.w2(32'h3a43d013),
	.w3(32'h39b0762f),
	.w4(32'h3a0e4dce),
	.w5(32'h3a3405df),
	.w6(32'hb86bc711),
	.w7(32'h3a08e904),
	.w8(32'hba08d3de),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38043e44),
	.w1(32'hb98fdee3),
	.w2(32'hba32e19b),
	.w3(32'hb68ba6ce),
	.w4(32'hb9b1f2e1),
	.w5(32'hba62c412),
	.w6(32'hbab16bed),
	.w7(32'hb7ed8d1c),
	.w8(32'hbaeb9e20),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57bcce),
	.w1(32'hb9e8aa31),
	.w2(32'hb9d534f8),
	.w3(32'hba248a8f),
	.w4(32'hba05a963),
	.w5(32'hba5c34a8),
	.w6(32'hba8ebd15),
	.w7(32'hba0ebc14),
	.w8(32'h3a12ecf6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac87078),
	.w1(32'hbaa68386),
	.w2(32'hba58b901),
	.w3(32'h3a4ec34c),
	.w4(32'hba00a100),
	.w5(32'hba35e288),
	.w6(32'h3a9b7e6f),
	.w7(32'h3a07683d),
	.w8(32'h3812a3f5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acfeaab),
	.w1(32'hba632322),
	.w2(32'hbac15d04),
	.w3(32'h3b225e99),
	.w4(32'h3a1cf0a7),
	.w5(32'hba8e5924),
	.w6(32'h3ad672a8),
	.w7(32'hbadd6bee),
	.w8(32'hba081929),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add14c9),
	.w1(32'hb983ff41),
	.w2(32'hbad5c7e6),
	.w3(32'h3ab31b0c),
	.w4(32'h3aba5ba0),
	.w5(32'hb9331f12),
	.w6(32'h38f87efd),
	.w7(32'hbb01ca5e),
	.w8(32'hbb2fcae5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1778ea),
	.w1(32'hbb463719),
	.w2(32'hbb2b2dee),
	.w3(32'hbb4ff8ce),
	.w4(32'hbb6168a0),
	.w5(32'hbb1435ea),
	.w6(32'hbb28b3b1),
	.w7(32'hbb1f6957),
	.w8(32'hbac42d7a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e9c6e),
	.w1(32'hbb1cafa7),
	.w2(32'hbaae8e3e),
	.w3(32'hbb1eaa15),
	.w4(32'hbaee6f0b),
	.w5(32'hbae89018),
	.w6(32'hbacd07fe),
	.w7(32'hba71e1fe),
	.w8(32'h3adb0a44),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60cfb3),
	.w1(32'hba21f5b7),
	.w2(32'hb922c4c8),
	.w3(32'h3aa49ebf),
	.w4(32'hb7cb09a4),
	.w5(32'hbac8bd32),
	.w6(32'h39bcc9f5),
	.w7(32'hbb05cd51),
	.w8(32'h3b55a7b8),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca3956),
	.w1(32'h39c8aea4),
	.w2(32'h3a2a99cc),
	.w3(32'h3adab9af),
	.w4(32'h39fa88a4),
	.w5(32'h3a00a67e),
	.w6(32'h3a92c446),
	.w7(32'h3aaf2068),
	.w8(32'h38e6da0d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f79a8),
	.w1(32'h3a2ea17c),
	.w2(32'hb93fc9f7),
	.w3(32'h391b0f62),
	.w4(32'h38e83dcf),
	.w5(32'h3a9e57e2),
	.w6(32'hb9e34f37),
	.w7(32'hba1c4089),
	.w8(32'hb82ff532),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b5620),
	.w1(32'h3a954fe9),
	.w2(32'hba960619),
	.w3(32'hbadf6758),
	.w4(32'hba3695ca),
	.w5(32'h3a6fe257),
	.w6(32'hbac2ad1b),
	.w7(32'hb986ea46),
	.w8(32'hb99f32bb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4b2c),
	.w1(32'hbb40427a),
	.w2(32'hbab4e205),
	.w3(32'hbab033c8),
	.w4(32'hba5531d3),
	.w5(32'hbadefd7c),
	.w6(32'hba5bed24),
	.w7(32'hba9d2299),
	.w8(32'hbb4528d1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accd99c),
	.w1(32'h3a104e5c),
	.w2(32'hba91b3fc),
	.w3(32'h3a917777),
	.w4(32'hb7faf174),
	.w5(32'hbab6da24),
	.w6(32'h3a301bec),
	.w7(32'h39c17140),
	.w8(32'hb9f5a41b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfb9d4),
	.w1(32'hbb9fe9dd),
	.w2(32'hbaf8748c),
	.w3(32'hbb166142),
	.w4(32'hbb79469e),
	.w5(32'hbb9960aa),
	.w6(32'h3afe4bd7),
	.w7(32'hba8a8572),
	.w8(32'hbb9b536e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule