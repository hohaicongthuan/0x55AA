module layer_10_featuremap_55(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ec787),
	.w1(32'hbb11c208),
	.w2(32'hbb0c3e55),
	.w3(32'hb9b60061),
	.w4(32'h3b27c486),
	.w5(32'hbc30bcc0),
	.w6(32'h3a9062b1),
	.w7(32'h3c1183fc),
	.w8(32'hbc7e75e3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dd073),
	.w1(32'hbb5bba13),
	.w2(32'h3b9a34ab),
	.w3(32'hbc5c10be),
	.w4(32'hbb246f67),
	.w5(32'hbb1d3979),
	.w6(32'hbbc28cde),
	.w7(32'h3b8a8ea0),
	.w8(32'h3ba52dd2),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbd9ae),
	.w1(32'h3c141e89),
	.w2(32'hbb0496e2),
	.w3(32'hbc2686ff),
	.w4(32'hbc04c58a),
	.w5(32'hbb4825de),
	.w6(32'h3c3b076d),
	.w7(32'h3b7f6ca4),
	.w8(32'hbbda20c2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8888c8),
	.w1(32'hbafe715b),
	.w2(32'hbb922980),
	.w3(32'h3a39af65),
	.w4(32'h3b120721),
	.w5(32'h3b5981aa),
	.w6(32'hbc402385),
	.w7(32'hbc2daef4),
	.w8(32'h3baa11f1),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4029bf),
	.w1(32'hbc1f29ee),
	.w2(32'hbbee5d9d),
	.w3(32'hb68e5f74),
	.w4(32'hbb067c31),
	.w5(32'hbbb498fd),
	.w6(32'h3b2daab8),
	.w7(32'h3b0196d8),
	.w8(32'hbc10ebc8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cde22),
	.w1(32'h399f5e81),
	.w2(32'hbb934792),
	.w3(32'hbc06652c),
	.w4(32'h3a09334c),
	.w5(32'hbbaa0755),
	.w6(32'hba849a92),
	.w7(32'h3aefcc85),
	.w8(32'hbb5b7245),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33c3b3),
	.w1(32'hbb29bbe2),
	.w2(32'h3bf68ea5),
	.w3(32'hba130b5f),
	.w4(32'hbb2861f1),
	.w5(32'h3b9fbcb6),
	.w6(32'h3a5e50ac),
	.w7(32'h3ac4eecb),
	.w8(32'hba2ec4ef),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6ecff),
	.w1(32'hbbb78257),
	.w2(32'hbba696d1),
	.w3(32'h3b7b6f9f),
	.w4(32'h3b38ab49),
	.w5(32'hbc17b412),
	.w6(32'hbc69741a),
	.w7(32'hbc3629d6),
	.w8(32'hbbdf900f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba36842),
	.w1(32'h3b7f2c08),
	.w2(32'h3b555887),
	.w3(32'hbbac4aa2),
	.w4(32'h3b79a535),
	.w5(32'hbb866552),
	.w6(32'hbb555262),
	.w7(32'hbba78f39),
	.w8(32'hbbcffaea),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b2655),
	.w1(32'h3c483970),
	.w2(32'h3b5bbac3),
	.w3(32'h3b06e845),
	.w4(32'h3c469304),
	.w5(32'hba920520),
	.w6(32'hbbdfeb7a),
	.w7(32'hbb616385),
	.w8(32'h3b56e9f3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c405),
	.w1(32'h3b29393f),
	.w2(32'hbbcfb459),
	.w3(32'h3980e6a9),
	.w4(32'h3a6e96a7),
	.w5(32'hbbaaff05),
	.w6(32'h3b521dfa),
	.w7(32'h3b57a237),
	.w8(32'hbc254f13),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aa4ad),
	.w1(32'h3ac5cc9a),
	.w2(32'hbadc548d),
	.w3(32'h3b7ac34a),
	.w4(32'h3bb0e7c0),
	.w5(32'hbb5be812),
	.w6(32'hbc1d3ccf),
	.w7(32'hbc30696f),
	.w8(32'hbb1e09d8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d236),
	.w1(32'h38bfcbf9),
	.w2(32'hbbcbe8e7),
	.w3(32'hbacf0770),
	.w4(32'hb988e4a4),
	.w5(32'hbbea0b0f),
	.w6(32'hbb359f1b),
	.w7(32'hbb2bd8e7),
	.w8(32'hbb49d8a0),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58a958),
	.w1(32'hbbb7bd04),
	.w2(32'hbb0d5683),
	.w3(32'hba65bdaf),
	.w4(32'hbb40cfc4),
	.w5(32'hbb8ae3be),
	.w6(32'h3b25f6a5),
	.w7(32'h3ab9334a),
	.w8(32'hbbc85025),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba18962),
	.w1(32'h3a87c7bd),
	.w2(32'h3b73b334),
	.w3(32'h3a1046d3),
	.w4(32'h3b724bc4),
	.w5(32'hbb08e214),
	.w6(32'hbb60b662),
	.w7(32'hbad2d399),
	.w8(32'hbb2e51fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3952fae7),
	.w1(32'h3ac4b38e),
	.w2(32'h3a7bd3d5),
	.w3(32'hbaa5d286),
	.w4(32'h3afa44cb),
	.w5(32'hb9fdf7a8),
	.w6(32'hbbb8a336),
	.w7(32'hbbc9fb3a),
	.w8(32'h3b1d597d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b394bbb),
	.w1(32'h3b81f206),
	.w2(32'hbac60bc5),
	.w3(32'hb901e353),
	.w4(32'hb995d3ac),
	.w5(32'hbae02377),
	.w6(32'h3b415ce3),
	.w7(32'h3ae78fe0),
	.w8(32'hbb8beae5),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ee590),
	.w1(32'hbbf4d580),
	.w2(32'hbc299210),
	.w3(32'hbc4636b2),
	.w4(32'hbc2691e3),
	.w5(32'hbc81c936),
	.w6(32'hbc79ea36),
	.w7(32'hbc309275),
	.w8(32'hbc4b27f6),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42e1b4),
	.w1(32'hba66c45d),
	.w2(32'hba80f8b3),
	.w3(32'hbb1813d8),
	.w4(32'hbb461e17),
	.w5(32'hbb9a3056),
	.w6(32'hbbc1cdd4),
	.w7(32'hbc1e4320),
	.w8(32'hbc1587f2),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c1568),
	.w1(32'hbc1208c8),
	.w2(32'hbb347064),
	.w3(32'h3b0078ba),
	.w4(32'h3b77d69d),
	.w5(32'h3b87828f),
	.w6(32'hbbe80d1c),
	.w7(32'hbbf79d82),
	.w8(32'hbaf0ef29),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab50eb0),
	.w1(32'hbb17ed67),
	.w2(32'h3b028266),
	.w3(32'h3b9fa36c),
	.w4(32'h3a90ad47),
	.w5(32'hba1f2d76),
	.w6(32'hbb060c42),
	.w7(32'h39b2e878),
	.w8(32'hbb646933),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f1236d),
	.w1(32'hbb1c858c),
	.w2(32'h3a30a76b),
	.w3(32'hbb9b37dd),
	.w4(32'hbc0cf329),
	.w5(32'hbafafa1e),
	.w6(32'hbb3e736b),
	.w7(32'hbb2c6b6f),
	.w8(32'h3a3908d1),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bc022),
	.w1(32'hbc8819c3),
	.w2(32'hbc46bcb3),
	.w3(32'hbc0c612c),
	.w4(32'hbc2e03b2),
	.w5(32'hbc2b27d9),
	.w6(32'hbc2affb0),
	.w7(32'hbc032f22),
	.w8(32'hbc3972a0),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07698f),
	.w1(32'h3b30d78a),
	.w2(32'h3b20c545),
	.w3(32'h3bbe64b6),
	.w4(32'h3c04d553),
	.w5(32'h3a3cd820),
	.w6(32'h3ba01803),
	.w7(32'h3bd78251),
	.w8(32'h3b127ac5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba64b737),
	.w1(32'hbba0df2e),
	.w2(32'h3c14b31a),
	.w3(32'h3b4d45f0),
	.w4(32'hbafc7362),
	.w5(32'hbbae5f7e),
	.w6(32'h3b9838b1),
	.w7(32'hbb0505c0),
	.w8(32'hbc06c568),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1106b8),
	.w1(32'h3a1953b1),
	.w2(32'h3b0b5a53),
	.w3(32'hbbbc5b82),
	.w4(32'hbb955f37),
	.w5(32'h3c53ea85),
	.w6(32'hbc18373e),
	.w7(32'hbbc9475d),
	.w8(32'h3c81ea99),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd3d828),
	.w1(32'hbc849eac),
	.w2(32'hb9633393),
	.w3(32'h3b7418bb),
	.w4(32'h3a92017b),
	.w5(32'hb9796e25),
	.w6(32'h3bf3d56b),
	.w7(32'h3ba66f29),
	.w8(32'hb81fbad5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab253b6),
	.w1(32'h3a4edb74),
	.w2(32'h3969ffc6),
	.w3(32'h3a3d465f),
	.w4(32'h3ad6eb76),
	.w5(32'h38c4f48f),
	.w6(32'h3b177bab),
	.w7(32'h3acf2494),
	.w8(32'h39c2fc1d),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23ecaf),
	.w1(32'hb9c899b1),
	.w2(32'hbadecb07),
	.w3(32'hbac5a028),
	.w4(32'hbaa397ee),
	.w5(32'hbafdd2fb),
	.w6(32'hbab59995),
	.w7(32'hbac5415e),
	.w8(32'hbaaac158),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4179eb),
	.w1(32'h3af8d25c),
	.w2(32'h3ae1d634),
	.w3(32'h3b263c95),
	.w4(32'h3b48fcb5),
	.w5(32'h3a24404d),
	.w6(32'h3b6981b0),
	.w7(32'h3b3d714c),
	.w8(32'h3b2f4edc),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391787a1),
	.w1(32'hb7cd5a7d),
	.w2(32'h3a2708d0),
	.w3(32'hb9991dfc),
	.w4(32'hb9c4cc38),
	.w5(32'h39b2d725),
	.w6(32'hb9d4e6e9),
	.w7(32'hba05d993),
	.w8(32'h39e799d4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3d749),
	.w1(32'h3a48e5b6),
	.w2(32'hba8f94de),
	.w3(32'h3a6859f3),
	.w4(32'h39f4ca2b),
	.w5(32'hb9997bd3),
	.w6(32'h3ae49dbd),
	.w7(32'h3abb4a5e),
	.w8(32'hba4d6756),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba523a26),
	.w1(32'hb9489d07),
	.w2(32'h3a68b487),
	.w3(32'h3a5e7600),
	.w4(32'h39d7f413),
	.w5(32'h3991bbf3),
	.w6(32'hba84a6a0),
	.w7(32'hba894714),
	.w8(32'h39cd9453),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b11a3b),
	.w1(32'h3b002c4c),
	.w2(32'h3af6ad2a),
	.w3(32'h3b046a31),
	.w4(32'h3b184743),
	.w5(32'h3b286aa3),
	.w6(32'h3abc8648),
	.w7(32'h3ad082f2),
	.w8(32'h3b36a756),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4710d0),
	.w1(32'h3984e59e),
	.w2(32'hb98a73bd),
	.w3(32'h3ad0eb3c),
	.w4(32'h38930970),
	.w5(32'hb98fca89),
	.w6(32'hb9835fab),
	.w7(32'hb99dd538),
	.w8(32'hb9fc5a95),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0353bd),
	.w1(32'hb9cc01b4),
	.w2(32'h394666c5),
	.w3(32'hb9b6bdb3),
	.w4(32'hba37afd6),
	.w5(32'h3a579a2a),
	.w6(32'hba7129b5),
	.w7(32'hba01543a),
	.w8(32'h3aa5be00),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeacef2),
	.w1(32'hbae808c9),
	.w2(32'hbac75872),
	.w3(32'h36b3c952),
	.w4(32'hbb05fe1d),
	.w5(32'h3a945a40),
	.w6(32'hbb00ae5c),
	.w7(32'hba191fb6),
	.w8(32'hba9b4041),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb405f),
	.w1(32'h3c12e4e2),
	.w2(32'h3ba95986),
	.w3(32'h3b490531),
	.w4(32'h3bc8d58c),
	.w5(32'h3b457f96),
	.w6(32'h3b9b53ac),
	.w7(32'h3ba198c6),
	.w8(32'h3b8f7896),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9050bcd),
	.w1(32'h3bc89dcf),
	.w2(32'h3bf2ac32),
	.w3(32'h3b4cb0e9),
	.w4(32'h3b96b656),
	.w5(32'h3b4c9e5d),
	.w6(32'h3bcddc6f),
	.w7(32'h3bb1bdcd),
	.w8(32'h3b9e9c08),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6d965),
	.w1(32'h3aeb725b),
	.w2(32'h3afbd35e),
	.w3(32'h3ab8c8b3),
	.w4(32'h3a09d2fd),
	.w5(32'h3a7cbf09),
	.w6(32'h3aa264ca),
	.w7(32'h3a2d0478),
	.w8(32'h3a9df763),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e7e74),
	.w1(32'h39dcd5b5),
	.w2(32'hbaa59c98),
	.w3(32'hb9c81185),
	.w4(32'h3994d934),
	.w5(32'hbaf7604f),
	.w6(32'hba065a94),
	.w7(32'hb89c8943),
	.w8(32'hbab43172),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf767c7),
	.w1(32'hbaa9ea6b),
	.w2(32'h39fcb29e),
	.w3(32'hbb21f02d),
	.w4(32'hbb05ada9),
	.w5(32'hb8b1a43b),
	.w6(32'hbb006408),
	.w7(32'hbad61d85),
	.w8(32'h39c34d2e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b5845),
	.w1(32'h3a9b808c),
	.w2(32'h3a1c781f),
	.w3(32'hb9918004),
	.w4(32'h3a383554),
	.w5(32'hb97d215e),
	.w6(32'h3a79d2ff),
	.w7(32'h3afd9e8f),
	.w8(32'hb996168b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ccf2d),
	.w1(32'hbaa7189d),
	.w2(32'hb8c30869),
	.w3(32'hbb0bca62),
	.w4(32'hbb0c32e3),
	.w5(32'hbb69ef12),
	.w6(32'hbb72a753),
	.w7(32'hbb637b0a),
	.w8(32'hbb1266b8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f463a4),
	.w1(32'h3b61bb80),
	.w2(32'h3b377fea),
	.w3(32'h3abb972d),
	.w4(32'h3b8fad4c),
	.w5(32'h3acb1e1d),
	.w6(32'h3a848301),
	.w7(32'h3b27c0a9),
	.w8(32'h3b64138d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917a150),
	.w1(32'h3b54f0d3),
	.w2(32'h3b01df77),
	.w3(32'h3ba614f9),
	.w4(32'h3b96c56c),
	.w5(32'hbb0f4d2d),
	.w6(32'h3b66df82),
	.w7(32'h3b1a1109),
	.w8(32'h3a88b91b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff3070),
	.w1(32'hba7de9a1),
	.w2(32'h398a41a4),
	.w3(32'h39f14e00),
	.w4(32'h391d8f5d),
	.w5(32'h3b24bcd7),
	.w6(32'hbbad825d),
	.w7(32'hbab3f407),
	.w8(32'h3b0cfda6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2ec23),
	.w1(32'hbc44a0d7),
	.w2(32'hbc2effab),
	.w3(32'hbc45b4e0),
	.w4(32'hbc5d7321),
	.w5(32'hbc594ea8),
	.w6(32'hbc931ceb),
	.w7(32'hbc5f4df7),
	.w8(32'hbc3b26ee),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22571),
	.w1(32'hbac33ba4),
	.w2(32'hba8d2de0),
	.w3(32'hbabcd54e),
	.w4(32'hbaefeb61),
	.w5(32'h37537dd9),
	.w6(32'hbac182e4),
	.w7(32'hbae753fc),
	.w8(32'hba8b85e4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984f830),
	.w1(32'hba2f53b0),
	.w2(32'h3a7d5f8e),
	.w3(32'h39985494),
	.w4(32'hb8c38a9e),
	.w5(32'h3979b349),
	.w6(32'hb885a8f8),
	.w7(32'hb9e6dc81),
	.w8(32'h39fc54eb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fb4b42),
	.w1(32'hb9e3af2a),
	.w2(32'h3936b08a),
	.w3(32'hba4976b9),
	.w4(32'hba0a7928),
	.w5(32'hbab9164c),
	.w6(32'hba985d90),
	.w7(32'hba5a3cea),
	.w8(32'hbaa28e39),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e3ebd),
	.w1(32'hbb0e97f6),
	.w2(32'hba8925f2),
	.w3(32'hbb35e6f8),
	.w4(32'hb9417e77),
	.w5(32'hba5219e9),
	.w6(32'hbaf6ffd4),
	.w7(32'hbab6f43e),
	.w8(32'hbaa467f8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c70119),
	.w1(32'hbabfa4ea),
	.w2(32'hba2fb95f),
	.w3(32'h392ba92c),
	.w4(32'hb98119c3),
	.w5(32'h3a2599ac),
	.w6(32'hbad83beb),
	.w7(32'hba14cf1c),
	.w8(32'h38950a15),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02588e),
	.w1(32'hbbc323da),
	.w2(32'hbbae639d),
	.w3(32'hbb8a0195),
	.w4(32'hbbb57806),
	.w5(32'hbbd9f3c7),
	.w6(32'hbc00173e),
	.w7(32'hbbd76712),
	.w8(32'hbbac3840),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae20f39),
	.w1(32'hbabb2d64),
	.w2(32'hbafd5efc),
	.w3(32'hbac07842),
	.w4(32'hba332dbc),
	.w5(32'hba6bf380),
	.w6(32'hba1cbbac),
	.w7(32'hb8d2fd80),
	.w8(32'hba746c8c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba193bf0),
	.w1(32'hb979c925),
	.w2(32'hba364d90),
	.w3(32'h3963cea6),
	.w4(32'hb984197d),
	.w5(32'hba49a490),
	.w6(32'h382f6462),
	.w7(32'hba58606a),
	.w8(32'hba637743),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab804b4),
	.w1(32'hba6f2997),
	.w2(32'h3b120b59),
	.w3(32'hbae664a8),
	.w4(32'hba75716c),
	.w5(32'h3a9ac900),
	.w6(32'hba71e2a4),
	.w7(32'hbaa0afa8),
	.w8(32'h3a9379b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91ffe0),
	.w1(32'h3a59815d),
	.w2(32'hb7aedd36),
	.w3(32'h3996ab3f),
	.w4(32'hb8da83df),
	.w5(32'hb95d0de7),
	.w6(32'h3943980c),
	.w7(32'hb98b5121),
	.w8(32'hba7c0004),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0c1fd),
	.w1(32'hba867ea3),
	.w2(32'h3a5f1fd9),
	.w3(32'hb9cc923e),
	.w4(32'hba79990a),
	.w5(32'h3a68294d),
	.w6(32'hbaa4e285),
	.w7(32'hbafd39f8),
	.w8(32'h398762ad),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f41b8),
	.w1(32'h3a37685d),
	.w2(32'h3a8de145),
	.w3(32'h3a805f77),
	.w4(32'h39a12ba5),
	.w5(32'hba2c5865),
	.w6(32'h3a8538e1),
	.w7(32'h39567482),
	.w8(32'hb93a6d92),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc0598),
	.w1(32'hbb5a7759),
	.w2(32'hbb864c4c),
	.w3(32'hbb283e5e),
	.w4(32'hbb5c904e),
	.w5(32'hbb683559),
	.w6(32'hbb8cb779),
	.w7(32'hbb810c7d),
	.w8(32'hbb6aa454),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8de610),
	.w1(32'hbbc013a3),
	.w2(32'hbaf12335),
	.w3(32'hbbc8cfbd),
	.w4(32'hbb4f9ce1),
	.w5(32'hbb60e419),
	.w6(32'hbb90cd6f),
	.w7(32'hbb8e2cf3),
	.w8(32'hbb33ec71),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac982c9),
	.w1(32'h3a99a2b5),
	.w2(32'hba78f552),
	.w3(32'h3b258f68),
	.w4(32'h3b048790),
	.w5(32'hbace5b7c),
	.w6(32'h3b0b2af5),
	.w7(32'h3b04124d),
	.w8(32'hba4a2370),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6907dc),
	.w1(32'hba369d47),
	.w2(32'h399ee4c6),
	.w3(32'hbadf7e01),
	.w4(32'hbacadd0a),
	.w5(32'hb8a18a67),
	.w6(32'hba35a064),
	.w7(32'hba54aec6),
	.w8(32'h3a0a5e66),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e2831),
	.w1(32'h3a1d358a),
	.w2(32'h3a15fb23),
	.w3(32'h39cbc255),
	.w4(32'hba668192),
	.w5(32'h3a0a4dc9),
	.w6(32'h3a46e7c0),
	.w7(32'h39d3669e),
	.w8(32'h3a072590),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a84b2),
	.w1(32'h3a1a1ed6),
	.w2(32'hb9db59f8),
	.w3(32'h3a0c922a),
	.w4(32'h3a03336b),
	.w5(32'hba33e88c),
	.w6(32'h3a27b31d),
	.w7(32'h3a14f3f3),
	.w8(32'hba500b2f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e3213),
	.w1(32'hbaefabc8),
	.w2(32'hbaf969fe),
	.w3(32'hbb2d74cd),
	.w4(32'hbb3c210d),
	.w5(32'hbafafe0a),
	.w6(32'hbb6d26be),
	.w7(32'hbb5d012c),
	.w8(32'hbb5b6570),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41aba9),
	.w1(32'hb9f98c09),
	.w2(32'h3af06e06),
	.w3(32'hb94f9ccd),
	.w4(32'h3ac17f5d),
	.w5(32'h3ad542c4),
	.w6(32'hbb2e4d3b),
	.w7(32'hb97549ec),
	.w8(32'h3af6ed04),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2b0f0),
	.w1(32'hbb722187),
	.w2(32'hbbae329f),
	.w3(32'hbb5923b6),
	.w4(32'hb9d6194f),
	.w5(32'hbbf386e1),
	.w6(32'hbb9f3cd1),
	.w7(32'hbb3bf5a5),
	.w8(32'hbba24b39),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b05b1),
	.w1(32'h3bcafa8d),
	.w2(32'h3c0b256f),
	.w3(32'h3b85496d),
	.w4(32'h3c01f17b),
	.w5(32'h3b8139ae),
	.w6(32'h3b2e324f),
	.w7(32'h3b83bff0),
	.w8(32'h3bebf9ea),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc169b),
	.w1(32'h39185999),
	.w2(32'h3a324e74),
	.w3(32'hbadcc856),
	.w4(32'hba3c507b),
	.w5(32'h3978a5fc),
	.w6(32'hbb082b10),
	.w7(32'hba86cdbe),
	.w8(32'h39eea4d9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c726a4),
	.w1(32'h39549521),
	.w2(32'hb9b44e35),
	.w3(32'h39c8405d),
	.w4(32'h399fa07b),
	.w5(32'hba7c92e0),
	.w6(32'h39ef341b),
	.w7(32'h39eb7d78),
	.w8(32'hb98f184f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55078f),
	.w1(32'hb944d5af),
	.w2(32'hba634576),
	.w3(32'hbb033c51),
	.w4(32'hba670a02),
	.w5(32'hba5d6949),
	.w6(32'hbaa1b46c),
	.w7(32'hba2edc9b),
	.w8(32'hba80aeca),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa19ee5),
	.w1(32'hbb148ec5),
	.w2(32'hbb0a0701),
	.w3(32'hbb076bd5),
	.w4(32'hbb78f713),
	.w5(32'hbb0deb77),
	.w6(32'hbb2cbcb3),
	.w7(32'hbb31018a),
	.w8(32'hbaf5f938),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba409dd9),
	.w1(32'hba860993),
	.w2(32'h3964a526),
	.w3(32'hba3336e6),
	.w4(32'hba8fa111),
	.w5(32'hb9dd13fa),
	.w6(32'hba5b0c00),
	.w7(32'hba9423b7),
	.w8(32'hb9f65e98),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba104855),
	.w1(32'hbbc0f449),
	.w2(32'hbb614f95),
	.w3(32'hbb80fa55),
	.w4(32'hbc0e2569),
	.w5(32'hbb14eeca),
	.w6(32'hbbfa8278),
	.w7(32'hbbba120b),
	.w8(32'hbb092e9c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b4ab4),
	.w1(32'hbba5ac6e),
	.w2(32'hbbd8e251),
	.w3(32'hbb52eb33),
	.w4(32'hbc3ab213),
	.w5(32'hbb9cf2eb),
	.w6(32'hbc2ad929),
	.w7(32'hbc08ed99),
	.w8(32'hbb9de118),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba884968),
	.w1(32'h3b3fa052),
	.w2(32'h3a9901e1),
	.w3(32'h3aacc8fe),
	.w4(32'h3b018a71),
	.w5(32'hbab0f195),
	.w6(32'h3b25b238),
	.w7(32'h3afd4db7),
	.w8(32'h3a8cb367),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42079e),
	.w1(32'h38f978d1),
	.w2(32'hba6e4dc6),
	.w3(32'hbae6688d),
	.w4(32'hba391e6a),
	.w5(32'hba7058ff),
	.w6(32'hbb0652bd),
	.w7(32'hba617f7d),
	.w8(32'h3896f7e6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a5281),
	.w1(32'hba91b9d5),
	.w2(32'hba839164),
	.w3(32'hb9dbbd47),
	.w4(32'h39b76abf),
	.w5(32'hba02797f),
	.w6(32'hbad892ca),
	.w7(32'h39193dcb),
	.w8(32'hb9b3f4d5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f90e),
	.w1(32'hb93cf345),
	.w2(32'hba1682b9),
	.w3(32'hb9b264cf),
	.w4(32'h3aad382f),
	.w5(32'hba8f571c),
	.w6(32'hb9dd526c),
	.w7(32'h39e99723),
	.w8(32'hb957e902),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d9dbf),
	.w1(32'hbbaa38b4),
	.w2(32'hbb99ec6b),
	.w3(32'hbbb16a65),
	.w4(32'hbbbb5c34),
	.w5(32'hbb7fae94),
	.w6(32'hbba69119),
	.w7(32'hbb80de04),
	.w8(32'hbb164625),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb5cd0),
	.w1(32'hba513df5),
	.w2(32'hba9c3e30),
	.w3(32'hba99240b),
	.w4(32'hba5d3ea3),
	.w5(32'hbab0024b),
	.w6(32'hba23010f),
	.w7(32'hbaa1857c),
	.w8(32'hb9d302a5),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa231c),
	.w1(32'hbae3ade0),
	.w2(32'hba3a8c4e),
	.w3(32'hbab653eb),
	.w4(32'hbb008991),
	.w5(32'hba7b45db),
	.w6(32'hbaa5a47f),
	.w7(32'hba64bfa6),
	.w8(32'hba53a50f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba948969),
	.w1(32'h39a3d3c6),
	.w2(32'h39eabbd8),
	.w3(32'hbacfd982),
	.w4(32'hba1425b7),
	.w5(32'h39018fec),
	.w6(32'hba1dbaf8),
	.w7(32'hb907ec60),
	.w8(32'h396dfaa0),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c1b02e),
	.w1(32'hb9be2b35),
	.w2(32'h3a26ff5a),
	.w3(32'hba0daef0),
	.w4(32'hb940142d),
	.w5(32'h3a1d7307),
	.w6(32'hba1bb175),
	.w7(32'hb806d5bf),
	.w8(32'h39edc24c),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0da9cf),
	.w1(32'h3b41fb13),
	.w2(32'h3b2cb080),
	.w3(32'h3b1ae5f2),
	.w4(32'h3b5f3f2a),
	.w5(32'h3ad31559),
	.w6(32'h3a85ddf8),
	.w7(32'h3aad7d9f),
	.w8(32'h3b073f10),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d11bd),
	.w1(32'hba848adc),
	.w2(32'h3a271fdd),
	.w3(32'hba403389),
	.w4(32'hb9f732d7),
	.w5(32'h39f96bd0),
	.w6(32'hba63e08e),
	.w7(32'hba2ebab5),
	.w8(32'hb6d8d8e9),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6981b5),
	.w1(32'h3a5f6793),
	.w2(32'h3a2a5426),
	.w3(32'h3a814911),
	.w4(32'h3a2f66a1),
	.w5(32'hb9844ec6),
	.w6(32'hbaaf954b),
	.w7(32'h3afc7117),
	.w8(32'h388362ac),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2269f),
	.w1(32'hbc44e6c5),
	.w2(32'hbbfe0a72),
	.w3(32'hbc32c4fa),
	.w4(32'hbc4004d1),
	.w5(32'hbbcd1387),
	.w6(32'hbc80cf54),
	.w7(32'hbc4dec34),
	.w8(32'hbbed2ca6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a96fb),
	.w1(32'h3ae0f785),
	.w2(32'h3b28f807),
	.w3(32'h3b05a087),
	.w4(32'h39e3f5ad),
	.w5(32'h3b25bba3),
	.w6(32'h3af3dcc2),
	.w7(32'h3ab68ae5),
	.w8(32'h3b5d08a8),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a5870),
	.w1(32'h3aa5a9ba),
	.w2(32'h3ad85b5e),
	.w3(32'h3a01c130),
	.w4(32'h3a0c1cca),
	.w5(32'h374d4ab0),
	.w6(32'h38075475),
	.w7(32'h39e1da91),
	.w8(32'hbb11221e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38480e),
	.w1(32'hb9a47437),
	.w2(32'h3a955876),
	.w3(32'hbabb8051),
	.w4(32'hb9ebeb14),
	.w5(32'h39cdf489),
	.w6(32'hba47155b),
	.w7(32'hb9e857b4),
	.w8(32'h39bcd5a5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3f0840),
	.w1(32'h38ffd8d4),
	.w2(32'h3a27f66a),
	.w3(32'hba60207f),
	.w4(32'h39bc887f),
	.w5(32'h3a5ebb54),
	.w6(32'hbad843cf),
	.w7(32'hba571749),
	.w8(32'h3a04f612),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8c7df),
	.w1(32'h3b1af360),
	.w2(32'h39097316),
	.w3(32'h3b4d892d),
	.w4(32'h3b8df669),
	.w5(32'h39fbdf68),
	.w6(32'h3b1d054b),
	.w7(32'h3b671867),
	.w8(32'hbad3114c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d3e7e),
	.w1(32'h3b3378f5),
	.w2(32'h3aecd2a5),
	.w3(32'h3a9eb3e7),
	.w4(32'h3ae53f8d),
	.w5(32'h3a6466d9),
	.w6(32'h3b09fc4f),
	.w7(32'h3a8f67bf),
	.w8(32'h3b2e4394),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96db99),
	.w1(32'hba97895d),
	.w2(32'h3a978280),
	.w3(32'hbb10dca8),
	.w4(32'hbb118e72),
	.w5(32'h3a9e4f12),
	.w6(32'hbac0a1ba),
	.w7(32'hbaa2c342),
	.w8(32'h3a63eaa2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3d754),
	.w1(32'h3a917770),
	.w2(32'hbaf0a6cd),
	.w3(32'h39c7360d),
	.w4(32'h3a9fe8a2),
	.w5(32'hbb0a230e),
	.w6(32'hbaa48f0b),
	.w7(32'hb9d19a9d),
	.w8(32'hbb03e559),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07626b),
	.w1(32'hbb2f0673),
	.w2(32'hbaf66110),
	.w3(32'hba965fbc),
	.w4(32'h3a0ed8d1),
	.w5(32'hb9ef2ecc),
	.w6(32'hba148278),
	.w7(32'h38f7a0bd),
	.w8(32'hba69d871),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9084ce),
	.w1(32'hbc3fccd6),
	.w2(32'hbbfe317e),
	.w3(32'hbc2544ff),
	.w4(32'hbc62e3ce),
	.w5(32'hbc011ee8),
	.w6(32'hbc62467b),
	.w7(32'hbc485f80),
	.w8(32'hbc084c45),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc47968),
	.w1(32'h3c3829ca),
	.w2(32'h3c16b57c),
	.w3(32'h3c2a98c8),
	.w4(32'h3c243ca3),
	.w5(32'h3bd1b73a),
	.w6(32'h3c15e249),
	.w7(32'h3bfa864e),
	.w8(32'h3b7619d0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26ae3e),
	.w1(32'h3b66a046),
	.w2(32'h3b826813),
	.w3(32'h3b98826d),
	.w4(32'h3b443468),
	.w5(32'h3a0992ee),
	.w6(32'h3b25654c),
	.w7(32'h3b04d075),
	.w8(32'h3b8cfe05),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f869c),
	.w1(32'hbb1e360f),
	.w2(32'hbad1c034),
	.w3(32'hb9c6fc55),
	.w4(32'hb7fad609),
	.w5(32'h392abc73),
	.w6(32'hbb02cb8b),
	.w7(32'hb87472e0),
	.w8(32'hbb0de70e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985d6ff),
	.w1(32'h3a701bc5),
	.w2(32'hbabb67b4),
	.w3(32'h38e998d3),
	.w4(32'h3970e43f),
	.w5(32'hbb2b9e19),
	.w6(32'hba2360b0),
	.w7(32'hb86ecf95),
	.w8(32'hbb367816),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f51f8),
	.w1(32'hbc549d4b),
	.w2(32'hbc569880),
	.w3(32'hbbbc55dd),
	.w4(32'hbc63afe8),
	.w5(32'hbbdee7a6),
	.w6(32'hbc63433a),
	.w7(32'hbc3b8ef5),
	.w8(32'hbbdcc398),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a843d8d),
	.w1(32'h3a8b963c),
	.w2(32'hba49a104),
	.w3(32'h3b08ba55),
	.w4(32'h3a83ca6d),
	.w5(32'hbaa039e2),
	.w6(32'h3b1bdfd8),
	.w7(32'h3a6cb654),
	.w8(32'hb9ed8bfd),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5afd18),
	.w1(32'hb9b53983),
	.w2(32'h39edf77f),
	.w3(32'hbaa1dd2e),
	.w4(32'hba0302e1),
	.w5(32'hb90582f2),
	.w6(32'hbaadfb13),
	.w7(32'hb9f1dfc4),
	.w8(32'h3941d6b3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdfdda),
	.w1(32'h3a360b9f),
	.w2(32'hb9fda33f),
	.w3(32'hba980023),
	.w4(32'h3972466e),
	.w5(32'hbaacef76),
	.w6(32'hb9e59a9f),
	.w7(32'h3a16820c),
	.w8(32'hb981613a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb912dff),
	.w1(32'hb9e19eef),
	.w2(32'h3a3677ac),
	.w3(32'hbb05687c),
	.w4(32'h39c1de5a),
	.w5(32'hba0862ae),
	.w6(32'hbb405a6c),
	.w7(32'hbb04b583),
	.w8(32'h3a981642),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4169b),
	.w1(32'h3b162be1),
	.w2(32'h3b44140b),
	.w3(32'h3b288bfd),
	.w4(32'h3b2c9ecc),
	.w5(32'h3b35bf21),
	.w6(32'h3b40e656),
	.w7(32'h3b23affe),
	.w8(32'h3b94d1e8),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2d073),
	.w1(32'h3b2663f3),
	.w2(32'hbb4897e3),
	.w3(32'h3af0a8b9),
	.w4(32'h3a8e5640),
	.w5(32'hba792bcd),
	.w6(32'h3b3977d1),
	.w7(32'hba62c5dc),
	.w8(32'hbb5f51f7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10f36d),
	.w1(32'h3a08ea41),
	.w2(32'h3a92dab8),
	.w3(32'hb91f904d),
	.w4(32'h3abf8c45),
	.w5(32'h3aac0b30),
	.w6(32'hb95a79dc),
	.w7(32'hb9ecf322),
	.w8(32'h3a4ffc89),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e658a),
	.w1(32'hba363e9d),
	.w2(32'hbadebf23),
	.w3(32'hba81a508),
	.w4(32'hbabec40c),
	.w5(32'hbae04ce7),
	.w6(32'hbb1175bc),
	.w7(32'hba928711),
	.w8(32'hba5d2371),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a4e12),
	.w1(32'hbb20a1f9),
	.w2(32'hbaff2f67),
	.w3(32'hbacdea34),
	.w4(32'hbac7a9f2),
	.w5(32'hbabeb847),
	.w6(32'hba2ed8ec),
	.w7(32'hba78ba35),
	.w8(32'hbaf63ad2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb133630),
	.w1(32'hb913a015),
	.w2(32'h3a22bafa),
	.w3(32'h3b05ccd5),
	.w4(32'h3af18388),
	.w5(32'hb929f6b7),
	.w6(32'h3a89d362),
	.w7(32'h3a24f885),
	.w8(32'h3a1535af),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a292b72),
	.w1(32'h39cbd6b3),
	.w2(32'h3af13950),
	.w3(32'h39b7b38f),
	.w4(32'h38d6ad1d),
	.w5(32'h3a731861),
	.w6(32'h3a11ac95),
	.w7(32'h392ac1a9),
	.w8(32'h3adc287c),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e2bbf),
	.w1(32'h3a389c7c),
	.w2(32'h397a718b),
	.w3(32'h39922a84),
	.w4(32'h394f4576),
	.w5(32'h3963f5c0),
	.w6(32'h3abc5a2d),
	.w7(32'h3a9c71f9),
	.w8(32'h39b4475c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0a7658),
	.w1(32'h39fc7611),
	.w2(32'h398a275f),
	.w3(32'h39ab5edc),
	.w4(32'h39526a98),
	.w5(32'hb9940c4b),
	.w6(32'h3a5b0829),
	.w7(32'h3a33de2c),
	.w8(32'h3a514fef),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace566c),
	.w1(32'h3a83bbe4),
	.w2(32'hba82a4f1),
	.w3(32'h3a94f9ce),
	.w4(32'hb9905eb9),
	.w5(32'hbac557c2),
	.w6(32'h3ac959b3),
	.w7(32'h3a82cb3d),
	.w8(32'hba4db92f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada6318),
	.w1(32'h3aa710cc),
	.w2(32'h3b52a550),
	.w3(32'h3ac0be6f),
	.w4(32'h3ac93195),
	.w5(32'h3a59e0c0),
	.w6(32'h3aad61ee),
	.w7(32'h3a12eab0),
	.w8(32'h3b3fea38),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b4a6),
	.w1(32'h3ad6d6ea),
	.w2(32'h3a768b4c),
	.w3(32'h3b2b710d),
	.w4(32'h3aef2c98),
	.w5(32'h3a302627),
	.w6(32'h3b12954b),
	.w7(32'h3aa06f43),
	.w8(32'h39ace29b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f8b763),
	.w1(32'hbaf2e145),
	.w2(32'hbade79f3),
	.w3(32'h3a94137a),
	.w4(32'hba9bdcd8),
	.w5(32'hbabafc02),
	.w6(32'hbb17853f),
	.w7(32'hbafd97ce),
	.w8(32'hbacf1c00),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb851e5a0),
	.w1(32'h3babeda7),
	.w2(32'h3b92ebd0),
	.w3(32'h3ad957c3),
	.w4(32'h3b39f54f),
	.w5(32'h3b20dd73),
	.w6(32'h3b7a4ada),
	.w7(32'h3b6dd630),
	.w8(32'h3b7d5a8c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9a9e0),
	.w1(32'h3a87abdf),
	.w2(32'h3a1b2722),
	.w3(32'h3a8b7c17),
	.w4(32'h39c7e9b6),
	.w5(32'h39c7e375),
	.w6(32'h3971e587),
	.w7(32'hb83120f9),
	.w8(32'h3a1ffecc),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ddab43),
	.w1(32'h3a6396d2),
	.w2(32'h3a23689e),
	.w3(32'h3855a910),
	.w4(32'h3a309093),
	.w5(32'hb89bc4fd),
	.w6(32'h39a4d701),
	.w7(32'h3a5f671e),
	.w8(32'hb967e96e),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81d3f4c),
	.w1(32'hb986bc15),
	.w2(32'h39700796),
	.w3(32'hba2ba0db),
	.w4(32'hba50389a),
	.w5(32'hb9ca15db),
	.w6(32'hbac34876),
	.w7(32'hba8be130),
	.w8(32'hb99cf4e9),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41751d),
	.w1(32'h3ab87d9b),
	.w2(32'h39f0427b),
	.w3(32'hba293b8a),
	.w4(32'h3a562418),
	.w5(32'hbac94b53),
	.w6(32'hbab4fdf0),
	.w7(32'h39f0f7af),
	.w8(32'hba6f9e08),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a63c6),
	.w1(32'hbb786862),
	.w2(32'hbaeb2568),
	.w3(32'hbb66dbe5),
	.w4(32'hbb2f4657),
	.w5(32'hbb8d25f1),
	.w6(32'hbb7866b5),
	.w7(32'hbb101f28),
	.w8(32'hbb622e07),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b0a4a),
	.w1(32'h38ebee3a),
	.w2(32'hb9140895),
	.w3(32'hb93ac08f),
	.w4(32'hb973ae0a),
	.w5(32'hb978e26b),
	.w6(32'hbb0af61e),
	.w7(32'hba9c5695),
	.w8(32'hba9d2eca),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376eb1d3),
	.w1(32'hbaf321c5),
	.w2(32'hbab0fcc8),
	.w3(32'hba00e3ce),
	.w4(32'hbaa2ec67),
	.w5(32'hba6b2c1d),
	.w6(32'hba3d5e82),
	.w7(32'hba031759),
	.w8(32'hb8f5d7c2),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0643ee),
	.w1(32'hbaf550d0),
	.w2(32'h39e3f909),
	.w3(32'hb7af02a3),
	.w4(32'hba84838a),
	.w5(32'h3a35231b),
	.w6(32'hbaa654bd),
	.w7(32'hba87c547),
	.w8(32'h3a4e43c2),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f5b4),
	.w1(32'h3ae1357e),
	.w2(32'h3ac42088),
	.w3(32'h3ab42f62),
	.w4(32'h3acc7052),
	.w5(32'h3a997fb6),
	.w6(32'h3ab326da),
	.w7(32'h3b3d3ddf),
	.w8(32'h3acc855f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43d974),
	.w1(32'hb8b45705),
	.w2(32'hb96a5f68),
	.w3(32'h3913e03a),
	.w4(32'h3a9529dc),
	.w5(32'hba40ec5e),
	.w6(32'h3a4ed51c),
	.w7(32'h39cd3526),
	.w8(32'hba80b790),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a351e60),
	.w1(32'h3b022bc8),
	.w2(32'h3b411548),
	.w3(32'h3a96930d),
	.w4(32'h3b399195),
	.w5(32'h3b02fc19),
	.w6(32'h3a9416d6),
	.w7(32'h3abe649a),
	.w8(32'h3b03b52e),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb047be5),
	.w1(32'hbbcb7e81),
	.w2(32'hbba9d46a),
	.w3(32'hbbfcc87c),
	.w4(32'hbbf15942),
	.w5(32'hbbca6026),
	.w6(32'hbc0a781c),
	.w7(32'hbbc6cace),
	.w8(32'hbbc0ee23),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1320e),
	.w1(32'h3b35e51e),
	.w2(32'h3ae2a123),
	.w3(32'h3b3d1061),
	.w4(32'h3b4aee28),
	.w5(32'h3ac22c9d),
	.w6(32'h3b3da134),
	.w7(32'h3b382a36),
	.w8(32'h3b7fcde0),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba840bfa),
	.w1(32'h399a9b7a),
	.w2(32'h3af0269c),
	.w3(32'h3a2385e7),
	.w4(32'h3a9624f8),
	.w5(32'h3aa620ff),
	.w6(32'h3ac45354),
	.w7(32'h3ad6d202),
	.w8(32'h3ab0b3df),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03ad18),
	.w1(32'hba1dd627),
	.w2(32'hbb216018),
	.w3(32'hbb5e4b3a),
	.w4(32'hba6da59f),
	.w5(32'hbb44a1ec),
	.w6(32'hbb7a4c0a),
	.w7(32'hbabf5a36),
	.w8(32'hbb621664),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83a1dab),
	.w1(32'h3b22387d),
	.w2(32'h3aff26f5),
	.w3(32'h3a0718cb),
	.w4(32'h3ae57c79),
	.w5(32'h3abd6719),
	.w6(32'hbab12493),
	.w7(32'h3a0e27d7),
	.w8(32'h3b10cda5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5285e9),
	.w1(32'h39ecc3ac),
	.w2(32'hb9f75ea3),
	.w3(32'h3ad5a6f6),
	.w4(32'h3a71bd21),
	.w5(32'hbacc2cad),
	.w6(32'h385c073b),
	.w7(32'hb928d9eb),
	.w8(32'hbada5cc1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a283f),
	.w1(32'hb8d01047),
	.w2(32'h3a398a12),
	.w3(32'hba03c40e),
	.w4(32'hb97a9763),
	.w5(32'hb9ef2a47),
	.w6(32'hba62a4f1),
	.w7(32'hba28ec21),
	.w8(32'h38594098),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba321d91),
	.w1(32'h3baeaf7c),
	.w2(32'h3b45ae98),
	.w3(32'h3b82c544),
	.w4(32'h3bd466d6),
	.w5(32'h3b3562f9),
	.w6(32'h3baefa0c),
	.w7(32'h3b831938),
	.w8(32'h3badc5d8),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1dd644),
	.w1(32'hbac2b854),
	.w2(32'hb99d1e09),
	.w3(32'hba9eba6c),
	.w4(32'hbad6ef7a),
	.w5(32'hba87a6a3),
	.w6(32'hba29bf81),
	.w7(32'hbac322a4),
	.w8(32'hba9afdc0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58f91e),
	.w1(32'h3a850331),
	.w2(32'hb9863b5e),
	.w3(32'h3a399c08),
	.w4(32'h3a6e21f4),
	.w5(32'hba1bb1f3),
	.w6(32'h3a44f121),
	.w7(32'h3a67e747),
	.w8(32'hba02cb02),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c88e),
	.w1(32'hb9809933),
	.w2(32'h39ee4279),
	.w3(32'hba4c32a2),
	.w4(32'hb9dc075d),
	.w5(32'h39bc3445),
	.w6(32'hba483e59),
	.w7(32'hb9f5628c),
	.w8(32'hb9a279b5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915b279),
	.w1(32'h3a90dcbb),
	.w2(32'h39b54047),
	.w3(32'h39b7254a),
	.w4(32'h390b4b12),
	.w5(32'h395137ea),
	.w6(32'hb9fa1120),
	.w7(32'h399fa9e4),
	.w8(32'h3a4ca697),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5180cc),
	.w1(32'h3b9d7544),
	.w2(32'hba2cb716),
	.w3(32'h3b7d4c17),
	.w4(32'h3b736b55),
	.w5(32'h3a977805),
	.w6(32'h3b0fd415),
	.w7(32'h3b13f767),
	.w8(32'h3b125c1b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbd3af),
	.w1(32'hbb0206b5),
	.w2(32'h3a119772),
	.w3(32'hbb845561),
	.w4(32'hbaf949ca),
	.w5(32'hb9deaf80),
	.w6(32'hbb1a45fc),
	.w7(32'hbabc4b7c),
	.w8(32'h39d55a39),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57bb0c),
	.w1(32'h3a2dfea4),
	.w2(32'h3a497b92),
	.w3(32'h39f977ad),
	.w4(32'h3a2ca2ac),
	.w5(32'h3a167c57),
	.w6(32'h39cfbebe),
	.w7(32'h3a0d2884),
	.w8(32'h3a721a76),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba103d99),
	.w1(32'h3af93406),
	.w2(32'hba2cef95),
	.w3(32'h3acae709),
	.w4(32'h3b834a6d),
	.w5(32'hbaedd70a),
	.w6(32'hba67abff),
	.w7(32'h3af1c1b4),
	.w8(32'hba6d10e2),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14fe49),
	.w1(32'hb96d4ee4),
	.w2(32'h3b33a2b8),
	.w3(32'hba55de54),
	.w4(32'hb98e607c),
	.w5(32'h3aa2cf3b),
	.w6(32'hba48ed84),
	.w7(32'hba243942),
	.w8(32'h3b373ce8),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad06963),
	.w1(32'hbb152cd2),
	.w2(32'hbb91027b),
	.w3(32'hba939cf7),
	.w4(32'hbae99a1b),
	.w5(32'hbb75848f),
	.w6(32'hbae9b9e6),
	.w7(32'hbabaace5),
	.w8(32'hbb44e417),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bc09f),
	.w1(32'h3ab4821d),
	.w2(32'h3b08d370),
	.w3(32'h387c0ab5),
	.w4(32'h3b4fe838),
	.w5(32'h38f4c119),
	.w6(32'h3a5e4d3d),
	.w7(32'h3b18c21f),
	.w8(32'h3aceb3b3),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae528ef),
	.w1(32'h3b0bd717),
	.w2(32'h3b374b82),
	.w3(32'h3acbc8e8),
	.w4(32'h3ad7f35d),
	.w5(32'h3b0d9394),
	.w6(32'h3ae1108b),
	.w7(32'h3b13697a),
	.w8(32'h3b05c46d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b6618),
	.w1(32'h3a909c7d),
	.w2(32'h3a35c635),
	.w3(32'h3a8cbc09),
	.w4(32'h398e3db3),
	.w5(32'hba459897),
	.w6(32'h3a888d2d),
	.w7(32'h385839c5),
	.w8(32'hba407868),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d7607),
	.w1(32'h3aeeba47),
	.w2(32'h3b57d6a7),
	.w3(32'h3acc3af0),
	.w4(32'h3b88f83d),
	.w5(32'h3b77ddeb),
	.w6(32'h3b0f5332),
	.w7(32'h3b837c3d),
	.w8(32'hbb020934),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4185a),
	.w1(32'h3bb6f992),
	.w2(32'h3c0a74ea),
	.w3(32'h3b29f424),
	.w4(32'h3be5b266),
	.w5(32'h3ad7315c),
	.w6(32'hbba8d6b9),
	.w7(32'h3bb57dec),
	.w8(32'hbc6141c7),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b07f3),
	.w1(32'h3c03b72c),
	.w2(32'hbabed830),
	.w3(32'h3c23f702),
	.w4(32'h3c680709),
	.w5(32'h38a81a81),
	.w6(32'hbd08df8b),
	.w7(32'hbc9c39d0),
	.w8(32'hbb7aeac6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b20a6),
	.w1(32'hbbc422b8),
	.w2(32'hbc1a1925),
	.w3(32'h3a0be067),
	.w4(32'hbb380980),
	.w5(32'hbba26fb1),
	.w6(32'hbaeca802),
	.w7(32'hbb11f122),
	.w8(32'hbc16c771),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e60c9d),
	.w1(32'hbb5e8ba3),
	.w2(32'h3aead835),
	.w3(32'h3bc0b452),
	.w4(32'h3b49120c),
	.w5(32'hbaecfe15),
	.w6(32'hbbb5a300),
	.w7(32'hbb2c4442),
	.w8(32'hbb950673),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab552be),
	.w1(32'hbb0f86eb),
	.w2(32'h3953f9ea),
	.w3(32'h3b1c7410),
	.w4(32'h3a66e998),
	.w5(32'hbb0505de),
	.w6(32'hbc3bd443),
	.w7(32'hbc135f64),
	.w8(32'hbb9a95ff),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b182846),
	.w1(32'h3a59c78b),
	.w2(32'hba98252b),
	.w3(32'h3a3bd147),
	.w4(32'hb9a2a86c),
	.w5(32'hbbb47bd0),
	.w6(32'hb94edd94),
	.w7(32'h3aeda6c0),
	.w8(32'h3b8963d2),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6b49a),
	.w1(32'hbc3ef087),
	.w2(32'hbac64686),
	.w3(32'hbb9a7e9f),
	.w4(32'hbc5f5c22),
	.w5(32'hb83dc1e2),
	.w6(32'h3cc57ad9),
	.w7(32'h3c92b925),
	.w8(32'hb7e5abd5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf369e2),
	.w1(32'hba816dfe),
	.w2(32'h3c85e113),
	.w3(32'hbb06462e),
	.w4(32'hbaffc4c3),
	.w5(32'hbccb741d),
	.w6(32'hbb5459bd),
	.w7(32'hbad4044c),
	.w8(32'hbbf6874d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3095a0),
	.w1(32'h3ccf0499),
	.w2(32'hb9801458),
	.w3(32'hbb935272),
	.w4(32'h3c848547),
	.w5(32'h3b9b7aff),
	.w6(32'hbce1ae69),
	.w7(32'hbccb2761),
	.w8(32'hbad43336),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993e2dd),
	.w1(32'hbb08109f),
	.w2(32'hbc2d1b3d),
	.w3(32'h3b0c52c6),
	.w4(32'hbaf6b294),
	.w5(32'h3b0bdec2),
	.w6(32'hbaac29c2),
	.w7(32'hb99f9eca),
	.w8(32'h3ba89adb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bd3a0),
	.w1(32'hbc21d328),
	.w2(32'hbb9ed324),
	.w3(32'hbc141842),
	.w4(32'hbc92b558),
	.w5(32'h3c07794c),
	.w6(32'h3c9ce41e),
	.w7(32'h3c93a3ea),
	.w8(32'h3bfdfde4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb739c58),
	.w1(32'h3b40971e),
	.w2(32'hba0f3a9b),
	.w3(32'h3c0a3bbb),
	.w4(32'h3b677fba),
	.w5(32'hba617f7f),
	.w6(32'h3bc8ccfc),
	.w7(32'h3bb76f21),
	.w8(32'hbb840f0d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0feca),
	.w1(32'hbbdb8456),
	.w2(32'hbbe85354),
	.w3(32'h3af3c99a),
	.w4(32'hbb581aff),
	.w5(32'hbb6f82a8),
	.w6(32'hbc00a0c6),
	.w7(32'hbbd8f72d),
	.w8(32'h3b30fc03),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc989315),
	.w1(32'hbbdcaa68),
	.w2(32'hbb76b3b9),
	.w3(32'hbc379596),
	.w4(32'hbc4942d4),
	.w5(32'hbc09a43f),
	.w6(32'hbaf07ae1),
	.w7(32'hbbf3060a),
	.w8(32'hbbfb8e61),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca40a),
	.w1(32'hbc4468ea),
	.w2(32'h3aebcaf1),
	.w3(32'hbb0ce242),
	.w4(32'hbb9551d4),
	.w5(32'h3ab3329e),
	.w6(32'h3ba7df13),
	.w7(32'h3c23aa76),
	.w8(32'h3b5c6be7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387c6ce5),
	.w1(32'h3b38d2fc),
	.w2(32'hbb48414e),
	.w3(32'hbaeef337),
	.w4(32'h3a1debbf),
	.w5(32'h3cf4af5b),
	.w6(32'h3b19a06a),
	.w7(32'h3b474361),
	.w8(32'h3a64b76d),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccaea26),
	.w1(32'hbbbad33d),
	.w2(32'h3bd7d9c0),
	.w3(32'h3c793b5d),
	.w4(32'hbb9e7bd2),
	.w5(32'h3c9ed42b),
	.w6(32'h3995adfe),
	.w7(32'h3c28c52d),
	.w8(32'h3c4a8d21),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5498c3),
	.w1(32'hbc2a47d5),
	.w2(32'h3bb95d7e),
	.w3(32'h3c32cbaf),
	.w4(32'hbc73cc0a),
	.w5(32'h3be4cfe0),
	.w6(32'h3c9a5dfd),
	.w7(32'h3c6fdf65),
	.w8(32'hbc953b8c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c951948),
	.w1(32'hbae94310),
	.w2(32'hbc38fcae),
	.w3(32'h3ca2939d),
	.w4(32'h3cb418a4),
	.w5(32'hbc148d75),
	.w6(32'hbd049895),
	.w7(32'hbcb32af7),
	.w8(32'hbb433b6e),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde3a48),
	.w1(32'h3ba93436),
	.w2(32'h3a9206b6),
	.w3(32'hbc1484ec),
	.w4(32'h3c03ae8d),
	.w5(32'h3adbb995),
	.w6(32'hbb1edca8),
	.w7(32'h3a4ba352),
	.w8(32'h3b831fa8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d25a6),
	.w1(32'hb81750d4),
	.w2(32'h3bfba054),
	.w3(32'h3a32f0cf),
	.w4(32'h392d7688),
	.w5(32'h3b7c17ca),
	.w6(32'h3b839a9a),
	.w7(32'h3a8285fe),
	.w8(32'h3c69cc5b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b16d5),
	.w1(32'hbba9033c),
	.w2(32'hbbeef5f8),
	.w3(32'hbc01f495),
	.w4(32'hbbb97390),
	.w5(32'hbb8d3dc4),
	.w6(32'h3b9199f9),
	.w7(32'h3bd091b1),
	.w8(32'h3c947749),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf2fa94),
	.w1(32'hbcef35c6),
	.w2(32'h3a6ab64b),
	.w3(32'hbc8d0855),
	.w4(32'hbcfb4da5),
	.w5(32'hbb334516),
	.w6(32'h3cf0b66d),
	.w7(32'h3c63d66f),
	.w8(32'h3b0d3661),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f2af5),
	.w1(32'hbbea83a8),
	.w2(32'hbbe6ad62),
	.w3(32'hbbe22948),
	.w4(32'hbc5bff23),
	.w5(32'h3b26c3bd),
	.w6(32'h3c16f528),
	.w7(32'hbac095dd),
	.w8(32'h3cda94ae),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfdb5f1),
	.w1(32'hbc76a269),
	.w2(32'hbb195863),
	.w3(32'hbc8a3780),
	.w4(32'hbcdfdde9),
	.w5(32'hbb55f87d),
	.w6(32'h3cd5143e),
	.w7(32'h3beef892),
	.w8(32'hbb603aed),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c004e20),
	.w1(32'h3c61ea71),
	.w2(32'h39753606),
	.w3(32'hba31c0d9),
	.w4(32'h3b715715),
	.w5(32'hbca0f5ea),
	.w6(32'h3af0fba2),
	.w7(32'h39d2e595),
	.w8(32'hba50782b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70ecd7),
	.w1(32'h3c4bafc4),
	.w2(32'h3c7b0c5a),
	.w3(32'hbcbfd6a1),
	.w4(32'hbc0c325c),
	.w5(32'h3c1b5390),
	.w6(32'hbc23cfc7),
	.w7(32'hbbfe0244),
	.w8(32'hbbcd28af),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cadb500),
	.w1(32'h3c62b703),
	.w2(32'hba7c763b),
	.w3(32'h3cbbfd15),
	.w4(32'h3cb10502),
	.w5(32'h3c3c233b),
	.w6(32'hbcaf32e1),
	.w7(32'hbc8114ed),
	.w8(32'hbc1852ae),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8f72b),
	.w1(32'hbb79ed91),
	.w2(32'h3a9a842b),
	.w3(32'h3c4d5b6d),
	.w4(32'h3b3e80ed),
	.w5(32'h3bd0cd32),
	.w6(32'hbc6e2829),
	.w7(32'hbc0e4040),
	.w8(32'h3b86f9f5),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc17baa),
	.w1(32'hbbc72876),
	.w2(32'h3aad5f66),
	.w3(32'h3b345933),
	.w4(32'hba42ce1a),
	.w5(32'hbab77aa0),
	.w6(32'h38f07440),
	.w7(32'h3afc96f8),
	.w8(32'h3b557235),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd00c),
	.w1(32'hbc193af5),
	.w2(32'h3b8b3a1e),
	.w3(32'hbc239a48),
	.w4(32'hbc0133a3),
	.w5(32'h3bafe731),
	.w6(32'h3ad83540),
	.w7(32'h3b007af1),
	.w8(32'hb8a6d324),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c6ae2),
	.w1(32'hb97621c0),
	.w2(32'hbc34ca34),
	.w3(32'hbb80faea),
	.w4(32'hbb3df25f),
	.w5(32'hbbec07eb),
	.w6(32'hbc00f7dc),
	.w7(32'hbabc79c0),
	.w8(32'hba9f9e65),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ff264),
	.w1(32'h389f11e0),
	.w2(32'h3c636ea9),
	.w3(32'h3ae83a6f),
	.w4(32'h3b96dcba),
	.w5(32'h3a772862),
	.w6(32'h3c173c7d),
	.w7(32'h3c028bd2),
	.w8(32'hbbc83700),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10f10e),
	.w1(32'h3be6e801),
	.w2(32'h3b99fa55),
	.w3(32'h3bf6affd),
	.w4(32'h3b6623b9),
	.w5(32'hba37e23a),
	.w6(32'hbcbb9cb8),
	.w7(32'hbc7f9645),
	.w8(32'hbb06d599),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b943f50),
	.w1(32'h3bc6fa2f),
	.w2(32'h3944dfaa),
	.w3(32'hbc4a3f0d),
	.w4(32'hbbf668d6),
	.w5(32'hbbb64e92),
	.w6(32'hbb9ab5a9),
	.w7(32'hbbf356f7),
	.w8(32'hbb1c3e6e),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba492eda),
	.w1(32'hbb0b3b9b),
	.w2(32'h3a8030e9),
	.w3(32'hbbb4b613),
	.w4(32'h3acdcac3),
	.w5(32'hbb6cd4dc),
	.w6(32'h3ac10757),
	.w7(32'h3b1aa569),
	.w8(32'hbb32ac36),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad4c3),
	.w1(32'h3c37c96c),
	.w2(32'h3a39050b),
	.w3(32'h3c16785f),
	.w4(32'h3c9dd0cd),
	.w5(32'h3b3cc526),
	.w6(32'hbb454ed0),
	.w7(32'hbb0f36ac),
	.w8(32'h3bb5cf3c),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dd7b8),
	.w1(32'hba5a369c),
	.w2(32'hbb3c74ef),
	.w3(32'hba847f4b),
	.w4(32'hbb6e3c18),
	.w5(32'hbbb5e6f4),
	.w6(32'h3b9b99ae),
	.w7(32'h38274f74),
	.w8(32'hbb8c1fd7),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a539abc),
	.w1(32'h3bc75814),
	.w2(32'hbc662954),
	.w3(32'h3b10e2b2),
	.w4(32'h3becfe67),
	.w5(32'h3be337ad),
	.w6(32'h3b15c300),
	.w7(32'h3c1bca83),
	.w8(32'h387b0d24),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdc1880),
	.w1(32'hbd115412),
	.w2(32'hbba913a4),
	.w3(32'h3c50e076),
	.w4(32'hbacfb797),
	.w5(32'hbaaa220e),
	.w6(32'h3cbac8c8),
	.w7(32'h3c430a61),
	.w8(32'h3c21d01d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc739e13),
	.w1(32'hbb1b9e80),
	.w2(32'h38af9386),
	.w3(32'hbccedca5),
	.w4(32'hbcbbe365),
	.w5(32'hbb2c6719),
	.w6(32'hbb11af2c),
	.w7(32'hb9d1d595),
	.w8(32'hba9354f0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e15f6),
	.w1(32'h3b09affc),
	.w2(32'h3b3dc083),
	.w3(32'hbb66a291),
	.w4(32'h3b1043be),
	.w5(32'h3aff0072),
	.w6(32'hbb3dc7c8),
	.w7(32'h3a1892b8),
	.w8(32'hba340412),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1604af),
	.w1(32'hbbcca92d),
	.w2(32'h3b922f61),
	.w3(32'hbac5b85e),
	.w4(32'hba6ac5ff),
	.w5(32'h3b7606e6),
	.w6(32'hbaed9818),
	.w7(32'h3abf0ddb),
	.w8(32'h3b6f6eb9),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341d56),
	.w1(32'hbbdab9e8),
	.w2(32'h3c2d912d),
	.w3(32'h3c109b3a),
	.w4(32'h3ac9f647),
	.w5(32'h3badcd47),
	.w6(32'h3b24ae98),
	.w7(32'hba52e3f0),
	.w8(32'hbd016782),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c476444),
	.w1(32'h3bf28a7e),
	.w2(32'hbb4c2f08),
	.w3(32'h3ceb141a),
	.w4(32'h3ce43e4d),
	.w5(32'hbb31677b),
	.w6(32'hbd0e2114),
	.w7(32'hbc54b834),
	.w8(32'h3cbcded0),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2976ac),
	.w1(32'h3b91974c),
	.w2(32'hba7cf3f8),
	.w3(32'hbcfd6bc2),
	.w4(32'hbcefbda6),
	.w5(32'h3a99d6eb),
	.w6(32'h3cbecfa4),
	.w7(32'h3bc2a3f1),
	.w8(32'hba20f7ec),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb30a65),
	.w1(32'hbbb9c615),
	.w2(32'hba8282de),
	.w3(32'hbbe0347e),
	.w4(32'hbc015157),
	.w5(32'hba2c8665),
	.w6(32'hbbdf4ae8),
	.w7(32'hbc0e6d23),
	.w8(32'hbb64a2b7),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18060d),
	.w1(32'hbc2800ba),
	.w2(32'h3b1a320d),
	.w3(32'hbbd6ba70),
	.w4(32'hbc72d1ca),
	.w5(32'h3b273452),
	.w6(32'hbb17e635),
	.w7(32'hbb9602df),
	.w8(32'h3c82582f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c018f23),
	.w1(32'h3d07b2ae),
	.w2(32'hbac7dfa6),
	.w3(32'hbc2d3e10),
	.w4(32'hbc43e192),
	.w5(32'hbc4f299c),
	.w6(32'h3aa49953),
	.w7(32'hbc0d2b09),
	.w8(32'h3c06ca15),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d7f5c),
	.w1(32'h3cddd43e),
	.w2(32'h3b93c594),
	.w3(32'hbc96faec),
	.w4(32'hbc076e0b),
	.w5(32'h3b564ae2),
	.w6(32'h3b5be01a),
	.w7(32'hbc382ee9),
	.w8(32'hbc3adde0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf25d0e),
	.w1(32'h3c191dec),
	.w2(32'h3b280e52),
	.w3(32'h3b9e5b86),
	.w4(32'h3c1246e0),
	.w5(32'h3b420efb),
	.w6(32'hbc735792),
	.w7(32'hbb110d20),
	.w8(32'h3b037d79),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43e83f),
	.w1(32'h3b13de39),
	.w2(32'hbb355bf7),
	.w3(32'h3b37a98d),
	.w4(32'h3b282f50),
	.w5(32'hbb7edfc7),
	.w6(32'h3b037159),
	.w7(32'h3a311c18),
	.w8(32'h3b02eaa3),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e2bd1),
	.w1(32'hbbf0d93c),
	.w2(32'hbb84a630),
	.w3(32'h3a8780d9),
	.w4(32'h3a90673b),
	.w5(32'hbbe83cf0),
	.w6(32'h3b26ed06),
	.w7(32'h3ba23e34),
	.w8(32'hbbd605af),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb508905),
	.w1(32'hbb950280),
	.w2(32'h3adaa470),
	.w3(32'hbb1549d8),
	.w4(32'hbb52df4f),
	.w5(32'hbbae133a),
	.w6(32'hbb99cc35),
	.w7(32'hbb1c6b01),
	.w8(32'h3bcbf7a0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b5662),
	.w1(32'hbba1fb64),
	.w2(32'h3b320c7e),
	.w3(32'h3c87c624),
	.w4(32'h3cd14d4b),
	.w5(32'hbbc932c7),
	.w6(32'h3c526868),
	.w7(32'h3c352049),
	.w8(32'hbc37600d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd4c0e),
	.w1(32'h3bff28d6),
	.w2(32'h3c86d842),
	.w3(32'hbae73391),
	.w4(32'hbb04c018),
	.w5(32'hbb0bbccf),
	.w6(32'hbc382ea6),
	.w7(32'hbba91c61),
	.w8(32'hbc93bfec),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c746b0a),
	.w1(32'h3bc3469d),
	.w2(32'hbbacd87b),
	.w3(32'hbb8cd9df),
	.w4(32'h3c142d8f),
	.w5(32'h3ad2824a),
	.w6(32'hbd675369),
	.w7(32'hbd01f7bb),
	.w8(32'hbb966c5d),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3eff33),
	.w1(32'hbc3af9b4),
	.w2(32'h3c459eca),
	.w3(32'h3c824798),
	.w4(32'h3bbc5e4f),
	.w5(32'h3c13b66f),
	.w6(32'h3c0a596c),
	.w7(32'h3c2c37b0),
	.w8(32'h3c2bb317),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9026eac),
	.w1(32'hba04dbec),
	.w2(32'hbb92e747),
	.w3(32'hba556e28),
	.w4(32'hb960eb91),
	.w5(32'hbb3b0e88),
	.w6(32'h3a2959a2),
	.w7(32'h3aa78bd6),
	.w8(32'hbaa47146),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba93106),
	.w1(32'hb9f8808d),
	.w2(32'hbbae973e),
	.w3(32'hb941a8de),
	.w4(32'h398b8cfc),
	.w5(32'hbb1b38ef),
	.w6(32'h3b210b92),
	.w7(32'h3b5cc441),
	.w8(32'h3cba7d94),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce68d6a),
	.w1(32'hbc8b1d3c),
	.w2(32'hbb22a417),
	.w3(32'hbcd5c5b7),
	.w4(32'hbd12d491),
	.w5(32'h3ba7bbe9),
	.w6(32'h3cf69073),
	.w7(32'h3bb58e04),
	.w8(32'hba8c4871),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3e344),
	.w1(32'hbc2e3a74),
	.w2(32'h3b040fcd),
	.w3(32'hba880675),
	.w4(32'hbc1817f4),
	.w5(32'hba89e3ff),
	.w6(32'hbad18658),
	.w7(32'hbc55feaa),
	.w8(32'hbc187051),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb296d48),
	.w1(32'hbb525ec1),
	.w2(32'hbc4eba2e),
	.w3(32'hbc0446b9),
	.w4(32'hbc6a1f34),
	.w5(32'hbc1bd67e),
	.w6(32'hbc59f1bf),
	.w7(32'hbc222431),
	.w8(32'hbb849424),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaffbfa),
	.w1(32'hbb2a402f),
	.w2(32'hbbb127a8),
	.w3(32'hbc520d1b),
	.w4(32'hbc06d535),
	.w5(32'hbc1145d2),
	.w6(32'hbc7598bf),
	.w7(32'hbc140920),
	.w8(32'hbc08c980),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f0ff),
	.w1(32'hbb1e0b88),
	.w2(32'h3acb018c),
	.w3(32'hbb5e6859),
	.w4(32'hbb4dffcb),
	.w5(32'h3ad21217),
	.w6(32'hbb7db845),
	.w7(32'hbbeb1824),
	.w8(32'h3b4c086a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ce32d),
	.w1(32'h3abf3a98),
	.w2(32'hba8c5ec5),
	.w3(32'h3a06d784),
	.w4(32'h3b67254d),
	.w5(32'hbc0830f8),
	.w6(32'h3b15e8fb),
	.w7(32'h3ae107b3),
	.w8(32'h3c820561),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a2737),
	.w1(32'h3ba33c15),
	.w2(32'h3b2dc2f1),
	.w3(32'hbcff2ae8),
	.w4(32'hbc9c62db),
	.w5(32'hbb144d25),
	.w6(32'hbb2805b0),
	.w7(32'hbc23f85d),
	.w8(32'h3bdf7df9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70b442),
	.w1(32'h393c2419),
	.w2(32'hbba4d506),
	.w3(32'hbcc49585),
	.w4(32'hbc60bb4c),
	.w5(32'hb9c9f68e),
	.w6(32'h3c193182),
	.w7(32'h3c45f033),
	.w8(32'h38e6907f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c6f4c),
	.w1(32'hbc11d19c),
	.w2(32'h3bd44b2b),
	.w3(32'hbc8a36fb),
	.w4(32'hbc9cd1ae),
	.w5(32'hbbee50a0),
	.w6(32'hbc159196),
	.w7(32'hbc3eda37),
	.w8(32'hba7a4249),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5aadc2),
	.w1(32'h3bfcdc44),
	.w2(32'h3a10e662),
	.w3(32'hbc815fd7),
	.w4(32'hbb836e8c),
	.w5(32'hbbc3975b),
	.w6(32'hbc55e599),
	.w7(32'hbc62394e),
	.w8(32'h3bb0911e),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda9eb8),
	.w1(32'h3c3ea6c8),
	.w2(32'hbbea9392),
	.w3(32'hbbfbcaae),
	.w4(32'hbbef0e3d),
	.w5(32'hbb0dd1d9),
	.w6(32'h3c18c3a2),
	.w7(32'hbaf4e4e7),
	.w8(32'hba9edec4),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c7756),
	.w1(32'hba8b2f07),
	.w2(32'hbaf72d7d),
	.w3(32'hbb47e64e),
	.w4(32'hbbb0542b),
	.w5(32'h3b4b5a11),
	.w6(32'h39438656),
	.w7(32'hbbba79c5),
	.w8(32'h3a0ecf45),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cc5b2),
	.w1(32'hbbd09780),
	.w2(32'hb9afd322),
	.w3(32'h3c07b74b),
	.w4(32'h3c5f5b4f),
	.w5(32'hbb7dd418),
	.w6(32'h3b92a2d3),
	.w7(32'h3c42905f),
	.w8(32'h3a01fea0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77faee),
	.w1(32'h37a6dacd),
	.w2(32'hbaf3213b),
	.w3(32'h3b8f4c13),
	.w4(32'h3c66961d),
	.w5(32'h3c07d04a),
	.w6(32'hbb98f3e7),
	.w7(32'hb963a507),
	.w8(32'h3be16933),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe62d84),
	.w1(32'hbbe73536),
	.w2(32'hbc2f6525),
	.w3(32'hbbfd542f),
	.w4(32'hbbfc6f66),
	.w5(32'hbaa96eb6),
	.w6(32'hbc469cca),
	.w7(32'hba3f9fd4),
	.w8(32'hbbf5b534),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad51f2),
	.w1(32'hbac90140),
	.w2(32'hbc046dda),
	.w3(32'h3b78c46a),
	.w4(32'h3b1ff663),
	.w5(32'h3b7c364d),
	.w6(32'hba93bcee),
	.w7(32'h3b8aa886),
	.w8(32'hbc14fcf3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90579a),
	.w1(32'hbca713bb),
	.w2(32'hbba06b46),
	.w3(32'h3be998fc),
	.w4(32'h3b012c24),
	.w5(32'h389874b4),
	.w6(32'h3b967b4d),
	.w7(32'h3b4d24c8),
	.w8(32'h3bae62ae),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a26d),
	.w1(32'hbc4f8b64),
	.w2(32'h3b0b9fc3),
	.w3(32'hbb0fd81b),
	.w4(32'hbbe85e92),
	.w5(32'h392941ed),
	.w6(32'hbb118e7b),
	.w7(32'hbb95b184),
	.w8(32'hbb5a7445),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2e6b3),
	.w1(32'hbba36069),
	.w2(32'hb962449b),
	.w3(32'h3aba394d),
	.w4(32'h3abc9120),
	.w5(32'h3b4656bc),
	.w6(32'hb99f147b),
	.w7(32'h3b7f87d3),
	.w8(32'h3a6d6a34),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d605),
	.w1(32'h3b1ba43f),
	.w2(32'h3c19b109),
	.w3(32'h3af5f3fa),
	.w4(32'h3a3dc3d6),
	.w5(32'h3a88cdae),
	.w6(32'h3b188a8e),
	.w7(32'hbbd07c00),
	.w8(32'hbcbc0f93),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88747e),
	.w1(32'h3c37b59c),
	.w2(32'h3b02d316),
	.w3(32'h3bb0bac4),
	.w4(32'h3b6073fd),
	.w5(32'hbaac2ab4),
	.w6(32'hbd0507d8),
	.w7(32'hbc97a4c8),
	.w8(32'hbaf8dbf4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5c9e9),
	.w1(32'hba8e4609),
	.w2(32'h3bca17dd),
	.w3(32'hbbb79636),
	.w4(32'h3b840a9d),
	.w5(32'hba8778a8),
	.w6(32'hbb01140f),
	.w7(32'h3a7c2b52),
	.w8(32'hba22344b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1da561),
	.w1(32'h3b267f37),
	.w2(32'h3ace0d08),
	.w3(32'hbbcada8a),
	.w4(32'hba5ef240),
	.w5(32'h3c04c8c5),
	.w6(32'h3bd4dd49),
	.w7(32'h3b9a0dfc),
	.w8(32'h3ba780dc),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4154e9),
	.w1(32'hbbfaec6d),
	.w2(32'hbbbb9b29),
	.w3(32'h3c8e889d),
	.w4(32'h3c3f9612),
	.w5(32'hbbe4a6b5),
	.w6(32'h3c1094e5),
	.w7(32'h3cb09b6d),
	.w8(32'h3b80216e),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf16b57),
	.w1(32'hbc874f9c),
	.w2(32'hba039c8e),
	.w3(32'hbaaf5551),
	.w4(32'hbbda02aa),
	.w5(32'hb9531e34),
	.w6(32'h3cd05630),
	.w7(32'h3ca27897),
	.w8(32'hbba7c87f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d1530),
	.w1(32'hbbe420de),
	.w2(32'h3b43096e),
	.w3(32'h3c0b5d90),
	.w4(32'hb889d985),
	.w5(32'hbbb030e3),
	.w6(32'hba05cb2d),
	.w7(32'h3b583653),
	.w8(32'hbc0c2266),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41910a),
	.w1(32'h3c0e7981),
	.w2(32'h3952879d),
	.w3(32'hbc08abdd),
	.w4(32'hbc39fbe6),
	.w5(32'h3bbfee98),
	.w6(32'hbc6c25a0),
	.w7(32'hbc855b7c),
	.w8(32'h3b230782),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a01f),
	.w1(32'h3b257e5d),
	.w2(32'hbb108977),
	.w3(32'h3bc3709c),
	.w4(32'hbad2aed1),
	.w5(32'h3a97cc4e),
	.w6(32'h3b987d48),
	.w7(32'hb98080b7),
	.w8(32'h3bf0cfb3),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08ad11),
	.w1(32'h3c1a25c1),
	.w2(32'h3aa830c3),
	.w3(32'hbb32adf8),
	.w4(32'h3b926e1a),
	.w5(32'h3b487c3f),
	.w6(32'hbb9235e3),
	.w7(32'hbbfef1c0),
	.w8(32'hbb089b33),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87fc8e),
	.w1(32'h3c0b1e65),
	.w2(32'hbb07dca8),
	.w3(32'hbaa842e1),
	.w4(32'hbac7261e),
	.w5(32'hbc2b527b),
	.w6(32'hba9f85ce),
	.w7(32'h3888f803),
	.w8(32'hbb502ce6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed2f2),
	.w1(32'h3c65102e),
	.w2(32'hbb654271),
	.w3(32'hbc09ac06),
	.w4(32'hbad033b4),
	.w5(32'h3a16862b),
	.w6(32'hbb937eba),
	.w7(32'hbc1abed8),
	.w8(32'hbc710a39),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7db23),
	.w1(32'hbbee3ec0),
	.w2(32'hba37610b),
	.w3(32'h3c4ee6b1),
	.w4(32'h3ccc306b),
	.w5(32'hba845177),
	.w6(32'hbb9aa9f8),
	.w7(32'h3b9761a7),
	.w8(32'hbbad9310),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cb250),
	.w1(32'h3ad7753c),
	.w2(32'hba8920e9),
	.w3(32'hbb75847b),
	.w4(32'hbc252779),
	.w5(32'hbb0811bd),
	.w6(32'hbb5a3a8c),
	.w7(32'hb876d2f6),
	.w8(32'hba05428c),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1eb5b8),
	.w1(32'hbae70c81),
	.w2(32'hb8c73274),
	.w3(32'hba40b85e),
	.w4(32'hbb068ab2),
	.w5(32'h3b0901cc),
	.w6(32'h3a34ae7a),
	.w7(32'hb84663a3),
	.w8(32'hb9b681f3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c81dc),
	.w1(32'hbb6180b6),
	.w2(32'h3a05c457),
	.w3(32'h3b41da79),
	.w4(32'hbb824cbe),
	.w5(32'hbc2e7aa7),
	.w6(32'h3631d990),
	.w7(32'hbb10d9ff),
	.w8(32'hbbacdec2),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e4620),
	.w1(32'h3806964b),
	.w2(32'h3b144bf8),
	.w3(32'h3c28cc29),
	.w4(32'h3c982f24),
	.w5(32'h3b69f2c9),
	.w6(32'h3a55cba4),
	.w7(32'hbb86e907),
	.w8(32'hbb837807),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea37da),
	.w1(32'h3b8d01a7),
	.w2(32'hbbe7678f),
	.w3(32'h3b32c94d),
	.w4(32'h3b550a94),
	.w5(32'hbad838c6),
	.w6(32'hbbd342ae),
	.w7(32'h3a1885d4),
	.w8(32'h3c03b519),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bf487),
	.w1(32'hbc8c70e8),
	.w2(32'hbb9eac5d),
	.w3(32'hbbbbe25b),
	.w4(32'hbc4d4bb0),
	.w5(32'h3c312e9b),
	.w6(32'h3c09d2d5),
	.w7(32'h3c129712),
	.w8(32'h3b0fa42c),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab3289),
	.w1(32'hbcc7028e),
	.w2(32'h3af4b7f1),
	.w3(32'h3cc62e24),
	.w4(32'h3c72d647),
	.w5(32'h3c88dfdd),
	.w6(32'h3c8eb479),
	.w7(32'h3c94c41e),
	.w8(32'hbbbb5ef0),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca87359),
	.w1(32'hbca7bef0),
	.w2(32'h3b8caf39),
	.w3(32'h3d02cc21),
	.w4(32'h3ce7a0c2),
	.w5(32'h3b49bb7c),
	.w6(32'h3c1d86b2),
	.w7(32'h3cb3824e),
	.w8(32'hbbe5660b),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule