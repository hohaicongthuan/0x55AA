module layer_8_featuremap_100(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8038e5),
	.w1(32'h3bc58e90),
	.w2(32'h3baa7e51),
	.w3(32'hbc10dcc5),
	.w4(32'h3bdcae13),
	.w5(32'h3c347e92),
	.w6(32'hbb3b3f05),
	.w7(32'h3a762509),
	.w8(32'h3c10bc72),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafa48f),
	.w1(32'hb99b776b),
	.w2(32'h3ad9b818),
	.w3(32'h3b81cd4b),
	.w4(32'hbb136a2a),
	.w5(32'h3c23a65a),
	.w6(32'h3bff0639),
	.w7(32'h3bf7811d),
	.w8(32'h3c8ea189),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdb0f5f),
	.w1(32'hbb5ebc13),
	.w2(32'h3ba8fa6e),
	.w3(32'hbb30bafd),
	.w4(32'hbbd00b32),
	.w5(32'hbafa2966),
	.w6(32'h3b5193c6),
	.w7(32'h3ba8b660),
	.w8(32'h3c9937ce),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d2cca),
	.w1(32'h3c0ce835),
	.w2(32'h3c055876),
	.w3(32'h3bf155e5),
	.w4(32'h3bbf98a1),
	.w5(32'h3c21611b),
	.w6(32'h3c8d0841),
	.w7(32'hbaeb6805),
	.w8(32'h3a40229e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f0fd8),
	.w1(32'h3c8e3458),
	.w2(32'h3c86e20f),
	.w3(32'h3c41e74f),
	.w4(32'h3c17a322),
	.w5(32'h3cbec59c),
	.w6(32'h3b868eb2),
	.w7(32'h3c27a45c),
	.w8(32'h3cae637d),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce806da),
	.w1(32'h3c3c66ed),
	.w2(32'h3cf4ebce),
	.w3(32'h3cb900bb),
	.w4(32'h3c68b0a5),
	.w5(32'h3c4b8e87),
	.w6(32'h3c801b7d),
	.w7(32'h3bc59e1f),
	.w8(32'h3baedee4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032930),
	.w1(32'h3bcbd130),
	.w2(32'hbb0cf0a3),
	.w3(32'h3bc9e404),
	.w4(32'hba8f6c7c),
	.w5(32'hbae7d801),
	.w6(32'h3aed5f6f),
	.w7(32'hb9edd7d5),
	.w8(32'hbb5072fd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1cea0),
	.w1(32'h3c092fde),
	.w2(32'h3cedbbed),
	.w3(32'h3c14e3f0),
	.w4(32'h3c3cff49),
	.w5(32'h3c05ef1c),
	.w6(32'h3cb714e6),
	.w7(32'h3cbb75a6),
	.w8(32'h3bc7cae8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51f6cf),
	.w1(32'hbc01dadf),
	.w2(32'hbc17bdbc),
	.w3(32'h3c67233d),
	.w4(32'h3c99592b),
	.w5(32'h3ca656e0),
	.w6(32'h3be25d28),
	.w7(32'h3c4b3ff4),
	.w8(32'h3c89555a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa0d0),
	.w1(32'hbb914568),
	.w2(32'h3a981c17),
	.w3(32'h3c09e647),
	.w4(32'hba704c45),
	.w5(32'h3b865502),
	.w6(32'hbbb967c3),
	.w7(32'h3b37e910),
	.w8(32'h3bf03173),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2148e8),
	.w1(32'hbc583c9c),
	.w2(32'h3b5491e0),
	.w3(32'hbbce0db2),
	.w4(32'h3b527679),
	.w5(32'h38094a05),
	.w6(32'hbc80fd4d),
	.w7(32'h3b744be3),
	.w8(32'h3aef4665),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50250f),
	.w1(32'hbc2e2f30),
	.w2(32'h3c32e02c),
	.w3(32'h3aa0cb89),
	.w4(32'h3b7b6930),
	.w5(32'h3c095b8b),
	.w6(32'hbc56defb),
	.w7(32'h3bb3b70d),
	.w8(32'h3c3f88ba),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b886b96),
	.w1(32'h3bcef748),
	.w2(32'h3be42acb),
	.w3(32'h3cbcc2da),
	.w4(32'h3badca61),
	.w5(32'h3c56f8a5),
	.w6(32'h3cc8b8d3),
	.w7(32'h3c042fad),
	.w8(32'h3c96ffb6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4e1a7),
	.w1(32'hbac51475),
	.w2(32'h3b1440e0),
	.w3(32'h3a0ddd75),
	.w4(32'h39370434),
	.w5(32'h3ad59524),
	.w6(32'h3c16a781),
	.w7(32'h3adb93ee),
	.w8(32'h3b8b1bb5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeaa687),
	.w1(32'h3b6377b7),
	.w2(32'h3a8951a2),
	.w3(32'h3c0ba887),
	.w4(32'h3b342a2e),
	.w5(32'hb7f96e0c),
	.w6(32'h3ba668d4),
	.w7(32'h3afc1936),
	.w8(32'h3a0b8b7b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e39ae8),
	.w1(32'h3bb1b01f),
	.w2(32'hb937f3dd),
	.w3(32'h3ba1d6f7),
	.w4(32'h3bd4826d),
	.w5(32'hbb4b7a6a),
	.w6(32'h3bb62f6f),
	.w7(32'h3b11b4d1),
	.w8(32'hbb0e076b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa167b2),
	.w1(32'h3b88bb94),
	.w2(32'h39b8b88f),
	.w3(32'hbaa5a766),
	.w4(32'hbc063afa),
	.w5(32'hbc4cb0c9),
	.w6(32'hbaf3bfa0),
	.w7(32'hbaad11ec),
	.w8(32'hbc9e548a),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ac81a),
	.w1(32'hbb3ea501),
	.w2(32'h39888712),
	.w3(32'hbbeaee07),
	.w4(32'h3b92826b),
	.w5(32'h3c4f81a1),
	.w6(32'h3b4270d7),
	.w7(32'hbb619d73),
	.w8(32'h3c258cd9),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e3831),
	.w1(32'h39f3f352),
	.w2(32'h3c56f91b),
	.w3(32'hbb27ac20),
	.w4(32'h3c19afd0),
	.w5(32'hbc055e90),
	.w6(32'h3bef3806),
	.w7(32'h3c1ae507),
	.w8(32'h3ba1f3ae),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5eed2c),
	.w1(32'h3b9ed593),
	.w2(32'h3d02df01),
	.w3(32'h3ccd6dc0),
	.w4(32'h3a967145),
	.w5(32'h3c69a407),
	.w6(32'h3cf68413),
	.w7(32'h3d6abcc1),
	.w8(32'h3d9ea2a0),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c678db7),
	.w1(32'h399eff02),
	.w2(32'hbb0402c3),
	.w3(32'hbaf74db2),
	.w4(32'hbb9a99d5),
	.w5(32'h3c93e8e7),
	.w6(32'h3a831975),
	.w7(32'hbc9ecd3e),
	.w8(32'hbbb02c6c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65a0c9),
	.w1(32'hbc593beb),
	.w2(32'hbbb29684),
	.w3(32'h3bd7ffdc),
	.w4(32'h3adba69b),
	.w5(32'h3c4cc241),
	.w6(32'h3c197e68),
	.w7(32'h3b93c51f),
	.w8(32'h3bcb6e98),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb581db1),
	.w1(32'h3c91a003),
	.w2(32'h3cc38ce1),
	.w3(32'h3b336b7e),
	.w4(32'h3d1677c6),
	.w5(32'h3cfd8ddf),
	.w6(32'h3beecba4),
	.w7(32'h3d169028),
	.w8(32'h3d142976),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3044ca),
	.w1(32'hbc1dd118),
	.w2(32'h3bb6ae09),
	.w3(32'hbb716d97),
	.w4(32'h3ba31f6d),
	.w5(32'h3c205398),
	.w6(32'hbc0ab543),
	.w7(32'h3bb03802),
	.w8(32'h3c1bf155),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0acac),
	.w1(32'h3b11223b),
	.w2(32'h3b86f8b4),
	.w3(32'h3b5d900b),
	.w4(32'h3a7a341b),
	.w5(32'hbabad314),
	.w6(32'h3b7cb2d0),
	.w7(32'hbbdde68d),
	.w8(32'hbc503b6c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ca23e),
	.w1(32'h3c2b113b),
	.w2(32'h3cf98687),
	.w3(32'h3c22cefc),
	.w4(32'h3ac62640),
	.w5(32'h3b92638f),
	.w6(32'h3c0d3fec),
	.w7(32'h3d19f327),
	.w8(32'h3d3ec9c9),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4df78),
	.w1(32'h3b2bda0d),
	.w2(32'hbafda6c8),
	.w3(32'h3c0b0b66),
	.w4(32'hb9a24de3),
	.w5(32'hbc09c33b),
	.w6(32'h3b1678db),
	.w7(32'hbc062f0e),
	.w8(32'hbc206530),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6ea052),
	.w1(32'h3c098680),
	.w2(32'h3c6ad90f),
	.w3(32'hbc6695c2),
	.w4(32'h3d55ec88),
	.w5(32'h3da8a62f),
	.w6(32'hbd23a9c8),
	.w7(32'h3c853674),
	.w8(32'h3ccd522a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9bd259),
	.w1(32'hb9e575e6),
	.w2(32'h3c246fe5),
	.w3(32'hbbe3153a),
	.w4(32'hb94541c1),
	.w5(32'h3bb407cb),
	.w6(32'hbbbbe3f6),
	.w7(32'h3c19ced7),
	.w8(32'h3c62356e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac85433),
	.w1(32'hbbad0fc6),
	.w2(32'hbbe90d0e),
	.w3(32'hba7a8ff3),
	.w4(32'h3b8bd801),
	.w5(32'h3c0dc706),
	.w6(32'hbb805748),
	.w7(32'h3b940d0f),
	.w8(32'h3ca926f3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb806378),
	.w1(32'h3b15081c),
	.w2(32'hbaef3b0e),
	.w3(32'h3c69bd2b),
	.w4(32'hbb3fad00),
	.w5(32'hbb8d644e),
	.w6(32'h3b828c5b),
	.w7(32'hbc455d98),
	.w8(32'hbc46abeb),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d14dc),
	.w1(32'h3ba6367c),
	.w2(32'hbbc00b97),
	.w3(32'h3b8bec0b),
	.w4(32'hbbfa5813),
	.w5(32'h3be108e9),
	.w6(32'h3c1293f1),
	.w7(32'h3b94f684),
	.w8(32'h3c9cd562),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fd84c),
	.w1(32'hbc2c6a68),
	.w2(32'hbbdc28c5),
	.w3(32'hbc0a5225),
	.w4(32'hbb8e9e1a),
	.w5(32'h3cac4d59),
	.w6(32'h3b050355),
	.w7(32'h3b984b40),
	.w8(32'h3d6b34e8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47f0ae),
	.w1(32'hbc4e191d),
	.w2(32'h3aea19fa),
	.w3(32'hbad01828),
	.w4(32'hbbabcfd9),
	.w5(32'hbbe17060),
	.w6(32'h3bcffa2d),
	.w7(32'h39bc677b),
	.w8(32'h3bbd920e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5c82c),
	.w1(32'hbc0f1b11),
	.w2(32'h3bd18bd9),
	.w3(32'h3c1d7dd9),
	.w4(32'hbca314b1),
	.w5(32'hbc1f9475),
	.w6(32'h3c3b0e7f),
	.w7(32'hbc1e5512),
	.w8(32'h3c00b234),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a9908),
	.w1(32'h3c16c2d9),
	.w2(32'hbbe9f8d3),
	.w3(32'h3b8a800d),
	.w4(32'h3c87257a),
	.w5(32'h3c203bcc),
	.w6(32'h3c00664e),
	.w7(32'hbbd461ef),
	.w8(32'h3b071f2d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23492c),
	.w1(32'hbb354489),
	.w2(32'h3ab45019),
	.w3(32'hbab964ee),
	.w4(32'hbc654c04),
	.w5(32'hbbf024b0),
	.w6(32'hbbb3a41d),
	.w7(32'hbc946456),
	.w8(32'hbc877708),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a3c5f),
	.w1(32'hbcbb135e),
	.w2(32'h3c27c708),
	.w3(32'hbbbeece4),
	.w4(32'h3bc88ac2),
	.w5(32'h3b99961d),
	.w6(32'hbc84ab3a),
	.w7(32'h3c9bf6cd),
	.w8(32'h3c0fd926),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb9c2f),
	.w1(32'hbaa89c72),
	.w2(32'h3bb86784),
	.w3(32'h3b48ad20),
	.w4(32'h3adc0cff),
	.w5(32'hbc8c9492),
	.w6(32'hbb60fa83),
	.w7(32'h3c03e050),
	.w8(32'h39d1cb24),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbde3a),
	.w1(32'hbb9522f3),
	.w2(32'hbad5da52),
	.w3(32'hbc82acd2),
	.w4(32'hbb5d2bd2),
	.w5(32'hbb9328a7),
	.w6(32'hbbc85006),
	.w7(32'hbb63981f),
	.w8(32'hbbaa791d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c2d6f),
	.w1(32'h3c80dee3),
	.w2(32'h3cf8dbb5),
	.w3(32'h3d0abf58),
	.w4(32'h3ca9d3bc),
	.w5(32'h3c9b45f7),
	.w6(32'h3d17c11b),
	.w7(32'h3d04c0c8),
	.w8(32'h3d5dbfcf),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3bd3f),
	.w1(32'hbba388d8),
	.w2(32'hbc6537ac),
	.w3(32'h3c1ecc8d),
	.w4(32'h3c62e99b),
	.w5(32'h3a67ffa4),
	.w6(32'h3c92e773),
	.w7(32'hbbea648d),
	.w8(32'h3a71bea4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4ae0),
	.w1(32'h3ba6717e),
	.w2(32'hbb72e18f),
	.w3(32'hbc00cae3),
	.w4(32'hbc0905a4),
	.w5(32'h3c49a4f6),
	.w6(32'h3b45f53f),
	.w7(32'hbbcb3ec0),
	.w8(32'hbbf86361),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd1543),
	.w1(32'hbbb9c6c2),
	.w2(32'h3bf4f62c),
	.w3(32'h3c0f50b1),
	.w4(32'h3bc08c83),
	.w5(32'h3b5cc540),
	.w6(32'hbc890f70),
	.w7(32'h3c4dd4ef),
	.w8(32'h3c876ae9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd25d89),
	.w1(32'h3bacba63),
	.w2(32'h3c51c39c),
	.w3(32'h3bc4b3e6),
	.w4(32'h3bcf9c3a),
	.w5(32'h3bb50eae),
	.w6(32'h3c349cbe),
	.w7(32'h3c04be5e),
	.w8(32'hb9d18eaa),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf5698),
	.w1(32'hba2ec256),
	.w2(32'hbbe17963),
	.w3(32'h3c01d4c0),
	.w4(32'h3c3af247),
	.w5(32'h3b8b0c4a),
	.w6(32'h3beaaa4a),
	.w7(32'hbb8f32ad),
	.w8(32'h3af372a6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e2276),
	.w1(32'h3b51020c),
	.w2(32'h3be4da90),
	.w3(32'hbc998a3a),
	.w4(32'hbc33643c),
	.w5(32'hbc4c0f70),
	.w6(32'hbc529adb),
	.w7(32'hbb90dd04),
	.w8(32'hbb8acee2),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9921a80),
	.w1(32'h3c17ba59),
	.w2(32'h3d01c02a),
	.w3(32'hbba7145d),
	.w4(32'h3c47ece5),
	.w5(32'h3c9a9442),
	.w6(32'hbbf85c3d),
	.w7(32'h3ca175bd),
	.w8(32'h3c268660),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b335ba1),
	.w1(32'hbb9825e4),
	.w2(32'h3ad6cae8),
	.w3(32'h3c61930f),
	.w4(32'h3c52cabd),
	.w5(32'h3b6d4230),
	.w6(32'h3c36c2f4),
	.w7(32'hbc32c8c4),
	.w8(32'hbc89b5b0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabc707),
	.w1(32'hbbab2812),
	.w2(32'h3c074eb4),
	.w3(32'hbc8d116b),
	.w4(32'h3aeadae1),
	.w5(32'hbc18f1bb),
	.w6(32'hbc77ab65),
	.w7(32'hbb8891f5),
	.w8(32'hbc643a07),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4621a7),
	.w1(32'hba58f7d4),
	.w2(32'h3c45d0a9),
	.w3(32'hbbbefb9e),
	.w4(32'h3cbc9fab),
	.w5(32'h3c8a79d8),
	.w6(32'h3b6e8e06),
	.w7(32'h3d56b4d3),
	.w8(32'h3d48c75a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa393c),
	.w1(32'h3d51f172),
	.w2(32'h3d766cde),
	.w3(32'h3d00f255),
	.w4(32'h3c0c12ee),
	.w5(32'h3cb08a0c),
	.w6(32'h3d56a5fb),
	.w7(32'h3d20df1a),
	.w8(32'h3d585fef),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc912f5),
	.w1(32'h3c5ec68f),
	.w2(32'h3cd2fb5d),
	.w3(32'h3be095c8),
	.w4(32'h3bac14db),
	.w5(32'h3c94a083),
	.w6(32'h3c98a04a),
	.w7(32'h3cc9e0fa),
	.w8(32'h3cf5926d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc855fbd),
	.w1(32'hbc1c3944),
	.w2(32'h3a99d606),
	.w3(32'hbc20cf01),
	.w4(32'hbafdfbf9),
	.w5(32'hba46ecc6),
	.w6(32'hbc541462),
	.w7(32'hbbb5a844),
	.w8(32'h3c22b390),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a006bf7),
	.w1(32'hba1487f2),
	.w2(32'h3c2f3638),
	.w3(32'h3b2f9ea3),
	.w4(32'hbb50bc72),
	.w5(32'hbc3e3be5),
	.w6(32'h3b547017),
	.w7(32'hba19ce7d),
	.w8(32'hbc8bdec2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3890cf37),
	.w1(32'hb90033c3),
	.w2(32'h3c80ee06),
	.w3(32'hbc36126f),
	.w4(32'hbb2c146d),
	.w5(32'hbbe107f8),
	.w6(32'hbc98dd6d),
	.w7(32'h3c30a0aa),
	.w8(32'h3bed4b30),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e6d40),
	.w1(32'h39e58965),
	.w2(32'h3b577333),
	.w3(32'h3b51c083),
	.w4(32'h3bcce1da),
	.w5(32'h3a93f94b),
	.w6(32'hbbc6a8c3),
	.w7(32'hbbb10317),
	.w8(32'hbbfec893),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c875341),
	.w1(32'h3c13e5d5),
	.w2(32'h3c13ba8e),
	.w3(32'h3cf67707),
	.w4(32'h3bc12b9f),
	.w5(32'h3c1fb42e),
	.w6(32'h3cb05914),
	.w7(32'hbc1fdfd1),
	.w8(32'hbc14a203),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad07fd6),
	.w1(32'h3c897d85),
	.w2(32'h3afb1c46),
	.w3(32'h3c13a29c),
	.w4(32'h3acd92ce),
	.w5(32'h3b26ca28),
	.w6(32'hbb67da08),
	.w7(32'h3be5ac53),
	.w8(32'h3c0951eb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd66d1b),
	.w1(32'h3bd01270),
	.w2(32'h3c81df27),
	.w3(32'h3c106a1e),
	.w4(32'hbc1e9e57),
	.w5(32'h3ae1f8de),
	.w6(32'h3c4d62ea),
	.w7(32'hbb895027),
	.w8(32'h3ba52470),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65b0a2),
	.w1(32'h3c12d78c),
	.w2(32'hbd1325f2),
	.w3(32'hbb5cd1a8),
	.w4(32'hbb480931),
	.w5(32'hbc0791f0),
	.w6(32'hbc6729a6),
	.w7(32'hbc513076),
	.w8(32'h3bd5cedd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906ab08),
	.w1(32'h3bfbf7ee),
	.w2(32'h39ebb604),
	.w3(32'h3ace7b5a),
	.w4(32'h3bcdd80e),
	.w5(32'h39057a22),
	.w6(32'h3c855eba),
	.w7(32'h3aab49e5),
	.w8(32'hbba5c769),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b249412),
	.w1(32'h3b7ee5d0),
	.w2(32'h3cba4367),
	.w3(32'h3cb476bb),
	.w4(32'hbb039101),
	.w5(32'h3c038e12),
	.w6(32'h3c89fce4),
	.w7(32'hbb4cb5a9),
	.w8(32'h3cb327aa),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cf611),
	.w1(32'h3b9b28c6),
	.w2(32'h3c1f05e0),
	.w3(32'hbb45c7c6),
	.w4(32'hbc1a4d32),
	.w5(32'hbb8bafd9),
	.w6(32'h3b0f7ce1),
	.w7(32'h3c0f5eea),
	.w8(32'h3cc1eb7c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e578d),
	.w1(32'h3b5ef3d5),
	.w2(32'hba761ae1),
	.w3(32'hbbee381c),
	.w4(32'hba6282fa),
	.w5(32'h3a8ff191),
	.w6(32'h3bd8d84d),
	.w7(32'hb9524046),
	.w8(32'h3aa0fc43),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b8b93),
	.w1(32'h3b4c33f6),
	.w2(32'h3c2b7fd3),
	.w3(32'h3be5e6a9),
	.w4(32'h3c252ad7),
	.w5(32'h3c1cc951),
	.w6(32'h3a361a76),
	.w7(32'h3c6ac297),
	.w8(32'h3ca29a1d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14b7c8),
	.w1(32'h3b8f16ed),
	.w2(32'h3c8d9ca0),
	.w3(32'h3bae60f3),
	.w4(32'hbab65ca9),
	.w5(32'h3bbfcde8),
	.w6(32'h3c20933f),
	.w7(32'h3c40ab6b),
	.w8(32'h3ccd9285),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67ef51),
	.w1(32'h3b1096fc),
	.w2(32'h3baa7327),
	.w3(32'hbb72a270),
	.w4(32'h3c2fb7e4),
	.w5(32'h3d0bbce7),
	.w6(32'h3ae63fcd),
	.w7(32'h3ba775cd),
	.w8(32'h3d18dff4),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c799da5),
	.w1(32'hbaf62e34),
	.w2(32'h3bda99e9),
	.w3(32'hbbfc3be1),
	.w4(32'hbb980db0),
	.w5(32'hbc41fb63),
	.w6(32'hb8bb9843),
	.w7(32'hbc2d41df),
	.w8(32'hbc2484c6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983a089),
	.w1(32'h3acbe979),
	.w2(32'h3c6ea4e4),
	.w3(32'hbcd12f99),
	.w4(32'h3b947871),
	.w5(32'h3ca93647),
	.w6(32'hbcd12ba3),
	.w7(32'h3c78dc3f),
	.w8(32'h3cc793bd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c237c),
	.w1(32'hbb1f7caa),
	.w2(32'h3a569d07),
	.w3(32'hbb9d954e),
	.w4(32'h3bacced9),
	.w5(32'h3c639068),
	.w6(32'hb99d158a),
	.w7(32'hbaa6f4d6),
	.w8(32'h3c020588),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3eee),
	.w1(32'hbb89bc16),
	.w2(32'hbb89cbfd),
	.w3(32'h3aa61b7f),
	.w4(32'hbc256dd0),
	.w5(32'hbbd89ca8),
	.w6(32'h38b730ac),
	.w7(32'hbc469723),
	.w8(32'h3ba1dfce),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d562fd),
	.w1(32'h3aeb60c5),
	.w2(32'hbadaf8e7),
	.w3(32'hbc022c62),
	.w4(32'hbb121876),
	.w5(32'hb9dec6c2),
	.w6(32'h3aa897b2),
	.w7(32'hbb7eb385),
	.w8(32'hbb6a1762),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6d39f),
	.w1(32'hbc0edffe),
	.w2(32'h3c99ef56),
	.w3(32'hbc9946ef),
	.w4(32'hbcab2cd5),
	.w5(32'hbaa5f3e2),
	.w6(32'hbc5ef602),
	.w7(32'hbb17f168),
	.w8(32'h3ca9973e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca6f29d),
	.w1(32'hbc395d5e),
	.w2(32'hb9f5f56a),
	.w3(32'hbc4b551f),
	.w4(32'hbba2e04d),
	.w5(32'hbc3cb2cc),
	.w6(32'hbc4e1b06),
	.w7(32'hbca1a587),
	.w8(32'hbcff9d98),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69fb05),
	.w1(32'hb9172976),
	.w2(32'h3bc31490),
	.w3(32'h3c8f2a88),
	.w4(32'h3c5960e8),
	.w5(32'h3b8250fd),
	.w6(32'hbb8695b3),
	.w7(32'h3ae9512b),
	.w8(32'h3b91c063),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dce59),
	.w1(32'hbb52ce6e),
	.w2(32'hba3613ab),
	.w3(32'hbc1a6550),
	.w4(32'hbb7e9ae6),
	.w5(32'hbb20288c),
	.w6(32'hbb83f829),
	.w7(32'h3c27a795),
	.w8(32'hbab21ec0),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1b3a4),
	.w1(32'h3c2c4476),
	.w2(32'h3c6f23c5),
	.w3(32'h3ba4fc45),
	.w4(32'h3ba62398),
	.w5(32'h3c6d110d),
	.w6(32'hbbadcee8),
	.w7(32'h3bd9f7d5),
	.w8(32'h3c8ee907),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37449f),
	.w1(32'h3bbf1f00),
	.w2(32'h3c019517),
	.w3(32'h3b9a8619),
	.w4(32'h3a5bad92),
	.w5(32'hb9284dfc),
	.w6(32'h3c23e09f),
	.w7(32'h3bb72d21),
	.w8(32'h3bf4e414),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b4556),
	.w1(32'h3a350d8d),
	.w2(32'hbbb0b81a),
	.w3(32'h3b392a8a),
	.w4(32'h3b9a4032),
	.w5(32'h3c302005),
	.w6(32'h3b81f660),
	.w7(32'hbb731597),
	.w8(32'hbca669b1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba376c),
	.w1(32'h38d74112),
	.w2(32'hbbbe222f),
	.w3(32'h3a0762f7),
	.w4(32'h3ba66267),
	.w5(32'h3b985bb7),
	.w6(32'hbbe34c70),
	.w7(32'hba9eb267),
	.w8(32'hbc3216f2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6102f8),
	.w1(32'hbb918256),
	.w2(32'hbc506130),
	.w3(32'hb9b9ab8f),
	.w4(32'hbc5be482),
	.w5(32'hbbc9edc6),
	.w6(32'h3b37c34e),
	.w7(32'h3bb03ac5),
	.w8(32'hbc11607f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cff480f),
	.w1(32'h3cb1be27),
	.w2(32'h3ca577d6),
	.w3(32'h3bdb2274),
	.w4(32'h3c6a5746),
	.w5(32'h3cc482cf),
	.w6(32'h3bd416d7),
	.w7(32'h3d33a153),
	.w8(32'h3ce64330),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f250b),
	.w1(32'h3ce88e96),
	.w2(32'h3d2240cb),
	.w3(32'h3d21efbc),
	.w4(32'h3d0e5e00),
	.w5(32'h3d101de1),
	.w6(32'h3d128127),
	.w7(32'h3ccb8715),
	.w8(32'h3db98760),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6f063),
	.w1(32'h3b04d783),
	.w2(32'h3cf64d79),
	.w3(32'h3ca0a27d),
	.w4(32'h3c5dd5fc),
	.w5(32'h3d0b047a),
	.w6(32'hbb89f5c8),
	.w7(32'h3d68b7d9),
	.w8(32'h3dc089ba),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc47c),
	.w1(32'h3ce60a32),
	.w2(32'h3c7bc6dd),
	.w3(32'hbc41347e),
	.w4(32'hbb59ae31),
	.w5(32'h3b4134f2),
	.w6(32'hbc137c53),
	.w7(32'hbc08ed7e),
	.w8(32'h3cf5744d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf952d9),
	.w1(32'hbc86b06c),
	.w2(32'hbb1baf3d),
	.w3(32'h3c0380dd),
	.w4(32'h3c42f787),
	.w5(32'h3baef4b5),
	.w6(32'hba170f8f),
	.w7(32'hba64bce9),
	.w8(32'hbafa05c6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28f18d),
	.w1(32'hbc9be48c),
	.w2(32'hba2288ea),
	.w3(32'h3c5626ad),
	.w4(32'h3bd17249),
	.w5(32'h3c15f3b1),
	.w6(32'h3bfc2071),
	.w7(32'hbbf412c3),
	.w8(32'hbb3a8453),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9478ed),
	.w1(32'hbb5e5f42),
	.w2(32'hbaad796f),
	.w3(32'hbb065b80),
	.w4(32'hba2042ec),
	.w5(32'hbb8af0a0),
	.w6(32'hbb153fc6),
	.w7(32'h3a1e62ae),
	.w8(32'h3a7bd21a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89cc85),
	.w1(32'h3b1bd73b),
	.w2(32'h3c4d7cf3),
	.w3(32'h3baf308e),
	.w4(32'h39b8a7b2),
	.w5(32'h3be8bc65),
	.w6(32'hbb53c9b6),
	.w7(32'hbcf07c4f),
	.w8(32'h3c101ee2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5afc0),
	.w1(32'hbcb0d056),
	.w2(32'h3c6e8baa),
	.w3(32'h3c95ca59),
	.w4(32'hbc746271),
	.w5(32'hba525c82),
	.w6(32'h3d4487f8),
	.w7(32'h3be5ade3),
	.w8(32'h3c8b8c48),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fe8b1),
	.w1(32'h3cb4b638),
	.w2(32'hbb8d1fb5),
	.w3(32'hbb84579a),
	.w4(32'hbbde0087),
	.w5(32'h3cbe7537),
	.w6(32'hbbae782e),
	.w7(32'hbcfe0a31),
	.w8(32'hb9dee2c0),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc72b7ab),
	.w1(32'hbcf04182),
	.w2(32'h3cd7ffee),
	.w3(32'h3c6fd2e0),
	.w4(32'hbce71c32),
	.w5(32'h3c1c3717),
	.w6(32'h3d1ed8f5),
	.w7(32'h3bbb9d13),
	.w8(32'h3cf0efec),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc255f16),
	.w1(32'hb9b231f7),
	.w2(32'h3c1b42f1),
	.w3(32'hbc0debee),
	.w4(32'h3b0f0c75),
	.w5(32'h3b783013),
	.w6(32'h3ae3e233),
	.w7(32'h3cb02a02),
	.w8(32'h3d67da4a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07d63c),
	.w1(32'hbb8c06e6),
	.w2(32'h3c3e43d6),
	.w3(32'h3c6a1b61),
	.w4(32'h3b851eda),
	.w5(32'h3c277ffe),
	.w6(32'h3c4da0e6),
	.w7(32'h3c3ca3a6),
	.w8(32'h3c8ba83d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69cc72),
	.w1(32'hbb10b78e),
	.w2(32'hbc4b4070),
	.w3(32'h3b42f011),
	.w4(32'h3938e2fe),
	.w5(32'h3c0991ee),
	.w6(32'h3aecc11b),
	.w7(32'h3b9b4b90),
	.w8(32'hbc2f90ed),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41c526),
	.w1(32'h3d0930f1),
	.w2(32'h3d4d8d7a),
	.w3(32'h3d20a1bb),
	.w4(32'h3d0b2261),
	.w5(32'h3cdc14db),
	.w6(32'hbc97ceba),
	.w7(32'h3d9ff103),
	.w8(32'h3da09755),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d01cc97),
	.w1(32'h3ca6c844),
	.w2(32'hbad9a9e0),
	.w3(32'hbbfb8ccb),
	.w4(32'hbc177987),
	.w5(32'h3a4118ff),
	.w6(32'hbc5a6ead),
	.w7(32'h3c66df6c),
	.w8(32'hbc620f85),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c121f1f),
	.w1(32'h3cb187bf),
	.w2(32'hbbbadd7e),
	.w3(32'h3c5393cb),
	.w4(32'h3b6efa54),
	.w5(32'hbae333ca),
	.w6(32'hbced9615),
	.w7(32'h3c2aa64a),
	.w8(32'h3b857a09),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3ed60),
	.w1(32'h3bee0e49),
	.w2(32'hbc9283b4),
	.w3(32'h3b8e2f61),
	.w4(32'h3c6cbc9b),
	.w5(32'hbbed51a2),
	.w6(32'h3c0017bf),
	.w7(32'h3c192fc6),
	.w8(32'hbc5430c9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc344cde),
	.w1(32'hbcd8e40a),
	.w2(32'hbc9d57d6),
	.w3(32'h3ca12e76),
	.w4(32'hbc9e0ff8),
	.w5(32'hbc265e42),
	.w6(32'hbca9b607),
	.w7(32'h3c465348),
	.w8(32'h3c5c70e4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3c190),
	.w1(32'h3b9385d6),
	.w2(32'h3c5467ab),
	.w3(32'hb9258a60),
	.w4(32'h3b98e7d0),
	.w5(32'h3c5e802c),
	.w6(32'hbcd68a0c),
	.w7(32'h3b8fe1b9),
	.w8(32'h3891fac3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4e09da),
	.w1(32'h3c62400d),
	.w2(32'hbc9dc88d),
	.w3(32'h3ab9d8c0),
	.w4(32'h3b995f8f),
	.w5(32'h391bbf71),
	.w6(32'h3b2cc498),
	.w7(32'h3bb1970e),
	.w8(32'h3c917c8c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b708c66),
	.w1(32'h3cda02ac),
	.w2(32'h3c767e85),
	.w3(32'h3ccb3a3d),
	.w4(32'hbc83a649),
	.w5(32'h3be9bf6a),
	.w6(32'hb921bd1e),
	.w7(32'h3c3d9954),
	.w8(32'h3cb42b84),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d62a9),
	.w1(32'hbc30308f),
	.w2(32'hb9ab3159),
	.w3(32'h3bf56558),
	.w4(32'hba2776f8),
	.w5(32'h3c71c869),
	.w6(32'h3a550bcc),
	.w7(32'h3b2706bd),
	.w8(32'hbcadf828),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80ff8),
	.w1(32'h3c6b9ade),
	.w2(32'h3cedbd2c),
	.w3(32'h3c0e6a5c),
	.w4(32'h3c5ad209),
	.w5(32'h3c5a43db),
	.w6(32'hb92ef785),
	.w7(32'hbcb5b4b9),
	.w8(32'h3d2f3404),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81a58c),
	.w1(32'hbba7a97f),
	.w2(32'h3c41df0b),
	.w3(32'h3c137ee3),
	.w4(32'h3a7d824d),
	.w5(32'hb9d42a3b),
	.w6(32'h3d5f9a59),
	.w7(32'h3d7239e4),
	.w8(32'h3ca8a727),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c945a6f),
	.w1(32'h3c8016d7),
	.w2(32'h3b7ee1bb),
	.w3(32'h3c07f630),
	.w4(32'hbb9f52c2),
	.w5(32'h3ba93db3),
	.w6(32'hbcc29c72),
	.w7(32'h3c54898f),
	.w8(32'h3be53371),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037948),
	.w1(32'h3a5aa24d),
	.w2(32'hbc232981),
	.w3(32'h3b84e648),
	.w4(32'hbc66c748),
	.w5(32'h3c019295),
	.w6(32'hbc0e17c3),
	.w7(32'hbd27a7f0),
	.w8(32'hbc677603),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0e47f7),
	.w1(32'hbc6ad628),
	.w2(32'hbbd1950e),
	.w3(32'h3cb7886e),
	.w4(32'h3d0aa604),
	.w5(32'h3cf907c8),
	.w6(32'h3d07ffea),
	.w7(32'h3be609c8),
	.w8(32'h3c83f935),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8979fd),
	.w1(32'hbca47eeb),
	.w2(32'hbc7adb4f),
	.w3(32'h3c6d84fc),
	.w4(32'hbc947e42),
	.w5(32'h3c4e94e9),
	.w6(32'hbbb3787f),
	.w7(32'h3c4321c7),
	.w8(32'h3d95cd41),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2f549c),
	.w1(32'hbc836d97),
	.w2(32'hbaafe7a7),
	.w3(32'h3cd4c3e6),
	.w4(32'hbbb9a0df),
	.w5(32'h3c9ef859),
	.w6(32'h3c5ba665),
	.w7(32'h3bc08303),
	.w8(32'hbbe7f153),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c865028),
	.w1(32'hbcb81411),
	.w2(32'h3cbee6ee),
	.w3(32'hbbde759d),
	.w4(32'hbd20c6ac),
	.w5(32'hbc597874),
	.w6(32'hbaa9c62b),
	.w7(32'hbcceba3c),
	.w8(32'hbc19b75c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0d8329),
	.w1(32'hbba675fe),
	.w2(32'hbc88fb2c),
	.w3(32'hbc8a8208),
	.w4(32'hbd01c61d),
	.w5(32'hbc8ec502),
	.w6(32'hba99fbae),
	.w7(32'hbd12fc2a),
	.w8(32'hbd0a55c4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39484e14),
	.w1(32'hbc8f6f08),
	.w2(32'h3c98336f),
	.w3(32'hbcc8f133),
	.w4(32'h3c0c36b3),
	.w5(32'h3caa00bc),
	.w6(32'hbd05cb18),
	.w7(32'hbd141860),
	.w8(32'hbc5928cf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7df9fc),
	.w1(32'hbc8a01bc),
	.w2(32'h3ce98138),
	.w3(32'h3c3bbe54),
	.w4(32'hbca90e01),
	.w5(32'hbc039932),
	.w6(32'h3d95a7cb),
	.w7(32'hbaed23d5),
	.w8(32'h39936563),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae869d),
	.w1(32'h3b898485),
	.w2(32'h3bea8521),
	.w3(32'hbc05dc2b),
	.w4(32'hba39268b),
	.w5(32'h3ca54e40),
	.w6(32'h3c6407b3),
	.w7(32'hbcdf31a9),
	.w8(32'hbc9a3b8b),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ffd12),
	.w1(32'h3b2f966c),
	.w2(32'h3bca1c34),
	.w3(32'h3c10d666),
	.w4(32'h3a696a6f),
	.w5(32'h3c0aea40),
	.w6(32'h3c172443),
	.w7(32'h3bb7f660),
	.w8(32'h3c015cbf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb971c62c),
	.w1(32'h3a56cf68),
	.w2(32'hbc931c8d),
	.w3(32'hb98f78a0),
	.w4(32'hbc6f139f),
	.w5(32'hbc66c658),
	.w6(32'hbb236bc2),
	.w7(32'hbc88c78a),
	.w8(32'hbc9c6d16),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa16460),
	.w1(32'h3c4ada8c),
	.w2(32'hbaffc38e),
	.w3(32'hbc60efc9),
	.w4(32'h3b25c39c),
	.w5(32'h3c48461a),
	.w6(32'h3c314bf6),
	.w7(32'hbb858985),
	.w8(32'hbd0a2a08),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cab0a7e),
	.w1(32'h3b279987),
	.w2(32'h3ba024da),
	.w3(32'hbb92c890),
	.w4(32'hbb716dc6),
	.w5(32'h3b080543),
	.w6(32'h3b8a53f6),
	.w7(32'hbb6a9e0d),
	.w8(32'h3b579ca5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c627d9f),
	.w1(32'h3b84e8f1),
	.w2(32'h3b9013d6),
	.w3(32'h3c9a2a07),
	.w4(32'h3d0d5f53),
	.w5(32'h3cef1206),
	.w6(32'h3bdf0e47),
	.w7(32'h3c139cfd),
	.w8(32'h3ce6b672),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d5f72),
	.w1(32'h38b23282),
	.w2(32'hbb380e0f),
	.w3(32'hbaf12150),
	.w4(32'hbbc9b86e),
	.w5(32'hbb65eda4),
	.w6(32'h3ce09d44),
	.w7(32'h3a8bbdb1),
	.w8(32'hbbd5ca98),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6de812),
	.w1(32'h3b577703),
	.w2(32'h3c12acb3),
	.w3(32'h3c59e9c9),
	.w4(32'h3bfc2110),
	.w5(32'h3ca38fa3),
	.w6(32'h3ab0ea5a),
	.w7(32'hbccfef49),
	.w8(32'hbdb09735),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc06140),
	.w1(32'h3bd5da4f),
	.w2(32'hbc491765),
	.w3(32'h3b2bdd25),
	.w4(32'h3b52e438),
	.w5(32'h3b7e5241),
	.w6(32'hbc72619a),
	.w7(32'hbb960aca),
	.w8(32'h3c23ce0c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0adef0),
	.w1(32'hbc848d29),
	.w2(32'h3c0169cd),
	.w3(32'hbbdf90ba),
	.w4(32'h3b837b20),
	.w5(32'h3bd332f4),
	.w6(32'h3d2c6269),
	.w7(32'h3bba5892),
	.w8(32'h3c11d722),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b882d36),
	.w1(32'hbadd0404),
	.w2(32'h3c5fa8ca),
	.w3(32'h3c92c670),
	.w4(32'hbbf7c00f),
	.w5(32'hbb98f4e9),
	.w6(32'h3c1672af),
	.w7(32'h3a1266b7),
	.w8(32'hbc8f6c0c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc02a99),
	.w1(32'h3a738705),
	.w2(32'hbba03351),
	.w3(32'h3aee175c),
	.w4(32'h398fc885),
	.w5(32'h3b65ce79),
	.w6(32'hbc0041c9),
	.w7(32'h3c911830),
	.w8(32'h3ca4879e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule