module layer_8_featuremap_230(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59378b),
	.w1(32'hbc788775),
	.w2(32'h3d04b5e3),
	.w3(32'hbc25403a),
	.w4(32'hbcacbc21),
	.w5(32'h3c9fb6ff),
	.w6(32'hbc92e57a),
	.w7(32'h3cb6fbe3),
	.w8(32'h3cc351ed),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb0254),
	.w1(32'hba500cc1),
	.w2(32'hbb9e80ed),
	.w3(32'hbb98bf28),
	.w4(32'h3b61d845),
	.w5(32'hbbc218e6),
	.w6(32'hbba8d6c9),
	.w7(32'hbab96d71),
	.w8(32'hbc076a01),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f2b6f),
	.w1(32'h3c431b74),
	.w2(32'h3c351a2b),
	.w3(32'hb9ced057),
	.w4(32'h3bff2121),
	.w5(32'h3c44e976),
	.w6(32'h3c1b83a0),
	.w7(32'h3c1c1814),
	.w8(32'hbbeb2c80),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c4597),
	.w1(32'h3c2fb590),
	.w2(32'hbb83a188),
	.w3(32'hbced1b9a),
	.w4(32'hba4ff110),
	.w5(32'h3b7943f0),
	.w6(32'h3a81616e),
	.w7(32'hbbcf8890),
	.w8(32'hbbe2f8ea),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8d5899),
	.w1(32'hb9ac18c4),
	.w2(32'hbc240d73),
	.w3(32'hbcaf05b9),
	.w4(32'h3b5df7d2),
	.w5(32'hbb902683),
	.w6(32'h3bdca728),
	.w7(32'hbbb873ae),
	.w8(32'hbc058961),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f218),
	.w1(32'hbbb86844),
	.w2(32'hbb5380ac),
	.w3(32'h3bc804e4),
	.w4(32'hbcac2f66),
	.w5(32'hbc7b9c34),
	.w6(32'hbbe90ef2),
	.w7(32'h3b16154a),
	.w8(32'hbcdfce52),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6506f6),
	.w1(32'hbacf4747),
	.w2(32'hbb8adb0f),
	.w3(32'h3b50f8c2),
	.w4(32'hbb4afb0c),
	.w5(32'hbb39efb7),
	.w6(32'hbbe5bd1a),
	.w7(32'hbbc29e3a),
	.w8(32'hbb85c439),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3af482),
	.w1(32'h3c683e98),
	.w2(32'hbc8a8a88),
	.w3(32'hbc303696),
	.w4(32'h3c5c3456),
	.w5(32'hbb93265d),
	.w6(32'hbc1ba9ef),
	.w7(32'hbd0194b7),
	.w8(32'h3bbf1f88),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946f35),
	.w1(32'h3b59be63),
	.w2(32'hbc59d21e),
	.w3(32'h3b94848f),
	.w4(32'h3c2ba49c),
	.w5(32'hbb0d5443),
	.w6(32'hbba91933),
	.w7(32'hbc562848),
	.w8(32'h3a73722d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3849f7),
	.w1(32'h3b1fa5f1),
	.w2(32'h3ccfaac3),
	.w3(32'hbc265824),
	.w4(32'h3c3bdd2a),
	.w5(32'h3cf61f4c),
	.w6(32'hbbdc39b2),
	.w7(32'h3cd5f014),
	.w8(32'hbc4604b9),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc66e86),
	.w1(32'h3cfb3481),
	.w2(32'h3d3abb35),
	.w3(32'hbcc385be),
	.w4(32'h3b384cdc),
	.w5(32'h3d038641),
	.w6(32'h3c0942fd),
	.w7(32'h3c48387e),
	.w8(32'h3bea6d48),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9f3d9),
	.w1(32'hbbe8d7e5),
	.w2(32'h3c86fb40),
	.w3(32'hbca06f50),
	.w4(32'hbba03bdf),
	.w5(32'h3b9e362f),
	.w6(32'hb9186c66),
	.w7(32'h3c554b9d),
	.w8(32'hbbd25d04),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedec07),
	.w1(32'hbc4b9c74),
	.w2(32'h3b895324),
	.w3(32'h394edb36),
	.w4(32'hb9d1f28b),
	.w5(32'hbb0bab87),
	.w6(32'hbb9a3803),
	.w7(32'hb936f8a6),
	.w8(32'hbb9a428a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae16623),
	.w1(32'h3b5ba1e8),
	.w2(32'h3aa61a4c),
	.w3(32'hbb760bb5),
	.w4(32'hba93e81e),
	.w5(32'hba4f9449),
	.w6(32'h3c2f0386),
	.w7(32'h3bf2c507),
	.w8(32'hbc303a5a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb010a7),
	.w1(32'hba34f0ed),
	.w2(32'h398ea7a5),
	.w3(32'hbc5cc86b),
	.w4(32'h3ad46105),
	.w5(32'h3ba509b8),
	.w6(32'hbc0d1d18),
	.w7(32'hbb98923a),
	.w8(32'hbb119934),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d135a),
	.w1(32'hbc28f158),
	.w2(32'h3cfd01a3),
	.w3(32'h3b5aa5e9),
	.w4(32'hbc8ef8e6),
	.w5(32'h3cc0abd5),
	.w6(32'hbbec54ca),
	.w7(32'h3d025b96),
	.w8(32'h3cce0bf3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cefbcad),
	.w1(32'hbc7f852b),
	.w2(32'h3b2b8470),
	.w3(32'h3c94eb43),
	.w4(32'hbc24f656),
	.w5(32'hba2cfad8),
	.w6(32'hbb744058),
	.w7(32'hbc0d47cb),
	.w8(32'hb9c00f51),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd99ad5),
	.w1(32'h3b803b34),
	.w2(32'h3c5a7460),
	.w3(32'hbc765573),
	.w4(32'hbb91875e),
	.w5(32'h39d94292),
	.w6(32'hbc134551),
	.w7(32'h3c29b330),
	.w8(32'h3ba59d4e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd03c2d5),
	.w1(32'hbccfc0ba),
	.w2(32'h3dd2032b),
	.w3(32'hbd1d13a6),
	.w4(32'hbd8fc4e4),
	.w5(32'h3d867271),
	.w6(32'hbcd3304c),
	.w7(32'h3d8c3b52),
	.w8(32'h3da79c58),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc30149),
	.w1(32'hbc461ce9),
	.w2(32'hbbe6cc9a),
	.w3(32'h3bc12827),
	.w4(32'h3a93b6a9),
	.w5(32'h398381c6),
	.w6(32'hbc4215f2),
	.w7(32'hbbf12fc8),
	.w8(32'hbc9dc1e9),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a1c3e),
	.w1(32'hbc29479c),
	.w2(32'hbc47f169),
	.w3(32'h3c1041a0),
	.w4(32'hbc4494c0),
	.w5(32'hbc7c1fef),
	.w6(32'h3c34d1a1),
	.w7(32'hbc4fdac6),
	.w8(32'hbc80e7f8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5c2d),
	.w1(32'hbc24de7e),
	.w2(32'hbc17f9b9),
	.w3(32'h3aafc0c0),
	.w4(32'hbc473aef),
	.w5(32'hbc8a776e),
	.w6(32'hbc21dcff),
	.w7(32'h3aab559a),
	.w8(32'hbc520a8d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd28a977),
	.w1(32'h3cb3bd73),
	.w2(32'h3db8a19e),
	.w3(32'hbd20f4aa),
	.w4(32'hbbfd28f3),
	.w5(32'h3d7638db),
	.w6(32'hbc5264be),
	.w7(32'h3cf7dcdc),
	.w8(32'h3d081eca),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc570a7),
	.w1(32'hbb9d3288),
	.w2(32'hbc33270e),
	.w3(32'hbca8b1a5),
	.w4(32'h3b8e71e9),
	.w5(32'hbc5f56ba),
	.w6(32'h3aa20143),
	.w7(32'hbbf0f769),
	.w8(32'hbca70614),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36fb77),
	.w1(32'h3bcbb6bf),
	.w2(32'h3c0ef8ab),
	.w3(32'hbc42d533),
	.w4(32'hbb198786),
	.w5(32'h3b632b05),
	.w6(32'h3c0c9c28),
	.w7(32'h3aa611b5),
	.w8(32'hbc62f046),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd97ee6),
	.w1(32'hbb33213c),
	.w2(32'hbba843b8),
	.w3(32'hbcc14d82),
	.w4(32'hbca13795),
	.w5(32'hbc5135c4),
	.w6(32'hbc763065),
	.w7(32'h3ba57a5c),
	.w8(32'hbc46d0fb),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbefe4df),
	.w1(32'h3ba5af79),
	.w2(32'h3c4f8cb7),
	.w3(32'hbc1bd96e),
	.w4(32'hbb82ee8f),
	.w5(32'h3baab131),
	.w6(32'hbb7bc1c8),
	.w7(32'h3c5eb6a1),
	.w8(32'hbb7d68f3),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe2f563f),
	.w1(32'h3d8b4927),
	.w2(32'h3d92d195),
	.w3(32'hbd82e6ca),
	.w4(32'h3c9fe2ce),
	.w5(32'hbe037520),
	.w6(32'hbe00a200),
	.w7(32'hbd45b5f6),
	.w8(32'h3db1370c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09f003),
	.w1(32'hbbb55fff),
	.w2(32'h3c5a1316),
	.w3(32'hbc880fb7),
	.w4(32'hbc0a4730),
	.w5(32'h3b9c0705),
	.w6(32'hbcc349b1),
	.w7(32'hbba18e53),
	.w8(32'h3c35ad49),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd222d9),
	.w1(32'h3b895bba),
	.w2(32'h39a9839b),
	.w3(32'h3bf59b0c),
	.w4(32'h3c7fe28a),
	.w5(32'h3ca69ffe),
	.w6(32'hbaf48e44),
	.w7(32'hb8c50e86),
	.w8(32'h3c93533d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ad9cd),
	.w1(32'h3c14a2e0),
	.w2(32'h3b93a1e8),
	.w3(32'h3d03916f),
	.w4(32'h3a09f55b),
	.w5(32'h3929856d),
	.w6(32'hbbcb12c6),
	.w7(32'hbc0aa47b),
	.w8(32'hbbaf5bc4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12c987),
	.w1(32'hbcbce5e9),
	.w2(32'hbc6fd43d),
	.w3(32'h3b78fb68),
	.w4(32'hbbd37745),
	.w5(32'hbc2253b9),
	.w6(32'hbbf18d50),
	.w7(32'hbbd9cc53),
	.w8(32'hbcb58fe7),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5919e3),
	.w1(32'h3bbe869f),
	.w2(32'h3c4e3d1a),
	.w3(32'h3a8379e4),
	.w4(32'hbb820c3a),
	.w5(32'hbb90823c),
	.w6(32'h3c071422),
	.w7(32'h3c864d63),
	.w8(32'hbbf55111),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc64e796),
	.w1(32'h3c026a5d),
	.w2(32'h398dff8d),
	.w3(32'hbc868fd5),
	.w4(32'h3bf45efc),
	.w5(32'h3a1cf8c6),
	.w6(32'h3b53b116),
	.w7(32'h3ba0aa72),
	.w8(32'h3ba86b6a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb659dd4),
	.w1(32'hbbeed4cd),
	.w2(32'hbca7b52a),
	.w3(32'h3c192ee8),
	.w4(32'h3c5975f4),
	.w5(32'h39a6b850),
	.w6(32'h3aaaed92),
	.w7(32'hbb6cdf76),
	.w8(32'hbb8b7062),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3d2aa),
	.w1(32'hbc2e3bfa),
	.w2(32'h3c6e3203),
	.w3(32'hbc8d2323),
	.w4(32'hbc77cb59),
	.w5(32'h3c0967de),
	.w6(32'hbc977370),
	.w7(32'hbad7274c),
	.w8(32'h3acad7b2),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae44484),
	.w1(32'h3c098a91),
	.w2(32'hbbef07b9),
	.w3(32'hbc3307e4),
	.w4(32'h3c2396e1),
	.w5(32'hbb24c10e),
	.w6(32'h3b66a91a),
	.w7(32'hbc1952b0),
	.w8(32'hbc1abf5b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2705c2),
	.w1(32'h3a2dd54b),
	.w2(32'hbbd20425),
	.w3(32'hbbb9f9af),
	.w4(32'h3b919353),
	.w5(32'h3a0d8336),
	.w6(32'hbc23ef63),
	.w7(32'hbc0dce7f),
	.w8(32'hbb57adeb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4b4a),
	.w1(32'hbcb248fd),
	.w2(32'hbc112c1a),
	.w3(32'h3ba9a8ea),
	.w4(32'hbc7fb68b),
	.w5(32'hbc37f482),
	.w6(32'hbc08db43),
	.w7(32'hbc55ca24),
	.w8(32'hbbfb75d4),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32ace8),
	.w1(32'h3b5e9715),
	.w2(32'h3bb47d0d),
	.w3(32'hbbfbc164),
	.w4(32'hbbc37a11),
	.w5(32'h3aee0b38),
	.w6(32'h3b9da487),
	.w7(32'hb9b67927),
	.w8(32'h3968c73a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e3b27),
	.w1(32'hbc9db189),
	.w2(32'hbcb45840),
	.w3(32'hbd69fd7f),
	.w4(32'hbbf3667c),
	.w5(32'hbc926a1d),
	.w6(32'hbd10154a),
	.w7(32'hbbaa0a98),
	.w8(32'hbd07306b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc126158),
	.w1(32'hbc5ce327),
	.w2(32'h3c4c45b9),
	.w3(32'hbbf0bc42),
	.w4(32'hbc7c652d),
	.w5(32'h3c0397ed),
	.w6(32'hbc896163),
	.w7(32'hbb693a27),
	.w8(32'hbb8e9445),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a700),
	.w1(32'h3c7189cb),
	.w2(32'hbb6fba8b),
	.w3(32'h3a41cfa9),
	.w4(32'h3c24aae7),
	.w5(32'hbb915831),
	.w6(32'h3c47a6db),
	.w7(32'hbb4a1092),
	.w8(32'hbc5ac3dc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceeb94d),
	.w1(32'hbbed0525),
	.w2(32'h3c74c669),
	.w3(32'hbca9b65b),
	.w4(32'hbc648751),
	.w5(32'h39512774),
	.w6(32'hbc8740b2),
	.w7(32'h3a9c8267),
	.w8(32'hbb15136f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc71cf27),
	.w1(32'h3c023117),
	.w2(32'h3d0aceec),
	.w3(32'hbc4e6592),
	.w4(32'hbc21cd89),
	.w5(32'h3d0dc11c),
	.w6(32'hba1d4fcd),
	.w7(32'h3cc3c986),
	.w8(32'h3cc06b5a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcceec64),
	.w1(32'hbc053f45),
	.w2(32'h3c57e5fc),
	.w3(32'hbc68a9cf),
	.w4(32'hbc00fc05),
	.w5(32'h3ca3918e),
	.w6(32'hbbcc8a59),
	.w7(32'h3c012942),
	.w8(32'h3c87cce3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4de1a),
	.w1(32'hba3d6300),
	.w2(32'h3c2da189),
	.w3(32'h3bc251d0),
	.w4(32'hbb53b2f2),
	.w5(32'h3bb1aa9d),
	.w6(32'hbb8cda59),
	.w7(32'h3b71924c),
	.w8(32'hbbc0c684),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0a96b),
	.w1(32'hbc7112bf),
	.w2(32'h3cce791b),
	.w3(32'hbc4ab3be),
	.w4(32'hbcb779f4),
	.w5(32'h3b5c7da2),
	.w6(32'hb9aaa5cf),
	.w7(32'h3c574864),
	.w8(32'h3c96300d),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a8ad2),
	.w1(32'h3bf9d2c9),
	.w2(32'h3c21aef0),
	.w3(32'hbc111911),
	.w4(32'hbb347b1f),
	.w5(32'hb77c1ed3),
	.w6(32'hbba458c4),
	.w7(32'h3bc36971),
	.w8(32'hbbabae61),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb959efc),
	.w1(32'hbaf526c0),
	.w2(32'h3d19099a),
	.w3(32'hbcb479b3),
	.w4(32'hbccf258c),
	.w5(32'h3c8c65f9),
	.w6(32'h3ab4ecb7),
	.w7(32'h3cd25cc0),
	.w8(32'h3c0ca499),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca77407),
	.w1(32'h3c04ed8f),
	.w2(32'hbcd59084),
	.w3(32'h3c6aa066),
	.w4(32'h3bf2ac4f),
	.w5(32'hbd1cc084),
	.w6(32'h3c8051b1),
	.w7(32'h3b818824),
	.w8(32'hbcdff63c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a870e9a),
	.w1(32'h3b48e61c),
	.w2(32'h3d11fc8c),
	.w3(32'hbd08581f),
	.w4(32'hbcd3ee46),
	.w5(32'h3cff9e78),
	.w6(32'hbd1a0227),
	.w7(32'hbbe11c8a),
	.w8(32'h3d122dbe),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a3ef8),
	.w1(32'h3b6633ae),
	.w2(32'h3b61d694),
	.w3(32'hbc024c55),
	.w4(32'h3a8b4010),
	.w5(32'h3c0ae74c),
	.w6(32'h3aa72b89),
	.w7(32'hbbdfee1d),
	.w8(32'h3b3142a0),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc379698),
	.w1(32'hbc837d85),
	.w2(32'hbc5d3b77),
	.w3(32'hbc142d84),
	.w4(32'h3bb97c1e),
	.w5(32'h3caac51c),
	.w6(32'hbbe4320c),
	.w7(32'hbbff4808),
	.w8(32'h3ce89e20),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd87555),
	.w1(32'h3c1feb0c),
	.w2(32'h3c368464),
	.w3(32'h3b194c1a),
	.w4(32'hbb12f705),
	.w5(32'h3ab18bf1),
	.w6(32'h3ba659f2),
	.w7(32'h3c0d5dc4),
	.w8(32'h3be5f337),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c1260),
	.w1(32'hbd29bb7e),
	.w2(32'h3c125bc4),
	.w3(32'hbcea2438),
	.w4(32'hbc9ecf0b),
	.w5(32'h3b2a3f46),
	.w6(32'hbcb1310c),
	.w7(32'h3c8f3ed1),
	.w8(32'h3d181bbe),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b77963),
	.w1(32'h3cca063a),
	.w2(32'hbaf04475),
	.w3(32'hbb964f7f),
	.w4(32'h3c8a4711),
	.w5(32'h3ad8d318),
	.w6(32'h3b91a20b),
	.w7(32'hbb5eac72),
	.w8(32'hbaa7f57f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafe699),
	.w1(32'h3c771f77),
	.w2(32'h3aee9d72),
	.w3(32'hbd007eba),
	.w4(32'hbbd511c3),
	.w5(32'h3a718e4d),
	.w6(32'hbc697758),
	.w7(32'hbc29f5e1),
	.w8(32'h3b8636f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc92022f),
	.w1(32'hbb9bd335),
	.w2(32'h3c2dbf2e),
	.w3(32'hbca7a780),
	.w4(32'hbc522ad0),
	.w5(32'hb9dfeb22),
	.w6(32'hbb980267),
	.w7(32'hbbee83da),
	.w8(32'h3bfe6226),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7a36c),
	.w1(32'h3b06bf8f),
	.w2(32'hbbb06cf8),
	.w3(32'hbb310935),
	.w4(32'hbc6e5968),
	.w5(32'hbc669e3e),
	.w6(32'hbbd503e2),
	.w7(32'hbc272f22),
	.w8(32'hbc8d3a85),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9431ba),
	.w1(32'h3c1dd2b1),
	.w2(32'h3c8391ee),
	.w3(32'hbc1e28bc),
	.w4(32'hbc06c0f2),
	.w5(32'h3b963ae6),
	.w6(32'h3bdb11bb),
	.w7(32'h3c3a89ec),
	.w8(32'hb926957c),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d5581),
	.w1(32'h3a848f72),
	.w2(32'h3b234ffc),
	.w3(32'hbbcf7919),
	.w4(32'hbb26b7b4),
	.w5(32'h3c57898e),
	.w6(32'h3b916b17),
	.w7(32'hbba2bc61),
	.w8(32'hbbcc280e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7125e9),
	.w1(32'hbbb00bf6),
	.w2(32'hbc4dfcbd),
	.w3(32'hbc8bff32),
	.w4(32'h3c5d5ab1),
	.w5(32'h3c6f5cd6),
	.w6(32'hbc70ea2a),
	.w7(32'hbb554212),
	.w8(32'h3a01badd),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3a0d34),
	.w1(32'h3c18ce74),
	.w2(32'h3c1497f0),
	.w3(32'h3cace64d),
	.w4(32'h3c04e077),
	.w5(32'h3bba63cb),
	.w6(32'h3b6296f0),
	.w7(32'h3b8e0ca0),
	.w8(32'h3b98ec00),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b213d7b),
	.w1(32'hba09dfc4),
	.w2(32'h3bdaaa87),
	.w3(32'h3b5c2a98),
	.w4(32'hbb4bd6d7),
	.w5(32'h3aaf4e88),
	.w6(32'hbb7d8ffd),
	.w7(32'hba4d286d),
	.w8(32'hbb9ab67f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeec8d3),
	.w1(32'h3c3633eb),
	.w2(32'h3c82059d),
	.w3(32'hbbbc86ab),
	.w4(32'hbb4c4593),
	.w5(32'hb8e79ec9),
	.w6(32'h3b0ebba3),
	.w7(32'hb9f4d3ee),
	.w8(32'hbbd373b4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeccc17),
	.w1(32'h3b9bfa87),
	.w2(32'h3c596b96),
	.w3(32'hbc009b75),
	.w4(32'hbc2a947a),
	.w5(32'h3cd9393b),
	.w6(32'h3c1cad5e),
	.w7(32'h3bdcd9c5),
	.w8(32'hbc499193),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f7adc),
	.w1(32'hbc4b1cc3),
	.w2(32'hb8e7bc9a),
	.w3(32'hbbe518ea),
	.w4(32'hbc134244),
	.w5(32'h3b55a2e5),
	.w6(32'h3bb45597),
	.w7(32'h3c2fafe0),
	.w8(32'h3b447b41),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe700ed),
	.w1(32'h3824c606),
	.w2(32'hbc266631),
	.w3(32'h3b045762),
	.w4(32'hbba20d05),
	.w5(32'hbc30b4f2),
	.w6(32'h3bcaae10),
	.w7(32'hbb195538),
	.w8(32'hbc9e66c3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd214bbd),
	.w1(32'h3c096a50),
	.w2(32'h3d1e98ee),
	.w3(32'hbca5bd58),
	.w4(32'hbd225004),
	.w5(32'h3b0776e0),
	.w6(32'hbceb99d0),
	.w7(32'hbc003385),
	.w8(32'h3cfa5180),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96f800),
	.w1(32'hbc64fbf1),
	.w2(32'hbb46bed3),
	.w3(32'hbc8990bf),
	.w4(32'hbbf03ad1),
	.w5(32'hbaf95b3e),
	.w6(32'hbc13213f),
	.w7(32'h3aba39c6),
	.w8(32'h3c6eeb52),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cce78e6),
	.w1(32'h3b2b40ef),
	.w2(32'hbbf5d5a1),
	.w3(32'h3c879e5c),
	.w4(32'hbbd6aa70),
	.w5(32'h3a1570b2),
	.w6(32'h3a9e0190),
	.w7(32'hbbe288bc),
	.w8(32'hbcde586b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccae0e8),
	.w1(32'hbb08ba30),
	.w2(32'h3b3f7faf),
	.w3(32'hbc4827cf),
	.w4(32'hbbdd20b0),
	.w5(32'hbb28f503),
	.w6(32'hbb4231a0),
	.w7(32'hbbad45cb),
	.w8(32'hbc568658),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd003597),
	.w1(32'h3bc54837),
	.w2(32'h3c098ca2),
	.w3(32'hbc6aaed2),
	.w4(32'h3c2f8279),
	.w5(32'h3b8249d5),
	.w6(32'hbb9dcf41),
	.w7(32'h3bb66290),
	.w8(32'hbbf7b867),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4276),
	.w1(32'hbc230c25),
	.w2(32'h3bac86c8),
	.w3(32'hbbd0e8e8),
	.w4(32'hbc771460),
	.w5(32'hbbcd5b87),
	.w6(32'hbc2925eb),
	.w7(32'h3a3b48f3),
	.w8(32'hbbc5bca1),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5517ed),
	.w1(32'h3cc3f206),
	.w2(32'h3cf25888),
	.w3(32'hbc01736d),
	.w4(32'h394b8efe),
	.w5(32'h3c2ffa74),
	.w6(32'h3be3bcd6),
	.w7(32'h3c0c614d),
	.w8(32'h3c56b53a),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd58158),
	.w1(32'h3bd6bf1a),
	.w2(32'hbb740a99),
	.w3(32'h3c50350b),
	.w4(32'hbb12772a),
	.w5(32'hbc25d9f3),
	.w6(32'h3b79df62),
	.w7(32'hbbdc82e6),
	.w8(32'hbb95f822),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc994db8),
	.w1(32'h3cc17ec9),
	.w2(32'h3cc60c2a),
	.w3(32'hbc6a2b48),
	.w4(32'hbb8f5b85),
	.w5(32'h3a1b3ec1),
	.w6(32'h399d7bc4),
	.w7(32'h3bb63d75),
	.w8(32'h3c3e2e05),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca3652a),
	.w1(32'hbc55871b),
	.w2(32'h3c3c68e7),
	.w3(32'hbcb315af),
	.w4(32'hbc709a62),
	.w5(32'h3c1bf830),
	.w6(32'hbc8938d0),
	.w7(32'h3c3acf8a),
	.w8(32'h3ce88b62),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13291e),
	.w1(32'hbc11d958),
	.w2(32'h3b777bb1),
	.w3(32'hbbf2d401),
	.w4(32'hbbecd2cf),
	.w5(32'hbc174330),
	.w6(32'hbc14dbc5),
	.w7(32'h3c1be5f1),
	.w8(32'hbaee37ae),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0c004),
	.w1(32'h3841ad44),
	.w2(32'h39bcfbaf),
	.w3(32'hbc66ae2e),
	.w4(32'h3b35f848),
	.w5(32'hbb43ec76),
	.w6(32'h3bbefdb8),
	.w7(32'hb9d3d818),
	.w8(32'hbc52bcf1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ee293),
	.w1(32'h3b2090f5),
	.w2(32'hbab24abf),
	.w3(32'hbc9a3415),
	.w4(32'h3bd8ac19),
	.w5(32'hbb826e72),
	.w6(32'hbbade330),
	.w7(32'hbc9153ef),
	.w8(32'hbc2eb17d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc47074),
	.w1(32'hbb0f3951),
	.w2(32'h3cd069ed),
	.w3(32'hbce475ec),
	.w4(32'hbbc43d6b),
	.w5(32'h3cbf50dc),
	.w6(32'hbc4a6e8b),
	.w7(32'h3c0db412),
	.w8(32'hbbbd560e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51555b),
	.w1(32'hbcb7ef25),
	.w2(32'hbd78bc65),
	.w3(32'hbd1a1ca2),
	.w4(32'hbc77ae98),
	.w5(32'hbd0200cc),
	.w6(32'hbc4b6c0f),
	.w7(32'h3bda5c1b),
	.w8(32'hbd1fac9b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bf95c),
	.w1(32'hba581f8f),
	.w2(32'h3cb0c9cc),
	.w3(32'hbcffb1a7),
	.w4(32'hbcca1c45),
	.w5(32'h3c68a000),
	.w6(32'hbc0880a2),
	.w7(32'h3c5add33),
	.w8(32'h3be6be9f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc562f70),
	.w1(32'h3c819ed0),
	.w2(32'h3c1c79d7),
	.w3(32'hbcc47ce6),
	.w4(32'hbc0009de),
	.w5(32'h3c0df7e1),
	.w6(32'hbc3d2f17),
	.w7(32'hbc36b7b2),
	.w8(32'hbb9d4a5a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7ebd3),
	.w1(32'hbbe6b56d),
	.w2(32'hbb042912),
	.w3(32'h3b31433c),
	.w4(32'hbb81d4c1),
	.w5(32'h3b330a46),
	.w6(32'hbb1dce36),
	.w7(32'h3b88b9fb),
	.w8(32'h3c0d4e59),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8e501),
	.w1(32'hbad53b2f),
	.w2(32'h3bb064f1),
	.w3(32'h3c0a8c39),
	.w4(32'hbaa1968a),
	.w5(32'h3b1d0f15),
	.w6(32'hbb125436),
	.w7(32'h3ada38f5),
	.w8(32'hbb45e545),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5ef87),
	.w1(32'hba59b56b),
	.w2(32'hbbd4317f),
	.w3(32'h39a32491),
	.w4(32'hb95d8671),
	.w5(32'hb9c29512),
	.w6(32'hbb24fb80),
	.w7(32'hba9b66b0),
	.w8(32'hbb19726b),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20e566),
	.w1(32'h3c0c5619),
	.w2(32'h3cea9e03),
	.w3(32'hbbe4ef01),
	.w4(32'h3c036df6),
	.w5(32'h3c8f404b),
	.w6(32'h3c2ba445),
	.w7(32'h3c50b9fb),
	.w8(32'hbc0cc367),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb513a3),
	.w1(32'hbb6156d5),
	.w2(32'hbb9abcd7),
	.w3(32'hbc91746a),
	.w4(32'hbc228962),
	.w5(32'hbba57b59),
	.w6(32'hbb4104a0),
	.w7(32'hbc1e920b),
	.w8(32'hbc9ec880),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c9d6a),
	.w1(32'h3c4eb2c3),
	.w2(32'h3c6252e6),
	.w3(32'hbbb33abc),
	.w4(32'h3be23db4),
	.w5(32'h3c38d614),
	.w6(32'h3aa122ec),
	.w7(32'h3bf376fd),
	.w8(32'h3b1baa9c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c820d80),
	.w1(32'h3b866c8e),
	.w2(32'hbc5652e8),
	.w3(32'hba4d041f),
	.w4(32'hb9adaf70),
	.w5(32'hbbda39b1),
	.w6(32'hbbf4d2dd),
	.w7(32'hbbc732ee),
	.w8(32'hbba52092),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa65c4),
	.w1(32'hbac38725),
	.w2(32'h3bb99b0b),
	.w3(32'hbc2eacab),
	.w4(32'hbbb87c0b),
	.w5(32'h3b18954d),
	.w6(32'hbbbe33e1),
	.w7(32'h3b3e5b8a),
	.w8(32'hba19c42e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc250eb9),
	.w1(32'h3c06d508),
	.w2(32'h3c68e175),
	.w3(32'hbbee50fc),
	.w4(32'h3b884ae9),
	.w5(32'h3bdc8df0),
	.w6(32'h3bf99be0),
	.w7(32'h3c38c93e),
	.w8(32'h3b8bba1b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af86f6e),
	.w1(32'hbba99450),
	.w2(32'hbc6bc7e5),
	.w3(32'hbbcbe01e),
	.w4(32'hbbd24f7e),
	.w5(32'hbbf97279),
	.w6(32'h3ae5d1eb),
	.w7(32'hbc89cc91),
	.w8(32'h3b9af00b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c1d2b),
	.w1(32'h3be9bb26),
	.w2(32'h3c8288e2),
	.w3(32'hbcda46dc),
	.w4(32'hbb6c4dcf),
	.w5(32'h3c046b5e),
	.w6(32'hbc779fa4),
	.w7(32'hbb8a9529),
	.w8(32'hbc97cf01),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0f6f2),
	.w1(32'hb87d97b2),
	.w2(32'h3cbe8787),
	.w3(32'hbc59dfe0),
	.w4(32'hbc661ec3),
	.w5(32'h3b01521a),
	.w6(32'h3b308ebd),
	.w7(32'h3c700a3e),
	.w8(32'h3bdd33ed),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27f352),
	.w1(32'hbc391955),
	.w2(32'h3bd379b4),
	.w3(32'hbbb34352),
	.w4(32'hbc2c7cc9),
	.w5(32'hbc8092c1),
	.w6(32'hbb8d4980),
	.w7(32'h3bc9afcb),
	.w8(32'hb933f504),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13db51),
	.w1(32'h3cd3b791),
	.w2(32'h3c22502c),
	.w3(32'hbbbd98c3),
	.w4(32'h3c592c02),
	.w5(32'hbb8367cc),
	.w6(32'h3d03d830),
	.w7(32'h3bb5295a),
	.w8(32'hbca7ce11),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf62196),
	.w1(32'h3c2a9a43),
	.w2(32'h3b4d52b4),
	.w3(32'hbcd8f2ba),
	.w4(32'h3c9039cd),
	.w5(32'h3c13a942),
	.w6(32'h3bf59a10),
	.w7(32'hbb29c94a),
	.w8(32'hbb9f26fa),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4cad),
	.w1(32'hbb866db2),
	.w2(32'hbc698e4c),
	.w3(32'hbc5db9a2),
	.w4(32'hbb213b9f),
	.w5(32'hbc5d7763),
	.w6(32'hbb3f34af),
	.w7(32'hbc01a3f3),
	.w8(32'h3bee6ae1),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53278e),
	.w1(32'hba019006),
	.w2(32'h3c3545c4),
	.w3(32'h3b8ad37c),
	.w4(32'hbbc738fb),
	.w5(32'h3bcc9f46),
	.w6(32'h3b7b3ba5),
	.w7(32'h3bc07dd7),
	.w8(32'hbb243ba1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a868909),
	.w1(32'h3c557eb4),
	.w2(32'hbc550ebc),
	.w3(32'h3b8b8699),
	.w4(32'h3bf187c9),
	.w5(32'hbc3e0bb5),
	.w6(32'h3c7965e3),
	.w7(32'hbbb1edd6),
	.w8(32'hbc95585e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02aff8),
	.w1(32'hbbb060b3),
	.w2(32'h3c0ec502),
	.w3(32'hbc198044),
	.w4(32'hbbc6f9e1),
	.w5(32'hbc7be2a9),
	.w6(32'hbaa1cdb7),
	.w7(32'h3b98c524),
	.w8(32'hbc30533e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7beb5),
	.w1(32'h3bb381f4),
	.w2(32'h3ca50032),
	.w3(32'hbc6638ae),
	.w4(32'hbc78d587),
	.w5(32'h3c09d66b),
	.w6(32'hbc761763),
	.w7(32'hbae5852f),
	.w8(32'h3c92db7b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e0c9d),
	.w1(32'h3c0e8b99),
	.w2(32'hbadf9712),
	.w3(32'h3baaf70e),
	.w4(32'hbac11b38),
	.w5(32'hbb924434),
	.w6(32'h3bba9c22),
	.w7(32'h39a90baa),
	.w8(32'hbc63a8dc),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51dbe9),
	.w1(32'h3c8edd41),
	.w2(32'hbc1feb9d),
	.w3(32'hbc49c99d),
	.w4(32'h3c518682),
	.w5(32'hbbe8afbc),
	.w6(32'h3c7d86eb),
	.w7(32'hbc0e6cb7),
	.w8(32'hbca61ef0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc990a8c),
	.w1(32'h3bcd11d8),
	.w2(32'hbc1bdbf9),
	.w3(32'hbba9094e),
	.w4(32'h3c3cdee8),
	.w5(32'h3bac76df),
	.w6(32'h3c0d8639),
	.w7(32'hbb5a4b6d),
	.w8(32'h3b5d0e88),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b868554),
	.w1(32'h3c032dd9),
	.w2(32'h3bb0132e),
	.w3(32'h3c4dcfb4),
	.w4(32'h3b55cd49),
	.w5(32'h3c003786),
	.w6(32'hbb4c066f),
	.w7(32'hbba3939d),
	.w8(32'hba1b3995),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9efec),
	.w1(32'hbb50624c),
	.w2(32'hba352d90),
	.w3(32'hbb72c911),
	.w4(32'hbb34f78a),
	.w5(32'hbb2cf506),
	.w6(32'h3b8817b1),
	.w7(32'h3aa5acf6),
	.w8(32'hbbe4ca0c),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc239571),
	.w1(32'hba8d5f8c),
	.w2(32'hbb9915af),
	.w3(32'hbc11d130),
	.w4(32'hbbc1d0c5),
	.w5(32'hbc51b668),
	.w6(32'h3aa871e2),
	.w7(32'h3b43197b),
	.w8(32'hbc4b7e0a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b543a8b),
	.w1(32'h3bc8393f),
	.w2(32'h376aa088),
	.w3(32'h3be64029),
	.w4(32'h3c014659),
	.w5(32'h3b253625),
	.w6(32'hba942743),
	.w7(32'h3ba5d2fd),
	.w8(32'h3b842e4e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf5a61),
	.w1(32'h3ad93b19),
	.w2(32'h3a80b651),
	.w3(32'hbb2bdf64),
	.w4(32'hbbade005),
	.w5(32'hbc1d376d),
	.w6(32'h3c198c67),
	.w7(32'h3bdde7d4),
	.w8(32'hbc3b332e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc78cb02),
	.w1(32'hbc56f3ce),
	.w2(32'hbba80f4c),
	.w3(32'hbc8c723a),
	.w4(32'hbc03a0db),
	.w5(32'h3ac0ca44),
	.w6(32'hbc4d5728),
	.w7(32'hbb6b19a4),
	.w8(32'h3aa98161),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4c6b2),
	.w1(32'hbaeafb8c),
	.w2(32'hb9e04d2f),
	.w3(32'h3ba047a3),
	.w4(32'hbb4d821f),
	.w5(32'hbb0ae52f),
	.w6(32'hbb974b16),
	.w7(32'hbbc6c1cf),
	.w8(32'hbbca8082),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49c6f8),
	.w1(32'h3ab5dbde),
	.w2(32'h3bb2a3c6),
	.w3(32'hbaf509f0),
	.w4(32'h3b4a48c1),
	.w5(32'h3be69edb),
	.w6(32'hbab3e1b2),
	.w7(32'hbb1cdee2),
	.w8(32'h3be3d585),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7cb76),
	.w1(32'hbbbab2a8),
	.w2(32'h3b60c3eb),
	.w3(32'h3be9f567),
	.w4(32'hbc32e3d7),
	.w5(32'hbb232329),
	.w6(32'hbc92068d),
	.w7(32'hbb2b9ca8),
	.w8(32'h3c28fe96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c1837),
	.w1(32'hbb0a5e58),
	.w2(32'h3c48517a),
	.w3(32'hbac21a02),
	.w4(32'hbc490077),
	.w5(32'hbb6c8484),
	.w6(32'h3b86193d),
	.w7(32'h3c34babd),
	.w8(32'h389bc375),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc755744),
	.w1(32'hbc1f5a67),
	.w2(32'hb8de8f82),
	.w3(32'hbc942a28),
	.w4(32'hbc317a1a),
	.w5(32'hbbfa8149),
	.w6(32'hbbfe851e),
	.w7(32'hbb92a1c8),
	.w8(32'hbb95955f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba037d0),
	.w1(32'hbb9242c7),
	.w2(32'hbb3bbdbe),
	.w3(32'hbc2e10ef),
	.w4(32'h3bfeedbd),
	.w5(32'h3c43512c),
	.w6(32'hbb8384b3),
	.w7(32'hbbd2964b),
	.w8(32'h3b9984dc),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d7c14),
	.w1(32'h3b5a69e4),
	.w2(32'h3c9ced83),
	.w3(32'hbc930427),
	.w4(32'h3bb72968),
	.w5(32'h3c120d27),
	.w6(32'hbae3fc00),
	.w7(32'h3c4c48c2),
	.w8(32'hbc42ff01),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc423b90),
	.w1(32'h3b258702),
	.w2(32'h3ad95f8c),
	.w3(32'hbc378590),
	.w4(32'h3b8529de),
	.w5(32'h3ab40afe),
	.w6(32'h3b8a21ad),
	.w7(32'h3b7d0be8),
	.w8(32'hbb120de0),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c1b68),
	.w1(32'h3a9bcf50),
	.w2(32'hbb837d75),
	.w3(32'h3b0f5713),
	.w4(32'hbb80f6db),
	.w5(32'hbb4f144c),
	.w6(32'hbaf6a83e),
	.w7(32'h3aa226c0),
	.w8(32'h3b17c6e9),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae0c259),
	.w1(32'h3bda513f),
	.w2(32'h3abce5e7),
	.w3(32'hbb9987c7),
	.w4(32'h3c0e27cf),
	.w5(32'hbb42620d),
	.w6(32'h3c1514fc),
	.w7(32'h3b69c156),
	.w8(32'hbc60c9a9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b9171),
	.w1(32'hbc07a365),
	.w2(32'hbb27aa5a),
	.w3(32'hbc83fc3a),
	.w4(32'hbc8cfcf8),
	.w5(32'hbc797023),
	.w6(32'hbbc56b96),
	.w7(32'h3a9bcb26),
	.w8(32'h3b8af295),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc61843b),
	.w1(32'hbb1c78f8),
	.w2(32'h3b2431b1),
	.w3(32'hbbd7411d),
	.w4(32'h3b394c2e),
	.w5(32'h3b307df4),
	.w6(32'hbba4d24f),
	.w7(32'hbae9937d),
	.w8(32'hbac6136f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dd26c),
	.w1(32'hbc43b30d),
	.w2(32'h3bfe7db6),
	.w3(32'hbbeede73),
	.w4(32'hbc206f64),
	.w5(32'h3c649837),
	.w6(32'hbc3eb353),
	.w7(32'hbc8a06be),
	.w8(32'h3bdfe528),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule