module layer_10_featuremap_209(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a43cb1),
	.w1(32'hb992d1dc),
	.w2(32'h39252f10),
	.w3(32'h384b81ff),
	.w4(32'h380740b1),
	.w5(32'h3793fc36),
	.w6(32'hb99be6ad),
	.w7(32'h3889c92b),
	.w8(32'hb9abc490),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0da426),
	.w1(32'h3b54892d),
	.w2(32'h3bbe11bd),
	.w3(32'h3bbfc704),
	.w4(32'hba972dd4),
	.w5(32'h3a893931),
	.w6(32'h3b8687e4),
	.w7(32'hbb4dcdb5),
	.w8(32'h3a9203eb),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96aca9b),
	.w1(32'hb888db6f),
	.w2(32'hb9a480d1),
	.w3(32'hb920dfc4),
	.w4(32'h37e28e2f),
	.w5(32'hb93bdb9a),
	.w6(32'hb908b3fd),
	.w7(32'hb967b5ac),
	.w8(32'hb9aa5429),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe8c8b),
	.w1(32'hbaa8a593),
	.w2(32'hbafa90c5),
	.w3(32'hb9f53759),
	.w4(32'h392b83ab),
	.w5(32'hb88601c8),
	.w6(32'hba6b9ef7),
	.w7(32'hba3bd35c),
	.w8(32'hb9fb89ac),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93853e),
	.w1(32'h384bbc40),
	.w2(32'h3a3ad762),
	.w3(32'hba8880b7),
	.w4(32'hb9823193),
	.w5(32'h38e3a101),
	.w6(32'hba140c83),
	.w7(32'hb9fb6c15),
	.w8(32'hb8f801a9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de6797),
	.w1(32'h39930d03),
	.w2(32'h398b3264),
	.w3(32'h38571243),
	.w4(32'h399e9267),
	.w5(32'h395cbec4),
	.w6(32'h393d8ad8),
	.w7(32'h39a8527c),
	.w8(32'h38f9f64a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b4748),
	.w1(32'h3b3ae2b4),
	.w2(32'h3bf0173e),
	.w3(32'hb93eac1e),
	.w4(32'h3bc4e72a),
	.w5(32'h3c2f6e4b),
	.w6(32'hbb366eb0),
	.w7(32'h3b4cf796),
	.w8(32'h3c18c4a2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0495),
	.w1(32'h3c2f857a),
	.w2(32'h3c2aac6f),
	.w3(32'h3c83aac0),
	.w4(32'h3c4feb7b),
	.w5(32'h3bdb6613),
	.w6(32'h3c51821a),
	.w7(32'h3b9c6780),
	.w8(32'h3bde06b8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a3ea9),
	.w1(32'hba569ad7),
	.w2(32'h3a747160),
	.w3(32'hb845ee04),
	.w4(32'hbaa9a75d),
	.w5(32'h3a8e1f1f),
	.w6(32'h3993bebe),
	.w7(32'hb9c1cedd),
	.w8(32'h3a50c052),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c652e64),
	.w1(32'h3b1d5e38),
	.w2(32'h3c9a4cd8),
	.w3(32'h3c49da91),
	.w4(32'hba9e5135),
	.w5(32'h3c284a20),
	.w6(32'h3c0e8a74),
	.w7(32'hbb9a3a4b),
	.w8(32'h3bb0bd6d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9616f3),
	.w1(32'h3addfca7),
	.w2(32'h3a8c2d09),
	.w3(32'h3a9470f8),
	.w4(32'h3a13daae),
	.w5(32'h3a0c0fa5),
	.w6(32'h3a98ca38),
	.w7(32'h3961c357),
	.w8(32'hb9719e61),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a340ed2),
	.w1(32'hbbf89797),
	.w2(32'hb9cbdbbd),
	.w3(32'h3bb7abff),
	.w4(32'hbb1fe566),
	.w5(32'h3b53c084),
	.w6(32'h3b0bfc16),
	.w7(32'hbbbf4083),
	.w8(32'h3bfead5d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a705a),
	.w1(32'h3ba1f400),
	.w2(32'h3c9f72b6),
	.w3(32'h3bd01ce0),
	.w4(32'h3ad91174),
	.w5(32'h3c6ca7e4),
	.w6(32'h3b53fa71),
	.w7(32'hbad2b389),
	.w8(32'h3c08c035),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1d9d1),
	.w1(32'h3be9600c),
	.w2(32'h3c05a65c),
	.w3(32'h3b6db4d3),
	.w4(32'h3b879141),
	.w5(32'h3b832e20),
	.w6(32'h3b8f7a44),
	.w7(32'h3b599a37),
	.w8(32'h3b3d65c7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9aef2),
	.w1(32'hb9f501b6),
	.w2(32'h3bb1dacb),
	.w3(32'h3b639131),
	.w4(32'hbbb6f0c9),
	.w5(32'hba5d0819),
	.w6(32'h3bc009fc),
	.w7(32'hbb964bb7),
	.w8(32'h3a76a3bf),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c434a68),
	.w1(32'h3b87f56e),
	.w2(32'h3c6e0253),
	.w3(32'h3bd53099),
	.w4(32'hbaf129ad),
	.w5(32'h3bd5927a),
	.w6(32'h3c0d3473),
	.w7(32'h3a3461bd),
	.w8(32'h3b8e18a9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944a29d),
	.w1(32'hb98c5dab),
	.w2(32'hb9f624f8),
	.w3(32'h3a1d7bb0),
	.w4(32'hb89fb589),
	.w5(32'hba32853e),
	.w6(32'h396700f8),
	.w7(32'hb90d47dd),
	.w8(32'hba96c573),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a18a3),
	.w1(32'h3b4abda0),
	.w2(32'h3c4f24bb),
	.w3(32'h3c1b040b),
	.w4(32'h3a6faf63),
	.w5(32'h3c58685d),
	.w6(32'h3c119c5d),
	.w7(32'hba281440),
	.w8(32'h3c19211e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ad651),
	.w1(32'h3b221e54),
	.w2(32'h3c32bfa4),
	.w3(32'h3b10c59f),
	.w4(32'h3ae1443d),
	.w5(32'h3c19db4d),
	.w6(32'h3a64ae7c),
	.w7(32'h39a8eaa0),
	.w8(32'h3bcd1387),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9015592),
	.w1(32'hb911ec64),
	.w2(32'h389af10b),
	.w3(32'hb93af577),
	.w4(32'hb9587de5),
	.w5(32'hb6902fb6),
	.w6(32'hb94e6352),
	.w7(32'hb97492fd),
	.w8(32'h38db8db2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982d993),
	.w1(32'h391651f5),
	.w2(32'hb88ce062),
	.w3(32'hb96edd22),
	.w4(32'h39820ece),
	.w5(32'h38f3d89c),
	.w6(32'hb8a2d202),
	.w7(32'h38c23727),
	.w8(32'hb88f3f36),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4952d0),
	.w1(32'hbb64ee86),
	.w2(32'h3a59a441),
	.w3(32'hb9a791b3),
	.w4(32'hbbb330d0),
	.w5(32'h39b47d39),
	.w6(32'hb90cdf84),
	.w7(32'hbbbbd081),
	.w8(32'hbab8a7f7),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbb3682),
	.w1(32'hba56577c),
	.w2(32'h3c248ed7),
	.w3(32'h3c95d7e7),
	.w4(32'hbb9c83ec),
	.w5(32'h3c16a01e),
	.w6(32'h3c98ab70),
	.w7(32'hbb346861),
	.w8(32'h3c837146),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86a10a),
	.w1(32'h3a871f22),
	.w2(32'h3c70fee4),
	.w3(32'h3c1adf1d),
	.w4(32'hbbc1b95a),
	.w5(32'h3bcfc6bb),
	.w6(32'h3c184d1d),
	.w7(32'hbc0617da),
	.w8(32'h3b3a07cf),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbed535),
	.w1(32'h38e03ee3),
	.w2(32'h3c3d0521),
	.w3(32'h3c7e9ae8),
	.w4(32'hbbd90614),
	.w5(32'h3b5801a7),
	.w6(32'h3c81e077),
	.w7(32'hbc1e3deb),
	.w8(32'h3a149218),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eb51e3),
	.w1(32'hb847ba74),
	.w2(32'h398eb0e7),
	.w3(32'hb95f362d),
	.w4(32'h394a51e6),
	.w5(32'h3a0a0b63),
	.w6(32'hb92062de),
	.w7(32'hb8951caf),
	.w8(32'hb846e03b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5333c),
	.w1(32'hb998f66b),
	.w2(32'hb9e96790),
	.w3(32'hba96a9f6),
	.w4(32'hb901fff4),
	.w5(32'hb9a9d374),
	.w6(32'hb9dc8c13),
	.w7(32'hb952dff0),
	.w8(32'hb9b79383),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c61a),
	.w1(32'hbba31a57),
	.w2(32'h3b846530),
	.w3(32'hbb042faa),
	.w4(32'hbbc6f26c),
	.w5(32'hbbdd0c45),
	.w6(32'hbac90b63),
	.w7(32'hbb89b397),
	.w8(32'hbb957134),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb5a9),
	.w1(32'hbaf3198d),
	.w2(32'hbac936e5),
	.w3(32'h3b9c974a),
	.w4(32'hbb170752),
	.w5(32'hbab2eb61),
	.w6(32'h3bf427a9),
	.w7(32'hbb0ec0bf),
	.w8(32'hbabcc512),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0e8bd),
	.w1(32'hbb6dade3),
	.w2(32'h3c28f2b3),
	.w3(32'h3ae3deac),
	.w4(32'hbb919917),
	.w5(32'h3b4845d9),
	.w6(32'h3b6bdcc8),
	.w7(32'hbbb682b0),
	.w8(32'h393d4124),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955d347),
	.w1(32'h381cc9c9),
	.w2(32'hb8adcee4),
	.w3(32'hb9ee3c4a),
	.w4(32'h389b3039),
	.w5(32'hb7a9a62b),
	.w6(32'h3708d309),
	.w7(32'hb86702e5),
	.w8(32'hb872ed90),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38066139),
	.w1(32'h39525918),
	.w2(32'h38c3cc97),
	.w3(32'h3926b8e5),
	.w4(32'h395163c4),
	.w5(32'hb898db01),
	.w6(32'h398842c5),
	.w7(32'h36e7b786),
	.w8(32'hb9a3b9f1),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4f04a),
	.w1(32'h390378ca),
	.w2(32'h3bdfecee),
	.w3(32'h3b310c6b),
	.w4(32'hbb27b64a),
	.w5(32'h3b451889),
	.w6(32'h3b131ac4),
	.w7(32'hbb59e7bb),
	.w8(32'h3ac3161c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc596b4),
	.w1(32'h3757df0e),
	.w2(32'h3af9f313),
	.w3(32'h3bac0152),
	.w4(32'hba404e30),
	.w5(32'h39e5ec14),
	.w6(32'h3bb1376f),
	.w7(32'hbaec1fed),
	.w8(32'h3a1f95c1),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6aa535),
	.w1(32'h3a0534d2),
	.w2(32'hb99c5a79),
	.w3(32'h3a957b63),
	.w4(32'h3a90c9b4),
	.w5(32'hb9c42c06),
	.w6(32'h3a837814),
	.w7(32'h3a807fa8),
	.w8(32'h3a7aeedd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba486f4f),
	.w1(32'h3abfde8e),
	.w2(32'h3b7582db),
	.w3(32'h39ba04b6),
	.w4(32'h3b2d2f5d),
	.w5(32'h3b90979b),
	.w6(32'hbaf5b763),
	.w7(32'h3741de08),
	.w8(32'h3b5c847d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26c8f0),
	.w1(32'hbb8339b8),
	.w2(32'h3c692077),
	.w3(32'h3c139e20),
	.w4(32'hbb7d66b6),
	.w5(32'h3bc0c118),
	.w6(32'h3b0634a5),
	.w7(32'hbc3881cc),
	.w8(32'h3c04c2c6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0914b7),
	.w1(32'hbc318e4b),
	.w2(32'hbb7b2202),
	.w3(32'h3cb89300),
	.w4(32'hbc93058c),
	.w5(32'hbc463cad),
	.w6(32'h3cd56959),
	.w7(32'hbc84ce0b),
	.w8(32'hbbaee784),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca261f0),
	.w1(32'hbc31a078),
	.w2(32'hbbd73372),
	.w3(32'h3c984d5d),
	.w4(32'hbc541e0e),
	.w5(32'hbc19ab6b),
	.w6(32'h3ccd66cf),
	.w7(32'hbc293015),
	.w8(32'hbb12535c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd020b5),
	.w1(32'hba3c58b5),
	.w2(32'hba60be53),
	.w3(32'h3b92309f),
	.w4(32'hbb07be6a),
	.w5(32'hbb2da998),
	.w6(32'h3b8ecbe7),
	.w7(32'hbb0441e8),
	.w8(32'hba9754c8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce058b),
	.w1(32'h390dd917),
	.w2(32'h38e6f779),
	.w3(32'hb9d0566a),
	.w4(32'h3903b2c4),
	.w5(32'h389a2369),
	.w6(32'hb98b1590),
	.w7(32'h39c648c9),
	.w8(32'hb8e7e137),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6df60e),
	.w1(32'hba15f1e6),
	.w2(32'hba49faad),
	.w3(32'hba7977c2),
	.w4(32'hb9a65c61),
	.w5(32'hba2d9873),
	.w6(32'hba6bdaa5),
	.w7(32'hb9dba585),
	.w8(32'hb9fc9ab4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc176),
	.w1(32'hbb0a85c4),
	.w2(32'h39e719eb),
	.w3(32'h3bb95f87),
	.w4(32'hbacf5343),
	.w5(32'h3ad36c91),
	.w6(32'h3ba1c871),
	.w7(32'hba0ba74e),
	.w8(32'h3abe98a8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7acf82),
	.w1(32'h3a9b8233),
	.w2(32'h3c60e016),
	.w3(32'h3c3f6b51),
	.w4(32'hba4d0fc7),
	.w5(32'h3bd51ddf),
	.w6(32'h3c3e0a9a),
	.w7(32'h3b3188d1),
	.w8(32'h3beb38c1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c709ca7),
	.w1(32'hbaaf11b2),
	.w2(32'h3c5e6968),
	.w3(32'h3bf3c460),
	.w4(32'hbc05fc07),
	.w5(32'h3ba13930),
	.w6(32'h3c00c757),
	.w7(32'hbc2770a3),
	.w8(32'h3a98fc3c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9f3af6),
	.w1(32'h3a9d8a50),
	.w2(32'h3c79e91d),
	.w3(32'h3c36e4b8),
	.w4(32'hbbcaad71),
	.w5(32'h3bd010bb),
	.w6(32'h3c1f7a36),
	.w7(32'hbc28e7b9),
	.w8(32'h3ae845ab),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77972c),
	.w1(32'hb9410f78),
	.w2(32'h3bea95cb),
	.w3(32'h3c526bd3),
	.w4(32'hbb510633),
	.w5(32'h3b15c1f2),
	.w6(32'h3c2dd1cc),
	.w7(32'hbb72c4b5),
	.w8(32'h3b4f2d55),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11525b),
	.w1(32'h3c06aeb8),
	.w2(32'h3c8f850f),
	.w3(32'h3bb486f7),
	.w4(32'h3c127f74),
	.w5(32'h3c82ed61),
	.w6(32'hbafe5ee7),
	.w7(32'h3b00083e),
	.w8(32'h3c108501),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20565f),
	.w1(32'hb872ddab),
	.w2(32'h39863ebb),
	.w3(32'hba63cc83),
	.w4(32'hb87b39b6),
	.w5(32'h370ea697),
	.w6(32'hb9415536),
	.w7(32'hb86038d3),
	.w8(32'h38e0fa8c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7c4b7),
	.w1(32'hba62ab1a),
	.w2(32'hba8b0c0d),
	.w3(32'hb9c7a731),
	.w4(32'hb9ad5d6a),
	.w5(32'hba0fabbb),
	.w6(32'h39bcd085),
	.w7(32'h3a2c7fad),
	.w8(32'h3a7707a4),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b03da5),
	.w1(32'h379de1ae),
	.w2(32'hb9d26b4a),
	.w3(32'hba81f9c9),
	.w4(32'hb969306c),
	.w5(32'hb9bb3a40),
	.w6(32'hba5b0db5),
	.w7(32'hba310848),
	.w8(32'hb980a7bc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c215368),
	.w1(32'h3abfbbd2),
	.w2(32'h3c274e6a),
	.w3(32'h3b9f18f9),
	.w4(32'hbb04e8ef),
	.w5(32'h3b86bc77),
	.w6(32'h3b44945a),
	.w7(32'hbba5acd5),
	.w8(32'h39d91fb7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b180c47),
	.w1(32'h3a71e6cd),
	.w2(32'h3b56c1be),
	.w3(32'h3acffcc8),
	.w4(32'h39b115d5),
	.w5(32'h3b2b7fc0),
	.w6(32'h3a6b8862),
	.w7(32'hb99befbc),
	.w8(32'h3b082541),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d0548),
	.w1(32'h3b359952),
	.w2(32'h3c7cdb49),
	.w3(32'h3bf2c640),
	.w4(32'h3a876779),
	.w5(32'h3c26980d),
	.w6(32'h3bb2b29b),
	.w7(32'hbad91128),
	.w8(32'h3c0740a4),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5bca7),
	.w1(32'hbaf20baa),
	.w2(32'hb8d49e92),
	.w3(32'h3afe39be),
	.w4(32'h370780d1),
	.w5(32'h3a3e4a69),
	.w6(32'h3aeb1430),
	.w7(32'hba1663ec),
	.w8(32'h3aa678d6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d40df),
	.w1(32'h3941dabd),
	.w2(32'h39ecb210),
	.w3(32'hb7665fd8),
	.w4(32'hb9510e8a),
	.w5(32'hb8c00856),
	.w6(32'hb8d39e9b),
	.w7(32'hb98fccc2),
	.w8(32'hba14ea66),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b337bf),
	.w1(32'hb9a4e986),
	.w2(32'hb9a259f7),
	.w3(32'hba016c93),
	.w4(32'hb9a3f92c),
	.w5(32'hb9b58c48),
	.w6(32'hb9acd7e1),
	.w7(32'hb9f491a0),
	.w8(32'hb9a039ac),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d64be),
	.w1(32'hba1e8f56),
	.w2(32'h382e7c28),
	.w3(32'hb985fffa),
	.w4(32'hb9942859),
	.w5(32'hb9bfbc14),
	.w6(32'h396e399c),
	.w7(32'hb9b9f0a8),
	.w8(32'h39a0cb1b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2787a),
	.w1(32'hbafe6fa9),
	.w2(32'hb9df322b),
	.w3(32'h3a63507b),
	.w4(32'hbb26eefa),
	.w5(32'hba52aec9),
	.w6(32'h3b0c84da),
	.w7(32'hbab02b94),
	.w8(32'hba0f77cf),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adad59f),
	.w1(32'h3a837d5a),
	.w2(32'h3a8e4e68),
	.w3(32'h3a1b5c3e),
	.w4(32'h391cdde4),
	.w5(32'h39926f8a),
	.w6(32'h3a8d7928),
	.w7(32'h3a362c9f),
	.w8(32'h3a32ee56),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28efab),
	.w1(32'h3b8b147d),
	.w2(32'h3bd58ceb),
	.w3(32'h3c1a70bc),
	.w4(32'h3b693e63),
	.w5(32'h3b9033b3),
	.w6(32'h3bbc10a1),
	.w7(32'h3a803e9d),
	.w8(32'h3ac207b8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a3fa),
	.w1(32'h3a43a45b),
	.w2(32'h3b7f04ca),
	.w3(32'h3bbe783a),
	.w4(32'h3b1a3c58),
	.w5(32'h3b348341),
	.w6(32'h3baeb9cd),
	.w7(32'h3b41df3c),
	.w8(32'h3b95e3dc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9e181),
	.w1(32'hb8943a3f),
	.w2(32'h398a4038),
	.w3(32'hb8afdbec),
	.w4(32'h38f3eb24),
	.w5(32'h39f478c5),
	.w6(32'hb965468e),
	.w7(32'h38ac1ff9),
	.w8(32'hb9134cb4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940c5d6),
	.w1(32'hb9a49c38),
	.w2(32'hb9ce9160),
	.w3(32'hb8dd32b7),
	.w4(32'hb96e2d95),
	.w5(32'hb9641bdc),
	.w6(32'hba1b1bca),
	.w7(32'hb9d55912),
	.w8(32'hb9cf534c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f24895),
	.w1(32'hb895beff),
	.w2(32'h38a118ad),
	.w3(32'hb9f32311),
	.w4(32'hb989fa08),
	.w5(32'hb9082013),
	.w6(32'hb9fdf22d),
	.w7(32'hb9c11f01),
	.w8(32'hb9957176),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a53ec1),
	.w1(32'h37e5621c),
	.w2(32'hb7f05ed4),
	.w3(32'hb962e26f),
	.w4(32'h398833e8),
	.w5(32'h36128a44),
	.w6(32'h3786e4ec),
	.w7(32'hb94f65ef),
	.w8(32'hb9463a58),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d8e41),
	.w1(32'h3bcc4737),
	.w2(32'h3c5c813b),
	.w3(32'h3c19c997),
	.w4(32'h3c00782b),
	.w5(32'h3b8b9ea0),
	.w6(32'h3bde494e),
	.w7(32'h3c0a07cb),
	.w8(32'h3c1b5de3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c977467),
	.w1(32'h3b492de0),
	.w2(32'h3c707304),
	.w3(32'h3c54f960),
	.w4(32'hb8a0de48),
	.w5(32'h3c5efb4b),
	.w6(32'h3c0cd974),
	.w7(32'hbbaab563),
	.w8(32'h3c1758cc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c883353),
	.w1(32'hbb578cc2),
	.w2(32'h3bb0f005),
	.w3(32'h3c5c2339),
	.w4(32'hbbdd05f0),
	.w5(32'h3b3da3c5),
	.w6(32'h3c58c41a),
	.w7(32'hbb385266),
	.w8(32'h3bbbb754),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccd8d24),
	.w1(32'hbc0555e6),
	.w2(32'h3c932a93),
	.w3(32'h3c49494f),
	.w4(32'hbc9a6678),
	.w5(32'hbadb078e),
	.w6(32'h3c927652),
	.w7(32'hbcbe7d78),
	.w8(32'hba2596c2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ef63d),
	.w1(32'h378d12d2),
	.w2(32'hb999cc6a),
	.w3(32'h38369092),
	.w4(32'h393cf101),
	.w5(32'hb9109873),
	.w6(32'hb9f72325),
	.w7(32'hb96fca7d),
	.w8(32'hb9adb971),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65b5f7),
	.w1(32'h391ec413),
	.w2(32'hb741b6f7),
	.w3(32'hba2e7e4e),
	.w4(32'h39901c46),
	.w5(32'h384d73f9),
	.w6(32'hb9bcd6e4),
	.w7(32'h3905f760),
	.w8(32'hb8e9a6d3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7786d),
	.w1(32'h39b22a72),
	.w2(32'h396b0237),
	.w3(32'hb9b6f720),
	.w4(32'h39dece69),
	.w5(32'h39530be8),
	.w6(32'hb9b582eb),
	.w7(32'h39ba33c4),
	.w8(32'h38002d1c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b208f2a),
	.w1(32'hb965ab13),
	.w2(32'h3aaeae13),
	.w3(32'h3b2e385c),
	.w4(32'h39fd1349),
	.w5(32'h3b07c0b1),
	.w6(32'h3b0b262d),
	.w7(32'hb84003f3),
	.w8(32'h3aa339fb),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba03a109),
	.w1(32'hb99ef122),
	.w2(32'hb983dca1),
	.w3(32'hb9a8502b),
	.w4(32'hb91cdfa2),
	.w5(32'hb91fd0eb),
	.w6(32'hba386803),
	.w7(32'hb98717ca),
	.w8(32'hb9b23eb7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b364a7b),
	.w1(32'h3b0c9ff0),
	.w2(32'h3b61bc74),
	.w3(32'h3b595b2d),
	.w4(32'h3b736032),
	.w5(32'h3b2222ba),
	.w6(32'h3a332ce9),
	.w7(32'h3ab38747),
	.w8(32'h3ac7d16f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c347a5a),
	.w1(32'h3b861a40),
	.w2(32'h3c15994e),
	.w3(32'h3c16a0b9),
	.w4(32'h3a770a14),
	.w5(32'h3b7af9cd),
	.w6(32'h3c1519c2),
	.w7(32'h3b13c4e3),
	.w8(32'h3ba305d7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c545462),
	.w1(32'h3bb4b2d9),
	.w2(32'h3c621a0f),
	.w3(32'h3c06a930),
	.w4(32'hb9736489),
	.w5(32'h3bc74720),
	.w6(32'h3b8b6007),
	.w7(32'hbbc128a3),
	.w8(32'h39b67b5e),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be27657),
	.w1(32'h3a34f101),
	.w2(32'h3bdd3443),
	.w3(32'h3bacf471),
	.w4(32'hbabc2d87),
	.w5(32'h3b46ed58),
	.w6(32'h3bad08bf),
	.w7(32'hbaf2b56e),
	.w8(32'h3b50f590),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa83327),
	.w1(32'hb8ebfa00),
	.w2(32'h3bc230d6),
	.w3(32'h3a6d4f08),
	.w4(32'h3add5859),
	.w5(32'h3b555921),
	.w6(32'hb8a5bb8f),
	.w7(32'hba5db0a0),
	.w8(32'h3b861c4d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd00918),
	.w1(32'hb8dfae75),
	.w2(32'h3ba7f3c5),
	.w3(32'h3b6974e1),
	.w4(32'hbaae9ad0),
	.w5(32'h3af0ce29),
	.w6(32'h3b78c689),
	.w7(32'hbafa0e2a),
	.w8(32'hb9409b19),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6692d),
	.w1(32'h3acb171c),
	.w2(32'h3bd3d71b),
	.w3(32'h3b0b82f1),
	.w4(32'h3b3455e3),
	.w5(32'h3bf7fc46),
	.w6(32'hb95cd741),
	.w7(32'hba8169e2),
	.w8(32'h3b5641b4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ba0f24),
	.w1(32'hb8713167),
	.w2(32'hb8fada8f),
	.w3(32'hb918f9da),
	.w4(32'hb912783b),
	.w5(32'hb9266359),
	.w6(32'hb96fcc4a),
	.w7(32'hb89272cf),
	.w8(32'hb943571f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99793d9),
	.w1(32'hb851af06),
	.w2(32'h37d709cb),
	.w3(32'hb9cd33b5),
	.w4(32'hb888de56),
	.w5(32'hb73bb5ff),
	.w6(32'hb7bfc354),
	.w7(32'hb8152b96),
	.w8(32'hb8ea12cf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9340133),
	.w1(32'h37e99507),
	.w2(32'hb8ca53c3),
	.w3(32'h3934ca39),
	.w4(32'h38d4797c),
	.w5(32'h38494b94),
	.w6(32'hb8eaca46),
	.w7(32'hb883a89d),
	.w8(32'hb98a03f8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a1687),
	.w1(32'hba3ca911),
	.w2(32'hb9d4faf7),
	.w3(32'hb99b71b4),
	.w4(32'hba5270dc),
	.w5(32'hba2132e9),
	.w6(32'hb982e199),
	.w7(32'hba8212dd),
	.w8(32'hba2504eb),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c888311),
	.w1(32'hbabda4a4),
	.w2(32'hbb181fb2),
	.w3(32'h3c647109),
	.w4(32'hbb2c0e96),
	.w5(32'hbb95ba49),
	.w6(32'h3c3c7cca),
	.w7(32'hbbd3b2e2),
	.w8(32'hbb64d8e4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c201b),
	.w1(32'hba52de40),
	.w2(32'hba5e0cbb),
	.w3(32'hbaddc57d),
	.w4(32'hbb1aa8f9),
	.w5(32'hbab5203c),
	.w6(32'h3a7dbf3f),
	.w7(32'hba6e19a0),
	.w8(32'hb9aae4a0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20472d),
	.w1(32'h3b4bc85a),
	.w2(32'h3c28637a),
	.w3(32'h3b994fd9),
	.w4(32'hba847a19),
	.w5(32'h3bd16c0b),
	.w6(32'h3b91265a),
	.w7(32'hbae92d09),
	.w8(32'h3b71a161),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39786e),
	.w1(32'h3b8598be),
	.w2(32'h3be4bba4),
	.w3(32'h3c80d4c6),
	.w4(32'h3baba1e8),
	.w5(32'h3ba95490),
	.w6(32'h3c709697),
	.w7(32'h3bb653ae),
	.w8(32'h3bb446c8),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb98f2b),
	.w1(32'hbbbb3568),
	.w2(32'hba562b69),
	.w3(32'h3bcc419d),
	.w4(32'hbbc11d82),
	.w5(32'hbb89a41b),
	.w6(32'h3be783d9),
	.w7(32'hbbb0b1ea),
	.w8(32'hbaf8da04),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0566e9),
	.w1(32'h3b9f1cb6),
	.w2(32'h3c399db1),
	.w3(32'h3be3ffc0),
	.w4(32'hb8ef50c3),
	.w5(32'h3b607a88),
	.w6(32'h3bbb76e7),
	.w7(32'h3afc3dc7),
	.w8(32'h3be41d02),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b343417),
	.w1(32'hbbc2ec13),
	.w2(32'hbaad5967),
	.w3(32'h3a9d9ef7),
	.w4(32'hbc09ee44),
	.w5(32'hbb82c85d),
	.w6(32'hb8cd7101),
	.w7(32'hbc23be4a),
	.w8(32'hbbc756a1),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c805056),
	.w1(32'h3b5ec963),
	.w2(32'h3c2adef5),
	.w3(32'h3c5b05df),
	.w4(32'h3a0b5e99),
	.w5(32'h3b919032),
	.w6(32'h3c72e392),
	.w7(32'hb9684b1c),
	.w8(32'h3bcdb3c1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c06275d),
	.w1(32'h35f91e34),
	.w2(32'h3b9e8791),
	.w3(32'h3bbac218),
	.w4(32'hbb27d6da),
	.w5(32'hbb224e41),
	.w6(32'h3b96f4d2),
	.w7(32'hbb394a12),
	.w8(32'hba82e77a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ec721),
	.w1(32'hbb1c4d61),
	.w2(32'h3b8b39f4),
	.w3(32'h3c0d3c02),
	.w4(32'hbbd1dd18),
	.w5(32'hb93a0bbd),
	.w6(32'h3c08aa71),
	.w7(32'hbc0132f2),
	.w8(32'hbb40b926),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d1c9d),
	.w1(32'hb9e901bf),
	.w2(32'hba8ef9b7),
	.w3(32'hb9b7e35e),
	.w4(32'hba40b785),
	.w5(32'hbabc0121),
	.w6(32'hba3da979),
	.w7(32'hba211da0),
	.w8(32'hbab1ec5b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2124a6),
	.w1(32'hb886cbee),
	.w2(32'h3c3f1e99),
	.w3(32'h3bd13ec4),
	.w4(32'hbb9e89d6),
	.w5(32'h3b8a9751),
	.w6(32'h3bf54de6),
	.w7(32'hbb1fda51),
	.w8(32'h3bd4374e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0f7c7),
	.w1(32'hbb07460e),
	.w2(32'h3b85e50b),
	.w3(32'h3bd9be71),
	.w4(32'hbb37fdb0),
	.w5(32'hb9a4cd67),
	.w6(32'h3b4966c7),
	.w7(32'hbac41494),
	.w8(32'h3bd8ba1c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c459734),
	.w1(32'h3b2ec2d4),
	.w2(32'h3c5ad5b9),
	.w3(32'h3c08b41b),
	.w4(32'hbae937cf),
	.w5(32'h3c156f32),
	.w6(32'hb8bd5041),
	.w7(32'hbc21d425),
	.w8(32'h3c0d122a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0636e6),
	.w1(32'hbc59895c),
	.w2(32'hbc890121),
	.w3(32'h3cc81bf8),
	.w4(32'hbcb1c7d2),
	.w5(32'hbc8e526b),
	.w6(32'h3cb32b87),
	.w7(32'hbc8f6c48),
	.w8(32'hbc14c2e4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38b322),
	.w1(32'h3880754b),
	.w2(32'h3c8511fb),
	.w3(32'h3b931b65),
	.w4(32'hbb94b072),
	.w5(32'h3c1569fb),
	.w6(32'h3bac7b77),
	.w7(32'hbbf78ef6),
	.w8(32'h3b3328c5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf504d9),
	.w1(32'h3b44fcc4),
	.w2(32'h3c150a8f),
	.w3(32'h3bed6f8b),
	.w4(32'h3b082526),
	.w5(32'h3bd486e8),
	.w6(32'hbb51e927),
	.w7(32'hbbaa2a21),
	.w8(32'h3c03dafb),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f2df0),
	.w1(32'h39bc54a3),
	.w2(32'hb9e32130),
	.w3(32'hb93565ad),
	.w4(32'hb9eaa8b3),
	.w5(32'hb9bf9ec8),
	.w6(32'h39637c81),
	.w7(32'hba6e1b96),
	.w8(32'hbac77940),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb06b5c),
	.w1(32'h3c43109a),
	.w2(32'h3c915d18),
	.w3(32'h3c3463de),
	.w4(32'h3b948eb0),
	.w5(32'h3c3e4d8d),
	.w6(32'hbb4880a3),
	.w7(32'hbbb4bcf2),
	.w8(32'h3b3db38e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86953b),
	.w1(32'hbbc87d90),
	.w2(32'h3aa3960c),
	.w3(32'h3ac69d37),
	.w4(32'hbb84fc44),
	.w5(32'h3b7f7216),
	.w6(32'hba9fcdec),
	.w7(32'hbb91e106),
	.w8(32'h3b60ff39),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed91d8),
	.w1(32'hb8f75ec9),
	.w2(32'h39643a55),
	.w3(32'h3971e819),
	.w4(32'hb9e8d00f),
	.w5(32'h38aad1ef),
	.w6(32'h382e9420),
	.w7(32'hba48972c),
	.w8(32'hb9df6975),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b725819),
	.w1(32'h3b248462),
	.w2(32'h3b4bffd3),
	.w3(32'h3aa59a8f),
	.w4(32'h3a70bdfe),
	.w5(32'h3ac193e6),
	.w6(32'h3b3e1019),
	.w7(32'h3a7f84aa),
	.w8(32'h3a770837),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5a5f5),
	.w1(32'h3b6d8b00),
	.w2(32'h3c344279),
	.w3(32'h3b946cd9),
	.w4(32'h3b3db67a),
	.w5(32'h3bf9a6b8),
	.w6(32'h3b7e928f),
	.w7(32'h3b16215f),
	.w8(32'h3beac18a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba67f26),
	.w1(32'hbae6678d),
	.w2(32'h3c012841),
	.w3(32'h3b01f47e),
	.w4(32'hbb870b99),
	.w5(32'h3b3a817d),
	.w6(32'h3b069f56),
	.w7(32'hbbd57129),
	.w8(32'h39081506),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb25c69),
	.w1(32'hba928411),
	.w2(32'h3af2cc5d),
	.w3(32'h3b84c234),
	.w4(32'hbb5cd951),
	.w5(32'h3881416c),
	.w6(32'h3bf57bfa),
	.w7(32'hbacc4040),
	.w8(32'h3ade9095),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11c192),
	.w1(32'h3a138ecb),
	.w2(32'h3bc622ef),
	.w3(32'h3b974dc2),
	.w4(32'hbb4d57b6),
	.w5(32'h3adf56df),
	.w6(32'h3b7f45a1),
	.w7(32'hbb67a461),
	.w8(32'h3b2269da),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94da56),
	.w1(32'hbb7d29c1),
	.w2(32'h3a79d70c),
	.w3(32'h3be09377),
	.w4(32'hbac82463),
	.w5(32'h3b332ee2),
	.w6(32'h3b9538e9),
	.w7(32'hbb881a4b),
	.w8(32'h3afcd375),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a6c03),
	.w1(32'h3b31c18d),
	.w2(32'h3c0ebeb0),
	.w3(32'h3bd6b026),
	.w4(32'hba96e827),
	.w5(32'h3b3a8a43),
	.w6(32'h3bb7a786),
	.w7(32'hb9e69881),
	.w8(32'h3b28d4ff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba9af5),
	.w1(32'hba9fbf3b),
	.w2(32'h3b72f349),
	.w3(32'h3b715e52),
	.w4(32'hbb140adc),
	.w5(32'h3af9cfee),
	.w6(32'h3b7eee56),
	.w7(32'hbb574ba8),
	.w8(32'h3a9cfd88),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c5daea),
	.w1(32'h39f45949),
	.w2(32'h39ea5e93),
	.w3(32'h3896e9d4),
	.w4(32'h39b042e6),
	.w5(32'h39b71e3f),
	.w6(32'h39bf9647),
	.w7(32'h39b83c45),
	.w8(32'hb67f98fc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91fcdf),
	.w1(32'h3a5bb3a0),
	.w2(32'h3a72d1e1),
	.w3(32'h3a0dfc93),
	.w4(32'h39980774),
	.w5(32'h39a7204a),
	.w6(32'h3a626cf7),
	.w7(32'h39a1df86),
	.w8(32'h39a14d5c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39352662),
	.w1(32'hb91df889),
	.w2(32'hb79591e5),
	.w3(32'h39adf3a2),
	.w4(32'hb8db1656),
	.w5(32'hb8013ab1),
	.w6(32'h39a3e8a8),
	.w7(32'h389ce4ec),
	.w8(32'h37fe8420),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2d877),
	.w1(32'hb9c33e21),
	.w2(32'hba1503d6),
	.w3(32'h38ec13a8),
	.w4(32'hba0e5b7a),
	.w5(32'hba2ca1f5),
	.w6(32'hb9e769d7),
	.w7(32'hba6431e3),
	.w8(32'hbacb5725),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05528a),
	.w1(32'hbb15892a),
	.w2(32'h3ba4f7dc),
	.w3(32'h3b8a4413),
	.w4(32'hbba892c6),
	.w5(32'h3af616e3),
	.w6(32'h3b933e96),
	.w7(32'hbbd96869),
	.w8(32'hba7916f8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a053d),
	.w1(32'h3b193a83),
	.w2(32'h3b493bc3),
	.w3(32'h3aa1dc80),
	.w4(32'h3a4686ae),
	.w5(32'h3ab6deba),
	.w6(32'h3a99a79d),
	.w7(32'hb839223d),
	.w8(32'h3a163706),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba30df94),
	.w1(32'h3a51d9be),
	.w2(32'h3bb4df50),
	.w3(32'h3a9408b9),
	.w4(32'h3aed4860),
	.w5(32'h3b7f6ac4),
	.w6(32'hbb6cd8c6),
	.w7(32'hba3729b0),
	.w8(32'h3b32122f),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c88ac62),
	.w1(32'h3b2c3a30),
	.w2(32'h3be83679),
	.w3(32'h3c34fa14),
	.w4(32'hbb186235),
	.w5(32'h3a9f8180),
	.w6(32'h3c21b05b),
	.w7(32'hbb663507),
	.w8(32'h3b438da3),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993a666),
	.w1(32'h38fdb54c),
	.w2(32'hb8d8c12b),
	.w3(32'hb9ac8fe2),
	.w4(32'h389934d4),
	.w5(32'h39af0950),
	.w6(32'hb9570ce9),
	.w7(32'hb9949609),
	.w8(32'hb98f5318),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cf05d),
	.w1(32'h392a3895),
	.w2(32'h3a6867a4),
	.w3(32'h396a3c60),
	.w4(32'hb9d03248),
	.w5(32'h3867a754),
	.w6(32'h36dec697),
	.w7(32'hb94b1615),
	.w8(32'h39878589),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959b49c),
	.w1(32'h38b259b7),
	.w2(32'h37d3bc5f),
	.w3(32'hb978530d),
	.w4(32'h38f73c43),
	.w5(32'h38680bef),
	.w6(32'h38cb0492),
	.w7(32'h3900b305),
	.w8(32'h39164629),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b52e1),
	.w1(32'h3a8fde15),
	.w2(32'h3a661e8b),
	.w3(32'h3b001758),
	.w4(32'h39d54c45),
	.w5(32'h391d5388),
	.w6(32'h3b2abde0),
	.w7(32'h3a8cbe1c),
	.w8(32'h3a96542d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b197453),
	.w1(32'h3be3df06),
	.w2(32'h3c09fdad),
	.w3(32'h3a864aac),
	.w4(32'h3c0508ca),
	.w5(32'h3c6ab9f3),
	.w6(32'h38f16dc5),
	.w7(32'h3b33f13c),
	.w8(32'h3c02792d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf32c4e),
	.w1(32'h3af773a8),
	.w2(32'h3c4338b8),
	.w3(32'h3bb0187a),
	.w4(32'h3ab6b7fe),
	.w5(32'h3c09c3bf),
	.w6(32'h3b8b3616),
	.w7(32'h39b86946),
	.w8(32'h3bedd581),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd93c7),
	.w1(32'h3a9d01dd),
	.w2(32'h3adb5692),
	.w3(32'h3a18ec20),
	.w4(32'h3a33020a),
	.w5(32'h3a39ae13),
	.w6(32'hba0a23e9),
	.w7(32'h39924d37),
	.w8(32'h3a245ff5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99dca8),
	.w1(32'h3a5ea5d1),
	.w2(32'h3b5a6ca7),
	.w3(32'h3bac0205),
	.w4(32'h3904d5b2),
	.w5(32'h3add8cd2),
	.w6(32'h3ba09f3e),
	.w7(32'h3ac66ea7),
	.w8(32'h3b62e25d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3f264),
	.w1(32'hbad35099),
	.w2(32'h39a7c6f3),
	.w3(32'h3b662730),
	.w4(32'hbb04512e),
	.w5(32'hba2216f0),
	.w6(32'h3b1bec98),
	.w7(32'hbb4ca6b3),
	.w8(32'h3a24d6e6),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2da43),
	.w1(32'h3b0b4382),
	.w2(32'h3b80cb28),
	.w3(32'h3aa3ab4a),
	.w4(32'h3a7cc4e3),
	.w5(32'h3aecffb1),
	.w6(32'h3bb73a06),
	.w7(32'hba8a83fe),
	.w8(32'h3a4e4a64),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09bd63),
	.w1(32'h3b618036),
	.w2(32'h3c1d84da),
	.w3(32'h3ba7d963),
	.w4(32'h39d616ab),
	.w5(32'h3b33ddb2),
	.w6(32'h3b9bf6f8),
	.w7(32'hba8d73e1),
	.w8(32'h3b10d32a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be50d9b),
	.w1(32'h3b7c82c6),
	.w2(32'h3c3fcaac),
	.w3(32'h3bd76bea),
	.w4(32'h3aee571d),
	.w5(32'h3c225771),
	.w6(32'h3b9cdec1),
	.w7(32'h3aec2630),
	.w8(32'h3c155239),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26cb23),
	.w1(32'h3a9775f7),
	.w2(32'h3bbe6974),
	.w3(32'h3bfa165f),
	.w4(32'hbae4ff59),
	.w5(32'h3ac32562),
	.w6(32'h3bfd7061),
	.w7(32'hbb1a4cf3),
	.w8(32'h3b5219e8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f7613),
	.w1(32'h3b34add9),
	.w2(32'h3bf4b3b6),
	.w3(32'h3bb16b0f),
	.w4(32'hbb1050b0),
	.w5(32'h3b0fe9f9),
	.w6(32'h3b279624),
	.w7(32'hbb0199c6),
	.w8(32'h3b91c34a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd849e6),
	.w1(32'h3a200dfe),
	.w2(32'h3bea3071),
	.w3(32'h3ba4dd8b),
	.w4(32'h3967b5b4),
	.w5(32'h3bdc4a22),
	.w6(32'h398ff43d),
	.w7(32'hbb814a3a),
	.w8(32'h3b919428),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ec376),
	.w1(32'h3a53b26a),
	.w2(32'h3b1859bc),
	.w3(32'h3bb216e7),
	.w4(32'hbb15a7c5),
	.w5(32'hbabd708f),
	.w6(32'h3b996edf),
	.w7(32'hbb911992),
	.w8(32'hbb09eac8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb73924),
	.w1(32'h3a89b499),
	.w2(32'h3bddf935),
	.w3(32'h3b11743e),
	.w4(32'hb9de149f),
	.w5(32'h3b9f98c7),
	.w6(32'h3bad6a21),
	.w7(32'h3b0cfa3f),
	.w8(32'h3be92e43),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1ac52),
	.w1(32'hb91a11b4),
	.w2(32'h3b3af99f),
	.w3(32'h3b0d31ea),
	.w4(32'hbac85862),
	.w5(32'h3a3b1791),
	.w6(32'h3aa8f112),
	.w7(32'hbae9c6a5),
	.w8(32'hb8e0c412),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26a86d),
	.w1(32'hbbdc9bc1),
	.w2(32'h3b88fa44),
	.w3(32'h3c137b4e),
	.w4(32'hbbbf64a6),
	.w5(32'h3b7b3ac1),
	.w6(32'h3c271a5b),
	.w7(32'hbbf1c574),
	.w8(32'h3af03d60),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c143050),
	.w1(32'hba904b0f),
	.w2(32'hbb7ffe16),
	.w3(32'h3c0048fb),
	.w4(32'hb9a11315),
	.w5(32'hba9808e6),
	.w6(32'h3c12375d),
	.w7(32'hbb037a72),
	.w8(32'hba7974e5),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6e88f),
	.w1(32'h3a76353b),
	.w2(32'h3a9dbf6e),
	.w3(32'h3aea05e1),
	.w4(32'h3a575d71),
	.w5(32'h3a74654d),
	.w6(32'h3a5d3056),
	.w7(32'h3a6e8c12),
	.w8(32'h3a5452f5),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46ebb5),
	.w1(32'h3a33d063),
	.w2(32'hb8351678),
	.w3(32'h3a5baf39),
	.w4(32'h3abe17f5),
	.w5(32'h3a805557),
	.w6(32'h397f97b1),
	.w7(32'h390f2049),
	.w8(32'h3a1b6f3a),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b780427),
	.w1(32'h39bccab1),
	.w2(32'h3ac82ccb),
	.w3(32'h3ba9b650),
	.w4(32'hba528283),
	.w5(32'hbacceaba),
	.w6(32'h3b24fd77),
	.w7(32'hbac687cb),
	.w8(32'hb94a6557),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54173b),
	.w1(32'hb98ba1e6),
	.w2(32'h3b3c6e75),
	.w3(32'h3bf255a5),
	.w4(32'hbba025f5),
	.w5(32'hb9137482),
	.w6(32'h3bd917be),
	.w7(32'hbb95062d),
	.w8(32'h3a3adc8c),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c570af4),
	.w1(32'h3bb15d82),
	.w2(32'h3c721903),
	.w3(32'h3c3c1940),
	.w4(32'h3a42805b),
	.w5(32'h3c01ebd1),
	.w6(32'h3bc68dba),
	.w7(32'hbb7ad7ef),
	.w8(32'h3b895406),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba003be8),
	.w1(32'hb95c7f27),
	.w2(32'hb999e7cc),
	.w3(32'hb9309634),
	.w4(32'hb914c4cd),
	.w5(32'hb8e25de6),
	.w6(32'h36bf7e58),
	.w7(32'h398c6a13),
	.w8(32'h39346b9b),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131f3c),
	.w1(32'h3abac85a),
	.w2(32'h3c441103),
	.w3(32'h3bd5fd8e),
	.w4(32'hba80b678),
	.w5(32'h3bc10e27),
	.w6(32'h3b9d0cc2),
	.w7(32'hbac6d781),
	.w8(32'h3bbe2109),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf67118),
	.w1(32'hb96a4eb4),
	.w2(32'h3be4089c),
	.w3(32'h3ab20531),
	.w4(32'hbb2ce88e),
	.w5(32'h3b647d2a),
	.w6(32'h3b0f2a94),
	.w7(32'hba74645d),
	.w8(32'h3b69fb79),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3772a0f3),
	.w1(32'h3bad2e52),
	.w2(32'h3c669d12),
	.w3(32'h3af3f0c4),
	.w4(32'h3b9751ab),
	.w5(32'h3c2e38a2),
	.w6(32'hbb496935),
	.w7(32'h3867a3b7),
	.w8(32'h3c05b84f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d9250),
	.w1(32'hbbf6542c),
	.w2(32'h3c16553f),
	.w3(32'h3a03f077),
	.w4(32'hbc368357),
	.w5(32'h39ce2d1d),
	.w6(32'h39eb1981),
	.w7(32'hbc709797),
	.w8(32'hbb8bc59a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdd3e2),
	.w1(32'h39ead06d),
	.w2(32'h3a0ba2c8),
	.w3(32'h3b6742bf),
	.w4(32'hbac45b5f),
	.w5(32'hb90be887),
	.w6(32'h3b8a0efd),
	.w7(32'hba3f7813),
	.w8(32'h3b6315ee),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cb270),
	.w1(32'hba2ebf7c),
	.w2(32'hbae198ce),
	.w3(32'hba259550),
	.w4(32'hbab0de64),
	.w5(32'hbaed0d47),
	.w6(32'hbb154062),
	.w7(32'hbb18a716),
	.w8(32'hbaf54b25),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a5a9),
	.w1(32'hbb8dc002),
	.w2(32'hba99a65a),
	.w3(32'h3bac43d0),
	.w4(32'hbbb26ffe),
	.w5(32'hbb26bc14),
	.w6(32'h3be1fa35),
	.w7(32'hbbb71d22),
	.w8(32'hbb4186de),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4012f1),
	.w1(32'hbbcc0570),
	.w2(32'hbb94d02f),
	.w3(32'h3bf4877b),
	.w4(32'hbc1be11c),
	.w5(32'hbbc30c56),
	.w6(32'h3bd795e1),
	.w7(32'hbc091184),
	.w8(32'h3abaf023),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838a00),
	.w1(32'hbbb1411e),
	.w2(32'hb9c887d9),
	.w3(32'h3b809c1f),
	.w4(32'hbbc45f43),
	.w5(32'hba7cf684),
	.w6(32'h3bce4c4f),
	.w7(32'hbbc824c2),
	.w8(32'hbaa62d81),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0e15),
	.w1(32'h3967cb72),
	.w2(32'h3a9cfd6f),
	.w3(32'h3b2a197f),
	.w4(32'h3abaf057),
	.w5(32'h3ad4970e),
	.w6(32'hb9b2340c),
	.w7(32'h39741e04),
	.w8(32'h3ad4f981),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388a38f1),
	.w1(32'h3a0cdca9),
	.w2(32'h3a33010f),
	.w3(32'h39057f23),
	.w4(32'h391813c2),
	.w5(32'h39c16047),
	.w6(32'h39dd742d),
	.w7(32'h3a4acd5f),
	.w8(32'h3a8892f2),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea2b91),
	.w1(32'h3b77aa9c),
	.w2(32'h3b812f00),
	.w3(32'h3ba3061b),
	.w4(32'h398b3eb7),
	.w5(32'h3b182bb2),
	.w6(32'h3bb27683),
	.w7(32'hbab43a2f),
	.w8(32'h3b523b4f),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e851),
	.w1(32'hba98b751),
	.w2(32'h3894e5a4),
	.w3(32'hba8fbd48),
	.w4(32'hba9d9fd6),
	.w5(32'h38ba3540),
	.w6(32'hbb0ae552),
	.w7(32'hbac0d6d8),
	.w8(32'h3a4aca87),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f7139),
	.w1(32'hbb788207),
	.w2(32'h3b15d9dc),
	.w3(32'h3afa5b90),
	.w4(32'hbb88eb91),
	.w5(32'hb9bb17bd),
	.w6(32'h3af71d07),
	.w7(32'hbbbb999a),
	.w8(32'hbad7bba1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990313c),
	.w1(32'h36c8cf91),
	.w2(32'h3a05d649),
	.w3(32'hb9670e74),
	.w4(32'hb9e48ba2),
	.w5(32'hb9a77e7d),
	.w6(32'hb98274c6),
	.w7(32'hba0fcca1),
	.w8(32'hb9d95d27),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9bc67),
	.w1(32'h3b1b5d4b),
	.w2(32'h3bc85353),
	.w3(32'h3bc49d4e),
	.w4(32'h3b374fc8),
	.w5(32'h3b8345e7),
	.w6(32'h3baf6d45),
	.w7(32'hbabd4ad2),
	.w8(32'h3ab7a9d4),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c21fec),
	.w1(32'h3a0a9d52),
	.w2(32'h3a49a791),
	.w3(32'h392ad735),
	.w4(32'h38d26b66),
	.w5(32'h39d2fd63),
	.w6(32'h39c47833),
	.w7(32'h39cf134a),
	.w8(32'hb97c1646),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35a773),
	.w1(32'h3ad2c81d),
	.w2(32'h3af5a471),
	.w3(32'h38b102ef),
	.w4(32'h3ad15686),
	.w5(32'h3b02129e),
	.w6(32'h3ac48f87),
	.w7(32'h3acc2ade),
	.w8(32'h3ac9a090),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0afa75),
	.w1(32'h3a940407),
	.w2(32'h3b84dec7),
	.w3(32'h3be4ad80),
	.w4(32'hbab959ea),
	.w5(32'h3a9bb5e4),
	.w6(32'h3bf4be78),
	.w7(32'hbaadae65),
	.w8(32'h3acd77ac),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6059c1),
	.w1(32'h376c9942),
	.w2(32'h3c1b16a0),
	.w3(32'h3c578584),
	.w4(32'h3a7e53c5),
	.w5(32'h3c82b0d5),
	.w6(32'h3c1c65bb),
	.w7(32'hbb7723af),
	.w8(32'h3c16619a),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32cf18),
	.w1(32'hbb0636c6),
	.w2(32'h39b53f02),
	.w3(32'h3b6348fa),
	.w4(32'hbb5f11e1),
	.w5(32'hb717946d),
	.w6(32'h3be5ba50),
	.w7(32'hbaaacd1b),
	.w8(32'h39f89575),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23a2e7),
	.w1(32'h3a9d6a59),
	.w2(32'h3c1c3ec4),
	.w3(32'h3bdc5b55),
	.w4(32'hba86fcc6),
	.w5(32'h3bd25e9b),
	.w6(32'h3bb269ae),
	.w7(32'hbb55c56c),
	.w8(32'h3ba976b4),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a0919),
	.w1(32'hb982cfa8),
	.w2(32'h3ad40197),
	.w3(32'h3aaa26ba),
	.w4(32'hbac68779),
	.w5(32'hbb09c626),
	.w6(32'h3a33dd22),
	.w7(32'hbb1215c1),
	.w8(32'hbac22f9a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90c4d2),
	.w1(32'h3a93c106),
	.w2(32'h3c83d062),
	.w3(32'h3c1bf385),
	.w4(32'hbc07e867),
	.w5(32'h3b995377),
	.w6(32'h3c280bcb),
	.w7(32'hbb138430),
	.w8(32'h3c06a670),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bf68c),
	.w1(32'h3a7c2b7d),
	.w2(32'h3c135408),
	.w3(32'h3bd8d45e),
	.w4(32'hbba3d087),
	.w5(32'h3b039f45),
	.w6(32'h3bf8f0be),
	.w7(32'hbb72e184),
	.w8(32'h3b4ad7cf),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7b80),
	.w1(32'hb92b1fb4),
	.w2(32'h3c056578),
	.w3(32'h3b5d6fa1),
	.w4(32'h39a5cff1),
	.w5(32'h3c100a78),
	.w6(32'h3b8eb127),
	.w7(32'hba6dc3ce),
	.w8(32'h3baae81a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c847),
	.w1(32'hbab3ba53),
	.w2(32'hbb0f5b92),
	.w3(32'h3a9ea403),
	.w4(32'hbaeada40),
	.w5(32'hbb222ae7),
	.w6(32'hba246e2c),
	.w7(32'hbaeeaf25),
	.w8(32'hba788286),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38eed9),
	.w1(32'h3a34867e),
	.w2(32'h3bc7d388),
	.w3(32'h3b42d87a),
	.w4(32'hba424a62),
	.w5(32'h3b5cfd2f),
	.w6(32'h39830708),
	.w7(32'hbb1f7d1b),
	.w8(32'h3b085481),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91bbe77),
	.w1(32'h3aae06af),
	.w2(32'h3aa6d682),
	.w3(32'hb9907936),
	.w4(32'h3a8f73bc),
	.w5(32'h3aa215e7),
	.w6(32'h3a9fdb70),
	.w7(32'h3ac0aa7d),
	.w8(32'h3a9df95d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047d8b),
	.w1(32'h3a2a9fe1),
	.w2(32'h3ba75f1f),
	.w3(32'h3a83f7e9),
	.w4(32'hba6ec498),
	.w5(32'h3ad0cc3d),
	.w6(32'h3989ef44),
	.w7(32'hb820dbed),
	.w8(32'h3ade6009),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b162b50),
	.w1(32'h3aace45d),
	.w2(32'h3a484de3),
	.w3(32'h3b1c7c54),
	.w4(32'h39ee0fd0),
	.w5(32'h384e1b43),
	.w6(32'h3b4ecbdd),
	.w7(32'hbaa5b915),
	.w8(32'hb89386c8),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5f28b),
	.w1(32'h3aa51add),
	.w2(32'h3c12bcd0),
	.w3(32'h3bb5c7f8),
	.w4(32'hba78ba29),
	.w5(32'h3b6b5f85),
	.w6(32'h3bdef386),
	.w7(32'hba72666b),
	.w8(32'h3b8a0988),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4a556),
	.w1(32'h3b10f2d3),
	.w2(32'h3988b1f8),
	.w3(32'h3a33c9a4),
	.w4(32'h3afb9420),
	.w5(32'h3a255949),
	.w6(32'h3a476a63),
	.w7(32'hba11b79a),
	.w8(32'hb92e668f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0acca6),
	.w1(32'h3979d5c4),
	.w2(32'hb839c4fc),
	.w3(32'h39993ca7),
	.w4(32'h3a172720),
	.w5(32'hb8c63c5e),
	.w6(32'h39909dc9),
	.w7(32'h389d3e8b),
	.w8(32'hb9aa3725),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b952af0),
	.w1(32'hba2b5bbd),
	.w2(32'h39ccd515),
	.w3(32'h3b08aa50),
	.w4(32'hba7b87a6),
	.w5(32'hba14b9c8),
	.w6(32'h3ae81579),
	.w7(32'hbb598a7c),
	.w8(32'hbb2603e5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36d29a),
	.w1(32'h3a3f1888),
	.w2(32'h3bc77c3d),
	.w3(32'h3bff868d),
	.w4(32'hba0296ff),
	.w5(32'h3b502b3d),
	.w6(32'h3bcd881d),
	.w7(32'h3a16d512),
	.w8(32'h3bac26a2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b48d1),
	.w1(32'hb9f2af67),
	.w2(32'h3b742068),
	.w3(32'h3b9fc959),
	.w4(32'h3aa5c66e),
	.w5(32'h3b935985),
	.w6(32'h3a7304e1),
	.w7(32'hbb524190),
	.w8(32'h3ae8b1b0),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db4a9d),
	.w1(32'h3aa8e2c0),
	.w2(32'h3b1f720c),
	.w3(32'h3ab63273),
	.w4(32'h3ab4d981),
	.w5(32'h3b0d8387),
	.w6(32'h3b5879ae),
	.w7(32'h3ab65feb),
	.w8(32'h3b07745a),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbaaece),
	.w1(32'h3c1c499c),
	.w2(32'h3d05190f),
	.w3(32'h3c903e23),
	.w4(32'h3c1bacb6),
	.w5(32'h3ce20f0c),
	.w6(32'h3bd8406c),
	.w7(32'h3b8ad4cb),
	.w8(32'h3c4f912b),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce4845b),
	.w1(32'h3a42c1aa),
	.w2(32'h3c29940d),
	.w3(32'h3ca9e948),
	.w4(32'hbba0758d),
	.w5(32'hbae0c57c),
	.w6(32'h3c8a5a75),
	.w7(32'hbc220c28),
	.w8(32'hba12d89e),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07e8fa),
	.w1(32'h3a96d40e),
	.w2(32'h3acc3508),
	.w3(32'h395e20b2),
	.w4(32'h3b29a5b7),
	.w5(32'h3b01622b),
	.w6(32'h39b4961f),
	.w7(32'h3a9d2a2b),
	.w8(32'h3b19ecc6),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a79a8e),
	.w1(32'h3af8babb),
	.w2(32'hbb2bd168),
	.w3(32'h3a254203),
	.w4(32'h3b0cf684),
	.w5(32'hbaf5dd44),
	.w6(32'h398f024f),
	.w7(32'hbb4c2e05),
	.w8(32'hbace6e10),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59d876),
	.w1(32'hb9b52d68),
	.w2(32'hba60abfa),
	.w3(32'hbadd6a51),
	.w4(32'hba1e87e3),
	.w5(32'hbabd6160),
	.w6(32'hb9f9b2ce),
	.w7(32'hba82b55c),
	.w8(32'hba331578),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf60b9),
	.w1(32'hb91b7155),
	.w2(32'hb9ce15e7),
	.w3(32'hba8e9367),
	.w4(32'hba0c05e7),
	.w5(32'hba3acb27),
	.w6(32'hb96a2bf1),
	.w7(32'hb9d219b4),
	.w8(32'hb95bfafb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae8016),
	.w1(32'h3b146461),
	.w2(32'h3baf0961),
	.w3(32'h3997a0d3),
	.w4(32'h3b3e5170),
	.w5(32'h3bbd8214),
	.w6(32'hb8a546ba),
	.w7(32'h3b189760),
	.w8(32'h3b8ffc01),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20b4fb),
	.w1(32'h3a8da42a),
	.w2(32'h3b07f6d7),
	.w3(32'h3ba7d0d2),
	.w4(32'hbb3022b4),
	.w5(32'h3b09fa42),
	.w6(32'h3bb759a0),
	.w7(32'hba1fe390),
	.w8(32'h3b9c5644),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59cf6c),
	.w1(32'h3b9e368f),
	.w2(32'h3c655da9),
	.w3(32'h3c2bdc42),
	.w4(32'hbb345a36),
	.w5(32'h3bab000e),
	.w6(32'h3c03d384),
	.w7(32'hbbc7ce49),
	.w8(32'h392ff221),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa80dff),
	.w1(32'hba00d0bb),
	.w2(32'h3abc3341),
	.w3(32'h3accdb28),
	.w4(32'hba935f70),
	.w5(32'hb8d8d609),
	.w6(32'h3b82e0a2),
	.w7(32'h3aace1e1),
	.w8(32'h3b0ac245),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b8183),
	.w1(32'h3b91be05),
	.w2(32'h3c6f3de0),
	.w3(32'h3ba4a759),
	.w4(32'hbad9f7c5),
	.w5(32'h3c219408),
	.w6(32'h3b58dd53),
	.w7(32'hb99d76a6),
	.w8(32'h3bd520b9),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae220fb),
	.w1(32'hb996ec92),
	.w2(32'h3b3d84d3),
	.w3(32'hb886abf4),
	.w4(32'hb98efc82),
	.w5(32'h3b0e823c),
	.w6(32'h389c9853),
	.w7(32'hba7bb8b9),
	.w8(32'h3ae30a92),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390b3a37),
	.w1(32'h3a5b9146),
	.w2(32'h3a5e8108),
	.w3(32'hb99dad8b),
	.w4(32'h3a87d72f),
	.w5(32'h3a86a473),
	.w6(32'h3a4fa9b3),
	.w7(32'h3ab2dbd7),
	.w8(32'h3a6c5453),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459921),
	.w1(32'h3b6440ed),
	.w2(32'h3b1230e9),
	.w3(32'h3b2faf32),
	.w4(32'h3b4c23aa),
	.w5(32'h3b043520),
	.w6(32'h3b2921fa),
	.w7(32'h3ac3b3d3),
	.w8(32'h3a32dcf7),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b5cb1),
	.w1(32'hba1c22e0),
	.w2(32'hb9f707c8),
	.w3(32'h3a365942),
	.w4(32'hba3035df),
	.w5(32'hba220750),
	.w6(32'hbaa4eb34),
	.w7(32'hb9b76756),
	.w8(32'hba07f87f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33d18b),
	.w1(32'h3a01bc95),
	.w2(32'h3b58a1cc),
	.w3(32'h3c0173f8),
	.w4(32'hbb5d1bd8),
	.w5(32'hbb1d66b1),
	.w6(32'h3c0ec7c7),
	.w7(32'hbb5dd08f),
	.w8(32'h3a89d2db),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c70bf23),
	.w1(32'hbb660ac2),
	.w2(32'hbb3ced26),
	.w3(32'h3c0736ec),
	.w4(32'hbbdd4448),
	.w5(32'hbb66c13b),
	.w6(32'h3c621948),
	.w7(32'hbbbb096b),
	.w8(32'h3ab23b7f),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c486268),
	.w1(32'h3b248756),
	.w2(32'h3c0ac7ba),
	.w3(32'h3c03ebc0),
	.w4(32'hbb013b24),
	.w5(32'h3b6c8dd5),
	.w6(32'h3c178261),
	.w7(32'hbb125188),
	.w8(32'h3b99f236),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6124c4),
	.w1(32'h3a771ed8),
	.w2(32'hbaead4b0),
	.w3(32'h3b6c9b7d),
	.w4(32'h39d67f33),
	.w5(32'hbacc6a69),
	.w6(32'h3b9e0094),
	.w7(32'hb951050d),
	.w8(32'h3a479453),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5b8af9),
	.w1(32'h3aad5b6b),
	.w2(32'h3c21f63b),
	.w3(32'h3c0310e4),
	.w4(32'hbb48e3ff),
	.w5(32'h3b4ac3d8),
	.w6(32'h3c1ed838),
	.w7(32'hbb2e57b5),
	.w8(32'h3b93640c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8179a2),
	.w1(32'h3627d615),
	.w2(32'h3bb1ba97),
	.w3(32'h3b922f30),
	.w4(32'hba2dabb4),
	.w5(32'h3b329771),
	.w6(32'h3b81c618),
	.w7(32'hba134bcf),
	.w8(32'h3a9a1a63),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c882add),
	.w1(32'h3aa2cb22),
	.w2(32'h3c612c35),
	.w3(32'h3c604f46),
	.w4(32'hbb4592fc),
	.w5(32'h3c096b23),
	.w6(32'h3bebc1a3),
	.w7(32'hbbcb6cbe),
	.w8(32'h3b71d1bb),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61a339),
	.w1(32'h3ac8c404),
	.w2(32'h3abbf93b),
	.w3(32'hb9d3cbb1),
	.w4(32'h3a874c5f),
	.w5(32'h3a8d0a74),
	.w6(32'h3a647e8a),
	.w7(32'h3aae7630),
	.w8(32'h3aa23019),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a5a92),
	.w1(32'hba13ed47),
	.w2(32'hb9b2a577),
	.w3(32'h3acff728),
	.w4(32'hba0c6dd0),
	.w5(32'hb9a083bc),
	.w6(32'hb7e5bf09),
	.w7(32'hb9331d0f),
	.w8(32'hba1120bd),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39ba98),
	.w1(32'h39b07dc4),
	.w2(32'h3beb0c31),
	.w3(32'h3bfc112a),
	.w4(32'hbae9ae7f),
	.w5(32'h3ba35557),
	.w6(32'h3be37a1f),
	.w7(32'hbb581f68),
	.w8(32'h3bc1b098),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d2b77),
	.w1(32'hbb78a49f),
	.w2(32'h3c0d7378),
	.w3(32'h3c2e0f55),
	.w4(32'hbb81bf15),
	.w5(32'h3c2024ec),
	.w6(32'h3bd6f914),
	.w7(32'hbbefa55c),
	.w8(32'h3b56859e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73fd83),
	.w1(32'h3b06414f),
	.w2(32'h3c2104a8),
	.w3(32'h3bfb596c),
	.w4(32'hbb841a1b),
	.w5(32'h3b5d1917),
	.w6(32'h3c083b59),
	.w7(32'hbbd22cc3),
	.w8(32'h390bcd83),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50a9b8),
	.w1(32'h3ac91484),
	.w2(32'h3acf7caa),
	.w3(32'h3bb7ed77),
	.w4(32'h3bf5d3ae),
	.w5(32'h3a9e1a70),
	.w6(32'hba8c04dc),
	.w7(32'h3a958959),
	.w8(32'h3bbcd058),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8f854),
	.w1(32'hb90881f4),
	.w2(32'h37629a68),
	.w3(32'h39cb3bee),
	.w4(32'h39eb842f),
	.w5(32'h395f818d),
	.w6(32'h38b2af92),
	.w7(32'h39c75e17),
	.w8(32'h39285de4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab14df0),
	.w1(32'h3abe7e1f),
	.w2(32'h3a0d4b9e),
	.w3(32'h3ab60dbc),
	.w4(32'h3ac79ec0),
	.w5(32'h3a2a9541),
	.w6(32'h3b077e81),
	.w7(32'h3a7bf878),
	.w8(32'h396044cf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ed960),
	.w1(32'hbb3059a5),
	.w2(32'h3bb82fac),
	.w3(32'h3a23b373),
	.w4(32'h3bb1f097),
	.w5(32'h3c3dc3b0),
	.w6(32'hbb7053c6),
	.w7(32'hbb3eed48),
	.w8(32'h3bf9f8e3),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a3931),
	.w1(32'h3baa6e24),
	.w2(32'h3c55e273),
	.w3(32'h3c46cd0e),
	.w4(32'h3b7fc784),
	.w5(32'h3c567582),
	.w6(32'h3bde52b6),
	.w7(32'h3b3c975b),
	.w8(32'h3c0e2b0e),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11db86),
	.w1(32'h3aa06284),
	.w2(32'h3bb3bac0),
	.w3(32'h3b89316b),
	.w4(32'h3b685b65),
	.w5(32'h3bc08fde),
	.w6(32'hbb67be46),
	.w7(32'hbaa6faf8),
	.w8(32'h3b950016),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf473f3),
	.w1(32'hbbe8e32a),
	.w2(32'hbb268a3a),
	.w3(32'h3bb76f2f),
	.w4(32'hbc0b3cd1),
	.w5(32'hbb869212),
	.w6(32'h3bf92f0b),
	.w7(32'hbbe1a1fe),
	.w8(32'hbae76812),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3de92f),
	.w1(32'h3984c6a6),
	.w2(32'h3bf5bc04),
	.w3(32'h3c0c0ee3),
	.w4(32'hbb8cec59),
	.w5(32'h3ab6a33c),
	.w6(32'h3c14d606),
	.w7(32'hbbaf21e1),
	.w8(32'h3aee0958),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d097d),
	.w1(32'h37f9c71e),
	.w2(32'h3a7ea19f),
	.w3(32'hb98a4a6c),
	.w4(32'hba20e93b),
	.w5(32'hb91260be),
	.w6(32'hb9c73953),
	.w7(32'h37d06ec1),
	.w8(32'hb90a618c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4552c),
	.w1(32'hb9ae9d18),
	.w2(32'hbaa6bbd8),
	.w3(32'hb98dc209),
	.w4(32'h3aa62481),
	.w5(32'hb7b281b6),
	.w6(32'hb9e06530),
	.w7(32'h3899bef3),
	.w8(32'h3a563cf2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7c184),
	.w1(32'hbae02b6d),
	.w2(32'h39549fa2),
	.w3(32'h3a6f31a3),
	.w4(32'h381fd932),
	.w5(32'h3aed418a),
	.w6(32'hba9909ac),
	.w7(32'h3b188632),
	.w8(32'hb981572f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7df9b8),
	.w1(32'h38cfc531),
	.w2(32'hbab1f44d),
	.w3(32'hba957346),
	.w4(32'hb9abe321),
	.w5(32'hba6d6e3a),
	.w6(32'hba87de8a),
	.w7(32'hbb072d91),
	.w8(32'hbae7483b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9228fb),
	.w1(32'h3b3bb7ba),
	.w2(32'h3b7c311a),
	.w3(32'hba8534aa),
	.w4(32'h3adeb8d4),
	.w5(32'h3b6a232e),
	.w6(32'h399fa3d1),
	.w7(32'h3b09559f),
	.w8(32'h3b665dd5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c221564),
	.w1(32'h38da1ac0),
	.w2(32'h3bda2ff0),
	.w3(32'h3bb78dfd),
	.w4(32'hbb28cd9a),
	.w5(32'h3bc082f2),
	.w6(32'h3b791c4b),
	.w7(32'hbb619807),
	.w8(32'h3b63d022),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c109a25),
	.w1(32'h3a56238c),
	.w2(32'h3bdb3e79),
	.w3(32'h3bfa4fe9),
	.w4(32'hba882ce3),
	.w5(32'h3b9935aa),
	.w6(32'h3ba030b7),
	.w7(32'h3a4ffa5f),
	.w8(32'h3ab34662),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15e932),
	.w1(32'h39ec6481),
	.w2(32'hba9a3761),
	.w3(32'hbaa0340e),
	.w4(32'h3a36a256),
	.w5(32'hb99a52a9),
	.w6(32'h3a405717),
	.w7(32'h3a91cd7f),
	.w8(32'h3a6d7300),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a836cd3),
	.w1(32'h3adf133b),
	.w2(32'h3c2957c5),
	.w3(32'h3b86e59f),
	.w4(32'h3b73f18c),
	.w5(32'h3c4bd162),
	.w6(32'hbaf16dc8),
	.w7(32'hbb4a6a7f),
	.w8(32'h3c2e72de),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25813e),
	.w1(32'h3ab0741c),
	.w2(32'h3b8bc048),
	.w3(32'h3b2a8bac),
	.w4(32'h3a8b25c8),
	.w5(32'h3b699401),
	.w6(32'h3a97459b),
	.w7(32'h39af78b0),
	.w8(32'h3b338efa),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f261c),
	.w1(32'h3a78b2cb),
	.w2(32'h38feb9e2),
	.w3(32'h3ab877c7),
	.w4(32'h3a9356fa),
	.w5(32'h39b80371),
	.w6(32'h3aad0ecf),
	.w7(32'h3a23f6ca),
	.w8(32'h3a433f72),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b142a60),
	.w1(32'h3abe64fb),
	.w2(32'h3b78bf78),
	.w3(32'h3b12a9a0),
	.w4(32'h3aaa96af),
	.w5(32'h3b680444),
	.w6(32'h3a8e4bbe),
	.w7(32'h39cf6453),
	.w8(32'h3b3f677e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f73da0),
	.w1(32'hb6f0aea6),
	.w2(32'h39decbfc),
	.w3(32'hb9e4771d),
	.w4(32'hba5ba700),
	.w5(32'hba612ea1),
	.w6(32'hb9816a37),
	.w7(32'hb9a253cb),
	.w8(32'h38455a2b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab91e53),
	.w1(32'hba940d4b),
	.w2(32'hba7da112),
	.w3(32'hb9056bfe),
	.w4(32'hba95d060),
	.w5(32'hba30de1a),
	.w6(32'h39a781d8),
	.w7(32'h3987b0f5),
	.w8(32'h3a1887dc),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b21ae),
	.w1(32'h3a537dc3),
	.w2(32'h39e04e53),
	.w3(32'hba1eb6a4),
	.w4(32'h3a5328c7),
	.w5(32'h3a39f268),
	.w6(32'h3a5adeb5),
	.w7(32'h3a319025),
	.w8(32'h3a4b8ba5),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e6d462),
	.w1(32'h3a904c04),
	.w2(32'h39b8f405),
	.w3(32'h3a1b4284),
	.w4(32'h397cb723),
	.w5(32'hb940cbce),
	.w6(32'h3a7c27a1),
	.w7(32'h3a01c96b),
	.w8(32'h3a305da1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2a4da),
	.w1(32'h3abd6b4a),
	.w2(32'h3b361037),
	.w3(32'h3ba00b15),
	.w4(32'h3a9834a0),
	.w5(32'h3b138ba2),
	.w6(32'h3be37b92),
	.w7(32'h3a743cf2),
	.w8(32'h3ae63ef6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2dfbb),
	.w1(32'h3bbb930d),
	.w2(32'h3c75d0ce),
	.w3(32'h3bcdb584),
	.w4(32'h3b4f7dd0),
	.w5(32'h3c00cb1e),
	.w6(32'h3be7dd90),
	.w7(32'hb96dd69c),
	.w8(32'h3bd85715),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d516b),
	.w1(32'h3abe066c),
	.w2(32'h3be127ab),
	.w3(32'h3b19880a),
	.w4(32'h398f56a8),
	.w5(32'h3bbd5539),
	.w6(32'h3acba26d),
	.w7(32'hbacd7011),
	.w8(32'h3b5c2fa0),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becee82),
	.w1(32'h3b5e4aa8),
	.w2(32'h3c57da5c),
	.w3(32'h3bed2c75),
	.w4(32'h3b35b3e1),
	.w5(32'h3c24773a),
	.w6(32'h3b9fbe2d),
	.w7(32'h3b7a9983),
	.w8(32'h3c17126d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b006546),
	.w1(32'h3a5e6584),
	.w2(32'h397d62a0),
	.w3(32'h3acf7c44),
	.w4(32'h39896051),
	.w5(32'hba1411fd),
	.w6(32'h3ac23e5a),
	.w7(32'hb774294a),
	.w8(32'h39b31aa7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3936357d),
	.w1(32'h3b15eaca),
	.w2(32'h3aa19f43),
	.w3(32'h39dbf8cf),
	.w4(32'h3b00ca39),
	.w5(32'h3aa0afa8),
	.w6(32'h3ac1dce8),
	.w7(32'h3ab171df),
	.w8(32'h3aa848a1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4fe884),
	.w1(32'h3a7e8673),
	.w2(32'h3a1cd75e),
	.w3(32'h3a775744),
	.w4(32'h3a910b08),
	.w5(32'h3a866d0e),
	.w6(32'h3a6d89aa),
	.w7(32'h3a64afc1),
	.w8(32'h3a8523c2),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3532ff),
	.w1(32'h3a4aa907),
	.w2(32'h39a4a9bb),
	.w3(32'h3a6e4aa5),
	.w4(32'h3a73229d),
	.w5(32'h3a44d65d),
	.w6(32'h3a42974f),
	.w7(32'h3a0f7923),
	.w8(32'h3a60b99e),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b118a),
	.w1(32'h3ab370e9),
	.w2(32'h3bf7e7a2),
	.w3(32'h3bfdb76e),
	.w4(32'hb9b52dd9),
	.w5(32'h3b937a93),
	.w6(32'h3bce904a),
	.w7(32'h3aaf5dca),
	.w8(32'h3bdb9925),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b183056),
	.w1(32'h3952307b),
	.w2(32'h3a86a49e),
	.w3(32'h3a3a5176),
	.w4(32'hb9990668),
	.w5(32'h3a96850d),
	.w6(32'hba022a3e),
	.w7(32'h3a62f991),
	.w8(32'hb99c3d05),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86fd7a),
	.w1(32'hbb2e475c),
	.w2(32'hb992e7d4),
	.w3(32'h3ae5e756),
	.w4(32'hbb6531ca),
	.w5(32'hbac804ba),
	.w6(32'h3b4a816a),
	.w7(32'hbb0112ab),
	.w8(32'h3a657702),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e4bf9),
	.w1(32'hb9a5b77c),
	.w2(32'h3a0a7626),
	.w3(32'h3b36a0c4),
	.w4(32'hba090c88),
	.w5(32'hba14a510),
	.w6(32'h3b1d967c),
	.w7(32'hba19b610),
	.w8(32'hba63ad24),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81a366),
	.w1(32'h3abda129),
	.w2(32'h3ad162ba),
	.w3(32'hba09a1a6),
	.w4(32'h3ab1ad6e),
	.w5(32'h3ad7df47),
	.w6(32'h3aba146d),
	.w7(32'h3ac6c7d7),
	.w8(32'h3ad29fc3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e03d6),
	.w1(32'h3a0ac2e2),
	.w2(32'h3a847659),
	.w3(32'h3b6a9fcd),
	.w4(32'h3b0f807d),
	.w5(32'h3b074906),
	.w6(32'h39c455bc),
	.w7(32'h3a9f467f),
	.w8(32'h3b406fc6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adf9be6),
	.w1(32'h3a8b4c8d),
	.w2(32'h3978b726),
	.w3(32'h3a8b5fd9),
	.w4(32'h3aad91d9),
	.w5(32'h39cfdafc),
	.w6(32'h3a91b607),
	.w7(32'h3a24f169),
	.w8(32'h3a802b04),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f8df9),
	.w1(32'h3bb0e799),
	.w2(32'h3c80222e),
	.w3(32'h3c0192e0),
	.w4(32'h3aff6886),
	.w5(32'h3bd834c2),
	.w6(32'h3c080602),
	.w7(32'h3adc34a9),
	.w8(32'h3baa3f13),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c1860),
	.w1(32'hba2ac75b),
	.w2(32'hb9f7081c),
	.w3(32'hb9beb589),
	.w4(32'hba210c7f),
	.w5(32'hb9d8bfc1),
	.w6(32'hba2ed3cc),
	.w7(32'hba2816cc),
	.w8(32'hb89b85fa),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04fbda),
	.w1(32'hbbbec4dd),
	.w2(32'hbbbfae2c),
	.w3(32'h3c06fe0e),
	.w4(32'hbb975bce),
	.w5(32'hbbe62938),
	.w6(32'h3c349eae),
	.w7(32'hbb78a462),
	.w8(32'hbb5cf96a),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule