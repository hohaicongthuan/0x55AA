module layer_10_featuremap_365(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd8a66),
	.w1(32'h3bd0fb7a),
	.w2(32'hb90de661),
	.w3(32'hbb28271e),
	.w4(32'hba5d6874),
	.w5(32'h3c4e2db6),
	.w6(32'hbc29e52a),
	.w7(32'h3ba3fea0),
	.w8(32'h3b69b123),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1496ae),
	.w1(32'hbc7695ba),
	.w2(32'hbc5402ee),
	.w3(32'h3b87301b),
	.w4(32'h3bb7b3b5),
	.w5(32'h3b669c34),
	.w6(32'h3c54c45c),
	.w7(32'h3b4eefdf),
	.w8(32'h3c0bb990),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4ac08),
	.w1(32'h3b4f811f),
	.w2(32'h3a0f8742),
	.w3(32'h3b72409f),
	.w4(32'h3c3ca209),
	.w5(32'hbbb1654c),
	.w6(32'hbd8a2aa6),
	.w7(32'h3b7b3056),
	.w8(32'h3be8df99),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53945c),
	.w1(32'hbd02c985),
	.w2(32'h3b2e55e7),
	.w3(32'h3cd5e02d),
	.w4(32'h3bbbf379),
	.w5(32'hbb206a86),
	.w6(32'hbb86d7fe),
	.w7(32'h3b9d665d),
	.w8(32'hbbc10c7e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e6ba1),
	.w1(32'hbc4c37b0),
	.w2(32'hbb178417),
	.w3(32'hbc8c04d8),
	.w4(32'h3bcb5b77),
	.w5(32'hb93a6f48),
	.w6(32'hbc2499f2),
	.w7(32'h39c828bf),
	.w8(32'hbd8b3620),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8abef),
	.w1(32'hb92961ef),
	.w2(32'hbb45e353),
	.w3(32'hbb6de12f),
	.w4(32'h3a10b923),
	.w5(32'h3bf12796),
	.w6(32'hbb2e7888),
	.w7(32'hbc812ac0),
	.w8(32'hbb5ee080),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1fedaf),
	.w1(32'hbc23f5d3),
	.w2(32'hbae5c233),
	.w3(32'h3cc4c2f5),
	.w4(32'h3ce1c74a),
	.w5(32'hbc5be722),
	.w6(32'h3a9dfb85),
	.w7(32'h3bda9fdc),
	.w8(32'hbbd12f11),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a61205c),
	.w1(32'h3b812459),
	.w2(32'hbb0ec6bd),
	.w3(32'h3be349d8),
	.w4(32'hbc000fd0),
	.w5(32'h3b8dd4d0),
	.w6(32'hbcb6455e),
	.w7(32'h3a95ec3c),
	.w8(32'h38b0c9f8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5f4a4),
	.w1(32'hbbb9c28f),
	.w2(32'h3ac6f911),
	.w3(32'hba841ffd),
	.w4(32'h39b7264f),
	.w5(32'h3b1f6f1f),
	.w6(32'h3b9f1f00),
	.w7(32'h3b0d8ef6),
	.w8(32'h3b8d337f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1ccc6b),
	.w1(32'hbb3a1df4),
	.w2(32'hb900d590),
	.w3(32'hbc5e029e),
	.w4(32'hbb11db98),
	.w5(32'h3b51a319),
	.w6(32'h3af1cbfa),
	.w7(32'h3b069a00),
	.w8(32'h3bb683db),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd29134),
	.w1(32'hbbc3be1c),
	.w2(32'hbb88d834),
	.w3(32'hb93c9697),
	.w4(32'h3a83db14),
	.w5(32'h3cdaaa26),
	.w6(32'h3bd19cd5),
	.w7(32'hbaa4b3a6),
	.w8(32'h3ae22f3f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84dfac),
	.w1(32'hbb89bb22),
	.w2(32'h3d4ff0a8),
	.w3(32'h3c5d6fbf),
	.w4(32'h3d3755b0),
	.w5(32'h3ab23d75),
	.w6(32'h3bbd9397),
	.w7(32'hb89f6f19),
	.w8(32'h3bd138f6),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35b770),
	.w1(32'h3bb584e4),
	.w2(32'hbbc2a936),
	.w3(32'h3af7f32e),
	.w4(32'hbb9c8f42),
	.w5(32'hbcad4738),
	.w6(32'hbc1c39ba),
	.w7(32'hbc003e9c),
	.w8(32'hbd041515),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26e59),
	.w1(32'h3d320a82),
	.w2(32'hbc0e0fef),
	.w3(32'hbbfa8412),
	.w4(32'hbd49dd50),
	.w5(32'h3c08db2e),
	.w6(32'h3c1aa456),
	.w7(32'h3b914811),
	.w8(32'h3ca7e820),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc91552f),
	.w1(32'hbb578cc0),
	.w2(32'hbbbe4972),
	.w3(32'h3ae95676),
	.w4(32'h3b7867fc),
	.w5(32'hbb4c51bf),
	.w6(32'hbb129624),
	.w7(32'h3bac0d89),
	.w8(32'hbad0958b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb06381),
	.w1(32'h3adfd8e0),
	.w2(32'hbba2df67),
	.w3(32'h3c9afff6),
	.w4(32'hbafe89bb),
	.w5(32'h3bda834e),
	.w6(32'hbc11c244),
	.w7(32'hbc037d76),
	.w8(32'h3b6d848a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8874af),
	.w1(32'h39825f2b),
	.w2(32'hbbccb053),
	.w3(32'hbacae459),
	.w4(32'h3a79fc87),
	.w5(32'h3b58ab84),
	.w6(32'hbb41b3bc),
	.w7(32'hb9ac46ec),
	.w8(32'h3b6df7c9),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e78b4),
	.w1(32'hbb0114f9),
	.w2(32'hbbfe0582),
	.w3(32'hbc737675),
	.w4(32'hbb2b5d67),
	.w5(32'h3ba153fb),
	.w6(32'hbb296cbe),
	.w7(32'hbc2422f5),
	.w8(32'hbaa3537f),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4360fc),
	.w1(32'hbbcbee97),
	.w2(32'h3a71320c),
	.w3(32'hbbcccb77),
	.w4(32'hba1ac189),
	.w5(32'hbd5a2815),
	.w6(32'hba0c43b8),
	.w7(32'h3bdecf0b),
	.w8(32'hba1809b7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7afbdd),
	.w1(32'h3c8af6f6),
	.w2(32'hbad68fcb),
	.w3(32'h3a9d63ff),
	.w4(32'h3d6225bd),
	.w5(32'hbb6516be),
	.w6(32'h3bffd9a6),
	.w7(32'hbbad4b24),
	.w8(32'h3c01eef6),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a1892),
	.w1(32'h3b86b0ea),
	.w2(32'h3c85b007),
	.w3(32'hbb212c40),
	.w4(32'hbb03d95c),
	.w5(32'h3ba7ae35),
	.w6(32'h3b88972e),
	.w7(32'hbc87d66d),
	.w8(32'h3bdae2c1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24ecb0),
	.w1(32'h3c2e9c0d),
	.w2(32'h3b832147),
	.w3(32'hb9a05795),
	.w4(32'h3b7a4854),
	.w5(32'hbc16ed4e),
	.w6(32'hbd3975ff),
	.w7(32'h3b727eb8),
	.w8(32'hbbb5ee6b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0cb3),
	.w1(32'h3ab1eb59),
	.w2(32'hbd942e96),
	.w3(32'h3c0b6e8c),
	.w4(32'h3b43b356),
	.w5(32'hbbe4bc8c),
	.w6(32'h3b3d9060),
	.w7(32'hbbe0ec5d),
	.w8(32'h3c80c0c8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093787),
	.w1(32'hbab68d93),
	.w2(32'h3b663cad),
	.w3(32'h3af2f7a3),
	.w4(32'hb9bc772b),
	.w5(32'h3b4e98ff),
	.w6(32'h3c09a00d),
	.w7(32'hbcd4d649),
	.w8(32'h3b1c8d54),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59e0e5),
	.w1(32'hb9bfbdef),
	.w2(32'h3c02cfa5),
	.w3(32'hbb16a64e),
	.w4(32'h3bc540f9),
	.w5(32'h3ba1abcc),
	.w6(32'hbb25130d),
	.w7(32'h3beb148c),
	.w8(32'h3c039fd1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb92780),
	.w1(32'hbb35c405),
	.w2(32'h399ef664),
	.w3(32'h3bd0fa9c),
	.w4(32'h3bfdaa75),
	.w5(32'h3be3e91e),
	.w6(32'hbb8fbd6a),
	.w7(32'h3a364a41),
	.w8(32'h3b3d1644),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d8d3d),
	.w1(32'hbcaddf90),
	.w2(32'h3b84592e),
	.w3(32'h3aa21740),
	.w4(32'hba124e87),
	.w5(32'hbb384038),
	.w6(32'h3bc83fbb),
	.w7(32'h3a99a5d8),
	.w8(32'h3b2d9d07),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21be78),
	.w1(32'hbb28e968),
	.w2(32'hbca700f1),
	.w3(32'hbc0b3b36),
	.w4(32'h3b40e945),
	.w5(32'hbb4864a5),
	.w6(32'hbbc737cf),
	.w7(32'hbca26f43),
	.w8(32'h3a5331d6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae9902),
	.w1(32'hba81817c),
	.w2(32'hbcd29879),
	.w3(32'hba819f3a),
	.w4(32'hbb47af12),
	.w5(32'hbb8fb568),
	.w6(32'hbb64ab55),
	.w7(32'hbb9b549b),
	.w8(32'h3aa0968f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384936),
	.w1(32'hba39ff2e),
	.w2(32'h3c41674d),
	.w3(32'h3a14d0fa),
	.w4(32'h3b1178c9),
	.w5(32'hbc72b76b),
	.w6(32'h3be93f55),
	.w7(32'hbc4c7ca8),
	.w8(32'h3a975007),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba779420),
	.w1(32'hba764689),
	.w2(32'hb92d7449),
	.w3(32'hbbacb2d9),
	.w4(32'h3ba8fa30),
	.w5(32'hb971a30b),
	.w6(32'h3aa34a29),
	.w7(32'h3b49a4b4),
	.w8(32'hb9998b8f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6a6b2),
	.w1(32'h3b91a339),
	.w2(32'hbb0c5806),
	.w3(32'hba8e780a),
	.w4(32'hbc17fe9a),
	.w5(32'hbd29439c),
	.w6(32'hbc18c341),
	.w7(32'h3b70cfda),
	.w8(32'hbc63ff8b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88e279),
	.w1(32'hbc1ce4f7),
	.w2(32'hbc345c58),
	.w3(32'h3bb822df),
	.w4(32'hbb3ce70f),
	.w5(32'hbc5a30b8),
	.w6(32'h3a1d1f98),
	.w7(32'hbd12f187),
	.w8(32'hba53b8e8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094a91),
	.w1(32'hbd44e3ca),
	.w2(32'hbb97653d),
	.w3(32'h3b93156e),
	.w4(32'h3be3c918),
	.w5(32'hba64b8a5),
	.w6(32'h3aaabae8),
	.w7(32'h3c0da8b3),
	.w8(32'hbb47ec4b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fd42a),
	.w1(32'h3bc539fe),
	.w2(32'h398a034b),
	.w3(32'h3b9b0715),
	.w4(32'hb91bd351),
	.w5(32'hbc119c63),
	.w6(32'h3c18cc64),
	.w7(32'hbc18f0f8),
	.w8(32'h3ca0a616),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23739b),
	.w1(32'hbc119374),
	.w2(32'h3c353399),
	.w3(32'hbb3d92fe),
	.w4(32'h39a1b0bc),
	.w5(32'h3b59478c),
	.w6(32'h3b4604e2),
	.w7(32'h3afad02a),
	.w8(32'hbc896b51),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f10b),
	.w1(32'h3abde881),
	.w2(32'hbc7fe14e),
	.w3(32'h3b9a3126),
	.w4(32'h39a92f19),
	.w5(32'h3ca4b934),
	.w6(32'hba34f468),
	.w7(32'hbabe6e9a),
	.w8(32'hbc5a9402),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc032346),
	.w1(32'h3b4a6565),
	.w2(32'hbd42ff3b),
	.w3(32'h3aaa42c8),
	.w4(32'hbb477ff7),
	.w5(32'hbb390261),
	.w6(32'hba8a3fde),
	.w7(32'h3c0d6bd1),
	.w8(32'h3981b3ad),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398f16fb),
	.w1(32'hb9dc8dfe),
	.w2(32'hbc0e473f),
	.w3(32'hbca0314a),
	.w4(32'hbac7ff15),
	.w5(32'hbc70859c),
	.w6(32'h3c163837),
	.w7(32'h3b40a34d),
	.w8(32'hbb604b76),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a810524),
	.w1(32'hbbc99e70),
	.w2(32'hbbd86304),
	.w3(32'hbb1cce3e),
	.w4(32'h3b7ae087),
	.w5(32'h3b890af9),
	.w6(32'hbc19356d),
	.w7(32'h3c2d4d50),
	.w8(32'h3ced7c8e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df9df9),
	.w1(32'h3c1eb13c),
	.w2(32'h3c512206),
	.w3(32'hbb3da422),
	.w4(32'hba7c2fa9),
	.w5(32'h3a783bfd),
	.w6(32'h3abdf932),
	.w7(32'h3ba44ceb),
	.w8(32'hbaf81200),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd587d1),
	.w1(32'h3b793a16),
	.w2(32'h3ab36dc9),
	.w3(32'h3b9fd00f),
	.w4(32'h3adda3a7),
	.w5(32'h3c0e56e0),
	.w6(32'hbbfacb78),
	.w7(32'h3c06565f),
	.w8(32'h3c2bf707),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02905e),
	.w1(32'h39aaa597),
	.w2(32'hbbba2154),
	.w3(32'h3b49a0c2),
	.w4(32'h3bea6191),
	.w5(32'h3ab3e0d8),
	.w6(32'hbbc7a834),
	.w7(32'h3a79ec4a),
	.w8(32'hb8fe8142),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd42514),
	.w1(32'hba0b74c4),
	.w2(32'h3a26521c),
	.w3(32'hb9a44197),
	.w4(32'h3bd0601f),
	.w5(32'hba848cbd),
	.w6(32'hbbd32c32),
	.w7(32'h3c899d7d),
	.w8(32'hb9a38398),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949b70a),
	.w1(32'hbd070954),
	.w2(32'h3b05fbc1),
	.w3(32'h3c235035),
	.w4(32'h3bafcd63),
	.w5(32'hbc38f104),
	.w6(32'h3b08ecec),
	.w7(32'h3b01a840),
	.w8(32'h39fc7080),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c9a9f),
	.w1(32'h3ac68e43),
	.w2(32'h3b9ce2d9),
	.w3(32'h3be2979c),
	.w4(32'h3b66c04a),
	.w5(32'h3b0e9a2f),
	.w6(32'h3b8ec3f1),
	.w7(32'hbb42d50d),
	.w8(32'hbcb32c51),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf9750c),
	.w1(32'h3ba501c7),
	.w2(32'hbb4a996a),
	.w3(32'hbd09f052),
	.w4(32'h38e6b729),
	.w5(32'h3af5dd35),
	.w6(32'hbad0cb9d),
	.w7(32'hbad0251b),
	.w8(32'h39aa11ec),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ff717),
	.w1(32'hba9eff20),
	.w2(32'h3c4a3b01),
	.w3(32'hba20441e),
	.w4(32'h3bd3930f),
	.w5(32'h3b4ff74f),
	.w6(32'h3b98e84b),
	.w7(32'h3b9b74ac),
	.w8(32'h3d2c84ea),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14aa04),
	.w1(32'hbbec5536),
	.w2(32'hbc1fa36c),
	.w3(32'h3a914445),
	.w4(32'hbb17fee7),
	.w5(32'h3c31309e),
	.w6(32'h3bc060e0),
	.w7(32'h3addf4d3),
	.w8(32'h3b9d38c4),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84bebc),
	.w1(32'hbb9259bb),
	.w2(32'hbd542c72),
	.w3(32'h3c890968),
	.w4(32'hbcdf8ed8),
	.w5(32'h3be577c5),
	.w6(32'h3bbe3f9f),
	.w7(32'hbb8c1b8d),
	.w8(32'hbabc9a4a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a662e01),
	.w1(32'h3bce8f1f),
	.w2(32'h3b4eb74d),
	.w3(32'h3b005ad5),
	.w4(32'hbb607262),
	.w5(32'hb95de75b),
	.w6(32'h3b907e43),
	.w7(32'hbb191f00),
	.w8(32'hbaeee790),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d35c6),
	.w1(32'hbc3c0915),
	.w2(32'h3b097485),
	.w3(32'hbd7f6f0c),
	.w4(32'hbd092903),
	.w5(32'hbb5ab821),
	.w6(32'h3cc25c73),
	.w7(32'h3bae52ee),
	.w8(32'h3b5a66cd),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cc64f),
	.w1(32'h3c0dcec8),
	.w2(32'h3bc935bd),
	.w3(32'h3c54fd2e),
	.w4(32'h3a17cf03),
	.w5(32'hbb896dc9),
	.w6(32'h3bc1a0dd),
	.w7(32'hbb02c2f9),
	.w8(32'hbb544f77),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09ce4e),
	.w1(32'hbd6e2938),
	.w2(32'hbb6b0ad2),
	.w3(32'h3c0ab5bd),
	.w4(32'hbc843e95),
	.w5(32'h3ae505cb),
	.w6(32'hba17188e),
	.w7(32'hbbefd38a),
	.w8(32'h3c258468),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f9205),
	.w1(32'h3b044f56),
	.w2(32'h3b027e4f),
	.w3(32'hbb37145e),
	.w4(32'h3998325a),
	.w5(32'h3b97d996),
	.w6(32'hbbe58e79),
	.w7(32'h3bbc6af0),
	.w8(32'hbadcbc5a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aaefa),
	.w1(32'hbc0d9608),
	.w2(32'h3b1f12b0),
	.w3(32'h3beec4fa),
	.w4(32'hbc23cc00),
	.w5(32'hbc2011c8),
	.w6(32'hbb0edff8),
	.w7(32'hbb218720),
	.w8(32'hbb1f3f32),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8649e3),
	.w1(32'hbaa066bb),
	.w2(32'h3d047835),
	.w3(32'hbb19a1cf),
	.w4(32'h3c755af3),
	.w5(32'hbbc3aff7),
	.w6(32'hba8d7c33),
	.w7(32'h3a4f6cc3),
	.w8(32'h3bece66e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09dfef),
	.w1(32'hbb0eb282),
	.w2(32'h3c0cf126),
	.w3(32'h3be334f8),
	.w4(32'h3c9ea775),
	.w5(32'h39c18f03),
	.w6(32'h3b114493),
	.w7(32'hbc038954),
	.w8(32'hbc2adee4),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b051331),
	.w1(32'h3bae3d48),
	.w2(32'hbab68685),
	.w3(32'hbb129a52),
	.w4(32'h3be36685),
	.w5(32'hbb553e72),
	.w6(32'h3c4e6bc8),
	.w7(32'hbae6d073),
	.w8(32'h3bec8994),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13fcfc),
	.w1(32'hbc51af0c),
	.w2(32'hbc6fd5d1),
	.w3(32'hbbb53aa6),
	.w4(32'h3aeef7ba),
	.w5(32'h39f78032),
	.w6(32'h3ab9e5e2),
	.w7(32'hbc90d089),
	.w8(32'hbb83bee5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3276d1),
	.w1(32'hba205e35),
	.w2(32'hbab678a9),
	.w3(32'hbbd3c14b),
	.w4(32'hbbae12b0),
	.w5(32'h39720ba9),
	.w6(32'h3b4a1321),
	.w7(32'hbc5c12e1),
	.w8(32'h3bed1afd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c380373),
	.w1(32'hbbc77d03),
	.w2(32'h3ab269a9),
	.w3(32'h3a9991ec),
	.w4(32'hbbd31b49),
	.w5(32'h3b0f55e0),
	.w6(32'h3c236363),
	.w7(32'hba00bb2d),
	.w8(32'hbc0a8240),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57987c),
	.w1(32'hba023b18),
	.w2(32'h3c75ca5b),
	.w3(32'hba61d216),
	.w4(32'hbbb1716f),
	.w5(32'h3bcbc421),
	.w6(32'hbc602af8),
	.w7(32'hbb241783),
	.w8(32'hbb377f6f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc782a34),
	.w1(32'h3ce61a8e),
	.w2(32'hbbe7f198),
	.w3(32'hbba8ed47),
	.w4(32'hbc6f9adb),
	.w5(32'hba091fb4),
	.w6(32'hbc7aebee),
	.w7(32'h3a68183d),
	.w8(32'hbc169eff),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf18e8f),
	.w1(32'h3b4d84cd),
	.w2(32'hbb8ce12e),
	.w3(32'h3b181f1f),
	.w4(32'hbc4f4dca),
	.w5(32'hbb178e3f),
	.w6(32'hba9c6ac0),
	.w7(32'hbb7ba90b),
	.w8(32'hbc31bcf0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a89d5),
	.w1(32'hbcb1aba3),
	.w2(32'h3c15cc99),
	.w3(32'hbb9d59ee),
	.w4(32'h3b3185fc),
	.w5(32'hbaf78aa6),
	.w6(32'h3ba2cf11),
	.w7(32'hba852a99),
	.w8(32'h3bd2a8a4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b6581),
	.w1(32'hbbeb7c28),
	.w2(32'h3b08600d),
	.w3(32'h3c358b4f),
	.w4(32'h3ab05a47),
	.w5(32'hba4ba6a7),
	.w6(32'hb9c134bc),
	.w7(32'hbbbcba8c),
	.w8(32'h3c705a24),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba08634),
	.w1(32'h3b09b3bf),
	.w2(32'hbbddc148),
	.w3(32'hbc26c25e),
	.w4(32'hbb117d3e),
	.w5(32'hbc07a43e),
	.w6(32'h3cdabfec),
	.w7(32'h3b199195),
	.w8(32'h3b98d68e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd196d),
	.w1(32'h3ca7ac03),
	.w2(32'h3ab3c7c2),
	.w3(32'hbb348502),
	.w4(32'hb8860372),
	.w5(32'h3b17e3dd),
	.w6(32'hbb673b14),
	.w7(32'hbc8cf9df),
	.w8(32'h390955fa),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8ee60),
	.w1(32'h3c1bfa6e),
	.w2(32'h3bedf37e),
	.w3(32'hbb082d43),
	.w4(32'hbbf655a1),
	.w5(32'h3b420bf9),
	.w6(32'h3c1c8a27),
	.w7(32'hbbb89bdb),
	.w8(32'h3a827b3f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddfcfc),
	.w1(32'hbb453ad1),
	.w2(32'hbc37bbb5),
	.w3(32'hbc755e5d),
	.w4(32'h3b1c37c2),
	.w5(32'h3b891ec9),
	.w6(32'hba8ac206),
	.w7(32'hbc8f53b0),
	.w8(32'hbc68275a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb5e2bd),
	.w1(32'hba605bc1),
	.w2(32'h3c57e4de),
	.w3(32'h3b0c182c),
	.w4(32'h3ba5cde8),
	.w5(32'h39379d09),
	.w6(32'hbb4c15a3),
	.w7(32'h3bbbfea8),
	.w8(32'hbc94ad6a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabe0d9),
	.w1(32'h3ac90b88),
	.w2(32'hbc24d9a4),
	.w3(32'hbb32f781),
	.w4(32'hbb3ac4bf),
	.w5(32'h3ab72992),
	.w6(32'h39aa216a),
	.w7(32'h39b54dde),
	.w8(32'h3bdbbc05),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d2165),
	.w1(32'h38eb4da0),
	.w2(32'h3c005e5a),
	.w3(32'h3ba507df),
	.w4(32'h3bb5cf68),
	.w5(32'hba941b50),
	.w6(32'hbb470c47),
	.w7(32'h3c3248e7),
	.w8(32'h3ae55465),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3e468b),
	.w1(32'hbbdc0b23),
	.w2(32'hb9b92e23),
	.w3(32'h3bc3913c),
	.w4(32'hbc125bbf),
	.w5(32'hbc0b94c6),
	.w6(32'h3ba40cac),
	.w7(32'h3bae74c5),
	.w8(32'h3a423992),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3f27e),
	.w1(32'h3ba40d09),
	.w2(32'h3b42d13e),
	.w3(32'hba6f73ab),
	.w4(32'h3c28e92c),
	.w5(32'hbab6bfc2),
	.w6(32'hbbf95289),
	.w7(32'hbaa366a6),
	.w8(32'hbc123941),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d76ad),
	.w1(32'hbbeae9eb),
	.w2(32'h3b6bf410),
	.w3(32'h3b6a2a98),
	.w4(32'hbaa21de8),
	.w5(32'hbc176ad3),
	.w6(32'hbad80859),
	.w7(32'hb9fcf821),
	.w8(32'h3c58b6c3),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0ab75),
	.w1(32'hbc32fe2c),
	.w2(32'hbc608042),
	.w3(32'h3ad8ed5e),
	.w4(32'h3bcd4189),
	.w5(32'hbc5440a1),
	.w6(32'hbb0a0e30),
	.w7(32'hbc39ae15),
	.w8(32'hb932f9ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750bd2),
	.w1(32'h3b88039c),
	.w2(32'hbc37aac4),
	.w3(32'h3c2fde8a),
	.w4(32'h3a77a645),
	.w5(32'hbc84c32d),
	.w6(32'hbc3ebe05),
	.w7(32'h3b57473b),
	.w8(32'hbbf540d6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be48bb9),
	.w1(32'hbb368807),
	.w2(32'h3ae593f9),
	.w3(32'h3b420e95),
	.w4(32'hbbdbf5dd),
	.w5(32'h3aedd695),
	.w6(32'hb8019b91),
	.w7(32'h3ba9f5a1),
	.w8(32'h3cb88160),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d7d8b),
	.w1(32'h3bc210a0),
	.w2(32'hbc1e41ed),
	.w3(32'hbbc72d76),
	.w4(32'h3adb8d68),
	.w5(32'hbc45ba84),
	.w6(32'h3c42736d),
	.w7(32'h3cbc11c8),
	.w8(32'hbc3ca411),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9924e5),
	.w1(32'hbc2d3d87),
	.w2(32'h3980eb13),
	.w3(32'h3bb23bfc),
	.w4(32'h3a4ce3d8),
	.w5(32'hbc01fb89),
	.w6(32'h3c421a65),
	.w7(32'hbaa72b12),
	.w8(32'hbb4292ae),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fb1ed),
	.w1(32'hbc523b4c),
	.w2(32'h3bdcfa75),
	.w3(32'h3a116457),
	.w4(32'h3c78e483),
	.w5(32'h3cd786e2),
	.w6(32'hba7a4cc5),
	.w7(32'hbbbac976),
	.w8(32'h3b635327),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23753f),
	.w1(32'hbc2889da),
	.w2(32'hbc474eec),
	.w3(32'h3b97915e),
	.w4(32'hbbeb0847),
	.w5(32'hbc99bdd8),
	.w6(32'hbbedab1f),
	.w7(32'hbb33db25),
	.w8(32'hbc81a33b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc780d03),
	.w1(32'hbba4cb86),
	.w2(32'hbba440ca),
	.w3(32'hbc000f6b),
	.w4(32'h3c87eb30),
	.w5(32'h3b8bc724),
	.w6(32'hbc1fad18),
	.w7(32'hbc761094),
	.w8(32'h38fa1722),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067e0a),
	.w1(32'h3bb8ade5),
	.w2(32'h3a3c9237),
	.w3(32'hbbc659ec),
	.w4(32'hbc9256a7),
	.w5(32'hbbed7965),
	.w6(32'hbc1b27c4),
	.w7(32'hbcadeb54),
	.w8(32'hbc926fcc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c4f25),
	.w1(32'hbb86b557),
	.w2(32'hbb0bcaca),
	.w3(32'h3d6d04f4),
	.w4(32'hbc860824),
	.w5(32'h3a08677d),
	.w6(32'hbb5f64f6),
	.w7(32'hbc63675f),
	.w8(32'hbbde867a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3d6cf4),
	.w1(32'hbb0b1009),
	.w2(32'h3b2089df),
	.w3(32'h3b079873),
	.w4(32'h3b3e7e85),
	.w5(32'h3c99f39c),
	.w6(32'h3c116d0d),
	.w7(32'h3b015d99),
	.w8(32'hbb358d22),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c319ca2),
	.w1(32'hbb89df4a),
	.w2(32'hbc6ed858),
	.w3(32'h3b197d41),
	.w4(32'hbc81e22d),
	.w5(32'hbbf448ae),
	.w6(32'hbb40ae57),
	.w7(32'h3b0584a4),
	.w8(32'h3b6a97d8),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4985e5),
	.w1(32'hba81d079),
	.w2(32'hbc295489),
	.w3(32'hbb0e91c1),
	.w4(32'hbd3f77a4),
	.w5(32'h3c7098c4),
	.w6(32'hb7621491),
	.w7(32'h3b4c2dcc),
	.w8(32'hbb7a20bd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d040),
	.w1(32'hbaf5b74e),
	.w2(32'hbcaefdf5),
	.w3(32'h3adee11b),
	.w4(32'h3b74b095),
	.w5(32'hbc568628),
	.w6(32'hbb51548b),
	.w7(32'hbc0ea9db),
	.w8(32'hbc41b773),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5325),
	.w1(32'hbc9d69a0),
	.w2(32'h3a1effbf),
	.w3(32'h3d06c231),
	.w4(32'hbc453f1b),
	.w5(32'hbc1c726d),
	.w6(32'hbba73e93),
	.w7(32'hbc48b23b),
	.w8(32'h3b8763e9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc482cba),
	.w1(32'hbc742c8f),
	.w2(32'h3bd4cca8),
	.w3(32'hba710947),
	.w4(32'h3c0a1833),
	.w5(32'hbc80fdcc),
	.w6(32'h3bef9869),
	.w7(32'hbd18ff51),
	.w8(32'h3cbfedd6),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38f4fb),
	.w1(32'hbc6b0cd6),
	.w2(32'hbd413138),
	.w3(32'h390efe94),
	.w4(32'h3b9c76e0),
	.w5(32'hb82c3ba2),
	.w6(32'h3c67eee0),
	.w7(32'hbb8fcff9),
	.w8(32'h3c04bfb4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9db086),
	.w1(32'h3b6806e0),
	.w2(32'hbc0434b1),
	.w3(32'hbc61724d),
	.w4(32'h3aaba622),
	.w5(32'h3a8f4ec0),
	.w6(32'h3bd14853),
	.w7(32'hbb818808),
	.w8(32'h3c1e5382),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9bfa),
	.w1(32'hbc466453),
	.w2(32'hbcd07b48),
	.w3(32'hbb862ed1),
	.w4(32'hb89ceb55),
	.w5(32'hbc9a8012),
	.w6(32'hbc300fd4),
	.w7(32'h3ae0edbb),
	.w8(32'hbc0d9c18),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89bb45),
	.w1(32'hbbff6331),
	.w2(32'hbc328057),
	.w3(32'h3c90812a),
	.w4(32'h3c5d57c2),
	.w5(32'hbcb0b5b3),
	.w6(32'hbbdce108),
	.w7(32'hbc2113c5),
	.w8(32'hba480dbd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63e440),
	.w1(32'hbb643693),
	.w2(32'h3bb4939b),
	.w3(32'hba525a4e),
	.w4(32'h3adc5188),
	.w5(32'hbafc50fd),
	.w6(32'hbb9a891e),
	.w7(32'h3c34069c),
	.w8(32'hbbdc7e56),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc890aee),
	.w1(32'hb9d32b59),
	.w2(32'h3c566e73),
	.w3(32'hbb90a908),
	.w4(32'h3adcce6d),
	.w5(32'hbbb4829f),
	.w6(32'hbd051bad),
	.w7(32'hbc2a3b5d),
	.w8(32'h3b5289bb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84e158),
	.w1(32'hbc18a149),
	.w2(32'h3bdddd44),
	.w3(32'hbcb92501),
	.w4(32'hbcc7000c),
	.w5(32'hbbb45291),
	.w6(32'hbbb4626f),
	.w7(32'hbd416e62),
	.w8(32'hba9c5994),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4200f),
	.w1(32'h3a168a85),
	.w2(32'hbba2a338),
	.w3(32'hbcc122cc),
	.w4(32'h3cc28432),
	.w5(32'hba1c14b8),
	.w6(32'hbc01316d),
	.w7(32'hbbaf14eb),
	.w8(32'h3ad3a5a4),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988f8fa),
	.w1(32'hbc4e8ee6),
	.w2(32'h3c50ea5f),
	.w3(32'hbbeb116d),
	.w4(32'h3bdd5603),
	.w5(32'hb95e7515),
	.w6(32'hbc4983b1),
	.w7(32'hbaf58630),
	.w8(32'hbc0b95d3),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb491ef7),
	.w1(32'h3c3a4bd0),
	.w2(32'hbceacb23),
	.w3(32'hbc8320fc),
	.w4(32'hbbfe8077),
	.w5(32'hbcd4a615),
	.w6(32'hbc0d8fcf),
	.w7(32'hbbf7969a),
	.w8(32'hbc86d7db),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0c0f61),
	.w1(32'hb7a6454a),
	.w2(32'hbc9bf4b8),
	.w3(32'hbb82dab6),
	.w4(32'h3c811377),
	.w5(32'hbc4fce5d),
	.w6(32'hba8836d9),
	.w7(32'hbb7cdbde),
	.w8(32'hbc36687e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21e6b0),
	.w1(32'hbb9a7885),
	.w2(32'h3a237032),
	.w3(32'hbb9662c5),
	.w4(32'h36af8ca0),
	.w5(32'h3bd30172),
	.w6(32'hbbe99751),
	.w7(32'h3b053298),
	.w8(32'hbb999514),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71bff2),
	.w1(32'hbb88c1c6),
	.w2(32'h3b084e87),
	.w3(32'h3b11a18f),
	.w4(32'hbc12f712),
	.w5(32'hbbb1c6c7),
	.w6(32'hbc7b5082),
	.w7(32'hbccc7159),
	.w8(32'hbb55af00),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb586f2),
	.w1(32'hbc7a798e),
	.w2(32'h3c1f15f6),
	.w3(32'h3cc177c7),
	.w4(32'hb95720b5),
	.w5(32'hba75ef7f),
	.w6(32'hbbd71c51),
	.w7(32'hbd804ce0),
	.w8(32'h3b56045c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40c741),
	.w1(32'hbc4e148c),
	.w2(32'hbae3f246),
	.w3(32'hbca040b7),
	.w4(32'hbaeeaf9d),
	.w5(32'h3bcdba29),
	.w6(32'hbbd99ece),
	.w7(32'h3bfabdcc),
	.w8(32'hbcc2e052),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08baec),
	.w1(32'hbcbd95cf),
	.w2(32'hbc8e88b6),
	.w3(32'h3d71e57a),
	.w4(32'h3bbd968e),
	.w5(32'hbcb5cf80),
	.w6(32'h3c522d98),
	.w7(32'h3b7ea6a4),
	.w8(32'hbc8a75b1),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc809616),
	.w1(32'hbc9bfd23),
	.w2(32'hba6ba0e2),
	.w3(32'hb99e6d51),
	.w4(32'h3bc05e5f),
	.w5(32'h3b53143c),
	.w6(32'h3bf44ae5),
	.w7(32'hbb8476c7),
	.w8(32'hbaada939),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9caf801),
	.w1(32'hb8274901),
	.w2(32'hbc16d05d),
	.w3(32'hbc97dc8b),
	.w4(32'hbb641720),
	.w5(32'hbd1e177b),
	.w6(32'hbd347afb),
	.w7(32'h3ba83d71),
	.w8(32'hbb373685),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cd1be),
	.w1(32'hbcbe1119),
	.w2(32'hbcdc43d4),
	.w3(32'hbb6574c5),
	.w4(32'hbb78e064),
	.w5(32'hbc768d03),
	.w6(32'hbb2d11b8),
	.w7(32'hba17dc7a),
	.w8(32'hbc00264d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9306ec),
	.w1(32'hbbb9324a),
	.w2(32'h3b7c392a),
	.w3(32'h3a93cb4a),
	.w4(32'hbc1d17a2),
	.w5(32'h3b38936d),
	.w6(32'hbb00ecd4),
	.w7(32'h3b9e04e2),
	.w8(32'h3c4ba7f5),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb3172e),
	.w1(32'h3b9d4eea),
	.w2(32'hbc6ac46f),
	.w3(32'h3bcd51fe),
	.w4(32'h3b23b0cb),
	.w5(32'hbb65ae52),
	.w6(32'h3a5b7e15),
	.w7(32'h3c235b99),
	.w8(32'h3ac0d06e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7893f4),
	.w1(32'hbb0f06db),
	.w2(32'hbaa81d05),
	.w3(32'h3b8f8144),
	.w4(32'hbc0297eb),
	.w5(32'h38c0ffa0),
	.w6(32'hbbb7ec65),
	.w7(32'h3c06d55f),
	.w8(32'hbba8d472),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c8b83),
	.w1(32'hbb8316a3),
	.w2(32'h3a8693d4),
	.w3(32'hbb96ffb8),
	.w4(32'h3afbdd60),
	.w5(32'hbbcd18bc),
	.w6(32'hbb420ce2),
	.w7(32'h3adf2e10),
	.w8(32'hbc408df6),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e277c),
	.w1(32'hbbdd5a3b),
	.w2(32'hbc118e3d),
	.w3(32'hbb0ba96d),
	.w4(32'h3bbb2137),
	.w5(32'hbb6ed928),
	.w6(32'h3b38d704),
	.w7(32'h3be02a54),
	.w8(32'hbbfcd5b2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5059c),
	.w1(32'h3c182b93),
	.w2(32'h3b9e7fe8),
	.w3(32'hbd3379c9),
	.w4(32'hbbe7096e),
	.w5(32'hb9bc50ef),
	.w6(32'h3c1056ad),
	.w7(32'hbc3cae34),
	.w8(32'hbbc4e1a7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3565f1),
	.w1(32'hbb3c13e5),
	.w2(32'hbb8c2db1),
	.w3(32'h3be749b6),
	.w4(32'hba86381c),
	.w5(32'hbad6630a),
	.w6(32'hbbbb1492),
	.w7(32'h39ebbd23),
	.w8(32'hbb7981de),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9929c),
	.w1(32'hb98e1b63),
	.w2(32'hbbbc763a),
	.w3(32'hbbfe1768),
	.w4(32'hbae713d9),
	.w5(32'h3a5bffd4),
	.w6(32'h3b652e15),
	.w7(32'hbb15b73d),
	.w8(32'h3c850ba0),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebb3cc),
	.w1(32'h3ba4d9de),
	.w2(32'hba775010),
	.w3(32'h3adcf008),
	.w4(32'hbc07162d),
	.w5(32'h3c08aef3),
	.w6(32'hbc7030b6),
	.w7(32'h3b81fb1c),
	.w8(32'h3b8638be),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62893d),
	.w1(32'h3b65deb3),
	.w2(32'hbc13aa25),
	.w3(32'h3ad4fd62),
	.w4(32'hbb37bace),
	.w5(32'h3ba30fb0),
	.w6(32'hbc97c6dc),
	.w7(32'hbb0b4541),
	.w8(32'h3c152953),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe46701),
	.w1(32'h3b04bf47),
	.w2(32'hba7b8869),
	.w3(32'h3c2d1e17),
	.w4(32'hbb60f376),
	.w5(32'hba411e24),
	.w6(32'h3c0503cc),
	.w7(32'h3a8b5538),
	.w8(32'h3ba7ca7f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e91b7),
	.w1(32'hbc1c5f6d),
	.w2(32'hbb91249f),
	.w3(32'hba3f6097),
	.w4(32'hbba59d54),
	.w5(32'hba743f97),
	.w6(32'h3b1a012d),
	.w7(32'hbbef3525),
	.w8(32'h3bf40f56),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8981b0),
	.w1(32'hbb14c84b),
	.w2(32'hbc8b78e9),
	.w3(32'hbbc1f4e6),
	.w4(32'h3bbc703f),
	.w5(32'h3c1d23d6),
	.w6(32'hb9a012ba),
	.w7(32'h3b65bcce),
	.w8(32'h3b8a46a1),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f811b),
	.w1(32'hb841aa3e),
	.w2(32'hbb8b2148),
	.w3(32'hba857f2f),
	.w4(32'h3c0d9e92),
	.w5(32'hbbfcf6fd),
	.w6(32'h3b8fac4e),
	.w7(32'hba45755c),
	.w8(32'hbb8cc2fe),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fcd71),
	.w1(32'hbbacf1a7),
	.w2(32'hbba29055),
	.w3(32'h3b722e43),
	.w4(32'h3bc94ba2),
	.w5(32'h3b96067b),
	.w6(32'h3b2a13a1),
	.w7(32'hbc40c3f5),
	.w8(32'hbbb2fd31),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0747d9),
	.w1(32'hbad8fef6),
	.w2(32'h3bb57eb7),
	.w3(32'h3a3bc5ae),
	.w4(32'h3bf000b8),
	.w5(32'hbc961618),
	.w6(32'h3b0cfe35),
	.w7(32'hbb851f0a),
	.w8(32'h39e2faed),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb254881),
	.w1(32'hb9711607),
	.w2(32'h3b3c37ae),
	.w3(32'hb88acc51),
	.w4(32'h3b509032),
	.w5(32'h3b815a10),
	.w6(32'hbae9cddd),
	.w7(32'hbbf0a90a),
	.w8(32'hbb8cb8d6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8c117),
	.w1(32'hbc2a0d3d),
	.w2(32'hbb830c3b),
	.w3(32'hbb701be6),
	.w4(32'h3bb9e87e),
	.w5(32'h3bd33e3a),
	.w6(32'hba5fcd86),
	.w7(32'h3a0e8956),
	.w8(32'h394782a5),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a2a95),
	.w1(32'h3b86af35),
	.w2(32'hbb23d549),
	.w3(32'h3c0c6fed),
	.w4(32'hbc6b4a72),
	.w5(32'h3c2c1d00),
	.w6(32'h39da9c21),
	.w7(32'hb9a7a4fc),
	.w8(32'h3ac56379),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6ec1a),
	.w1(32'h3c673ef3),
	.w2(32'h3b86f9e4),
	.w3(32'h3bd3bf4d),
	.w4(32'h3b076917),
	.w5(32'h3b05f121),
	.w6(32'h3c1d6320),
	.w7(32'h3bb61fbb),
	.w8(32'hb9c1d037),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8beb9b),
	.w1(32'hbb25ce68),
	.w2(32'hbb4477b0),
	.w3(32'hbbf074ee),
	.w4(32'hbbc33f99),
	.w5(32'hbb0bf049),
	.w6(32'hbb455c19),
	.w7(32'hbcdaeaba),
	.w8(32'h3b385f89),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5fd504),
	.w1(32'hb99a0e84),
	.w2(32'h3796f862),
	.w3(32'hbb785905),
	.w4(32'h3a999a80),
	.w5(32'h3c148a73),
	.w6(32'h3b4126bd),
	.w7(32'hbb38477b),
	.w8(32'hbbabe3c7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c038fbc),
	.w1(32'hbba2eeaf),
	.w2(32'hbac8ca25),
	.w3(32'hbb0c144c),
	.w4(32'hbb98867f),
	.w5(32'h3b8a2b73),
	.w6(32'hbb95abeb),
	.w7(32'h3bc7a059),
	.w8(32'h3b9b39f1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedc2f1),
	.w1(32'h39f1e1c6),
	.w2(32'hbb24e406),
	.w3(32'h3c266341),
	.w4(32'h3bb4ad45),
	.w5(32'h3b4ff53c),
	.w6(32'h3a73dae0),
	.w7(32'hbb964d9c),
	.w8(32'h39822d8d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fe4b4),
	.w1(32'hbbd9ebb6),
	.w2(32'hbc02bd97),
	.w3(32'h38d15006),
	.w4(32'h3c73f2ea),
	.w5(32'hbba03fc7),
	.w6(32'h3a05e4a8),
	.w7(32'hbbf9cda9),
	.w8(32'hbbb20dfb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b524257),
	.w1(32'hbc594ab0),
	.w2(32'h39a4c0f1),
	.w3(32'h3c4bb5b6),
	.w4(32'hbc68d5de),
	.w5(32'hbb8fdeb9),
	.w6(32'hbac466ce),
	.w7(32'h3b73c26b),
	.w8(32'hbb3aa45b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fb0e0),
	.w1(32'h3c0d3f20),
	.w2(32'h3c1ef703),
	.w3(32'hbc24ea3a),
	.w4(32'hbb931c5b),
	.w5(32'hbbda36b7),
	.w6(32'h3bc31a90),
	.w7(32'hbbfa04fc),
	.w8(32'hbb61a31d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba999af7),
	.w1(32'hbb915a36),
	.w2(32'h3b91f7a7),
	.w3(32'hbb917ca6),
	.w4(32'hbb94daa2),
	.w5(32'h3b28e39b),
	.w6(32'hbbdeb2a4),
	.w7(32'hbc02fb47),
	.w8(32'h3acee8a4),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad09e80),
	.w1(32'hbbddadac),
	.w2(32'h3afde4b2),
	.w3(32'h3b97ed5a),
	.w4(32'hbb6a9e8f),
	.w5(32'h3bc698bc),
	.w6(32'hbbad6a00),
	.w7(32'hbbb5ecfc),
	.w8(32'hbba5f7ba),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a998729),
	.w1(32'hbbb4fcc9),
	.w2(32'h3bfb2034),
	.w3(32'hbb86173c),
	.w4(32'h3c65695d),
	.w5(32'h3be1ce19),
	.w6(32'h3af964dd),
	.w7(32'hbc09c148),
	.w8(32'hbba42347),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffb2a5),
	.w1(32'hbbfd65fa),
	.w2(32'hbba6b83f),
	.w3(32'hbc505ae6),
	.w4(32'hbc429ac2),
	.w5(32'h3bc25122),
	.w6(32'hbb99509d),
	.w7(32'hbbbbd756),
	.w8(32'h3c2e4a1f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9536c),
	.w1(32'hba97ec99),
	.w2(32'hbaf375f6),
	.w3(32'h3b521095),
	.w4(32'hbaee09e1),
	.w5(32'hbb82448b),
	.w6(32'hbda5ed16),
	.w7(32'h3c1d2923),
	.w8(32'h3ba92e28),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7811e9),
	.w1(32'hbc303a34),
	.w2(32'hbc53687f),
	.w3(32'h3be58ffc),
	.w4(32'h3cb74405),
	.w5(32'h3c00126c),
	.w6(32'hb977103a),
	.w7(32'hbb0be57a),
	.w8(32'h3b85f43d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1372c4),
	.w1(32'hbccece65),
	.w2(32'h3c378d18),
	.w3(32'hbc0056e1),
	.w4(32'h3bc1258e),
	.w5(32'hba540ea9),
	.w6(32'hbb8c0956),
	.w7(32'h3bd6b17d),
	.w8(32'h3bc3a185),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4193b2),
	.w1(32'h3a71b013),
	.w2(32'h3c0fab36),
	.w3(32'hbb2fb4ae),
	.w4(32'h3abb1529),
	.w5(32'h3b626283),
	.w6(32'h3b753068),
	.w7(32'h3b3b4939),
	.w8(32'h3b0ecc34),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9721aa),
	.w1(32'h39c33ec5),
	.w2(32'hba9041b9),
	.w3(32'hbc7d220b),
	.w4(32'hbb13405f),
	.w5(32'h3b772e5c),
	.w6(32'h3c06e2d3),
	.w7(32'hbc7be258),
	.w8(32'h3b012c58),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8c171),
	.w1(32'hbb434665),
	.w2(32'h3c1fa018),
	.w3(32'h3b6eea83),
	.w4(32'hbb6ca1e1),
	.w5(32'hbc013bc0),
	.w6(32'hbba9c691),
	.w7(32'hbb619332),
	.w8(32'h3bd5edfd),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cdc62),
	.w1(32'hba5a2d68),
	.w2(32'hbb7065c6),
	.w3(32'hbc3ee1de),
	.w4(32'hbbceabe9),
	.w5(32'h3aec1cd6),
	.w6(32'hbb3486e3),
	.w7(32'hbb8be799),
	.w8(32'h3b29ee37),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e02c2d),
	.w1(32'h3b568ca2),
	.w2(32'hbb63a222),
	.w3(32'hbaf2346b),
	.w4(32'hba16a4a1),
	.w5(32'h3ab99afa),
	.w6(32'hbd72546a),
	.w7(32'hbcba4722),
	.w8(32'h39e31d42),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00a899),
	.w1(32'hbb742188),
	.w2(32'h3b866db0),
	.w3(32'hba2f536c),
	.w4(32'h3c388caf),
	.w5(32'h3c0fe390),
	.w6(32'hbbff3bf5),
	.w7(32'hbb0cc270),
	.w8(32'hbba848fb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac53e2),
	.w1(32'hbb7a9153),
	.w2(32'hbc04aa69),
	.w3(32'h3a8db662),
	.w4(32'h3bcb252d),
	.w5(32'hbbc9726b),
	.w6(32'h3ac4ddd0),
	.w7(32'h3a80272e),
	.w8(32'hba093263),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1414a),
	.w1(32'hbb0401ad),
	.w2(32'hbc48990c),
	.w3(32'hbb63e8e1),
	.w4(32'h3a6c815b),
	.w5(32'hb805858d),
	.w6(32'h3c00c5d2),
	.w7(32'h3ab6f08b),
	.w8(32'hbcefd1fb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26d666),
	.w1(32'h3b923e81),
	.w2(32'h3a870b9b),
	.w3(32'h3c2f2569),
	.w4(32'hbb1ff8b9),
	.w5(32'h3a0f3840),
	.w6(32'hbbc31130),
	.w7(32'h3bf1729f),
	.w8(32'hb920d0a1),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa5579),
	.w1(32'hbc41622a),
	.w2(32'hbb6e6299),
	.w3(32'hbbeaad8a),
	.w4(32'hbcc0eabb),
	.w5(32'h3b9db038),
	.w6(32'h3cf3863e),
	.w7(32'hbcccaa51),
	.w8(32'h3b0c8c52),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a0e2d),
	.w1(32'h3b7e0a70),
	.w2(32'hbb2d50c1),
	.w3(32'h3992ff52),
	.w4(32'hb9bee6b9),
	.w5(32'hbb4ecebf),
	.w6(32'hbd1a47d8),
	.w7(32'hbb41bf49),
	.w8(32'h3b3d851b),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f7c13),
	.w1(32'hbb991ab0),
	.w2(32'hba913706),
	.w3(32'hba9c1cc6),
	.w4(32'h3b7d5b76),
	.w5(32'h3b26b187),
	.w6(32'h3bf24621),
	.w7(32'h3af7464e),
	.w8(32'h3b794f2e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8563c),
	.w1(32'hbb3b02bf),
	.w2(32'hb90a3aac),
	.w3(32'h3baf1d26),
	.w4(32'h3b33c871),
	.w5(32'h39db2a63),
	.w6(32'h3af5b8b5),
	.w7(32'hbbf09797),
	.w8(32'hbc126168),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d3a68),
	.w1(32'hbb9de531),
	.w2(32'h3bef8bb7),
	.w3(32'hbb887f24),
	.w4(32'h3b3b3ba7),
	.w5(32'hbc180a71),
	.w6(32'hbae164f0),
	.w7(32'hbd150bbc),
	.w8(32'h3c3bd039),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a920c),
	.w1(32'hbbf98379),
	.w2(32'hbb739676),
	.w3(32'hbadfca3f),
	.w4(32'h3b9da876),
	.w5(32'h3bbb7718),
	.w6(32'h3b873cb9),
	.w7(32'h3aa6cd49),
	.w8(32'h3b2f1531),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5d2be),
	.w1(32'hbbc01d7b),
	.w2(32'h3c919fa7),
	.w3(32'h3b6b3407),
	.w4(32'h3ae0d611),
	.w5(32'h3ab933a1),
	.w6(32'h3d01ab7d),
	.w7(32'h3b710d2c),
	.w8(32'h3a15123d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96f8cb),
	.w1(32'h3b3fd614),
	.w2(32'hbb3b2cf2),
	.w3(32'hbb79bb74),
	.w4(32'h3925e7b2),
	.w5(32'hbbf8aa2c),
	.w6(32'h3af01cb8),
	.w7(32'h3b09adc7),
	.w8(32'h3c1ebdfa),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9df4f5),
	.w1(32'hbaed8e60),
	.w2(32'hb94f0b56),
	.w3(32'hba159bc6),
	.w4(32'hbc4d0e2a),
	.w5(32'h3ad97536),
	.w6(32'h3c1eee5a),
	.w7(32'h3c2ac38f),
	.w8(32'h3a9ff403),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda8dfd),
	.w1(32'h3b72b93b),
	.w2(32'h3b3b1beb),
	.w3(32'h3c26bcfb),
	.w4(32'h3b250260),
	.w5(32'h3b0fa8af),
	.w6(32'hbb5a3111),
	.w7(32'hb8ac6e1e),
	.w8(32'h3cf5e068),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a890bab),
	.w1(32'hbb35f33e),
	.w2(32'hbb432a30),
	.w3(32'hbccf530b),
	.w4(32'hbb03a94f),
	.w5(32'h3bc3f9eb),
	.w6(32'h3c0911c1),
	.w7(32'hbb87d67b),
	.w8(32'h3bc8bff5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb3a54),
	.w1(32'h3a3bd996),
	.w2(32'hbd038927),
	.w3(32'h38f3c53a),
	.w4(32'h3adf0d4f),
	.w5(32'hbc0cbbe6),
	.w6(32'h3a936eff),
	.w7(32'hbb02d44e),
	.w8(32'hbb18677d),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d43fe),
	.w1(32'hbbded980),
	.w2(32'hbbd5215d),
	.w3(32'h39921a8a),
	.w4(32'h3bd0cfc1),
	.w5(32'hbb431fb6),
	.w6(32'h3c762b3b),
	.w7(32'hbc4a2672),
	.w8(32'h3a3fb636),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4c20),
	.w1(32'h3b074bbb),
	.w2(32'h3b292d94),
	.w3(32'h3b19ec26),
	.w4(32'h3c0b04a8),
	.w5(32'hbb3ba703),
	.w6(32'hbb4ef02c),
	.w7(32'hbd7c9d33),
	.w8(32'hbc304797),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a750c35),
	.w1(32'h3b5072cf),
	.w2(32'hbbb46dbb),
	.w3(32'h3c8a5d63),
	.w4(32'h3b55c191),
	.w5(32'h3c5e09fb),
	.w6(32'hbc830301),
	.w7(32'h3be946e3),
	.w8(32'h3ba03f8b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ec5f7),
	.w1(32'h3b59ad52),
	.w2(32'hbae54b1e),
	.w3(32'h3a8927a1),
	.w4(32'hbc2a0b37),
	.w5(32'h3a835f3c),
	.w6(32'h3bc0730b),
	.w7(32'hbabdad78),
	.w8(32'h3c00a982),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc323832),
	.w1(32'h3cc2108e),
	.w2(32'h3a84ae2d),
	.w3(32'h3b954f2d),
	.w4(32'hbb8a4791),
	.w5(32'hbb07152e),
	.w6(32'h3bf5407d),
	.w7(32'h3918c52d),
	.w8(32'hbbc50d8a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ae512),
	.w1(32'hbc236511),
	.w2(32'hbc93681e),
	.w3(32'hbca1b668),
	.w4(32'hba16b351),
	.w5(32'h3c456dbe),
	.w6(32'h3c877af1),
	.w7(32'h3b22d248),
	.w8(32'h3b259788),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18b2bb),
	.w1(32'hbc0eac7a),
	.w2(32'hbbe0e9e8),
	.w3(32'h3b04602a),
	.w4(32'hbc22820f),
	.w5(32'hbcba7780),
	.w6(32'h3b6c1f9a),
	.w7(32'hbaaceece),
	.w8(32'h3a260a38),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c540400),
	.w1(32'hbc5ca712),
	.w2(32'h3bc0fee2),
	.w3(32'h3c56a32c),
	.w4(32'h3b7edff1),
	.w5(32'hbc5866d7),
	.w6(32'hbb9b1895),
	.w7(32'hba98a2d9),
	.w8(32'h3ad2ced0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44589f),
	.w1(32'hbc71d9ef),
	.w2(32'hbc6aacc5),
	.w3(32'hbcd6d194),
	.w4(32'hb94849eb),
	.w5(32'h3b25d345),
	.w6(32'h3c634ce3),
	.w7(32'hbc7de91d),
	.w8(32'h3c4fa8c6),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd76698),
	.w1(32'hbb9dd4c4),
	.w2(32'hbc46ccdd),
	.w3(32'h3a09e21c),
	.w4(32'h3c8cf004),
	.w5(32'h3cd4da75),
	.w6(32'h3a95c820),
	.w7(32'hbbf86314),
	.w8(32'h3bcb76ab),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1836c),
	.w1(32'h3c0147df),
	.w2(32'hbc84985f),
	.w3(32'hbc6be1a9),
	.w4(32'hb9fb81ae),
	.w5(32'hbd30434f),
	.w6(32'hbc1ec986),
	.w7(32'h3ae55268),
	.w8(32'h3aca74b5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007353),
	.w1(32'h3bdada30),
	.w2(32'hba821ad3),
	.w3(32'h3c19d5db),
	.w4(32'hbc187416),
	.w5(32'hbbd40e97),
	.w6(32'h3ab789b2),
	.w7(32'h3c05af2c),
	.w8(32'hbcce22f9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5224ab),
	.w1(32'hbb983ac1),
	.w2(32'h3a3bf90d),
	.w3(32'hbc585cf6),
	.w4(32'h3c239328),
	.w5(32'h3cfdf72e),
	.w6(32'hbb09f1fc),
	.w7(32'hbb4330d0),
	.w8(32'h3c42322c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba830b4a),
	.w1(32'hbb394978),
	.w2(32'hbc6639f4),
	.w3(32'h3c909a8a),
	.w4(32'hbcb502d2),
	.w5(32'h3aaee3db),
	.w6(32'h3babad42),
	.w7(32'hb94f2621),
	.w8(32'hbc3cf9bc),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c217ef1),
	.w1(32'h3c484b7e),
	.w2(32'hbaa26a47),
	.w3(32'hbbd98549),
	.w4(32'h3a6fa24c),
	.w5(32'h3940c1ad),
	.w6(32'hba9a48d7),
	.w7(32'hbb3c6b87),
	.w8(32'hbc108af5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2ef1),
	.w1(32'hbcc13f1e),
	.w2(32'h3c14c719),
	.w3(32'h3c455cee),
	.w4(32'hb8afdc95),
	.w5(32'hbc9d00d1),
	.w6(32'hb96f4710),
	.w7(32'hbd1932de),
	.w8(32'h3b1fad26),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a47a9e8),
	.w1(32'hbbcf8549),
	.w2(32'hb9f92f5b),
	.w3(32'h3be33c05),
	.w4(32'hbccb8d61),
	.w5(32'hbcf5a18f),
	.w6(32'hbaaacd33),
	.w7(32'hbc250909),
	.w8(32'hbd0d6c69),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2511ef),
	.w1(32'h394f9e32),
	.w2(32'hbc141735),
	.w3(32'h3c46292b),
	.w4(32'h3b88d444),
	.w5(32'h3b2a3300),
	.w6(32'h3c781510),
	.w7(32'h3af31663),
	.w8(32'hbd08dcc7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e9fb4),
	.w1(32'h3c3d475e),
	.w2(32'h3cc8df33),
	.w3(32'h3d358e2e),
	.w4(32'hbbe53552),
	.w5(32'h3c2f051c),
	.w6(32'h3b542fac),
	.w7(32'h3a225f12),
	.w8(32'h3baf9a04),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08825),
	.w1(32'hbc5e7269),
	.w2(32'h3c24e0ee),
	.w3(32'hba687b47),
	.w4(32'h3c22e0fa),
	.w5(32'h3bc71454),
	.w6(32'hbb8d9bf2),
	.w7(32'h3b96ad92),
	.w8(32'h3b9884fd),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba5359),
	.w1(32'hbcb4a550),
	.w2(32'h3b293796),
	.w3(32'hb959b26f),
	.w4(32'hbaf6c04a),
	.w5(32'h3b2b94b2),
	.w6(32'hbbc92251),
	.w7(32'h3a4bd85e),
	.w8(32'hbcbfdd75),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb210e31),
	.w1(32'hbc12ad28),
	.w2(32'hba848f5d),
	.w3(32'hbc81b339),
	.w4(32'h3bacf467),
	.w5(32'hbc0cd29d),
	.w6(32'h3c60601d),
	.w7(32'h3b0e4689),
	.w8(32'hbc5d1c68),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf3c08),
	.w1(32'hbc91a136),
	.w2(32'hbae59900),
	.w3(32'hbacb9769),
	.w4(32'hbb210663),
	.w5(32'hbc9903a1),
	.w6(32'h3aff58f0),
	.w7(32'h3b816a90),
	.w8(32'h3ad859ad),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcad08c),
	.w1(32'hbc07ea9a),
	.w2(32'h3c0fd948),
	.w3(32'h3c0ddf92),
	.w4(32'hbb67cc4a),
	.w5(32'hba5981ee),
	.w6(32'h3ba1c15d),
	.w7(32'h3b5a87c3),
	.w8(32'hbaeae234),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca87ff),
	.w1(32'h3b8e8ac3),
	.w2(32'hbc871ed8),
	.w3(32'hbae314ca),
	.w4(32'hbae5a7cd),
	.w5(32'h3aef3e91),
	.w6(32'hbc485d9a),
	.w7(32'hbb8341a7),
	.w8(32'hbbde18c2),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eabc6),
	.w1(32'h3bad5181),
	.w2(32'h3ca5adef),
	.w3(32'hbae06c3a),
	.w4(32'hbc83f37f),
	.w5(32'hbc5aa05e),
	.w6(32'hba33ce47),
	.w7(32'hbbdc7be5),
	.w8(32'h39c6b737),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03cf7b),
	.w1(32'hbbd63564),
	.w2(32'hbb568279),
	.w3(32'hbb78fffc),
	.w4(32'h3cd06c8a),
	.w5(32'hbab1d2ba),
	.w6(32'hbbccb018),
	.w7(32'hbb61b7fb),
	.w8(32'hbbfb1027),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd18258e),
	.w1(32'hbbe1c213),
	.w2(32'h3c6fc60b),
	.w3(32'hbb4884f4),
	.w4(32'h3c1dfa38),
	.w5(32'hba46870b),
	.w6(32'hbc8bcb05),
	.w7(32'h3c40659f),
	.w8(32'h3c44002e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc496067),
	.w1(32'hbb0b6aed),
	.w2(32'h39d9c2d8),
	.w3(32'hba2ff778),
	.w4(32'h3baa19fd),
	.w5(32'h39afdfad),
	.w6(32'h3c12b771),
	.w7(32'h3ca4436a),
	.w8(32'h3aabdda6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d6fd3),
	.w1(32'hbc5e165b),
	.w2(32'h3a52d173),
	.w3(32'hbc0aa8cd),
	.w4(32'hbc596a61),
	.w5(32'hbab67bc3),
	.w6(32'hbc346ba6),
	.w7(32'hbb88a8d0),
	.w8(32'h3a7a13f0),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94763b),
	.w1(32'hbbe0d0d0),
	.w2(32'h3ba1fdf6),
	.w3(32'hbc77f2d9),
	.w4(32'hbb2c3ae4),
	.w5(32'h3a125c1e),
	.w6(32'hbbecdc4b),
	.w7(32'hba34e3ed),
	.w8(32'h3b706f1e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3704b2),
	.w1(32'h3bf44539),
	.w2(32'hbb4ce07f),
	.w3(32'hbba67ba9),
	.w4(32'h3d0b213b),
	.w5(32'h3bd64b79),
	.w6(32'hbc344163),
	.w7(32'hbc0ff30c),
	.w8(32'h3bed5842),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24cd5c),
	.w1(32'hbcf756fb),
	.w2(32'hbbc3c5d0),
	.w3(32'hbba69a8a),
	.w4(32'h3b310d78),
	.w5(32'hbb7495e4),
	.w6(32'hba982fc2),
	.w7(32'hbb8af3d1),
	.w8(32'h3bb1f2e8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6898),
	.w1(32'h3b0721b5),
	.w2(32'h3a33d1df),
	.w3(32'hbcea3fa6),
	.w4(32'hbc2b4d5a),
	.w5(32'h3c2b8eed),
	.w6(32'h3b1c4452),
	.w7(32'hbbb2b975),
	.w8(32'h3a1897bc),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3d3c5),
	.w1(32'h3cd0c831),
	.w2(32'hbb693dc0),
	.w3(32'hb97d80ab),
	.w4(32'hbbd890af),
	.w5(32'h3cc24c9c),
	.w6(32'hbc043cad),
	.w7(32'hbab65d19),
	.w8(32'h3aa0f6c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996b2a3),
	.w1(32'hbbee8583),
	.w2(32'hbb261540),
	.w3(32'h3c8397dd),
	.w4(32'hbc7a30b4),
	.w5(32'hbafb9c8a),
	.w6(32'h3c53f045),
	.w7(32'hbbc74975),
	.w8(32'hbb101c4f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bfb95),
	.w1(32'hbbc15975),
	.w2(32'hbb5c0a4b),
	.w3(32'h3a4d0d79),
	.w4(32'hbc09d171),
	.w5(32'hba06b1ab),
	.w6(32'hbbcc2f9a),
	.w7(32'h3c11a502),
	.w8(32'hbaced488),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e4eaf),
	.w1(32'hb883606d),
	.w2(32'hbbb1d171),
	.w3(32'hbb104923),
	.w4(32'h3bb3330c),
	.w5(32'hbbb93803),
	.w6(32'hbb87ee9e),
	.w7(32'hbbbc7627),
	.w8(32'h3bb8f6b0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ea959),
	.w1(32'hbb29dee1),
	.w2(32'hbac9040c),
	.w3(32'h3a9c3e60),
	.w4(32'h3c846102),
	.w5(32'hbadb76f4),
	.w6(32'h3c9686d3),
	.w7(32'hbd139f48),
	.w8(32'hbc2c22e2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41db73),
	.w1(32'hbc64f7db),
	.w2(32'hbb9aeea1),
	.w3(32'hbc0195c8),
	.w4(32'hbba12558),
	.w5(32'hba7c0a4c),
	.w6(32'hba483efe),
	.w7(32'hbb6d64c3),
	.w8(32'hbb1cf032),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19f6ec),
	.w1(32'h3a9a3ed7),
	.w2(32'h3bb1bdc8),
	.w3(32'h3a368d2d),
	.w4(32'h3b822eca),
	.w5(32'hbb703929),
	.w6(32'hbb80d9df),
	.w7(32'hbbb07deb),
	.w8(32'h3b053b1d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3bafe7),
	.w1(32'hbc385e07),
	.w2(32'h3ac5ff3a),
	.w3(32'hbcb2ab38),
	.w4(32'hb920dc1b),
	.w5(32'hbc81c9e3),
	.w6(32'h3b345142),
	.w7(32'h3ad91e79),
	.w8(32'hbc169519),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba690b96),
	.w1(32'h3c707c43),
	.w2(32'hbb8f14c2),
	.w3(32'hba46ef4a),
	.w4(32'h3bc7e7f4),
	.w5(32'h3bfce39e),
	.w6(32'h3aef79ad),
	.w7(32'hbc6ffe21),
	.w8(32'h3cb4c1c1),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c494ee7),
	.w1(32'hbb389463),
	.w2(32'hba33de0f),
	.w3(32'h3b746c8c),
	.w4(32'hbb136650),
	.w5(32'hbbc93246),
	.w6(32'hbb7135cc),
	.w7(32'hbd2e06e9),
	.w8(32'h3acae252),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f65f),
	.w1(32'hbc2b4835),
	.w2(32'h3a13e631),
	.w3(32'hbc0c544d),
	.w4(32'h3bee5ea4),
	.w5(32'hbbfa61e3),
	.w6(32'hbb17893a),
	.w7(32'h38d7ae0d),
	.w8(32'hbcc20112),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb494038),
	.w1(32'hbc0cbf7d),
	.w2(32'hbc25c945),
	.w3(32'h3c16d438),
	.w4(32'h3b3331b6),
	.w5(32'h39a16e66),
	.w6(32'h3b773e62),
	.w7(32'h3cba68b1),
	.w8(32'h38da55b4),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac667d),
	.w1(32'hbc1b18af),
	.w2(32'h3bca924c),
	.w3(32'hbaaada97),
	.w4(32'hbb9e4eab),
	.w5(32'hbb9e0862),
	.w6(32'hba1d9887),
	.w7(32'h3ac33157),
	.w8(32'hb9ef4c0c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91a719),
	.w1(32'h3b528ae8),
	.w2(32'hbc16cb97),
	.w3(32'h3b822746),
	.w4(32'hba32da63),
	.w5(32'hbc10cf94),
	.w6(32'h3bef7272),
	.w7(32'hbae3e0cb),
	.w8(32'h39a6e84d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3123f8),
	.w1(32'hbc0d4bed),
	.w2(32'h3a124a33),
	.w3(32'h3b17c39c),
	.w4(32'h3a97e755),
	.w5(32'hbc05fd29),
	.w6(32'hbb90aad5),
	.w7(32'hb9189a93),
	.w8(32'h3b4ab8d1),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96b6017),
	.w1(32'hbbc927ec),
	.w2(32'h3d42749f),
	.w3(32'h3b3afdd1),
	.w4(32'h3cd60471),
	.w5(32'hbbef6dc0),
	.w6(32'hbb448d96),
	.w7(32'h3c82d06b),
	.w8(32'h3b8d6471),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb964a6d6),
	.w1(32'hbbd5dc77),
	.w2(32'h3b19edb8),
	.w3(32'hba720885),
	.w4(32'hbc15b57d),
	.w5(32'hb9a01adf),
	.w6(32'hbc22827d),
	.w7(32'hbb0760ab),
	.w8(32'hbce47453),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa92cf9),
	.w1(32'h3adbabca),
	.w2(32'hbc11588c),
	.w3(32'h3c564c75),
	.w4(32'hba0fbd9e),
	.w5(32'hbbf9b7e9),
	.w6(32'h3ba953d4),
	.w7(32'hbcb3069e),
	.w8(32'hbad01081),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd3303),
	.w1(32'h3c55fcec),
	.w2(32'hbb92acd4),
	.w3(32'hb9ca0cf2),
	.w4(32'hbb995f52),
	.w5(32'hbd1bf054),
	.w6(32'h3a0befd0),
	.w7(32'h3b1e0fff),
	.w8(32'h3b85b89b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8dfe42),
	.w1(32'hbc93bab9),
	.w2(32'h3b0a7d0c),
	.w3(32'hbb249df1),
	.w4(32'h3c6978c2),
	.w5(32'hbbfa9238),
	.w6(32'hbb5db555),
	.w7(32'hbaaccaeb),
	.w8(32'hbb8ca8fd),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b2e2fb),
	.w1(32'hbab638a6),
	.w2(32'hbc57f36f),
	.w3(32'h3c04d577),
	.w4(32'h388ae2ba),
	.w5(32'hbd0e5a36),
	.w6(32'hbb3d47bd),
	.w7(32'h3bb99cc4),
	.w8(32'h3b7aea61),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3242c6),
	.w1(32'h3bc7e324),
	.w2(32'h3b338072),
	.w3(32'hbbd04112),
	.w4(32'hbc07b97b),
	.w5(32'h39efc3db),
	.w6(32'h3bb1945a),
	.w7(32'hbae5ab2c),
	.w8(32'h3b8a3926),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd50273),
	.w1(32'h3bf3456e),
	.w2(32'h3b8e0f6b),
	.w3(32'hbb8fe8e2),
	.w4(32'hbaa3f4b6),
	.w5(32'hba2e2ca8),
	.w6(32'hbb31214e),
	.w7(32'h3c3dd3ee),
	.w8(32'hbbb81f1f),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0deed),
	.w1(32'hbc0474d9),
	.w2(32'h3be13cab),
	.w3(32'hba9b0b77),
	.w4(32'h3b824256),
	.w5(32'hba90417f),
	.w6(32'hbb8020ca),
	.w7(32'h3b260eb7),
	.w8(32'h398306cf),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c69c4),
	.w1(32'hbbd07819),
	.w2(32'hbc38b025),
	.w3(32'h3b2f67d9),
	.w4(32'hbc86d235),
	.w5(32'hba57ac1e),
	.w6(32'hbb6b09a4),
	.w7(32'h3ac507e4),
	.w8(32'hbabcd9d7),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67eaf8),
	.w1(32'hbbfe8280),
	.w2(32'h3bf13fcc),
	.w3(32'h3ac8b7bc),
	.w4(32'h3c4288a8),
	.w5(32'h3c23b5f2),
	.w6(32'h3be4a23c),
	.w7(32'hbc0f2f67),
	.w8(32'h3c8d26bf),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ebc0fb),
	.w1(32'h3c51111e),
	.w2(32'h3c40bd10),
	.w3(32'hbc30a4d8),
	.w4(32'h3c85a45c),
	.w5(32'h3a2acde5),
	.w6(32'hbc794541),
	.w7(32'hbc264d2e),
	.w8(32'h3bb81e37),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5abb6),
	.w1(32'hbc480d98),
	.w2(32'h3c0bd545),
	.w3(32'h3c272215),
	.w4(32'hbbc65b93),
	.w5(32'h3c22156d),
	.w6(32'h388c661c),
	.w7(32'h3b41445b),
	.w8(32'h3bb61fe9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1038ec),
	.w1(32'h3beedfc9),
	.w2(32'h3c661bee),
	.w3(32'hbc1f88d7),
	.w4(32'hbba281d7),
	.w5(32'h3cf783e0),
	.w6(32'hbc992971),
	.w7(32'h3c960e38),
	.w8(32'hbb58c62b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a280),
	.w1(32'h3c30f7fd),
	.w2(32'hbcef3d0d),
	.w3(32'hbcb217d3),
	.w4(32'h3973c244),
	.w5(32'hbc58a858),
	.w6(32'h3c7a4d24),
	.w7(32'hbc772890),
	.w8(32'hbd075e85),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc392d1),
	.w1(32'h3cdafc6e),
	.w2(32'hbb4d6312),
	.w3(32'h3b6caf04),
	.w4(32'h3bb41abd),
	.w5(32'hbd0660d8),
	.w6(32'h3c88d45e),
	.w7(32'hbc24868d),
	.w8(32'hbb8e4f71),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc0e1e9),
	.w1(32'hb97e43b1),
	.w2(32'hba70ef6a),
	.w3(32'h3b9ef13c),
	.w4(32'hbbdeda93),
	.w5(32'hbc1464c9),
	.w6(32'hbaadbb7f),
	.w7(32'hba2c77c9),
	.w8(32'h3c11ceb3),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2e5df),
	.w1(32'hba754464),
	.w2(32'hbc6242ef),
	.w3(32'h3c8ac907),
	.w4(32'h3bdfef2d),
	.w5(32'hbc40f4f7),
	.w6(32'h3b586e7f),
	.w7(32'hbc666bcb),
	.w8(32'hbb31cbdc),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c6a63),
	.w1(32'h3be6b191),
	.w2(32'hbc81c836),
	.w3(32'h3c53ffb1),
	.w4(32'hbbf18a02),
	.w5(32'h3c1dde7b),
	.w6(32'h3bd081e0),
	.w7(32'hbb272273),
	.w8(32'h3b3984a4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89c17b),
	.w1(32'hbc7765ab),
	.w2(32'hbcbd864c),
	.w3(32'h3b956230),
	.w4(32'hbbcf7d63),
	.w5(32'h3c873a5c),
	.w6(32'hbba3caeb),
	.w7(32'h3bd6df74),
	.w8(32'hbc5f2e06),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa616aa),
	.w1(32'h3b8a4777),
	.w2(32'hbbe8c06e),
	.w3(32'hb9a34013),
	.w4(32'hbc09aea6),
	.w5(32'h3b4e021a),
	.w6(32'h3cc1e081),
	.w7(32'h3ca3fcea),
	.w8(32'h3ae852d4),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87f3a2),
	.w1(32'h3b406b9b),
	.w2(32'hbc283c22),
	.w3(32'h3bc075cf),
	.w4(32'hbc043146),
	.w5(32'h3c01fd49),
	.w6(32'h39bdd29c),
	.w7(32'h3a6c4cf4),
	.w8(32'hbc181a1e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c010c6c),
	.w1(32'h3c0c094c),
	.w2(32'h3c1d46b2),
	.w3(32'h3b9e6330),
	.w4(32'h3b92790e),
	.w5(32'hbbd655fa),
	.w6(32'hbc206949),
	.w7(32'h3aed20ad),
	.w8(32'h3b6131db),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbeebab),
	.w1(32'hba6f6adb),
	.w2(32'hbc074507),
	.w3(32'h394c5307),
	.w4(32'h3a1a6384),
	.w5(32'hbc5084cd),
	.w6(32'hbc7f9e18),
	.w7(32'hbcd23ec6),
	.w8(32'h3b2409d0),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30b182),
	.w1(32'hbb9bf789),
	.w2(32'h3bc6e7cd),
	.w3(32'hbcc3b259),
	.w4(32'hbc58b958),
	.w5(32'h3c8595c9),
	.w6(32'hbc8c0155),
	.w7(32'hbc1b7af0),
	.w8(32'h3c1d4fc8),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a046f33),
	.w1(32'h3ba11246),
	.w2(32'h3a8357dd),
	.w3(32'h3b89c4f0),
	.w4(32'hbc6675af),
	.w5(32'h3c0e2a20),
	.w6(32'hbcebf720),
	.w7(32'h3bf43091),
	.w8(32'hbc1c0d41),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac07f1a),
	.w1(32'hb96b5144),
	.w2(32'h3afa6080),
	.w3(32'h3b8e81f0),
	.w4(32'hba9135c0),
	.w5(32'hbaf26e9e),
	.w6(32'h3b0fa600),
	.w7(32'h3c6346d8),
	.w8(32'hba3ec782),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e1ec1),
	.w1(32'h3b605b39),
	.w2(32'hbb039096),
	.w3(32'hbc092b27),
	.w4(32'h3b194a23),
	.w5(32'hbaadf27f),
	.w6(32'h3c8127dc),
	.w7(32'hbb81d650),
	.w8(32'hb8bc0273),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396b5c97),
	.w1(32'h3b494526),
	.w2(32'h3b3658e7),
	.w3(32'h3bbb0ab6),
	.w4(32'hbb7fab3b),
	.w5(32'h3c9a5a0d),
	.w6(32'h3c2155cd),
	.w7(32'h3c0b5f18),
	.w8(32'hbb5562be),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012f16),
	.w1(32'h3996f5c4),
	.w2(32'h3c27fff4),
	.w3(32'hbb8449d1),
	.w4(32'h3ab29ff9),
	.w5(32'hbc38e829),
	.w6(32'hbc46190d),
	.w7(32'h3b56546e),
	.w8(32'h3a8fb8ae),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b262653),
	.w1(32'hba6245e7),
	.w2(32'h3c171397),
	.w3(32'hbc0ae1b8),
	.w4(32'hba132ec4),
	.w5(32'h3b809e54),
	.w6(32'h3abfc45a),
	.w7(32'hbb38c8b4),
	.w8(32'hbc0582e7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb42d0383),
	.w1(32'hbb836677),
	.w2(32'h3b37cef2),
	.w3(32'h3c624971),
	.w4(32'hbb0d5ba3),
	.w5(32'hbbf21cac),
	.w6(32'h3b413d50),
	.w7(32'h3c5ec995),
	.w8(32'hbaa7a6da),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf936fb),
	.w1(32'h3c95412f),
	.w2(32'h3b15fe58),
	.w3(32'hbc532256),
	.w4(32'h3d143e8a),
	.w5(32'h3b7e10cb),
	.w6(32'h3ca4aa20),
	.w7(32'hbac7034f),
	.w8(32'h3c6633ac),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1d147),
	.w1(32'hbcac9aea),
	.w2(32'h3b4b8a94),
	.w3(32'h398e52e4),
	.w4(32'h3bf1e03a),
	.w5(32'h3b19d708),
	.w6(32'h3b9f2d45),
	.w7(32'h3a95e7d0),
	.w8(32'h3aa987a1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58ee65),
	.w1(32'hbbd732f5),
	.w2(32'h3b1adc27),
	.w3(32'h3b4fe8db),
	.w4(32'hbb0a9e71),
	.w5(32'hbc20df61),
	.w6(32'h3bd7a5fd),
	.w7(32'hbc6f2551),
	.w8(32'hbc298cd9),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9ba98),
	.w1(32'h3a0f5661),
	.w2(32'h3c136299),
	.w3(32'hbb663a0d),
	.w4(32'h3b7bf0f6),
	.w5(32'h3be225a8),
	.w6(32'h3ba025df),
	.w7(32'h3af969bd),
	.w8(32'hbcba1912),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcae5366),
	.w1(32'h3ce9a696),
	.w2(32'hbd08b757),
	.w3(32'hbc5dcdb7),
	.w4(32'hbbcb2450),
	.w5(32'h3b10ea76),
	.w6(32'h38a1c8f5),
	.w7(32'hbb4aa536),
	.w8(32'hbb22b68d),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b002d32),
	.w1(32'h3be66eb9),
	.w2(32'hbc87ae54),
	.w3(32'hbc171e48),
	.w4(32'hbb1a36a6),
	.w5(32'hbc49156b),
	.w6(32'h3a6ad862),
	.w7(32'h3bb82188),
	.w8(32'h3aed4453),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8e10f6),
	.w1(32'h3a7d9600),
	.w2(32'hbc25c712),
	.w3(32'h3b981fad),
	.w4(32'hbbf4da2e),
	.w5(32'hbba08339),
	.w6(32'h3c49b39a),
	.w7(32'hbba46ff2),
	.w8(32'h3c08b630),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb530c8d),
	.w1(32'h3b5876ec),
	.w2(32'hbb76311c),
	.w3(32'hbb20dd91),
	.w4(32'hbb997b62),
	.w5(32'hbb037910),
	.w6(32'hbcf8ddc7),
	.w7(32'hbb9ed0bd),
	.w8(32'h3a889ebd),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule