module layer_10_featuremap_455(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb525cf),
	.w1(32'hbb9a020b),
	.w2(32'hbb26837c),
	.w3(32'hbb9c30d5),
	.w4(32'hbc1b534e),
	.w5(32'hb9d52b67),
	.w6(32'hbad028ec),
	.w7(32'hbb4b22a6),
	.w8(32'hba884d22),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee4019),
	.w1(32'h3be7c6f0),
	.w2(32'h3b6b9540),
	.w3(32'hbaddbb2e),
	.w4(32'hbbcfd70e),
	.w5(32'hbc0f3b7c),
	.w6(32'hbba87d5b),
	.w7(32'h3ba394f2),
	.w8(32'hbbbcdcfa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9606f),
	.w1(32'hbc862353),
	.w2(32'hbc1b5b04),
	.w3(32'h3beaf60d),
	.w4(32'h3aaa9301),
	.w5(32'hbc63f68a),
	.w6(32'h3a5b683b),
	.w7(32'hbc4a7137),
	.w8(32'h3c88ced5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1eefde),
	.w1(32'h3b8e0721),
	.w2(32'h3ba34075),
	.w3(32'hbb8a91c4),
	.w4(32'h3bfc1f2b),
	.w5(32'hba352d41),
	.w6(32'hbc72c52d),
	.w7(32'h3bd789c9),
	.w8(32'h3caadb58),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c433b70),
	.w1(32'h3b51a8d9),
	.w2(32'hba6287e2),
	.w3(32'h3d11cb0e),
	.w4(32'hbaa895ee),
	.w5(32'h3c1f036d),
	.w6(32'h3c342230),
	.w7(32'h3b031ed8),
	.w8(32'h3aaa78db),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83d492),
	.w1(32'hbb8697ab),
	.w2(32'hbc5d6e4f),
	.w3(32'hbb9187b5),
	.w4(32'hbb21a8c1),
	.w5(32'h3c073998),
	.w6(32'hbaafee5e),
	.w7(32'hba536802),
	.w8(32'hbbcb3765),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42758f),
	.w1(32'h3b86c2ab),
	.w2(32'hbb8449b6),
	.w3(32'hbbbc3c49),
	.w4(32'hbb199ba3),
	.w5(32'hbc8f4dba),
	.w6(32'hbc05c6f7),
	.w7(32'hbbdf8044),
	.w8(32'h3b1a4e58),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92460d8),
	.w1(32'h3c2914df),
	.w2(32'hbc54d682),
	.w3(32'hbc1c683b),
	.w4(32'h3c6f5b4a),
	.w5(32'h3b992d0b),
	.w6(32'hba6c1eca),
	.w7(32'h3c0bb5a6),
	.w8(32'h3cb59c2c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11c18a),
	.w1(32'h3b20c74e),
	.w2(32'h3c78e438),
	.w3(32'h3a843c60),
	.w4(32'h3b5d84d1),
	.w5(32'h3c926047),
	.w6(32'h3b8c3d9f),
	.w7(32'h3c0b6806),
	.w8(32'h3ca999cc),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e2e4ae),
	.w1(32'hbaafb558),
	.w2(32'h3ad9f53f),
	.w3(32'h3d40341f),
	.w4(32'h3bbba670),
	.w5(32'h39d22a34),
	.w6(32'h3c1284ad),
	.w7(32'hba67ba77),
	.w8(32'hbbda99be),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc4a42),
	.w1(32'hbb084ad4),
	.w2(32'h3bff83be),
	.w3(32'hb9eb998d),
	.w4(32'hbbad6c69),
	.w5(32'hbbfe3763),
	.w6(32'hbc0c5a05),
	.w7(32'hbc794a2e),
	.w8(32'hbc2fc73e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14cd53),
	.w1(32'hbafb4dca),
	.w2(32'h3906bd01),
	.w3(32'hbb92955d),
	.w4(32'hbbab6baf),
	.w5(32'h3c9d9005),
	.w6(32'hbc384ba0),
	.w7(32'hbba0726d),
	.w8(32'h3b221c57),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb0fee),
	.w1(32'hbc270452),
	.w2(32'hbc7dac25),
	.w3(32'hbb00b37d),
	.w4(32'hbc12ddf6),
	.w5(32'hbc6b7056),
	.w6(32'hb9f884af),
	.w7(32'hbc47d051),
	.w8(32'hbc913f12),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3127c5),
	.w1(32'hbc8d770c),
	.w2(32'h3c711259),
	.w3(32'hbca5085a),
	.w4(32'hbc6b51a0),
	.w5(32'h3c93a91d),
	.w6(32'hbc8585c6),
	.w7(32'h3bc9906c),
	.w8(32'hbc5528fd),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a1c33),
	.w1(32'h3b23615b),
	.w2(32'hbb083928),
	.w3(32'h3bdc4b4c),
	.w4(32'h3cd361d7),
	.w5(32'h3cc1647b),
	.w6(32'hba4ecc06),
	.w7(32'hbb2ba54b),
	.w8(32'h3ce87951),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5eeafd),
	.w1(32'h3bd2e8ee),
	.w2(32'h3b7ee3d5),
	.w3(32'hbc09c494),
	.w4(32'h3c9395fa),
	.w5(32'hb919d846),
	.w6(32'h3bf18214),
	.w7(32'h388a821a),
	.w8(32'h3b6b38aa),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebaba4),
	.w1(32'hb9d36ea4),
	.w2(32'h3b0b53a4),
	.w3(32'hbc2fdd92),
	.w4(32'hbc01e27b),
	.w5(32'hbc150344),
	.w6(32'hba857151),
	.w7(32'hbc7828f9),
	.w8(32'hbc873ac0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb08cf),
	.w1(32'hbb2958c5),
	.w2(32'hbc086bc5),
	.w3(32'hbaac8aaa),
	.w4(32'hbbcaaf23),
	.w5(32'hbbc2125a),
	.w6(32'hbc324ca8),
	.w7(32'hbbd07dae),
	.w8(32'hbc2d7b43),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9c4c90),
	.w1(32'hbcd4b080),
	.w2(32'hbc8e9ba3),
	.w3(32'hbc656323),
	.w4(32'hbd04d99f),
	.w5(32'hbcaecf2d),
	.w6(32'hbc927f29),
	.w7(32'hbce904d4),
	.w8(32'hbc991ade),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07247a),
	.w1(32'h3b7e828f),
	.w2(32'h3b778101),
	.w3(32'hbc0c7598),
	.w4(32'hbad3e6b6),
	.w5(32'h3bba034d),
	.w6(32'hbc440a7b),
	.w7(32'hbc6be070),
	.w8(32'hbbdaf58b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02d804),
	.w1(32'h3c17b8c2),
	.w2(32'h3bd6d6bc),
	.w3(32'hbc256276),
	.w4(32'h3cbf87f9),
	.w5(32'h3c2070df),
	.w6(32'h3b72d537),
	.w7(32'h3baab6bf),
	.w8(32'hbc020a61),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0955b),
	.w1(32'hbba3c779),
	.w2(32'hbbf5b3b8),
	.w3(32'hbca53842),
	.w4(32'hbbacb8e7),
	.w5(32'hbb8074b9),
	.w6(32'hbc84892d),
	.w7(32'hbba32cc8),
	.w8(32'h3b73af69),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a812bed),
	.w1(32'h3ba8e024),
	.w2(32'h3b1fdea8),
	.w3(32'hbb80ecfc),
	.w4(32'h3be61ab4),
	.w5(32'h3aa1a072),
	.w6(32'h3b00a5b1),
	.w7(32'hbbbc6c3c),
	.w8(32'h3a89f616),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb83acb),
	.w1(32'h3bb818e5),
	.w2(32'hbb9b3226),
	.w3(32'h3bd64ed5),
	.w4(32'h3bd38fe6),
	.w5(32'hba8980a7),
	.w6(32'hbc062b73),
	.w7(32'hbaf76ebf),
	.w8(32'hbc08ae42),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7df73),
	.w1(32'h3bbafa9b),
	.w2(32'h3be0affa),
	.w3(32'hb907ffaa),
	.w4(32'h3c6f7354),
	.w5(32'hbb89e016),
	.w6(32'hbbbf7e47),
	.w7(32'h3bf2b82a),
	.w8(32'hbadf4955),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c085d),
	.w1(32'h3bd90aff),
	.w2(32'h389e8980),
	.w3(32'hbb365b2f),
	.w4(32'h3bd51783),
	.w5(32'hbbbb8aed),
	.w6(32'hbbefa211),
	.w7(32'h3a900773),
	.w8(32'h3a638730),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c59b8e5),
	.w1(32'h3a8af322),
	.w2(32'h3babf681),
	.w3(32'h3c7f212e),
	.w4(32'h3b9aed12),
	.w5(32'hbbff10e1),
	.w6(32'h3b695fd2),
	.w7(32'h3ae1e038),
	.w8(32'h3be93a8a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72f504),
	.w1(32'h3c2baab6),
	.w2(32'h3b20c868),
	.w3(32'hbadb0734),
	.w4(32'h3c074ac4),
	.w5(32'hbc31f52f),
	.w6(32'hbad693e0),
	.w7(32'h3ba0d510),
	.w8(32'h3b06e53a),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b959685),
	.w1(32'h3c92801f),
	.w2(32'h3bfa6b69),
	.w3(32'h3b8a4c81),
	.w4(32'h3b78d9c2),
	.w5(32'h3bb30a8c),
	.w6(32'h3bc681e8),
	.w7(32'hbb0bb804),
	.w8(32'hbaabe380),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c044a57),
	.w1(32'hbadb09f7),
	.w2(32'hba73b7eb),
	.w3(32'hba4c39f8),
	.w4(32'h3c2170d6),
	.w5(32'h3c19a4f0),
	.w6(32'hbc5b5715),
	.w7(32'h3baabf1a),
	.w8(32'h3baee5c2),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09988d),
	.w1(32'h3b8630ef),
	.w2(32'hbbd60e84),
	.w3(32'hbcdd689c),
	.w4(32'h3b4153c8),
	.w5(32'h3c8dab90),
	.w6(32'hbbca0d58),
	.w7(32'hbbd26d08),
	.w8(32'h3be0e76b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8db03d),
	.w1(32'h3b32b8fe),
	.w2(32'hbaba8cf7),
	.w3(32'h3c139e65),
	.w4(32'h3cd86273),
	.w5(32'h3c1e1d89),
	.w6(32'h3b8a4280),
	.w7(32'h3c1f3525),
	.w8(32'h3c3756b5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11a88d),
	.w1(32'h3835304a),
	.w2(32'h3c88df0a),
	.w3(32'hbbb7649b),
	.w4(32'hb9f19c73),
	.w5(32'h3a31dce6),
	.w6(32'hba99030f),
	.w7(32'hbac756a7),
	.w8(32'hbbeef7c5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9528f7),
	.w1(32'h3b995a9e),
	.w2(32'h3b0d5bfb),
	.w3(32'hbb76b0e9),
	.w4(32'h39f5783e),
	.w5(32'hbc3ca0a0),
	.w6(32'hbbb9ebb6),
	.w7(32'h3aa59218),
	.w8(32'hbbf20132),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5ec6),
	.w1(32'h3b9138e1),
	.w2(32'h3c5ddd81),
	.w3(32'hbbeb1bac),
	.w4(32'hbbf68c95),
	.w5(32'hb9591f6a),
	.w6(32'hbbbd58f3),
	.w7(32'hbb60abcb),
	.w8(32'hbca23789),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cf293),
	.w1(32'hbabb2847),
	.w2(32'hbb4835f5),
	.w3(32'hbc026647),
	.w4(32'hbb9d72ca),
	.w5(32'hbaeaec10),
	.w6(32'hbc576476),
	.w7(32'hbb0b0369),
	.w8(32'h3b350276),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81c9c79),
	.w1(32'h3b763dea),
	.w2(32'h3c3508b6),
	.w3(32'h3c61ff1e),
	.w4(32'h3bd0e295),
	.w5(32'hbc0f847b),
	.w6(32'h3b1c22e9),
	.w7(32'hbbd61f7f),
	.w8(32'hbbbd1fd9),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2cce47),
	.w1(32'hbc48d12a),
	.w2(32'hbc5e9cb8),
	.w3(32'h3ad48e45),
	.w4(32'hbc85b35b),
	.w5(32'hbb40a02a),
	.w6(32'hbbf8ac93),
	.w7(32'hbc4a4188),
	.w8(32'hbc190f27),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a12b1),
	.w1(32'hbb6f6c01),
	.w2(32'h39737bc1),
	.w3(32'hbc9b3415),
	.w4(32'hbc453ee5),
	.w5(32'hbc247e9b),
	.w6(32'hbc58ff95),
	.w7(32'hbac377c7),
	.w8(32'hbbb764c1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c20a1),
	.w1(32'hbb1888ff),
	.w2(32'h3915b14c),
	.w3(32'h3c07e438),
	.w4(32'hbc21a206),
	.w5(32'h3b2df628),
	.w6(32'hbc119bcc),
	.w7(32'hbb8d3774),
	.w8(32'h3ad0d5c6),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa938fd),
	.w1(32'hbc915445),
	.w2(32'hbb35de3f),
	.w3(32'h3c381c95),
	.w4(32'hbc8a4810),
	.w5(32'h3db93d6d),
	.w6(32'h3b8e4641),
	.w7(32'hbc5b8f66),
	.w8(32'hbc4bfeac),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99a712),
	.w1(32'hbb1e7bd6),
	.w2(32'h3c4e071d),
	.w3(32'hbcda7b3f),
	.w4(32'h3c28b742),
	.w5(32'h3d5970d8),
	.w6(32'hbb8c4dd0),
	.w7(32'hbc2e16f3),
	.w8(32'h3c83698d),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c279583),
	.w1(32'h3b04c463),
	.w2(32'hbb05859f),
	.w3(32'h3c5d5b3c),
	.w4(32'h3b24c56d),
	.w5(32'hbc1b4529),
	.w6(32'h3c82d246),
	.w7(32'hbb558adc),
	.w8(32'h39a95947),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d1698),
	.w1(32'hbba32abe),
	.w2(32'hbad26241),
	.w3(32'hbbbbc9d7),
	.w4(32'hbbbc0a49),
	.w5(32'hbbd96358),
	.w6(32'h3b7672f9),
	.w7(32'h3b12a5e7),
	.w8(32'h39e861cf),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393ab1bb),
	.w1(32'hbbb7fc3e),
	.w2(32'hbb9db152),
	.w3(32'h3bc2cd84),
	.w4(32'hbb6fa66a),
	.w5(32'hbc172d1a),
	.w6(32'h3b2b49b4),
	.w7(32'hbbd24958),
	.w8(32'hbc1ab56c),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2d036),
	.w1(32'hba1c2bfc),
	.w2(32'h3c0e9e5e),
	.w3(32'hbc42f595),
	.w4(32'h3bb9861b),
	.w5(32'hbc901082),
	.w6(32'hbb833131),
	.w7(32'h3ab5cde6),
	.w8(32'hbb8301b2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf801ed),
	.w1(32'hbbb156e8),
	.w2(32'h3ac8e5cd),
	.w3(32'hbacbb253),
	.w4(32'hba969489),
	.w5(32'hbc5faaa3),
	.w6(32'h3befbc44),
	.w7(32'hbc03fd63),
	.w8(32'hbc9537d5),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95acff),
	.w1(32'hbc0fa635),
	.w2(32'hbc3dcf32),
	.w3(32'hbc513e33),
	.w4(32'hbc93f331),
	.w5(32'hbc999bd3),
	.w6(32'hbc410c86),
	.w7(32'hbb23c0bd),
	.w8(32'hbc0edc2e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c74e6),
	.w1(32'hbc662ee5),
	.w2(32'h3acbe3a8),
	.w3(32'hbc3de200),
	.w4(32'hbcb2fb5b),
	.w5(32'h3b8b1d07),
	.w6(32'hbc6f2d8d),
	.w7(32'hbbe8db84),
	.w8(32'hbc0c923f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5488),
	.w1(32'h3c42d6ae),
	.w2(32'hbb95be5d),
	.w3(32'h3c55e18d),
	.w4(32'h3c98416f),
	.w5(32'h3c63469d),
	.w6(32'hb963a03c),
	.w7(32'h3c70be20),
	.w8(32'h3bbe6fff),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc701b27),
	.w1(32'hb9ff56bb),
	.w2(32'hbc2e8dd3),
	.w3(32'hbcb99094),
	.w4(32'hbbe69f18),
	.w5(32'h3c04c3ba),
	.w6(32'hbbd204bf),
	.w7(32'hba92fe06),
	.w8(32'hbba4d7d5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86325a),
	.w1(32'h3baf003b),
	.w2(32'h3aacafcf),
	.w3(32'h3b9c5be8),
	.w4(32'h3bb186fb),
	.w5(32'hbb85d7d0),
	.w6(32'hbbd673ab),
	.w7(32'h3bf70f73),
	.w8(32'hba464f85),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe45ca),
	.w1(32'h3b24b836),
	.w2(32'hbb4523a1),
	.w3(32'hbb2904b2),
	.w4(32'hbaad5faf),
	.w5(32'h3c30edf4),
	.w6(32'hba60a886),
	.w7(32'h3aec02b4),
	.w8(32'h3b4e0244),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdbe20),
	.w1(32'h3aa67f2c),
	.w2(32'h3c82fa32),
	.w3(32'h3c32b708),
	.w4(32'hbaca1d3a),
	.w5(32'h3ba55556),
	.w6(32'h390aec4b),
	.w7(32'hb9d91095),
	.w8(32'hbc8a03bc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19f897),
	.w1(32'hbb4da5f6),
	.w2(32'hba575e5b),
	.w3(32'h3c94321f),
	.w4(32'h3ba83140),
	.w5(32'h3befefa3),
	.w6(32'h3b967910),
	.w7(32'h3b21b643),
	.w8(32'h3c2bf32d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd18df),
	.w1(32'h390b7680),
	.w2(32'h3c8ceb34),
	.w3(32'hbbca689f),
	.w4(32'hba71dace),
	.w5(32'h3c0d832c),
	.w6(32'hbb68854a),
	.w7(32'h3c3c47fc),
	.w8(32'h3a5a5417),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ddbb4),
	.w1(32'hbae90825),
	.w2(32'hbbd06a54),
	.w3(32'h3cfcb277),
	.w4(32'h3b08dad8),
	.w5(32'h3a7cf8b4),
	.w6(32'h3bedf02e),
	.w7(32'h376bd366),
	.w8(32'h3a5d22e6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7eeec),
	.w1(32'hbbd622db),
	.w2(32'hbb4e8d4a),
	.w3(32'hbc6d79a8),
	.w4(32'h3b30edd3),
	.w5(32'hbb703073),
	.w6(32'hbc0d2184),
	.w7(32'hbbe3b820),
	.w8(32'hb9927e2c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcaae9a),
	.w1(32'h3b37c844),
	.w2(32'hbbd6e6db),
	.w3(32'h3b81558d),
	.w4(32'h3b6cdc10),
	.w5(32'h3ae5ac2b),
	.w6(32'hbb0f6200),
	.w7(32'h3aea4f3d),
	.w8(32'hbb3dd876),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb616c18),
	.w1(32'h3b7b3089),
	.w2(32'h3bbc053e),
	.w3(32'hbb86f5ac),
	.w4(32'h3ba42aad),
	.w5(32'hbb8f033d),
	.w6(32'hbb859100),
	.w7(32'h3c5d511f),
	.w8(32'h3bd5a57f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a973379),
	.w1(32'hbb5c6cfe),
	.w2(32'h3b9fc4d3),
	.w3(32'h3c19dd3f),
	.w4(32'h3c00f18b),
	.w5(32'hbb065c11),
	.w6(32'h38ec2ff7),
	.w7(32'h3b805b9c),
	.w8(32'hbb3148c6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b5272),
	.w1(32'h3c233ef8),
	.w2(32'hba4aebf1),
	.w3(32'h3b89880c),
	.w4(32'h3cc34c9b),
	.w5(32'h3c1c472e),
	.w6(32'hbbc91ffc),
	.w7(32'h3c130197),
	.w8(32'h3c1c7d68),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bbd97),
	.w1(32'h3b8c084d),
	.w2(32'hbbdaabff),
	.w3(32'hbc6c1e90),
	.w4(32'h3c20c1e9),
	.w5(32'hbbc26d73),
	.w6(32'h3a9ee649),
	.w7(32'hbbef1257),
	.w8(32'hbc5d7328),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb6a04c),
	.w1(32'hbb1ccc6a),
	.w2(32'h3b036b04),
	.w3(32'hbd0c4a34),
	.w4(32'hbbc3cd8d),
	.w5(32'h3c6b2297),
	.w6(32'hbcc08df0),
	.w7(32'hba405f4b),
	.w8(32'h3962c8c0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a2b7d),
	.w1(32'h3afe7647),
	.w2(32'h3b1525f1),
	.w3(32'h3b85aaa6),
	.w4(32'h3bcdb9c2),
	.w5(32'h3b6f209f),
	.w6(32'h3b372c81),
	.w7(32'h3b189cbd),
	.w8(32'hbbcca990),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810e17),
	.w1(32'hbae135b9),
	.w2(32'hba2ae7b9),
	.w3(32'hbb8c305d),
	.w4(32'hbc4e4ae9),
	.w5(32'hbc5297d0),
	.w6(32'hbc06bdfd),
	.w7(32'hbbb3e37a),
	.w8(32'hbc00c2b7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be024d5),
	.w1(32'hbc420e03),
	.w2(32'hbcaa268f),
	.w3(32'h3c23a26d),
	.w4(32'hbc817519),
	.w5(32'hbcc834bb),
	.w6(32'h3beff7d6),
	.w7(32'hbb59203b),
	.w8(32'hbc6d0c58),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1930e),
	.w1(32'hbac8a5c1),
	.w2(32'h3bae1b96),
	.w3(32'hbcc80aed),
	.w4(32'h3bcedbaf),
	.w5(32'hbca8a133),
	.w6(32'hbc82ec86),
	.w7(32'h3bf89abf),
	.w8(32'h3b150439),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5374c0),
	.w1(32'h3c03f59d),
	.w2(32'hbc16f466),
	.w3(32'hbc2684db),
	.w4(32'hbb5e2bb7),
	.w5(32'hbc939e27),
	.w6(32'h3981c9d9),
	.w7(32'h3b21570e),
	.w8(32'hbbb6f637),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc090dab),
	.w1(32'h3b86c4ed),
	.w2(32'h3a7aa067),
	.w3(32'h3ba74b27),
	.w4(32'h3a8393d1),
	.w5(32'h3b41a19f),
	.w6(32'hbbb19413),
	.w7(32'hbaa4be64),
	.w8(32'h3baea0d4),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a149b07),
	.w1(32'hbb53d427),
	.w2(32'hbacbe583),
	.w3(32'h3b2d1dfe),
	.w4(32'h3a9522f3),
	.w5(32'hba729f9d),
	.w6(32'h3bd91854),
	.w7(32'hba157da1),
	.w8(32'hba9a65ff),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf113b9),
	.w1(32'hbacdc8a2),
	.w2(32'hbba78f35),
	.w3(32'hbb91ead4),
	.w4(32'hbb4b659f),
	.w5(32'hbc84a31e),
	.w6(32'hbbe73ac7),
	.w7(32'h3b931f98),
	.w8(32'hbba6767d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f8972),
	.w1(32'hbba767ad),
	.w2(32'h3c79d3d0),
	.w3(32'hbb8a07f5),
	.w4(32'hb9c6c8de),
	.w5(32'h3c71a2c2),
	.w6(32'hbbd7fa04),
	.w7(32'hbb814e65),
	.w8(32'h3c3df283),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6fc72),
	.w1(32'hba849ca9),
	.w2(32'h3a3e53cb),
	.w3(32'h3a3a493b),
	.w4(32'hbac50c19),
	.w5(32'hbb7cb1df),
	.w6(32'h3acf1c32),
	.w7(32'hbaa22f15),
	.w8(32'hbb3bedb1),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42c643),
	.w1(32'hbb9a61a4),
	.w2(32'hbbc8d08f),
	.w3(32'h3abc7581),
	.w4(32'hbb4d3473),
	.w5(32'hbbbfd882),
	.w6(32'hbb159bd2),
	.w7(32'hb9a4838f),
	.w8(32'hbb306d7a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b03b92),
	.w1(32'h3a84fb29),
	.w2(32'hba8e872f),
	.w3(32'hbb5aaaf0),
	.w4(32'h3af2dad5),
	.w5(32'hbb8d281c),
	.w6(32'h39f69b98),
	.w7(32'hb9e92c24),
	.w8(32'hbb1cf56f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0f49c),
	.w1(32'h3b36d183),
	.w2(32'hbb87c4f0),
	.w3(32'hbb16d6c5),
	.w4(32'h3af5812b),
	.w5(32'hbbeab9fb),
	.w6(32'hbbab76f4),
	.w7(32'h3b0ed5b5),
	.w8(32'hbab81be2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6a03d9),
	.w1(32'h3a728cc3),
	.w2(32'h3b654598),
	.w3(32'hbb320da8),
	.w4(32'hb9ea4d2e),
	.w5(32'h3c85c728),
	.w6(32'hbb3f426e),
	.w7(32'hb6e8f62a),
	.w8(32'h3a8ab954),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbebd2bd),
	.w1(32'h3ab37b18),
	.w2(32'h3bb537d7),
	.w3(32'hbac780ac),
	.w4(32'h3b449401),
	.w5(32'h3c031a0d),
	.w6(32'h3ae109e4),
	.w7(32'h3a51397d),
	.w8(32'h3ababac5),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa902b9),
	.w1(32'h39c8c34d),
	.w2(32'hbb8a47a9),
	.w3(32'hba690337),
	.w4(32'h3abf8665),
	.w5(32'h3adbcc28),
	.w6(32'h38265833),
	.w7(32'h38b18ff4),
	.w8(32'h3ae02cb5),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3469d5),
	.w1(32'h3bd0ac13),
	.w2(32'h3b1c8530),
	.w3(32'hbb8deebb),
	.w4(32'h3c0c0bb5),
	.w5(32'hbbb7a692),
	.w6(32'hbac798fb),
	.w7(32'h3c14d2f6),
	.w8(32'h3b95954a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aa993),
	.w1(32'hb91e937c),
	.w2(32'h3a0b92a4),
	.w3(32'h3b8efe66),
	.w4(32'hbb0af13a),
	.w5(32'h39f5be1a),
	.w6(32'h3c12a664),
	.w7(32'hbb631bf2),
	.w8(32'hbb847917),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9496b83),
	.w1(32'h398e218e),
	.w2(32'hbb6b2e6f),
	.w3(32'hb74ebb2b),
	.w4(32'hb85afa5e),
	.w5(32'hbb84a7e8),
	.w6(32'hba4b9afe),
	.w7(32'h3a850ac1),
	.w8(32'h3b0e5e2c),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1ff42),
	.w1(32'h3a84c20e),
	.w2(32'hbaa105e2),
	.w3(32'h39976262),
	.w4(32'h3a3eda81),
	.w5(32'h3abaa662),
	.w6(32'h3aea70cf),
	.w7(32'hbaf7bc27),
	.w8(32'h3b8133ad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4b8d3),
	.w1(32'hbc0d86e8),
	.w2(32'h3b869946),
	.w3(32'hbb501eb7),
	.w4(32'hbbea7b5f),
	.w5(32'h3aed236c),
	.w6(32'hbbe9d811),
	.w7(32'hbb95cb6d),
	.w8(32'hbb06931a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff50a2),
	.w1(32'hb9bb9ede),
	.w2(32'h3c7263a5),
	.w3(32'hbc0b2019),
	.w4(32'hbb2a01c7),
	.w5(32'h3cc7d2df),
	.w6(32'hbb061874),
	.w7(32'hbc04be7f),
	.w8(32'h3c17bb13),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ed4a4),
	.w1(32'hbb01c4f7),
	.w2(32'hbbadf010),
	.w3(32'hba91ad60),
	.w4(32'h3b794fde),
	.w5(32'hbb343221),
	.w6(32'h3a9445e4),
	.w7(32'h3ba19db0),
	.w8(32'hbadb0944),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68546c),
	.w1(32'hbb642d03),
	.w2(32'hbb3dbe20),
	.w3(32'hba71191e),
	.w4(32'hba7204c9),
	.w5(32'hbc24ae51),
	.w6(32'hbb8030e3),
	.w7(32'h3ba7442c),
	.w8(32'hbbb5cd21),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07bb82),
	.w1(32'hba8ba2bb),
	.w2(32'hbbce4d68),
	.w3(32'hb98149ac),
	.w4(32'hbaa76bd4),
	.w5(32'hbc2c0d72),
	.w6(32'hba98474a),
	.w7(32'hbabbd0b8),
	.w8(32'hbc0a81ce),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb1f94),
	.w1(32'hbb559c08),
	.w2(32'hb9a84168),
	.w3(32'h3c591d2a),
	.w4(32'hbb956976),
	.w5(32'h3c10a888),
	.w6(32'h3b630d46),
	.w7(32'hbb439534),
	.w8(32'hbb2595c6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ad42a),
	.w1(32'hbadb2fa0),
	.w2(32'h3a92f529),
	.w3(32'hba5ae6bd),
	.w4(32'h3a378ddd),
	.w5(32'hbab9c3c8),
	.w6(32'hbada5928),
	.w7(32'h3b309d3a),
	.w8(32'hbbc054e3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a7613),
	.w1(32'hba49ee0e),
	.w2(32'hbc486eff),
	.w3(32'h3a8e6378),
	.w4(32'h3c0d2aef),
	.w5(32'hbbae26f5),
	.w6(32'h3a6de17b),
	.w7(32'hbb23f70a),
	.w8(32'hbc058bde),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895df93),
	.w1(32'h3b31bba7),
	.w2(32'h3b84cac1),
	.w3(32'hbaa29f94),
	.w4(32'h3b47bfa0),
	.w5(32'h3a2be7ca),
	.w6(32'hbb8cf1e7),
	.w7(32'h3a96d641),
	.w8(32'hbab7fc35),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba72bc),
	.w1(32'hba0beed1),
	.w2(32'hb9add28b),
	.w3(32'h3ac44095),
	.w4(32'h39e39af2),
	.w5(32'hbb640c40),
	.w6(32'hbab22b49),
	.w7(32'hba977c4a),
	.w8(32'hbb8e7ddd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45efb0),
	.w1(32'hbb826646),
	.w2(32'hbc11068b),
	.w3(32'hbad5f59f),
	.w4(32'hbacda57f),
	.w5(32'hbac51ab5),
	.w6(32'hbb450d9a),
	.w7(32'hbc01a0d3),
	.w8(32'hbbb8f8a4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebc7d6),
	.w1(32'h3b85ffca),
	.w2(32'hbbc4afba),
	.w3(32'hbbf06bdf),
	.w4(32'h3c2e81f5),
	.w5(32'hbbb4a96e),
	.w6(32'hbb1b06da),
	.w7(32'h3bc0677b),
	.w8(32'h3b6d92f8),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46801d),
	.w1(32'hbb7db089),
	.w2(32'h3ab7c961),
	.w3(32'h3ac90f88),
	.w4(32'hbb20a8f7),
	.w5(32'hbb8a1c19),
	.w6(32'hbadb5d4b),
	.w7(32'hbc09ea43),
	.w8(32'hbbeb945a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedd6e3),
	.w1(32'hb996f65f),
	.w2(32'h3b66fc17),
	.w3(32'hbbdc7bfd),
	.w4(32'hbb82025f),
	.w5(32'h3bd5f7fb),
	.w6(32'hbbcd0612),
	.w7(32'hbb0ef4db),
	.w8(32'h3b984077),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf58ea6),
	.w1(32'hbb68da1d),
	.w2(32'hbba43aae),
	.w3(32'hbc1e18e3),
	.w4(32'hbc166a93),
	.w5(32'hbbc30e66),
	.w6(32'hbc12b584),
	.w7(32'hbbcc4a3c),
	.w8(32'hbbac621e),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa8e64),
	.w1(32'hbb5cf513),
	.w2(32'hbbde8680),
	.w3(32'h3c026160),
	.w4(32'hba6f5a95),
	.w5(32'hbb9221c3),
	.w6(32'h3c1f068c),
	.w7(32'h3b42c25e),
	.w8(32'hbc7f4744),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2687ca),
	.w1(32'hbb8c2bf2),
	.w2(32'hbb8ce445),
	.w3(32'h3b5fcaab),
	.w4(32'hbab07e4e),
	.w5(32'hbbff0449),
	.w6(32'h3b6f1cb8),
	.w7(32'h3a939869),
	.w8(32'hbbe3e121),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5272),
	.w1(32'h3aa4f670),
	.w2(32'h3b18ca8c),
	.w3(32'hbbcf641a),
	.w4(32'h3a76e6ce),
	.w5(32'h3c1e310e),
	.w6(32'hbbd6589a),
	.w7(32'hba6ab3c6),
	.w8(32'h3b592538),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02e06a),
	.w1(32'h3a88b0e7),
	.w2(32'hbc02230b),
	.w3(32'hbc4a1d24),
	.w4(32'h3bce2cd2),
	.w5(32'hbc210e55),
	.w6(32'hbbd292a1),
	.w7(32'h3b91c01a),
	.w8(32'hbbe43a94),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fef1d),
	.w1(32'hbba4c783),
	.w2(32'h3ba8e24c),
	.w3(32'hba19f3f8),
	.w4(32'hbb2c48a9),
	.w5(32'h3c4b8110),
	.w6(32'h3b2c5fa2),
	.w7(32'hbb4912eb),
	.w8(32'h3b0c5fe9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93ec70),
	.w1(32'h3b029da5),
	.w2(32'hbbcb8d83),
	.w3(32'hbb96dd57),
	.w4(32'hbaa40c61),
	.w5(32'hbc26f274),
	.w6(32'hbaeaae10),
	.w7(32'hb9b8583b),
	.w8(32'hbb140477),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e7cb),
	.w1(32'h3acc21ef),
	.w2(32'h3bdfb8d1),
	.w3(32'h3a94df94),
	.w4(32'h3ab2df9e),
	.w5(32'h3b867bb3),
	.w6(32'hbbcf9571),
	.w7(32'h39eab619),
	.w8(32'h3b9a2a45),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5565a7),
	.w1(32'hbb02e0b7),
	.w2(32'hb9abf1b4),
	.w3(32'h3a442040),
	.w4(32'hbb70910c),
	.w5(32'h3bc0b814),
	.w6(32'h395b2ec2),
	.w7(32'hbb072d34),
	.w8(32'h3b348771),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0eba6e),
	.w1(32'hbace14e3),
	.w2(32'hbaa16286),
	.w3(32'hba846ed4),
	.w4(32'h39fae168),
	.w5(32'hb9a30de3),
	.w6(32'hb90eb695),
	.w7(32'hbaf81395),
	.w8(32'h3a9315c8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0adb6c),
	.w1(32'hba66cfda),
	.w2(32'hba669cb2),
	.w3(32'h3b6d4fd1),
	.w4(32'hbbd01df6),
	.w5(32'hbb9fc90e),
	.w6(32'h3a32ca4d),
	.w7(32'h3ade4b80),
	.w8(32'hb9bc105b),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f36efc),
	.w1(32'h3b953b13),
	.w2(32'hbba630b5),
	.w3(32'hbb33430c),
	.w4(32'h3b2cf6f6),
	.w5(32'hbba9553b),
	.w6(32'hb9c036a7),
	.w7(32'h3af2d5f3),
	.w8(32'hbaf0e27a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8e35),
	.w1(32'hbc0ccc73),
	.w2(32'hbb09ce0a),
	.w3(32'hbbf840bf),
	.w4(32'hbc08ae2b),
	.w5(32'hba250d0e),
	.w6(32'hbc38b882),
	.w7(32'hbc6cda77),
	.w8(32'hba1db938),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a9cf5),
	.w1(32'h3b0e0e75),
	.w2(32'h3afa892e),
	.w3(32'hbae52e4b),
	.w4(32'h3ab7758f),
	.w5(32'h3c1f00ca),
	.w6(32'hbb1ded31),
	.w7(32'h398adf22),
	.w8(32'h3c1a8be7),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb686720),
	.w1(32'hbc21735b),
	.w2(32'hb925a9a6),
	.w3(32'hbbe7c429),
	.w4(32'hbb5b10a6),
	.w5(32'hbb473e12),
	.w6(32'hbb2cc766),
	.w7(32'hbb8315e2),
	.w8(32'hba5bdff6),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b878316),
	.w1(32'hba98e466),
	.w2(32'h3a55f909),
	.w3(32'h3b66cfeb),
	.w4(32'hbb479ec0),
	.w5(32'hbbf3cd36),
	.w6(32'h3b66af4b),
	.w7(32'hbaadc05e),
	.w8(32'hbbe8044b),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d5e3d),
	.w1(32'h3a6c18b1),
	.w2(32'hba926a8c),
	.w3(32'h3b46477c),
	.w4(32'h3b523a8b),
	.w5(32'hbb48e036),
	.w6(32'hb9945471),
	.w7(32'hb971863b),
	.w8(32'hbc0b4812),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392a3eab),
	.w1(32'h3b1257cc),
	.w2(32'h3b00a691),
	.w3(32'h3b425355),
	.w4(32'h39fd2437),
	.w5(32'hbb7180b3),
	.w6(32'hbaa0c9e6),
	.w7(32'hba448916),
	.w8(32'h3a3a3aae),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90e85e2),
	.w1(32'h3bb95eb9),
	.w2(32'h3adbfadd),
	.w3(32'hb9f84d1d),
	.w4(32'h3bbb6170),
	.w5(32'hbb0559e7),
	.w6(32'hbaed3948),
	.w7(32'h3bd97b08),
	.w8(32'hbbbecf5a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43cbc3),
	.w1(32'h3ba0994c),
	.w2(32'h3b3db5b5),
	.w3(32'h3b8a5654),
	.w4(32'hbb8902cf),
	.w5(32'h39ab7a8d),
	.w6(32'h3bafc44d),
	.w7(32'hbaa99668),
	.w8(32'h3a5c7027),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0da04),
	.w1(32'h3a3de3e0),
	.w2(32'h3b066830),
	.w3(32'hbbe0881c),
	.w4(32'h39108574),
	.w5(32'hb9253642),
	.w6(32'hbc08fcda),
	.w7(32'hbaabb685),
	.w8(32'h3a8960fa),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39b67c),
	.w1(32'hbb231af0),
	.w2(32'hbbcaca1a),
	.w3(32'h3a477002),
	.w4(32'h3baf2d4a),
	.w5(32'hbbb260bc),
	.w6(32'h3b20ca6d),
	.w7(32'h3b8cadee),
	.w8(32'hbb1409d4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90ac91),
	.w1(32'h3b46956f),
	.w2(32'h39dcf296),
	.w3(32'hbc0b02e3),
	.w4(32'h3b3dcc9e),
	.w5(32'hbc004fb5),
	.w6(32'hbbdffb8c),
	.w7(32'hba200825),
	.w8(32'hbb9a9bee),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd85d2),
	.w1(32'hb9e4f8e1),
	.w2(32'hbbb8be93),
	.w3(32'h3c63bf86),
	.w4(32'hba1b03fd),
	.w5(32'hbc3d29ea),
	.w6(32'h3bff3169),
	.w7(32'hbb0e8cd2),
	.w8(32'hbbe4cab4),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91dd6d),
	.w1(32'h3b43e9e4),
	.w2(32'hbac3bb45),
	.w3(32'hbc10c357),
	.w4(32'h3ae3c392),
	.w5(32'hbc2391d0),
	.w6(32'h3acfa2b6),
	.w7(32'hb9ac18f7),
	.w8(32'hbc14053f),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b0dc7),
	.w1(32'hbb6e2c51),
	.w2(32'hbb0ea981),
	.w3(32'hbbf1717d),
	.w4(32'hbbaec7f8),
	.w5(32'hb95e4de2),
	.w6(32'hbb3bf843),
	.w7(32'hbbe13f60),
	.w8(32'h3b8c93b2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0758fd),
	.w1(32'h3a92d98f),
	.w2(32'h3a4a0e61),
	.w3(32'hbbd9c0cc),
	.w4(32'hba680832),
	.w5(32'hbb611afa),
	.w6(32'hbba90780),
	.w7(32'h3bbe0b64),
	.w8(32'h3b3c0b58),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3965626e),
	.w1(32'hba4b1ceb),
	.w2(32'h3b2f5865),
	.w3(32'hbbba5a52),
	.w4(32'hbb229fa9),
	.w5(32'hba56b762),
	.w6(32'hbacd853d),
	.w7(32'h39ee41df),
	.w8(32'h392d1810),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf12d9),
	.w1(32'hbb204668),
	.w2(32'h3c1dc51c),
	.w3(32'hbad5181b),
	.w4(32'hbb1c1f93),
	.w5(32'h3c44dd7c),
	.w6(32'hbba8831a),
	.w7(32'hba6a200a),
	.w8(32'hbbae900d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed6a02),
	.w1(32'h3a7caf9b),
	.w2(32'hbb3390b4),
	.w3(32'h3c1c60af),
	.w4(32'hbaed6e79),
	.w5(32'hbbbfbb57),
	.w6(32'h3b9c5b4a),
	.w7(32'hbb870d7e),
	.w8(32'hbc03733d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9860fa),
	.w1(32'hba879b2f),
	.w2(32'hbbbac405),
	.w3(32'hbafdbfbd),
	.w4(32'h3aa3d843),
	.w5(32'hbb6b0921),
	.w6(32'hbba642ab),
	.w7(32'h3ab6036d),
	.w8(32'hbaaa8daa),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a63778c),
	.w1(32'h3b436816),
	.w2(32'h3a9fbdaf),
	.w3(32'hba69b084),
	.w4(32'hbb02f37a),
	.w5(32'h3b79dc97),
	.w6(32'hbaa509f3),
	.w7(32'hbac52d76),
	.w8(32'hbb2cc748),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d3764),
	.w1(32'hbb0b20e4),
	.w2(32'hbb23234d),
	.w3(32'hbc15ea8d),
	.w4(32'hba9a71b4),
	.w5(32'hbb0fd85f),
	.w6(32'hbbe35f66),
	.w7(32'h3add7b7e),
	.w8(32'hbb972e99),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83fa40),
	.w1(32'hbac21f46),
	.w2(32'h3b5d907b),
	.w3(32'hbba49de1),
	.w4(32'hbac35acd),
	.w5(32'hbb93175f),
	.w6(32'hbba729be),
	.w7(32'hbb4b8cab),
	.w8(32'hbb18218a),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac2021),
	.w1(32'hbb03a03e),
	.w2(32'hbbd9e091),
	.w3(32'h3a41611b),
	.w4(32'hbb2174e0),
	.w5(32'hbbb73879),
	.w6(32'hbb35135f),
	.w7(32'hbb81c135),
	.w8(32'hbb4009de),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f981),
	.w1(32'h3b7ab0e0),
	.w2(32'h3b4fd703),
	.w3(32'hbbd42a59),
	.w4(32'hbb433842),
	.w5(32'h3c9e2338),
	.w6(32'hbba9cf6e),
	.w7(32'h3bca97ed),
	.w8(32'h38965fd1),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cc650),
	.w1(32'hba383c26),
	.w2(32'hbb132f74),
	.w3(32'h3ae78c27),
	.w4(32'h3aefd05a),
	.w5(32'hbbd20d65),
	.w6(32'h3b2efd01),
	.w7(32'h3ae12a9f),
	.w8(32'hbbd1f929),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0698d0),
	.w1(32'hb9a69f4b),
	.w2(32'hbacdb2cd),
	.w3(32'h3b4fcfe8),
	.w4(32'h3a971b95),
	.w5(32'h38bc10a0),
	.w6(32'h386d4e8f),
	.w7(32'h3aef805f),
	.w8(32'hba884a9e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec50ff),
	.w1(32'h3aa6316e),
	.w2(32'h3bb9d0b7),
	.w3(32'hbaf2a0c7),
	.w4(32'hbb4ab26e),
	.w5(32'h3add9fd1),
	.w6(32'hba68df52),
	.w7(32'hbbdee6f8),
	.w8(32'hbb9aacc4),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87f66e),
	.w1(32'hbba569bc),
	.w2(32'hbbb4d291),
	.w3(32'h3b09dfc5),
	.w4(32'hbb379a59),
	.w5(32'hbc16b1c7),
	.w6(32'hbb12e1f5),
	.w7(32'hbaf59393),
	.w8(32'hbc19b47e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d7544),
	.w1(32'hbb64ab87),
	.w2(32'hbb968d98),
	.w3(32'hba6ba391),
	.w4(32'hbbea58b9),
	.w5(32'hbb91246d),
	.w6(32'hbaae7cc8),
	.w7(32'hbba91c61),
	.w8(32'hbba3c0ff),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cc474),
	.w1(32'h3962c70e),
	.w2(32'h3b0569fb),
	.w3(32'h3b052ca2),
	.w4(32'h39932188),
	.w5(32'hbb69c123),
	.w6(32'h3aa2f2cc),
	.w7(32'hba753932),
	.w8(32'hbb05a848),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba11f11),
	.w1(32'h3bb14ac8),
	.w2(32'h3c7066f3),
	.w3(32'hbbddffbe),
	.w4(32'hbaff996f),
	.w5(32'h3c29e882),
	.w6(32'hbba160aa),
	.w7(32'hbb0a4061),
	.w8(32'h3bc4c154),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c2835e),
	.w1(32'hbbe71df8),
	.w2(32'h39f07a95),
	.w3(32'h3b8b5aee),
	.w4(32'hbb937cfd),
	.w5(32'h3a01ab98),
	.w6(32'h3b4a5c2a),
	.w7(32'h3981a5f6),
	.w8(32'hb8e48481),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b5f2f),
	.w1(32'hbb273d2c),
	.w2(32'h3ab8b448),
	.w3(32'hbaebfe80),
	.w4(32'h39c9b399),
	.w5(32'h3beeb082),
	.w6(32'hbb816447),
	.w7(32'h3afdaffc),
	.w8(32'h3a879950),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dce8f),
	.w1(32'h3a2a2e97),
	.w2(32'h3c121b24),
	.w3(32'hbbe913f0),
	.w4(32'h3b96aa35),
	.w5(32'h3c2fe737),
	.w6(32'hbb1b292a),
	.w7(32'h3b1ef1fe),
	.w8(32'h3bdcfdbc),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3e04b5),
	.w1(32'hbb49192f),
	.w2(32'hbba15848),
	.w3(32'hbb27324b),
	.w4(32'hbb3e92d0),
	.w5(32'hbbca0b7f),
	.w6(32'hba66417a),
	.w7(32'h3ac99110),
	.w8(32'h3a934682),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7898ed),
	.w1(32'hbba1d471),
	.w2(32'hbb7ff905),
	.w3(32'hbb960a71),
	.w4(32'hba73eef6),
	.w5(32'hbbacd860),
	.w6(32'hbbb5e3f1),
	.w7(32'h3b93df99),
	.w8(32'hbb231c0b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b58f4),
	.w1(32'hbad225e9),
	.w2(32'hbb2d65f5),
	.w3(32'hbb424585),
	.w4(32'hba9eb2ba),
	.w5(32'hbba9ebff),
	.w6(32'hbbab219d),
	.w7(32'hbb877926),
	.w8(32'hbb8e5ca7),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19c141),
	.w1(32'hbb8a00ec),
	.w2(32'h3b93ae45),
	.w3(32'hbba0b49c),
	.w4(32'hbab8b06c),
	.w5(32'hbb468b5e),
	.w6(32'hbb52877b),
	.w7(32'h3b3e0e23),
	.w8(32'hbbef6d9e),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2176c4),
	.w1(32'hba8e4173),
	.w2(32'h3b5cf842),
	.w3(32'h3bfe87bf),
	.w4(32'h3967096a),
	.w5(32'h3b993306),
	.w6(32'h3b5f6e76),
	.w7(32'hb912c60e),
	.w8(32'hbbd59efc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb247f),
	.w1(32'h3aa0c4fb),
	.w2(32'h3cc7c2f1),
	.w3(32'hbb18af4a),
	.w4(32'hb59172c9),
	.w5(32'h3caa5a31),
	.w6(32'h3b3fcb36),
	.w7(32'h3b14c024),
	.w8(32'h3b2a7a03),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b514ee2),
	.w1(32'hbaeebcbf),
	.w2(32'hb88e13ea),
	.w3(32'h3c270eed),
	.w4(32'h3b22e437),
	.w5(32'hbc043238),
	.w6(32'h3c9a83bc),
	.w7(32'hba9afcb9),
	.w8(32'hbb4f8886),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6b00d),
	.w1(32'h3b1fff96),
	.w2(32'hbbcf0f5d),
	.w3(32'h3c052c0b),
	.w4(32'h3b820faf),
	.w5(32'hbb4af2db),
	.w6(32'hbb461d47),
	.w7(32'hbb29bf4f),
	.w8(32'hbbf2d941),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea652e),
	.w1(32'hbad38312),
	.w2(32'hbbc369bb),
	.w3(32'h3b877fab),
	.w4(32'h3bdb74d1),
	.w5(32'hbc3e53a9),
	.w6(32'hb8f15e31),
	.w7(32'h3b687c93),
	.w8(32'hbc30faf5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2a02),
	.w1(32'hba4155ae),
	.w2(32'hbb52e5d6),
	.w3(32'hbac2223b),
	.w4(32'hb9a696aa),
	.w5(32'hba1f972f),
	.w6(32'hbbf9d937),
	.w7(32'hbb1f6155),
	.w8(32'hbb50bda4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b094ba1),
	.w1(32'hbb6c8f2e),
	.w2(32'hbb86bdd4),
	.w3(32'h3b755d7a),
	.w4(32'hbab1332f),
	.w5(32'hbc0c714e),
	.w6(32'h3b67677a),
	.w7(32'hbbaa9984),
	.w8(32'hbc1ab518),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b15fc),
	.w1(32'hbb95b234),
	.w2(32'hbabd8ba9),
	.w3(32'hbb80fbe1),
	.w4(32'h3ac4df41),
	.w5(32'hbb537ad6),
	.w6(32'hbb8e36a9),
	.w7(32'h3a2781bc),
	.w8(32'hbb16f109),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd47e5d),
	.w1(32'h3c26171e),
	.w2(32'h3a410237),
	.w3(32'hbab16804),
	.w4(32'h3abcd4bf),
	.w5(32'hbbddbdb4),
	.w6(32'h3a8d4a4c),
	.w7(32'h3b8a5463),
	.w8(32'hba9c0fbf),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76f723),
	.w1(32'hbb36fa30),
	.w2(32'h3c12be0c),
	.w3(32'h3b8aae85),
	.w4(32'hbbe65070),
	.w5(32'h3c5ce5c0),
	.w6(32'h3a71c2b8),
	.w7(32'hbb850bba),
	.w8(32'h3c00c9bf),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49076e),
	.w1(32'h3b5c66ac),
	.w2(32'h3bc29631),
	.w3(32'hbb632804),
	.w4(32'h3a8bf14b),
	.w5(32'h39a2e24b),
	.w6(32'h39ccc6e6),
	.w7(32'h3ac6a260),
	.w8(32'hbadaa8e4),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48b21f),
	.w1(32'hbb33b2df),
	.w2(32'h3b87d6fc),
	.w3(32'h3c05fc9d),
	.w4(32'hbac15d7a),
	.w5(32'h3b80ae3e),
	.w6(32'h3b931387),
	.w7(32'h3ac4fa76),
	.w8(32'hba9176fb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc8411),
	.w1(32'hbb790835),
	.w2(32'hbb8442ea),
	.w3(32'hbada0442),
	.w4(32'hbb4c297e),
	.w5(32'hbb394852),
	.w6(32'hb9d05b9f),
	.w7(32'h37de72c2),
	.w8(32'hbbba5f17),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaaad1),
	.w1(32'hba8b4d16),
	.w2(32'hbaa92ba3),
	.w3(32'hba268f78),
	.w4(32'hba6471b2),
	.w5(32'hbbd19460),
	.w6(32'hba898d08),
	.w7(32'hba62d763),
	.w8(32'hbb62933d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b351ca7),
	.w1(32'hbbf71f07),
	.w2(32'hbc18c811),
	.w3(32'h3b471194),
	.w4(32'hbba58240),
	.w5(32'hbb3be05a),
	.w6(32'h3b189a23),
	.w7(32'h3a7bea54),
	.w8(32'h3b0da93d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbf3b1),
	.w1(32'h3abe0066),
	.w2(32'hbb2e143d),
	.w3(32'hbbccb196),
	.w4(32'h3be0bd3e),
	.w5(32'hbbb270d3),
	.w6(32'hbb43847e),
	.w7(32'h3b7e4abc),
	.w8(32'hb9e02f18),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5af46),
	.w1(32'h3b7a9538),
	.w2(32'h3b34d229),
	.w3(32'hbb60819e),
	.w4(32'h39038727),
	.w5(32'h3abf359f),
	.w6(32'hbb1dc0ea),
	.w7(32'hbacd96f5),
	.w8(32'hbabbe70f),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c7ae7),
	.w1(32'h392d0cbc),
	.w2(32'hbabfcf1a),
	.w3(32'h3a990bf8),
	.w4(32'hbaa8ed54),
	.w5(32'hbb64cb7e),
	.w6(32'hbabe3761),
	.w7(32'hba8fd986),
	.w8(32'hbc0ef89a),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6667c6),
	.w1(32'h3b357a8f),
	.w2(32'hbbd4d4e8),
	.w3(32'h39d34463),
	.w4(32'h3bda61b7),
	.w5(32'hbbc9ff6f),
	.w6(32'hbb5d410c),
	.w7(32'h3b874c63),
	.w8(32'hb8987d3a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dcb8c),
	.w1(32'hbb5df8dc),
	.w2(32'hbb1f39a7),
	.w3(32'hbabc5442),
	.w4(32'h3b049d82),
	.w5(32'hbbd89810),
	.w6(32'hb9cf3920),
	.w7(32'hba90bbf2),
	.w8(32'hbbaaf885),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8a68d),
	.w1(32'h39928b50),
	.w2(32'hbb8aede8),
	.w3(32'h38b1a110),
	.w4(32'h3ba5d33c),
	.w5(32'hbc24d4d5),
	.w6(32'hbaffa740),
	.w7(32'hbad8f6b2),
	.w8(32'hbbb40cee),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ca231),
	.w1(32'hbafce36e),
	.w2(32'h3bbebb1d),
	.w3(32'h39447517),
	.w4(32'hbb46d469),
	.w5(32'h3be3e7d9),
	.w6(32'hbb94dfd7),
	.w7(32'hba8776db),
	.w8(32'hbae33292),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85d051),
	.w1(32'hbb61ad75),
	.w2(32'h3a64331c),
	.w3(32'hbbe29bf8),
	.w4(32'hbb64760e),
	.w5(32'hbaa8fa41),
	.w6(32'hbb62be8a),
	.w7(32'hbbdd9480),
	.w8(32'hbb1b3e9f),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b8fcd),
	.w1(32'h3b1ffe4c),
	.w2(32'hbbe23569),
	.w3(32'h3b03d0d5),
	.w4(32'h3b1a9bca),
	.w5(32'hbb5a0ea8),
	.w6(32'hbb7278c5),
	.w7(32'h3aa8cb67),
	.w8(32'hbbfc75c1),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f71f0),
	.w1(32'hbbbb3da2),
	.w2(32'hba76b13a),
	.w3(32'hba96b12a),
	.w4(32'hbb14d087),
	.w5(32'hbb549c3e),
	.w6(32'h3b75433d),
	.w7(32'hbb4a0dca),
	.w8(32'hbb2f0d96),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12717b),
	.w1(32'hbb1ad0a7),
	.w2(32'h3b8592c2),
	.w3(32'hbae013ae),
	.w4(32'hb9a377d7),
	.w5(32'h3c451a97),
	.w6(32'hba77cd63),
	.w7(32'h3a8ac4e3),
	.w8(32'h38e58660),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe57928),
	.w1(32'h3b2f6c99),
	.w2(32'h3a22999b),
	.w3(32'hbbd69850),
	.w4(32'h3ba2eeaf),
	.w5(32'hbb551d73),
	.w6(32'hbb7b8a78),
	.w7(32'h3a04c692),
	.w8(32'hbb7a255a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca9faa),
	.w1(32'hb982cc8d),
	.w2(32'hbaf72b3a),
	.w3(32'h3b1dbfaa),
	.w4(32'h3a22e9e4),
	.w5(32'hba711843),
	.w6(32'hb9851fc8),
	.w7(32'hb9dab347),
	.w8(32'h3a9ef4ac),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb405359),
	.w1(32'h3b230c6a),
	.w2(32'h3bf88447),
	.w3(32'hbb5195b6),
	.w4(32'h3a688100),
	.w5(32'h3aaa71c4),
	.w6(32'hba042309),
	.w7(32'hbb9bb8b3),
	.w8(32'h3b483a21),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa2a3c),
	.w1(32'h3c00922b),
	.w2(32'h3ae8aba6),
	.w3(32'hba33ce68),
	.w4(32'h3c3bf0b7),
	.w5(32'h3a9456e4),
	.w6(32'h3b8eeebf),
	.w7(32'h3c0b2571),
	.w8(32'h3b13c3d1),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb64c59),
	.w1(32'h3c41ce42),
	.w2(32'hbc1d90f7),
	.w3(32'hbbc97bc1),
	.w4(32'h3c14ecd1),
	.w5(32'hbbacf143),
	.w6(32'h390c9d84),
	.w7(32'h3a49e097),
	.w8(32'hbbca0e9a),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabec9a),
	.w1(32'hbab9d582),
	.w2(32'hbb099f68),
	.w3(32'hbc643cfd),
	.w4(32'hbb3a3729),
	.w5(32'hbb9169c5),
	.w6(32'hbc20f1c0),
	.w7(32'hba7d0f02),
	.w8(32'hbb8a34a6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb48210),
	.w1(32'h3aae0880),
	.w2(32'hb9ab3a1b),
	.w3(32'hbbc42f53),
	.w4(32'h3ac392ee),
	.w5(32'h3b2d85a0),
	.w6(32'hbbb196ca),
	.w7(32'h3b853790),
	.w8(32'h3b6e85f0),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa50f82),
	.w1(32'hbba82d1b),
	.w2(32'hbc16e284),
	.w3(32'h3b9082fe),
	.w4(32'hbb898db3),
	.w5(32'hbbcdd192),
	.w6(32'h3b853364),
	.w7(32'h372556fa),
	.w8(32'hbba261d4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b236d),
	.w1(32'hbbdf2c5e),
	.w2(32'hbb4e07d5),
	.w3(32'hba9e8817),
	.w4(32'hbbbb5600),
	.w5(32'hb9b56953),
	.w6(32'h3a9bac3a),
	.w7(32'hbaea8036),
	.w8(32'hbb653b7e),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09c96b),
	.w1(32'hbb9e1acc),
	.w2(32'h3a9d4d8d),
	.w3(32'h3b9b1765),
	.w4(32'hbb9f8ce4),
	.w5(32'h3c29c52e),
	.w6(32'h3ababbc5),
	.w7(32'hbba5467d),
	.w8(32'h3a863668),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f18b2),
	.w1(32'h3b0764fa),
	.w2(32'hbc549269),
	.w3(32'hbc011d7e),
	.w4(32'h3b3e094c),
	.w5(32'hbc4f1454),
	.w6(32'hbb7ca46f),
	.w7(32'hbac257c8),
	.w8(32'hbc276cf3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba995588),
	.w1(32'h3b3162c5),
	.w2(32'h3c6669f1),
	.w3(32'hbba01a87),
	.w4(32'hbb0786f7),
	.w5(32'h3d10bdc5),
	.w6(32'hbbc790ca),
	.w7(32'hbb2ecdb5),
	.w8(32'h3cafc131),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0ac08),
	.w1(32'h39142d49),
	.w2(32'hbc3102f0),
	.w3(32'h3b4776bc),
	.w4(32'hbaa92bdc),
	.w5(32'hbc1afed9),
	.w6(32'h3c1f6b2a),
	.w7(32'hbb708b2f),
	.w8(32'hbbf4ddc3),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb28631),
	.w1(32'hbb9c5d24),
	.w2(32'hbc6548c3),
	.w3(32'hbba05a8a),
	.w4(32'h3b95b7bf),
	.w5(32'hbc116a60),
	.w6(32'hbc14a4b9),
	.w7(32'hbaa02e0d),
	.w8(32'hbb5dfd29),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c32e5),
	.w1(32'hbb83e2f9),
	.w2(32'hbbd5b7f3),
	.w3(32'hbb92e86c),
	.w4(32'h38a3d341),
	.w5(32'hbb57aca0),
	.w6(32'hbbc30067),
	.w7(32'hbc071bd4),
	.w8(32'hbbc935ad),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f1897),
	.w1(32'hbbd74557),
	.w2(32'hba962418),
	.w3(32'h3bbb4dde),
	.w4(32'hbbfa6270),
	.w5(32'hbb42b076),
	.w6(32'h3b398be0),
	.w7(32'hbbc03010),
	.w8(32'hbb8ff46f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27e02a),
	.w1(32'hbae02852),
	.w2(32'hbbdbff35),
	.w3(32'h39a5f857),
	.w4(32'h3b80f9f2),
	.w5(32'hbb74599e),
	.w6(32'h3b2669ad),
	.w7(32'h3b86dcdf),
	.w8(32'hbb935c17),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d040),
	.w1(32'h3adc92c9),
	.w2(32'hba8900c6),
	.w3(32'hbaddef64),
	.w4(32'hbaf510a1),
	.w5(32'hbbe3216e),
	.w6(32'hbc011d64),
	.w7(32'hbb1a0685),
	.w8(32'hbb365dd9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6621e3),
	.w1(32'h3b8a7f94),
	.w2(32'h39972bf1),
	.w3(32'hb8719d68),
	.w4(32'h3bb927ee),
	.w5(32'hbae4f9c2),
	.w6(32'hbb45bce8),
	.w7(32'h3bb8e619),
	.w8(32'h3982b107),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68db70),
	.w1(32'h3b972cf3),
	.w2(32'hba31c550),
	.w3(32'h3b46e43f),
	.w4(32'h3bb55c15),
	.w5(32'hbabea8c4),
	.w6(32'h3bb3e783),
	.w7(32'h3bb138ab),
	.w8(32'h3b9ab73b),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c4d971),
	.w1(32'hba5a1953),
	.w2(32'h3b827d66),
	.w3(32'h3874b549),
	.w4(32'h37a3c1d1),
	.w5(32'hba159ad5),
	.w6(32'h3a102646),
	.w7(32'hbab8be9f),
	.w8(32'hbb90d959),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810d10),
	.w1(32'h3a49eace),
	.w2(32'hbacae13c),
	.w3(32'hb8d8042a),
	.w4(32'hbbd51493),
	.w5(32'h3b01071d),
	.w6(32'hbab50cc2),
	.w7(32'hba4a78cf),
	.w8(32'hba9584e2),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c2bec),
	.w1(32'h3bdf1000),
	.w2(32'hbb9e5f87),
	.w3(32'hbbb63453),
	.w4(32'h3c01b853),
	.w5(32'h3a030268),
	.w6(32'hbb94e14d),
	.w7(32'h3bf7c432),
	.w8(32'hbb32877c),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb777e3),
	.w1(32'hbb1e9935),
	.w2(32'hbaa12790),
	.w3(32'hbbb5444b),
	.w4(32'hbaf4c94b),
	.w5(32'hbac0b6d9),
	.w6(32'hbbe568fd),
	.w7(32'hbb3b5c60),
	.w8(32'hba86c487),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20c7a1),
	.w1(32'hba9e1c79),
	.w2(32'hba2ff481),
	.w3(32'hba32b3a8),
	.w4(32'hbae866fb),
	.w5(32'hba726a90),
	.w6(32'hbb052964),
	.w7(32'hbb37e0dd),
	.w8(32'hbb88aeaf),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f842c9),
	.w1(32'hbb131269),
	.w2(32'hbb3f14f0),
	.w3(32'hbaea3da2),
	.w4(32'hbb5341a5),
	.w5(32'hbad65516),
	.w6(32'hbb75cfa4),
	.w7(32'hba4074a7),
	.w8(32'h3a8685cc),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a1d3e),
	.w1(32'h3ab1e29c),
	.w2(32'h3aee50ec),
	.w3(32'hbae9b42e),
	.w4(32'h3b01798b),
	.w5(32'h3b1d0894),
	.w6(32'h38ba3548),
	.w7(32'h3b11f6ad),
	.w8(32'h3b854aac),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e5295),
	.w1(32'h3a1e6d61),
	.w2(32'hb9137640),
	.w3(32'h3a7ba0a9),
	.w4(32'hbacef7d5),
	.w5(32'hba98749f),
	.w6(32'h3afe0513),
	.w7(32'hbac65989),
	.w8(32'hbaa5da70),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3e9ab),
	.w1(32'h3abcca24),
	.w2(32'h3a877188),
	.w3(32'hba8b3586),
	.w4(32'h39803d04),
	.w5(32'hba86cb45),
	.w6(32'hba29bbe4),
	.w7(32'h3a0af260),
	.w8(32'hb965473e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d248cc),
	.w1(32'hb95deb7b),
	.w2(32'h39dc3e8f),
	.w3(32'hbb0d23a2),
	.w4(32'hba4c3ad5),
	.w5(32'h3a202ae3),
	.w6(32'hb92330e7),
	.w7(32'hba76d0f8),
	.w8(32'h398ba8c1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d4f89),
	.w1(32'h39bb2f1c),
	.w2(32'hb930a402),
	.w3(32'hba8991dc),
	.w4(32'h3a272b2c),
	.w5(32'hba008bf6),
	.w6(32'hb96952eb),
	.w7(32'h390eaf86),
	.w8(32'hb80bebec),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b19af),
	.w1(32'hbad8982a),
	.w2(32'hbad7038b),
	.w3(32'h3ac65bf1),
	.w4(32'hbb860c92),
	.w5(32'hba30488b),
	.w6(32'hb9c34c9c),
	.w7(32'hb90239de),
	.w8(32'hbac9bae0),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5932b3),
	.w1(32'hba47b2fd),
	.w2(32'hb969b802),
	.w3(32'hbb5adc27),
	.w4(32'hb91926aa),
	.w5(32'hb9c2d4de),
	.w6(32'hbb136bcd),
	.w7(32'h39a32915),
	.w8(32'h3990f62c),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abef51a),
	.w1(32'h399ab9da),
	.w2(32'hba051cdb),
	.w3(32'h3a8c4189),
	.w4(32'hb947af1c),
	.w5(32'hbae87576),
	.w6(32'h38e63887),
	.w7(32'hba8d32a0),
	.w8(32'hbab8a62a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178b53),
	.w1(32'h3b85b0bb),
	.w2(32'h3b27c73b),
	.w3(32'h3a9fd2b2),
	.w4(32'h3bb6562d),
	.w5(32'h3b918c7d),
	.w6(32'hb901826e),
	.w7(32'h3b985029),
	.w8(32'h3b762509),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f70c6),
	.w1(32'hba0ef4c8),
	.w2(32'h3a4718fc),
	.w3(32'h3bbef249),
	.w4(32'hba0255c4),
	.w5(32'h3aa51f5f),
	.w6(32'h3b8da3e5),
	.w7(32'hba44efe0),
	.w8(32'h39cd1d36),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfcd66),
	.w1(32'hb9255d72),
	.w2(32'hb99cc3a1),
	.w3(32'h3a0343b1),
	.w4(32'h3986824e),
	.w5(32'h395e94ba),
	.w6(32'h3a20f29f),
	.w7(32'h3a21cbcb),
	.w8(32'h3a4a1a58),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2421e),
	.w1(32'h3a8b0146),
	.w2(32'h3adebb78),
	.w3(32'h3a1c7d64),
	.w4(32'h3aa0a4e1),
	.w5(32'h3b7fa433),
	.w6(32'h3a5cd321),
	.w7(32'h3a433e67),
	.w8(32'h39904c57),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39abd46d),
	.w1(32'hbae1f1d1),
	.w2(32'hbb18a517),
	.w3(32'h3a69f743),
	.w4(32'hbb169405),
	.w5(32'hbb23a545),
	.w6(32'hba8a052c),
	.w7(32'hbb0f0348),
	.w8(32'hbb15bca7),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bf494),
	.w1(32'hbb096b3c),
	.w2(32'hbb79a9cd),
	.w3(32'hba8f63d2),
	.w4(32'hbb92438c),
	.w5(32'hbba07598),
	.w6(32'hba4e7edd),
	.w7(32'hbb85c52e),
	.w8(32'hbb9a7ee2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f4d33),
	.w1(32'hba01d25d),
	.w2(32'hbadc7d84),
	.w3(32'hba9a4a3e),
	.w4(32'hbb4dbc7b),
	.w5(32'hba8534fc),
	.w6(32'hba604df2),
	.w7(32'hbb27e15e),
	.w8(32'hbb3b27e0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982ccfc),
	.w1(32'hbb2b9428),
	.w2(32'hbb856db2),
	.w3(32'hbace7ef1),
	.w4(32'hbbaedca2),
	.w5(32'hbb5ffdd8),
	.w6(32'hbb443473),
	.w7(32'hbb8650c9),
	.w8(32'hbb991d9b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cf0a5),
	.w1(32'hbb0219b2),
	.w2(32'hba3b4679),
	.w3(32'hbb6f3358),
	.w4(32'hb84c1bf4),
	.w5(32'h3a9cc590),
	.w6(32'hbb713eb5),
	.w7(32'h39774537),
	.w8(32'h3a6883d0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bd5729),
	.w1(32'h39c5da4a),
	.w2(32'hbac16729),
	.w3(32'h3a60ee0e),
	.w4(32'h39ffdaba),
	.w5(32'hba4cfd43),
	.w6(32'hbac5fb86),
	.w7(32'hb9f2c986),
	.w8(32'hb890a22a),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41da58),
	.w1(32'hba80af6b),
	.w2(32'hb9b3d872),
	.w3(32'h3a9807e3),
	.w4(32'hba8ad5b1),
	.w5(32'hbaa4449f),
	.w6(32'hba5b323e),
	.w7(32'hba1e1b9b),
	.w8(32'hbb05af29),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74d7ee3),
	.w1(32'hbaadb44e),
	.w2(32'hbaa9250a),
	.w3(32'hbaaf0b3c),
	.w4(32'hba1527f1),
	.w5(32'h37e465eb),
	.w6(32'hb9acb34f),
	.w7(32'h39a2a97e),
	.w8(32'hba326bc6),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b02bb),
	.w1(32'hbaaae1b7),
	.w2(32'hbb0fcad0),
	.w3(32'hb9b7b06c),
	.w4(32'h38c0c5dd),
	.w5(32'hbaa9ed39),
	.w6(32'hb90a7112),
	.w7(32'h3abfd693),
	.w8(32'h3abd60ed),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb635a13),
	.w1(32'hbb0fac06),
	.w2(32'hbadcb1cb),
	.w3(32'hbb128347),
	.w4(32'hbad6f3b1),
	.w5(32'hba9334b9),
	.w6(32'h39a77dc8),
	.w7(32'hbaaeac75),
	.w8(32'hba763013),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38431cb5),
	.w1(32'hba98d922),
	.w2(32'h3975537e),
	.w3(32'h3a5b4897),
	.w4(32'h3a436f98),
	.w5(32'h3b5fbe06),
	.w6(32'h39938229),
	.w7(32'hba1c7545),
	.w8(32'hba2e3424),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a41243b),
	.w1(32'hba28afc7),
	.w2(32'hba86a904),
	.w3(32'h3b20ec28),
	.w4(32'hbb297973),
	.w5(32'hbad4a2ff),
	.w6(32'hb937a39d),
	.w7(32'hbb1f07c7),
	.w8(32'hba8dd150),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7eb0a),
	.w1(32'hbaf95352),
	.w2(32'hbb223a13),
	.w3(32'hbb0391d0),
	.w4(32'hbb95e9ba),
	.w5(32'hbb737022),
	.w6(32'hb9ef86c5),
	.w7(32'hbb9f9c93),
	.w8(32'hbb90c829),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0bc0d),
	.w1(32'hba902ed3),
	.w2(32'h39c43a24),
	.w3(32'hbb1d7e80),
	.w4(32'hba8a50ef),
	.w5(32'h3a84f9e8),
	.w6(32'hbaf37b3f),
	.w7(32'hbab7bc10),
	.w8(32'h3a71a0f8),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d9e12),
	.w1(32'h3a120b9a),
	.w2(32'hb99bd971),
	.w3(32'h3b13df4a),
	.w4(32'h3a71d8ba),
	.w5(32'h3a9f7e2c),
	.w6(32'h3a30d829),
	.w7(32'hb81fc0a9),
	.w8(32'hba7c5df5),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39529ff0),
	.w1(32'h38f41e9b),
	.w2(32'hb9fce4ed),
	.w3(32'h396fe851),
	.w4(32'h3a66fedd),
	.w5(32'hba4c8035),
	.w6(32'hb970064b),
	.w7(32'h3a7488f1),
	.w8(32'hba501f70),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93288f8),
	.w1(32'hba0d17d2),
	.w2(32'hb9959d15),
	.w3(32'hbab29309),
	.w4(32'hbaff87da),
	.w5(32'hb90dd7d1),
	.w6(32'h38d423f0),
	.w7(32'hbb0c9cf7),
	.w8(32'hbb1aef09),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8521d50),
	.w1(32'hbab247a2),
	.w2(32'hbacd1371),
	.w3(32'hb8596be0),
	.w4(32'hbb20cda6),
	.w5(32'hbb233d55),
	.w6(32'hba9fff6b),
	.w7(32'hbb1db4da),
	.w8(32'hbaf4e1eb),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb951dfba),
	.w1(32'h3b698b4d),
	.w2(32'hba827712),
	.w3(32'hbab199bc),
	.w4(32'h3a12af9a),
	.w5(32'hb9ba5cfa),
	.w6(32'hb9e91d27),
	.w7(32'hba5ddd2a),
	.w8(32'hbb27bd0c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5da0c8),
	.w1(32'hbb21c454),
	.w2(32'hbb35cf0a),
	.w3(32'hba8d7825),
	.w4(32'hbb6a92e1),
	.w5(32'hbb33ec84),
	.w6(32'hbb0316d1),
	.w7(32'hbb6169b9),
	.w8(32'hbb2671a8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23ac9a),
	.w1(32'hbaa8255f),
	.w2(32'hbabb2df7),
	.w3(32'hbb0bbb28),
	.w4(32'hba280cdc),
	.w5(32'hba207415),
	.w6(32'hbaf2f53f),
	.w7(32'hbad86225),
	.w8(32'hbb4568cc),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba058ebd),
	.w1(32'hb7d2dea7),
	.w2(32'hb8d51d95),
	.w3(32'hba2b31e6),
	.w4(32'h3a0976fc),
	.w5(32'h39a0f512),
	.w6(32'hbb05c338),
	.w7(32'hb75b7185),
	.w8(32'hba335228),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15178f),
	.w1(32'hb9ceea80),
	.w2(32'hb9e900c7),
	.w3(32'h3ac6cc68),
	.w4(32'h389ebf45),
	.w5(32'hb96c0bda),
	.w6(32'h3a7e28fa),
	.w7(32'hba5288e5),
	.w8(32'hbac8decd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00710e),
	.w1(32'hbb4ece08),
	.w2(32'hbb5bb300),
	.w3(32'hba2679a1),
	.w4(32'hbb2caed3),
	.w5(32'hbb1496ff),
	.w6(32'hbac1a5ff),
	.w7(32'hbaca873c),
	.w8(32'hbae4bb3d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0b27a),
	.w1(32'hba738415),
	.w2(32'hba8c1d43),
	.w3(32'hbb0e893e),
	.w4(32'h37b4a5b4),
	.w5(32'h3ae4b188),
	.w6(32'hbb0bc653),
	.w7(32'h3a278ce3),
	.w8(32'h3a608b6e),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f0d8),
	.w1(32'hbad151b2),
	.w2(32'hba5a2ae4),
	.w3(32'h385886eb),
	.w4(32'hbad8b854),
	.w5(32'hba363888),
	.w6(32'h39229907),
	.w7(32'hba162e17),
	.w8(32'hbaa23c96),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c5cf20),
	.w1(32'hbab1a490),
	.w2(32'hbaccbf17),
	.w3(32'hbaf06750),
	.w4(32'h39b3ef14),
	.w5(32'hba0029f8),
	.w6(32'hbab860e4),
	.w7(32'h393dbf82),
	.w8(32'hb98775c3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa64f2f),
	.w1(32'h3a265136),
	.w2(32'hba2090bb),
	.w3(32'h3a8d40b1),
	.w4(32'hba1850d4),
	.w5(32'hba81ef63),
	.w6(32'h3a2b44e7),
	.w7(32'hbab55e70),
	.w8(32'hbaae55ce),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cfd8df),
	.w1(32'h39ea1a2e),
	.w2(32'hbade80bb),
	.w3(32'h396efa78),
	.w4(32'h3955efb9),
	.w5(32'hba99ad61),
	.w6(32'h3a16c2e0),
	.w7(32'hb907e32c),
	.w8(32'hba978e30),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa00a97),
	.w1(32'hb9ab4d11),
	.w2(32'hbad011c9),
	.w3(32'h39b3d8a4),
	.w4(32'hb810fd27),
	.w5(32'hbb20fcf6),
	.w6(32'h39f3c23d),
	.w7(32'hbb09acd3),
	.w8(32'hba707266),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9952dad),
	.w1(32'h3a9ff64f),
	.w2(32'hba92ba47),
	.w3(32'h394c5acb),
	.w4(32'h3ac99660),
	.w5(32'h39525050),
	.w6(32'h3a2faccb),
	.w7(32'h390f0948),
	.w8(32'hb8aa4c76),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae969b3),
	.w1(32'h39ae0c63),
	.w2(32'h39f6e3ca),
	.w3(32'hba270548),
	.w4(32'h39d672be),
	.w5(32'h3a282fc0),
	.w6(32'hba1cf184),
	.w7(32'h36147024),
	.w8(32'h39557734),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392acfa3),
	.w1(32'h37dd0c23),
	.w2(32'h3ae2514c),
	.w3(32'h39d36f86),
	.w4(32'h3b10f5b7),
	.w5(32'h3afec9d8),
	.w6(32'h3a8a4a0f),
	.w7(32'h3ac45219),
	.w8(32'h3b0fe666),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d3578),
	.w1(32'hb9fabf07),
	.w2(32'hba4b8549),
	.w3(32'h3b0044d0),
	.w4(32'hb9e4791f),
	.w5(32'hba577edd),
	.w6(32'h3b219d80),
	.w7(32'hb930ae19),
	.w8(32'h3ad51320),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391363e2),
	.w1(32'h3a0e7d02),
	.w2(32'h3a577d15),
	.w3(32'h3b018af6),
	.w4(32'hbae23336),
	.w5(32'hbac9b6c4),
	.w6(32'h3b6036a4),
	.w7(32'hb91c07ea),
	.w8(32'hbace72fd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83f338),
	.w1(32'h38f50ce7),
	.w2(32'hbb0aad52),
	.w3(32'hbaddd1aa),
	.w4(32'hbabef8a6),
	.w5(32'hbb220599),
	.w6(32'hb9c13166),
	.w7(32'hbb29de51),
	.w8(32'hbb7b5b55),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb520c0e),
	.w1(32'hb9f9eda9),
	.w2(32'hb8a542e2),
	.w3(32'hbb5861c4),
	.w4(32'h399a273c),
	.w5(32'h39ea8cff),
	.w6(32'hbba32611),
	.w7(32'h39fee109),
	.w8(32'h389fcf1f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97b0549),
	.w1(32'h39bdc101),
	.w2(32'h39c28b4e),
	.w3(32'h39b5311d),
	.w4(32'h38660677),
	.w5(32'h3aad5582),
	.w6(32'hba9a167f),
	.w7(32'hba3dc1f3),
	.w8(32'hb9c6f7e9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dce02c),
	.w1(32'hbac9733a),
	.w2(32'hbafb54d1),
	.w3(32'h3a6fb247),
	.w4(32'hbb2b833c),
	.w5(32'hbacb5cd1),
	.w6(32'hbab86744),
	.w7(32'hbb6f006c),
	.w8(32'hbba292d4),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ebe2),
	.w1(32'h3a8657bd),
	.w2(32'h39869878),
	.w3(32'hbb202e9d),
	.w4(32'h3a9eaf6c),
	.w5(32'h3a5efdb5),
	.w6(32'hbb6c4993),
	.w7(32'hb9ce4ff5),
	.w8(32'hb9ef2ed2),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4479c),
	.w1(32'hbb17865c),
	.w2(32'hbae78599),
	.w3(32'hb91f641b),
	.w4(32'hbae16b7d),
	.w5(32'h3a283c05),
	.w6(32'hb9287dad),
	.w7(32'h39fed94e),
	.w8(32'h3ab49840),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf78a84),
	.w1(32'h3925f651),
	.w2(32'h38eacfa0),
	.w3(32'hb78cb830),
	.w4(32'hba277209),
	.w5(32'hb9f5cbb3),
	.w6(32'h3ae49786),
	.w7(32'hbae8e786),
	.w8(32'hbac6d236),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39acb091),
	.w1(32'hba95210e),
	.w2(32'hbb01dcde),
	.w3(32'hb9453676),
	.w4(32'hbb1d475c),
	.w5(32'hbb9205b5),
	.w6(32'h3601fe67),
	.w7(32'hbb57e17b),
	.w8(32'hbbd8a6e6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e4fec5),
	.w1(32'hba286319),
	.w2(32'hba9ce979),
	.w3(32'hbb3d62ca),
	.w4(32'hba961c1d),
	.w5(32'hbb092d7d),
	.w6(32'hbb70dd2c),
	.w7(32'hbadbc4cc),
	.w8(32'hbb08dbfa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule