module layer_8_featuremap_122(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b8477f),
	.w1(32'h3b2fa091),
	.w2(32'h3bf9c4c4),
	.w3(32'hb9ba719d),
	.w4(32'h3c8d1e50),
	.w5(32'hb97b3d50),
	.w6(32'hbb93da7a),
	.w7(32'h3c3b4da1),
	.w8(32'hbc177c05),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099411),
	.w1(32'h3c28b5a5),
	.w2(32'hba45d89c),
	.w3(32'h39376e26),
	.w4(32'hbc8be7c2),
	.w5(32'h3bc53d5c),
	.w6(32'h3c147463),
	.w7(32'hbc401b79),
	.w8(32'h3b57864f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14a524),
	.w1(32'hbb6cdd9e),
	.w2(32'hbc84c5cb),
	.w3(32'hbb8ca24f),
	.w4(32'hbc11f4be),
	.w5(32'h3c566cdb),
	.w6(32'h3bb17264),
	.w7(32'hbc016b54),
	.w8(32'h3bae26cd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b114070),
	.w1(32'h3c3464a6),
	.w2(32'h3c348789),
	.w3(32'hbae19c2c),
	.w4(32'hbc53701f),
	.w5(32'h3cee9fc3),
	.w6(32'hbcfe3ac8),
	.w7(32'h3bfd9f40),
	.w8(32'hbcecbd76),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf58c8d),
	.w1(32'h3cacfbfa),
	.w2(32'hbbbd2c67),
	.w3(32'hbc32407d),
	.w4(32'h3b3c85a8),
	.w5(32'hbbe3a0d3),
	.w6(32'h3bb081f8),
	.w7(32'h3bc389e9),
	.w8(32'hbca985b1),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9722196),
	.w1(32'hbb3ac5df),
	.w2(32'hbc20dcf2),
	.w3(32'hb8b5ee80),
	.w4(32'hbc93e63a),
	.w5(32'h3aa3c662),
	.w6(32'h3b524f1c),
	.w7(32'hbc62ac70),
	.w8(32'hbbd3b761),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b510891),
	.w1(32'h3ba3800e),
	.w2(32'hbacb00ba),
	.w3(32'h3b46205e),
	.w4(32'hbbadafd8),
	.w5(32'hb9ce7245),
	.w6(32'h3bba718f),
	.w7(32'h3c75afce),
	.w8(32'hbc4532e0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc017),
	.w1(32'h39ded0fc),
	.w2(32'h3c00a703),
	.w3(32'h3c327a29),
	.w4(32'h3a0b7893),
	.w5(32'hbb8b5ca0),
	.w6(32'h3c14a283),
	.w7(32'h3c2b6d30),
	.w8(32'hbc59543c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01b2d9),
	.w1(32'hbc744f23),
	.w2(32'h3b80ad9b),
	.w3(32'h3c149da9),
	.w4(32'h3b9de940),
	.w5(32'hbc8b501a),
	.w6(32'hbadb40b9),
	.w7(32'h3b2b0a02),
	.w8(32'hbc36cae7),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c962f5),
	.w1(32'h3b03e01b),
	.w2(32'hbc80dbd8),
	.w3(32'hbbabcd3e),
	.w4(32'hba9f15a3),
	.w5(32'hbc089f14),
	.w6(32'h3ba48a8e),
	.w7(32'hbd04c82b),
	.w8(32'h3d6897bf),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3e0b4f),
	.w1(32'hbd1ec0f3),
	.w2(32'hbcad18b9),
	.w3(32'h3c33499d),
	.w4(32'h3c169ab1),
	.w5(32'hbc560481),
	.w6(32'hbca61b93),
	.w7(32'hbc2272c3),
	.w8(32'hbcb0ceb3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c36a2dc),
	.w1(32'hbad525ee),
	.w2(32'h3c708dba),
	.w3(32'hbbdbaa8f),
	.w4(32'h3bad8fd9),
	.w5(32'hbc331adf),
	.w6(32'hbbf0f43d),
	.w7(32'h3b0db15b),
	.w8(32'hbc978366),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61c560),
	.w1(32'hba0642e0),
	.w2(32'hbc23423b),
	.w3(32'h3bcc82ed),
	.w4(32'hbb41cdd8),
	.w5(32'hbb53f3a9),
	.w6(32'h3cb7e06b),
	.w7(32'hbc1dfb4f),
	.w8(32'hbadb19c8),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b184096),
	.w1(32'h3b91f7ee),
	.w2(32'hbba7b27f),
	.w3(32'h3b69fe25),
	.w4(32'hbb89054e),
	.w5(32'hbc329288),
	.w6(32'h3c93b316),
	.w7(32'hbbb2f3a5),
	.w8(32'hb9d485c0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f6b94),
	.w1(32'h3c369778),
	.w2(32'hbb67a62b),
	.w3(32'h3b85fbae),
	.w4(32'hba97faa6),
	.w5(32'hbbb241ba),
	.w6(32'h3c497108),
	.w7(32'hbadead23),
	.w8(32'hbbbfeee0),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b6627),
	.w1(32'hbb612c93),
	.w2(32'hbb8a2d97),
	.w3(32'hbadf043f),
	.w4(32'hbc7cc201),
	.w5(32'hbc3f4e6e),
	.w6(32'hbb993609),
	.w7(32'hbb9d51d3),
	.w8(32'hbc6b9f65),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0721bb),
	.w1(32'hbcb5877c),
	.w2(32'hbbe7fd63),
	.w3(32'hb9b9f77c),
	.w4(32'hbc0c90a0),
	.w5(32'h3b2bf536),
	.w6(32'h3bbd3ed0),
	.w7(32'hbb6f07c8),
	.w8(32'h3b4db02b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf70d93),
	.w1(32'h3c8a75f4),
	.w2(32'hbbe0b2d5),
	.w3(32'h3c4c1f48),
	.w4(32'hbc69c14a),
	.w5(32'hbb52e589),
	.w6(32'h3c183467),
	.w7(32'hbba4d2b8),
	.w8(32'hbc50fd86),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7648d5),
	.w1(32'h3cd29e99),
	.w2(32'h3ca62333),
	.w3(32'h3c04233a),
	.w4(32'h3d046bc8),
	.w5(32'h3ceff25a),
	.w6(32'hbb236e1f),
	.w7(32'h3c209b19),
	.w8(32'h3c98096b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ddfbb),
	.w1(32'h3cf6185a),
	.w2(32'h3cc15804),
	.w3(32'h3c7514f6),
	.w4(32'h3bab796e),
	.w5(32'hbaba879b),
	.w6(32'h3d7e4cb8),
	.w7(32'hbc1ecb1d),
	.w8(32'hba147aac),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ca2e4),
	.w1(32'hbca26141),
	.w2(32'h3b2e4fdd),
	.w3(32'h3bc74976),
	.w4(32'h3a8fe746),
	.w5(32'h3ad075de),
	.w6(32'h3c493aae),
	.w7(32'h3c10106b),
	.w8(32'h3cdb8b7d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e09a7),
	.w1(32'hbb9e513a),
	.w2(32'hbd07db48),
	.w3(32'h3b1d4218),
	.w4(32'hbccedfcf),
	.w5(32'h3a70c1b8),
	.w6(32'hbd53e07e),
	.w7(32'hbcad17ff),
	.w8(32'hbc531f23),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241b30),
	.w1(32'h3c6456db),
	.w2(32'hbccc2953),
	.w3(32'h3c070702),
	.w4(32'hbc427ac5),
	.w5(32'hbcc5c4bc),
	.w6(32'hbc2ca3c1),
	.w7(32'hbc5a399f),
	.w8(32'h39558e0a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c6f3b),
	.w1(32'hbb48e5ef),
	.w2(32'hbb91e4c2),
	.w3(32'h388ac28c),
	.w4(32'hbbfdfe94),
	.w5(32'hbbd2f1fe),
	.w6(32'hbb3bcc6c),
	.w7(32'hbbf81dc7),
	.w8(32'hbb5cdef1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bb509),
	.w1(32'h3baeaee5),
	.w2(32'h3a068625),
	.w3(32'h3b6829b4),
	.w4(32'h3b86eecb),
	.w5(32'hbc9bed72),
	.w6(32'h3c0530e8),
	.w7(32'h3bccadf2),
	.w8(32'hbc80ce2d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85c6ae),
	.w1(32'hbc45e31e),
	.w2(32'h3c415bd7),
	.w3(32'hbb7adb8d),
	.w4(32'h3c31c075),
	.w5(32'hbb1030c4),
	.w6(32'hbc4699cd),
	.w7(32'hb852eb18),
	.w8(32'h3bcd785f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929a16),
	.w1(32'hbc0d0346),
	.w2(32'hbc0e4717),
	.w3(32'h3bb66d6f),
	.w4(32'hbbda2f38),
	.w5(32'hba3e7810),
	.w6(32'hbcedbab1),
	.w7(32'hbc2a01e9),
	.w8(32'hbc72f25a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e5698),
	.w1(32'h3d33f13a),
	.w2(32'h3c7a8b6a),
	.w3(32'h3db076b9),
	.w4(32'h3d6ac16c),
	.w5(32'h3c86b491),
	.w6(32'h3cf5065d),
	.w7(32'h3d69da4d),
	.w8(32'h3a3da0cb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e31e0),
	.w1(32'hbba41985),
	.w2(32'hbac15358),
	.w3(32'h3bcb299b),
	.w4(32'hbab2dadc),
	.w5(32'h3a1e69b3),
	.w6(32'hbca885fb),
	.w7(32'h3c810cea),
	.w8(32'hbb14b05c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda7c86),
	.w1(32'hbc86b8e6),
	.w2(32'h3b4290b3),
	.w3(32'hbc099e42),
	.w4(32'hbc0bc80b),
	.w5(32'hbc7f9343),
	.w6(32'hbbc4bbea),
	.w7(32'hbba73e22),
	.w8(32'h3b2f18a1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784c69),
	.w1(32'hbbedbf3e),
	.w2(32'hba04561b),
	.w3(32'h3abfbfec),
	.w4(32'h3b4a303c),
	.w5(32'h3ba281f3),
	.w6(32'hbc8e94ee),
	.w7(32'h3b0894eb),
	.w8(32'h3ba32be9),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0bc08),
	.w1(32'hbbc2f29f),
	.w2(32'hbc5ff768),
	.w3(32'h39f4ba5d),
	.w4(32'hbc8593f6),
	.w5(32'hbcae8cab),
	.w6(32'h3b2ece1b),
	.w7(32'hbc831386),
	.w8(32'hbd035019),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0acfb),
	.w1(32'h3c65a1c3),
	.w2(32'hbc600549),
	.w3(32'h3a75b90b),
	.w4(32'hbc47dca7),
	.w5(32'h3c998fc8),
	.w6(32'h3d243166),
	.w7(32'hbcc80089),
	.w8(32'h3d21b931),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32e0f2),
	.w1(32'h38747bc8),
	.w2(32'hb9989a6c),
	.w3(32'h3c3968bb),
	.w4(32'hbb2b2641),
	.w5(32'hbc42c64f),
	.w6(32'h3c2b1392),
	.w7(32'hbadbc87b),
	.w8(32'hbc62404b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f9d8e),
	.w1(32'hbb7e7663),
	.w2(32'h3b815b7d),
	.w3(32'h3c29155a),
	.w4(32'h3c0981aa),
	.w5(32'h3c5f0632),
	.w6(32'hbc45c958),
	.w7(32'h3b68cf8c),
	.w8(32'h3c85e529),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c873e7e),
	.w1(32'hbbc49cd7),
	.w2(32'hba7146e6),
	.w3(32'h3c171705),
	.w4(32'hbc7c6c76),
	.w5(32'hb81bbc79),
	.w6(32'hbc41d6ca),
	.w7(32'hbc5268ce),
	.w8(32'h3d7840ca),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c79421b),
	.w1(32'h3caa8c26),
	.w2(32'h3c545c9c),
	.w3(32'h3c467aca),
	.w4(32'hbc7aab3f),
	.w5(32'hbc828534),
	.w6(32'h3d00e360),
	.w7(32'hbb9b06f0),
	.w8(32'hbc868fa8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17899b),
	.w1(32'hbb788e29),
	.w2(32'hbb263614),
	.w3(32'h399eda43),
	.w4(32'hbb3185de),
	.w5(32'hbc948a96),
	.w6(32'h3b03569b),
	.w7(32'h3b9e4d03),
	.w8(32'hbb44a751),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc003c62),
	.w1(32'hbc2a8731),
	.w2(32'h3b19b525),
	.w3(32'hbc8e18f6),
	.w4(32'hbb145591),
	.w5(32'hbbdfad69),
	.w6(32'h3b926275),
	.w7(32'hbc47c381),
	.w8(32'hbc8ebd73),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f2d4),
	.w1(32'h3be2fd8d),
	.w2(32'h3ae4fafc),
	.w3(32'hbc018431),
	.w4(32'hbc035a71),
	.w5(32'h3a3a6fe5),
	.w6(32'h3c02c489),
	.w7(32'h3b899e97),
	.w8(32'hba3d30af),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0712ed),
	.w1(32'h3cae5698),
	.w2(32'h3c087657),
	.w3(32'h3d2a5223),
	.w4(32'h3c5d5b89),
	.w5(32'h3bddfc84),
	.w6(32'h3d187fb5),
	.w7(32'h3c0fb504),
	.w8(32'hbafb5f74),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6fc00a),
	.w1(32'hbbda88ca),
	.w2(32'h3c409e73),
	.w3(32'h3d2aac33),
	.w4(32'h3c8a6139),
	.w5(32'h3c44cca8),
	.w6(32'h3d47229b),
	.w7(32'h3c905238),
	.w8(32'h3ca0fc78),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f09b4),
	.w1(32'hbc55117e),
	.w2(32'hbc04124d),
	.w3(32'hbc85fd1b),
	.w4(32'h3a27f14a),
	.w5(32'h3b74df9b),
	.w6(32'hbc672500),
	.w7(32'hbb5097da),
	.w8(32'hba8247bf),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc929f3d),
	.w1(32'h3bb3349b),
	.w2(32'hbbbc5be4),
	.w3(32'h3c106278),
	.w4(32'h3ba67895),
	.w5(32'h3b4eb80c),
	.w6(32'h3c79da7a),
	.w7(32'hbbe1f5c0),
	.w8(32'h3b96182b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4c0049),
	.w1(32'h3c323542),
	.w2(32'hbb03192d),
	.w3(32'h3be64949),
	.w4(32'h3b998f1a),
	.w5(32'h3c1c586b),
	.w6(32'h3cc5de43),
	.w7(32'h3b826cd0),
	.w8(32'h3c4f8e47),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00f23e),
	.w1(32'hbc612faa),
	.w2(32'hba2a447b),
	.w3(32'hbc1d1a8d),
	.w4(32'hbafb8bb4),
	.w5(32'h3bf033a8),
	.w6(32'hbc9a4714),
	.w7(32'hbbc932d5),
	.w8(32'hbcc5b3a8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc199ff0),
	.w1(32'h3bc75c4f),
	.w2(32'hbaca68a4),
	.w3(32'hbb844fdf),
	.w4(32'h3c1f6b65),
	.w5(32'h3cc28827),
	.w6(32'h3b8487f0),
	.w7(32'h3c6011db),
	.w8(32'h3c382578),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81753a),
	.w1(32'hbc5eca41),
	.w2(32'h3b6dc106),
	.w3(32'h3a5af92f),
	.w4(32'hbc2a0aa1),
	.w5(32'hbc84d3bd),
	.w6(32'hbcc98105),
	.w7(32'hbb194700),
	.w8(32'hbb52dd9e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2a2b0),
	.w1(32'h3ca09e62),
	.w2(32'hbc86ba9d),
	.w3(32'hb993cfa6),
	.w4(32'hbca54f73),
	.w5(32'hbc787254),
	.w6(32'h3cc2d594),
	.w7(32'hbc07a200),
	.w8(32'hbc69fd76),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaaecaa),
	.w1(32'h3d215753),
	.w2(32'hbd13139f),
	.w3(32'hbb70a01c),
	.w4(32'hbd2d4c46),
	.w5(32'hbd3713b5),
	.w6(32'h392e090f),
	.w7(32'hbd09fc02),
	.w8(32'hbd07e028),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbebacf),
	.w1(32'h3cee19fb),
	.w2(32'hbc1bfd29),
	.w3(32'hbc5d4abc),
	.w4(32'hbcde12af),
	.w5(32'hbce274ee),
	.w6(32'h3d555778),
	.w7(32'hbc773946),
	.w8(32'h3b97d4de),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1df0dd),
	.w1(32'h3c183f6a),
	.w2(32'h3d242e4d),
	.w3(32'h3cab6312),
	.w4(32'h3d3727f5),
	.w5(32'h3d4b22f4),
	.w6(32'h3d23237b),
	.w7(32'h3d1a00c9),
	.w8(32'h3bded3ff),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc6b10),
	.w1(32'hbd8968d8),
	.w2(32'h39885b05),
	.w3(32'hbba8165d),
	.w4(32'h3c7184aa),
	.w5(32'h3b86c9da),
	.w6(32'hbda4bae8),
	.w7(32'h3babcaca),
	.w8(32'hbc87a42a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5425d0),
	.w1(32'h3c0f2eca),
	.w2(32'hbbca3ba6),
	.w3(32'h3b4a71bd),
	.w4(32'h3b7d825c),
	.w5(32'h3b6db54e),
	.w6(32'h3cbc8318),
	.w7(32'hbc3f7df2),
	.w8(32'h3b6d4ea0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2063cf),
	.w1(32'h3c0df7ec),
	.w2(32'h3994920a),
	.w3(32'hb870c81a),
	.w4(32'hbb7ea97a),
	.w5(32'h3c072a78),
	.w6(32'h3c857376),
	.w7(32'h3b523d3c),
	.w8(32'h3c85675b),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5affa0),
	.w1(32'hb97a9f6d),
	.w2(32'hbc6d21f3),
	.w3(32'h3b93bde2),
	.w4(32'hbb3b42ab),
	.w5(32'hbcf928df),
	.w6(32'hbcf74769),
	.w7(32'hbcac5c32),
	.w8(32'hbd1e677b),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5f6d4e),
	.w1(32'h3cbca396),
	.w2(32'hbbd3d0d2),
	.w3(32'h3c25e061),
	.w4(32'hbb93028d),
	.w5(32'hbb12d5c1),
	.w6(32'h3d29ae4c),
	.w7(32'h3a2903a1),
	.w8(32'h3b257d41),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d7776),
	.w1(32'hbbe985e7),
	.w2(32'h3bee77f7),
	.w3(32'h3b8d7e80),
	.w4(32'h3ba44c68),
	.w5(32'hbb727c6c),
	.w6(32'hbb384942),
	.w7(32'h3b221d5e),
	.w8(32'h3b55f6c7),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9453e2),
	.w1(32'hbc6cf6d1),
	.w2(32'hbc59560d),
	.w3(32'hbcd041af),
	.w4(32'hbb17ee3c),
	.w5(32'hbbae6aa4),
	.w6(32'hbd33da2a),
	.w7(32'hbc628255),
	.w8(32'hbb120287),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a8cb3),
	.w1(32'h3c4bcc91),
	.w2(32'h3c3dd766),
	.w3(32'h3b6660ca),
	.w4(32'h3c48eaf4),
	.w5(32'h3c3141ff),
	.w6(32'h3cd6ada6),
	.w7(32'h3c0c1a6d),
	.w8(32'hbc065b3a),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb781d7e),
	.w1(32'h3c98e48e),
	.w2(32'hbcabc9d4),
	.w3(32'hbbce8e5e),
	.w4(32'hbc84b617),
	.w5(32'hbd1ee18c),
	.w6(32'hbc519bbf),
	.w7(32'hbc5ebd7c),
	.w8(32'h39d9a505),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05481c),
	.w1(32'h3c237f96),
	.w2(32'h3bc96509),
	.w3(32'hba9ff36d),
	.w4(32'h3aeaf561),
	.w5(32'h3bc8811a),
	.w6(32'h3d0c51da),
	.w7(32'h3b16622a),
	.w8(32'h3b95d2a9),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0cdc9),
	.w1(32'h3af675b8),
	.w2(32'hbbb7723e),
	.w3(32'h3cfcd5cf),
	.w4(32'hbb50221c),
	.w5(32'hbbded775),
	.w6(32'h3c8ca029),
	.w7(32'hbc22a946),
	.w8(32'hbc8e3b52),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99f13d),
	.w1(32'h3ca5bc7b),
	.w2(32'hbb4e0533),
	.w3(32'h3c378d1b),
	.w4(32'h3aef9bc1),
	.w5(32'hbc0474b4),
	.w6(32'h3d06371b),
	.w7(32'hbbe33cec),
	.w8(32'hbc5f18f3),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38ac97),
	.w1(32'h3b5e5e1c),
	.w2(32'h3bebbeee),
	.w3(32'hbb393413),
	.w4(32'h3b3d567d),
	.w5(32'h3c76b7c2),
	.w6(32'h3c328470),
	.w7(32'h3c9f59b8),
	.w8(32'h3c8fa1c0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7a9bf),
	.w1(32'hbc9a8f8e),
	.w2(32'hbb2d749a),
	.w3(32'h3b2c097c),
	.w4(32'hbb68fd8e),
	.w5(32'hbc2954c8),
	.w6(32'hbcc7d652),
	.w7(32'h3adf2e21),
	.w8(32'h3bd87f21),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd80938),
	.w1(32'hbbb6f299),
	.w2(32'h3adc0d2b),
	.w3(32'hbcadff20),
	.w4(32'hbc176e24),
	.w5(32'hbb8bb386),
	.w6(32'h3c0376fb),
	.w7(32'hbbcba3bb),
	.w8(32'hbb3b5e94),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86baf3),
	.w1(32'hbc40153c),
	.w2(32'hbaa8182c),
	.w3(32'hbb62915b),
	.w4(32'h3bd10c3b),
	.w5(32'h3c9543ba),
	.w6(32'hbc33e35c),
	.w7(32'h38f89c42),
	.w8(32'hbc17105d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3baa6b),
	.w1(32'h3b142aa1),
	.w2(32'h3aca4c2e),
	.w3(32'h3b275e0f),
	.w4(32'hbbb42126),
	.w5(32'hbc090472),
	.w6(32'hbb269430),
	.w7(32'hbb65d189),
	.w8(32'hbc6a9166),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac7461),
	.w1(32'h3cfcb132),
	.w2(32'hbbd13bbd),
	.w3(32'h3c87bb5b),
	.w4(32'hba8d026a),
	.w5(32'h3a5085ee),
	.w6(32'h3d342120),
	.w7(32'h3c2d4321),
	.w8(32'hbaac8d23),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b8736),
	.w1(32'h3b1b49bb),
	.w2(32'hbc31bf4c),
	.w3(32'h3bc412ae),
	.w4(32'hbc240683),
	.w5(32'h3ae163ab),
	.w6(32'h3c00f7c4),
	.w7(32'h3ab0cdf6),
	.w8(32'hbb963f6f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0237bc),
	.w1(32'h3b34ca90),
	.w2(32'h3bd4f151),
	.w3(32'hbc804da6),
	.w4(32'h3b969791),
	.w5(32'hbbe86c87),
	.w6(32'h3c2987ad),
	.w7(32'h3c06e4a1),
	.w8(32'hbc945f06),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0be46),
	.w1(32'h3c15b230),
	.w2(32'h3c4ba15a),
	.w3(32'h3c3f15ba),
	.w4(32'hbaf9acc3),
	.w5(32'h3a7f0203),
	.w6(32'h3b23894b),
	.w7(32'hb94ce236),
	.w8(32'hbc531845),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca13cfa),
	.w1(32'hbc159858),
	.w2(32'hbc086840),
	.w3(32'hbb25b2f4),
	.w4(32'hbb4f0c12),
	.w5(32'h39947e81),
	.w6(32'hbaefa258),
	.w7(32'hbc28df31),
	.w8(32'h3adfd285),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc658fe8),
	.w1(32'hbbf08ee7),
	.w2(32'hbc925347),
	.w3(32'h3bd98f98),
	.w4(32'hbc1437cb),
	.w5(32'hbb52cfa9),
	.w6(32'hbac169a4),
	.w7(32'hbc97d216),
	.w8(32'hbcbe7044),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc5f106),
	.w1(32'h3ca11016),
	.w2(32'hbbdc3821),
	.w3(32'h3c298cc4),
	.w4(32'h390ea022),
	.w5(32'hbc822ddc),
	.w6(32'h3c8f3a50),
	.w7(32'h3b0d625c),
	.w8(32'hbcb00e31),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b0f9a),
	.w1(32'h3b076920),
	.w2(32'hbb261758),
	.w3(32'h3c4b570a),
	.w4(32'h3af3740b),
	.w5(32'h3bfe8c00),
	.w6(32'h3c99c3fb),
	.w7(32'hbbfd19d0),
	.w8(32'h3c1ec7b1),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fed03),
	.w1(32'h3c146c52),
	.w2(32'h3badad10),
	.w3(32'h3c850de1),
	.w4(32'h3c0f8363),
	.w5(32'h3be760fb),
	.w6(32'h3cc1ba98),
	.w7(32'h3b8c88f3),
	.w8(32'h3b38af60),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f939a),
	.w1(32'hbb66fca3),
	.w2(32'h3a64c270),
	.w3(32'h39eef8b3),
	.w4(32'h3b293242),
	.w5(32'h3b5a4510),
	.w6(32'hbba75546),
	.w7(32'hba167699),
	.w8(32'hb9b6dba1),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b160acf),
	.w1(32'hbae95845),
	.w2(32'hbaea91a3),
	.w3(32'hba7d49f6),
	.w4(32'hbafae953),
	.w5(32'h3a458b25),
	.w6(32'hbaa57735),
	.w7(32'h3ab7dae1),
	.w8(32'h3a4bba08),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac247b9),
	.w1(32'h3aed18ac),
	.w2(32'hbc25342e),
	.w3(32'h3bb0b92f),
	.w4(32'hbbb7fece),
	.w5(32'h3b932bc0),
	.w6(32'h3b0d4759),
	.w7(32'hbc765c7e),
	.w8(32'hb9cc3cdf),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6483ec),
	.w1(32'h3ba8cda7),
	.w2(32'h3b98059b),
	.w3(32'h3bea6197),
	.w4(32'h3bc95bb8),
	.w5(32'h3b682570),
	.w6(32'h3a731a85),
	.w7(32'h3bf744cf),
	.w8(32'hb931cfe4),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9d742),
	.w1(32'hbb0f3a8e),
	.w2(32'hbb4a0e28),
	.w3(32'h3c3b4bba),
	.w4(32'h389a043a),
	.w5(32'h3aec9454),
	.w6(32'h3c06243c),
	.w7(32'hbb161c22),
	.w8(32'hbb133c5e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caa62bd),
	.w1(32'h3b9df732),
	.w2(32'h3c443fce),
	.w3(32'h3cded08e),
	.w4(32'h3c778099),
	.w5(32'h3cc70ac1),
	.w6(32'h3ced647d),
	.w7(32'h3c2426a4),
	.w8(32'h3c6b4676),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c95e8d9),
	.w1(32'h3c42d8c6),
	.w2(32'h3a8fc504),
	.w3(32'h3cad0954),
	.w4(32'h3c175a81),
	.w5(32'h3adfb9d4),
	.w6(32'h3ca784e9),
	.w7(32'hbb953263),
	.w8(32'hbc1296dc),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c681c),
	.w1(32'h3c15cf83),
	.w2(32'h3c025a84),
	.w3(32'hbafa7daa),
	.w4(32'h3bd96024),
	.w5(32'h3b97d0bb),
	.w6(32'hba7fc410),
	.w7(32'hb9e54a32),
	.w8(32'h3b997c24),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2922c),
	.w1(32'hba9f0785),
	.w2(32'h3b0fa9c1),
	.w3(32'hbb6e3e73),
	.w4(32'hb93ed3ec),
	.w5(32'hbbf94995),
	.w6(32'h3ad39420),
	.w7(32'h3b9218bb),
	.w8(32'hbbda6d45),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292f6a),
	.w1(32'hbb1d54e8),
	.w2(32'h3b93260d),
	.w3(32'h3b824ade),
	.w4(32'h3bd8fb4e),
	.w5(32'h3d59b05a),
	.w6(32'h3ba098a0),
	.w7(32'h3c0234e4),
	.w8(32'h3d8712ba),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d75e191),
	.w1(32'h3bc6d322),
	.w2(32'hb8d72f61),
	.w3(32'h3b68c570),
	.w4(32'hbb5005ce),
	.w5(32'hbc3f358b),
	.w6(32'h3ad60f18),
	.w7(32'h3b139239),
	.w8(32'hbc158f31),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc51cde9),
	.w1(32'hba131dea),
	.w2(32'h3ab0aaad),
	.w3(32'hbb0aeea5),
	.w4(32'h3b993d89),
	.w5(32'h3abd834b),
	.w6(32'hba70427e),
	.w7(32'h3ad76b0d),
	.w8(32'h3c2ebfa6),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586b42),
	.w1(32'hbb64f599),
	.w2(32'h3ac7e02e),
	.w3(32'hba89cb35),
	.w4(32'h3b0354d1),
	.w5(32'h3b312725),
	.w6(32'hbbffc748),
	.w7(32'h3c05a732),
	.w8(32'h3b2c9a0d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4070ad),
	.w1(32'h3b085102),
	.w2(32'hbb8e471d),
	.w3(32'h3a8b6851),
	.w4(32'hbc087330),
	.w5(32'hbba36a58),
	.w6(32'hbb001d33),
	.w7(32'hbc047487),
	.w8(32'hbb16c8fc),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20f0c3),
	.w1(32'hbad511a8),
	.w2(32'hbb48f44f),
	.w3(32'h3c379e4c),
	.w4(32'h3bdaae20),
	.w5(32'hba826b21),
	.w6(32'h3c535332),
	.w7(32'h3b8c2f27),
	.w8(32'h3c2bd5b8),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149422),
	.w1(32'h3bac4d4d),
	.w2(32'hbbdcc782),
	.w3(32'hbac9a4c5),
	.w4(32'h3b5bd153),
	.w5(32'h3c01e0da),
	.w6(32'h3ba43d6b),
	.w7(32'h3a60bfab),
	.w8(32'h3c4e44d5),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11f013),
	.w1(32'hbbd1d81b),
	.w2(32'h3b76715e),
	.w3(32'hbba8a04c),
	.w4(32'h3b24145e),
	.w5(32'hbadc73bf),
	.w6(32'hbc0b06a6),
	.w7(32'hba89147e),
	.w8(32'hbb35ba1a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af21a70),
	.w1(32'hbb81cf4f),
	.w2(32'hbc8588d6),
	.w3(32'h3b4cb264),
	.w4(32'hbc18ef7d),
	.w5(32'h3ae3dd33),
	.w6(32'h3aac1038),
	.w7(32'hbc63116f),
	.w8(32'hbb1ea6d1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc73cdf),
	.w1(32'h3bf19512),
	.w2(32'hbc223733),
	.w3(32'h3c7d063b),
	.w4(32'hbaddac37),
	.w5(32'h3b4af6c2),
	.w6(32'h3ca95966),
	.w7(32'hbb75c55e),
	.w8(32'hba5144c7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedc35b),
	.w1(32'hbb433dc0),
	.w2(32'hbc341684),
	.w3(32'hba8d9c07),
	.w4(32'hbb988c21),
	.w5(32'h3bdb48dd),
	.w6(32'h3b0c6dbf),
	.w7(32'hbc43942a),
	.w8(32'hbad87ed3),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac41f3),
	.w1(32'hbad40ca8),
	.w2(32'h3c2a3c32),
	.w3(32'hbb00fe39),
	.w4(32'h3c1a553e),
	.w5(32'hbba1f24b),
	.w6(32'hbc833fc6),
	.w7(32'h3bbef961),
	.w8(32'hbc1de1ca),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b7af),
	.w1(32'hba8e65a8),
	.w2(32'hbb83ee48),
	.w3(32'hbada5fbd),
	.w4(32'h3b2df923),
	.w5(32'hbc812d65),
	.w6(32'hbaee5bfd),
	.w7(32'h3c05fba3),
	.w8(32'hbbc7c7ef),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb8105c),
	.w1(32'h3b0a2067),
	.w2(32'hbc4189e9),
	.w3(32'h3bcb0c13),
	.w4(32'hbbd90cdd),
	.w5(32'hbc0a8796),
	.w6(32'h3c835973),
	.w7(32'hbb602cde),
	.w8(32'hbb3c5055),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17c32e),
	.w1(32'h3b0786c9),
	.w2(32'h3b07afea),
	.w3(32'hbb2a85be),
	.w4(32'h3af3c6a0),
	.w5(32'hbc3b79f3),
	.w6(32'h3b090d94),
	.w7(32'h3bdee5eb),
	.w8(32'hbc115789),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d4763),
	.w1(32'hbc615945),
	.w2(32'h3a784b16),
	.w3(32'hbbf70319),
	.w4(32'hba9ce590),
	.w5(32'hbbb5dbf9),
	.w6(32'hbc0b6af1),
	.w7(32'hb9b53ae9),
	.w8(32'hbbb3c715),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacff34b),
	.w1(32'hb95f839e),
	.w2(32'h3bd600fc),
	.w3(32'hbb50f10d),
	.w4(32'hbb3a9a68),
	.w5(32'hbbccc6be),
	.w6(32'hb9eba7aa),
	.w7(32'h3a15d812),
	.w8(32'hbbb97f86),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb866636),
	.w1(32'hbb720c45),
	.w2(32'hbb87777b),
	.w3(32'h39d04263),
	.w4(32'hbc18273a),
	.w5(32'h3c1c4c43),
	.w6(32'hbb43eb2b),
	.w7(32'hbc3de885),
	.w8(32'h3c0ff54e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61c056),
	.w1(32'h3c681027),
	.w2(32'h3c69cc39),
	.w3(32'h3c789d26),
	.w4(32'h3c336ae0),
	.w5(32'h3bde556c),
	.w6(32'h3c555b9e),
	.w7(32'h3c5a2867),
	.w8(32'hbaa2695d),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7cfea),
	.w1(32'hba0b726d),
	.w2(32'hbbfd4dea),
	.w3(32'h3bc5e2b9),
	.w4(32'h3a3b0a22),
	.w5(32'h3c168dc4),
	.w6(32'h3ac713e0),
	.w7(32'hbb54a8b9),
	.w8(32'h3c1892d4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1f27b),
	.w1(32'h3a9a39ee),
	.w2(32'hbb8dbf24),
	.w3(32'hbbbac631),
	.w4(32'hbaa81e22),
	.w5(32'h3c595519),
	.w6(32'h3ba13ea3),
	.w7(32'hbc47e606),
	.w8(32'h3c6e4941),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb439f6f),
	.w1(32'hba5c6d55),
	.w2(32'hbbc1e8e3),
	.w3(32'h3ae672f9),
	.w4(32'hba1b140c),
	.w5(32'hbac00658),
	.w6(32'h3c6b71a8),
	.w7(32'hbc11b79f),
	.w8(32'h3bda035d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24445c),
	.w1(32'h3be69ace),
	.w2(32'h3b8a564f),
	.w3(32'hbb1021b3),
	.w4(32'hbabff3e3),
	.w5(32'h3b91fc44),
	.w6(32'hba41c7b4),
	.w7(32'h3b40fd6f),
	.w8(32'h3c26e976),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86d079),
	.w1(32'hbb4f0a01),
	.w2(32'hbbfd3b7f),
	.w3(32'h3c562d1b),
	.w4(32'hba248991),
	.w5(32'hbb8a7a82),
	.w6(32'h3c84755e),
	.w7(32'hbc46beb1),
	.w8(32'hbb999afb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ae5fc),
	.w1(32'hbc3e4dde),
	.w2(32'hbb449bfa),
	.w3(32'hb72ccf48),
	.w4(32'hbbc5c533),
	.w5(32'hbc5c6d98),
	.w6(32'h3be401d6),
	.w7(32'hbb3b5516),
	.w8(32'h3ae3c818),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be272f4),
	.w1(32'hbad784fc),
	.w2(32'hbbdb9ca4),
	.w3(32'hbbefc8ec),
	.w4(32'hbc33a21d),
	.w5(32'hbbd4e7c0),
	.w6(32'h3abdae5d),
	.w7(32'hbc7a591a),
	.w8(32'hbbee80d7),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc9a0c),
	.w1(32'hba104ac9),
	.w2(32'hbc8312db),
	.w3(32'hbafc39bc),
	.w4(32'hbc131192),
	.w5(32'h3bd19467),
	.w6(32'h3b20dfc6),
	.w7(32'hbbf49927),
	.w8(32'h3c3d65a2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c7bc1),
	.w1(32'hba772b07),
	.w2(32'h39cfbff5),
	.w3(32'hba6b85bb),
	.w4(32'hbab78e57),
	.w5(32'h3c6902e4),
	.w6(32'hb876817d),
	.w7(32'h3bcfd3e1),
	.w8(32'h3c3fdf73),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16c163),
	.w1(32'hbb995dbb),
	.w2(32'h3bf8b8ab),
	.w3(32'h3c4e5c7e),
	.w4(32'h3757743b),
	.w5(32'h3be23353),
	.w6(32'h3c071cf3),
	.w7(32'hbba408f7),
	.w8(32'hbbb74950),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c680719),
	.w1(32'hbc40e71f),
	.w2(32'hbb9d5e59),
	.w3(32'hbc0e1ba3),
	.w4(32'hbbdd3868),
	.w5(32'h3c3c0e0c),
	.w6(32'hbc5d6348),
	.w7(32'hbbaa9171),
	.w8(32'h3c26bbc4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39d358),
	.w1(32'hbbea27ac),
	.w2(32'hbb008047),
	.w3(32'h3b8c1745),
	.w4(32'h3b69c3a9),
	.w5(32'h3c09298b),
	.w6(32'h3b7e7a8e),
	.w7(32'hbb8bf694),
	.w8(32'h3c089989),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b3651b),
	.w1(32'h3b1db556),
	.w2(32'hbb85d240),
	.w3(32'h3b25b6cd),
	.w4(32'hba27d401),
	.w5(32'h3babc8ba),
	.w6(32'h3c13c0d7),
	.w7(32'h3bc0d07a),
	.w8(32'h3c0a9ff7),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b086c7e),
	.w1(32'h3b14d152),
	.w2(32'hbbad8bdb),
	.w3(32'h3bddea9d),
	.w4(32'hbb662e42),
	.w5(32'h3b688a6c),
	.w6(32'hbbb10dd0),
	.w7(32'hbb935c5d),
	.w8(32'h3bce58e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca467d),
	.w1(32'hb9b61e9a),
	.w2(32'h3c374fd0),
	.w3(32'h3b12fd65),
	.w4(32'h3bc4ef0f),
	.w5(32'h3c81dacb),
	.w6(32'h3bc4ae15),
	.w7(32'h3bd043f4),
	.w8(32'h3c47d2ec),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c664b75),
	.w1(32'h3bf605d4),
	.w2(32'hba6af900),
	.w3(32'h3a655c0a),
	.w4(32'hbaec323b),
	.w5(32'hbb745f91),
	.w6(32'h3b99027e),
	.w7(32'hbb3c6e32),
	.w8(32'hbb8c8edf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc728eb),
	.w1(32'hbbce0ba7),
	.w2(32'hbab9fcc9),
	.w3(32'h3a1b38bf),
	.w4(32'h3af9ab74),
	.w5(32'h3c2a8a28),
	.w6(32'hba58d2db),
	.w7(32'hbba9fdd2),
	.w8(32'h3c57218c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34f802),
	.w1(32'hb9d7ccef),
	.w2(32'hbb5a1ddf),
	.w3(32'h3a9cd68c),
	.w4(32'hbb9f8856),
	.w5(32'h3b171625),
	.w6(32'h3c2924a6),
	.w7(32'hbba24a2b),
	.w8(32'hb9827954),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6aa466),
	.w1(32'h3abe3e8f),
	.w2(32'h393e4957),
	.w3(32'hbb8814f0),
	.w4(32'hbb2efa36),
	.w5(32'h3c1b00b9),
	.w6(32'hbb1c447d),
	.w7(32'h3bf6d8d8),
	.w8(32'h3c8c35ac),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfdeb),
	.w1(32'hbbe74793),
	.w2(32'hba819ffe),
	.w3(32'h3adf7838),
	.w4(32'h3c5213ac),
	.w5(32'h3c532f55),
	.w6(32'hbb1e3fec),
	.w7(32'h3c1f272d),
	.w8(32'h3ccd9f97),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb362df),
	.w1(32'h3c75f0d3),
	.w2(32'hbc712b0a),
	.w3(32'h3b57f584),
	.w4(32'hbc46b2c1),
	.w5(32'hbbb31622),
	.w6(32'h3c16e54e),
	.w7(32'hbc609452),
	.w8(32'hba684beb),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73c318),
	.w1(32'hbb91d6ec),
	.w2(32'hbbb0dc66),
	.w3(32'hbbcfdddd),
	.w4(32'h3a933073),
	.w5(32'hba44994a),
	.w6(32'hbba82511),
	.w7(32'hbc35ca50),
	.w8(32'hbb30016b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule