module layer_10_featuremap_395(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac58e),
	.w1(32'hbb0c3d74),
	.w2(32'hbb3cdf02),
	.w3(32'hbb5f9f0e),
	.w4(32'hbb24517a),
	.w5(32'hbb4bb38f),
	.w6(32'hbb7bcd18),
	.w7(32'hb91ee1ae),
	.w8(32'hbaa92325),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9daf22d),
	.w1(32'h3b5fd268),
	.w2(32'h3b49904b),
	.w3(32'h3b8ffeee),
	.w4(32'h3bde339a),
	.w5(32'h3a44319f),
	.w6(32'h3b0f2a7c),
	.w7(32'hba446b0c),
	.w8(32'hb96a16c5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acde22a),
	.w1(32'h38000d98),
	.w2(32'h3b858efe),
	.w3(32'hbb1f643a),
	.w4(32'hbb91e7bd),
	.w5(32'hbc0f2988),
	.w6(32'h3b0821fa),
	.w7(32'hba826aaa),
	.w8(32'h3a8f817d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a52ee),
	.w1(32'hbafeefd9),
	.w2(32'h3a75a917),
	.w3(32'hbb23a4a4),
	.w4(32'h3b67a44f),
	.w5(32'h39d4929d),
	.w6(32'hbb7909e3),
	.w7(32'hba931207),
	.w8(32'h3bed469b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ee376),
	.w1(32'h379ff2fb),
	.w2(32'hbb804538),
	.w3(32'hbada9aa1),
	.w4(32'hb6cb2506),
	.w5(32'hb9fd3805),
	.w6(32'h3c09c973),
	.w7(32'hbb351929),
	.w8(32'hbb57763f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae3570),
	.w1(32'hbae86530),
	.w2(32'hbb564f34),
	.w3(32'h3974a02d),
	.w4(32'h3b1fa378),
	.w5(32'hbb83f7aa),
	.w6(32'hb9154897),
	.w7(32'hbb7d3960),
	.w8(32'hbb9f42e9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d23b8),
	.w1(32'hbaf4bdf2),
	.w2(32'hbbf82628),
	.w3(32'hbb66a0b6),
	.w4(32'hbb0439fb),
	.w5(32'h3c531117),
	.w6(32'h3b53e070),
	.w7(32'h3c041b31),
	.w8(32'hbb61cfa5),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc750467),
	.w1(32'hbb4d2288),
	.w2(32'hbc3c01eb),
	.w3(32'h3c4f576f),
	.w4(32'hbb5a4bb8),
	.w5(32'hbb089853),
	.w6(32'hbc4fded2),
	.w7(32'hbb5d1a30),
	.w8(32'hbbf81991),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeac8c8),
	.w1(32'h3abef962),
	.w2(32'h3a2c0b2a),
	.w3(32'hbb83ea72),
	.w4(32'hbb63f3c2),
	.w5(32'h3abfe24e),
	.w6(32'hbac32476),
	.w7(32'hbbb044c7),
	.w8(32'h3b2366d1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb147e33),
	.w1(32'hba1b18a5),
	.w2(32'h3b63c77a),
	.w3(32'h3b799a1c),
	.w4(32'hbab370f0),
	.w5(32'h3adbd7d5),
	.w6(32'hba4c4cc8),
	.w7(32'hbb325014),
	.w8(32'h3ad9224f),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913ccb),
	.w1(32'h39fe5fd5),
	.w2(32'h3b5b7265),
	.w3(32'hbb2a7b55),
	.w4(32'h3b7ce777),
	.w5(32'h3b8a33b5),
	.w6(32'h3ad5e57b),
	.w7(32'h3bbe05de),
	.w8(32'h3bdf715d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4e268),
	.w1(32'h3ba17acd),
	.w2(32'h3ab4ee54),
	.w3(32'h3be16da0),
	.w4(32'h3bdff6d2),
	.w5(32'h3b5be456),
	.w6(32'h3b7af9fb),
	.w7(32'h3b08a1cc),
	.w8(32'h39bef67e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a908b53),
	.w1(32'h3b542986),
	.w2(32'h3bd15c68),
	.w3(32'h3b2a8feb),
	.w4(32'h3bd4d9c2),
	.w5(32'hbaf9acda),
	.w6(32'h3b2d011f),
	.w7(32'hbb11f4f9),
	.w8(32'h3ba0ef5e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f17be8),
	.w1(32'h3aaff657),
	.w2(32'hb750d9fc),
	.w3(32'hbc14643a),
	.w4(32'hba1d31c7),
	.w5(32'hbb917c3c),
	.w6(32'h3bc52e30),
	.w7(32'h3b74408b),
	.w8(32'h3ba267f4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9874439),
	.w1(32'h3a4a6783),
	.w2(32'h3aff0a82),
	.w3(32'h3b7bbd25),
	.w4(32'hbb7fd415),
	.w5(32'hbb7e2b43),
	.w6(32'h3baf4f0f),
	.w7(32'hba51529b),
	.w8(32'hbb78625c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb840a),
	.w1(32'h39f6e10b),
	.w2(32'h3a6113a2),
	.w3(32'hbb52a45f),
	.w4(32'hbb93c9ae),
	.w5(32'h3adf4375),
	.w6(32'hba934a94),
	.w7(32'hbb2e37f4),
	.w8(32'hba8a609e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae93659),
	.w1(32'h3ac8c802),
	.w2(32'h3b343311),
	.w3(32'hba6e713a),
	.w4(32'h3931495b),
	.w5(32'h3a44a124),
	.w6(32'hba926e1e),
	.w7(32'h3ab61468),
	.w8(32'h3aba05ab),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd1e321),
	.w1(32'hbc1df11a),
	.w2(32'hbc4138d3),
	.w3(32'hbc619710),
	.w4(32'hbc2a18d8),
	.w5(32'hbc500321),
	.w6(32'hbc0cff69),
	.w7(32'hbc0095bd),
	.w8(32'hbbf1b70a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca6359),
	.w1(32'hbbd3008c),
	.w2(32'hbb8e925b),
	.w3(32'hbc110ce3),
	.w4(32'hbbee4c22),
	.w5(32'hbb95fa41),
	.w6(32'hbb2ca7c7),
	.w7(32'hbb579b0b),
	.w8(32'hbb260487),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb536459),
	.w1(32'h3a18a568),
	.w2(32'hbad92bab),
	.w3(32'h3a82f4ff),
	.w4(32'hbba8246b),
	.w5(32'hb97aba89),
	.w6(32'hbb1124f8),
	.w7(32'hb96d5a1b),
	.w8(32'hbb747c8f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedab01),
	.w1(32'h3b496998),
	.w2(32'h3ba22333),
	.w3(32'h3b805c17),
	.w4(32'h3b8cae9f),
	.w5(32'h3ae79bfa),
	.w6(32'h3a8dd655),
	.w7(32'hba169c08),
	.w8(32'hb9c51bfe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ea017),
	.w1(32'hb8bd4f29),
	.w2(32'h3a10495d),
	.w3(32'hbb075461),
	.w4(32'h3a5ced6e),
	.w5(32'h3bc8b8f7),
	.w6(32'h3b21e2c3),
	.w7(32'hba042327),
	.w8(32'h3b06f66c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35722f),
	.w1(32'hbccee649),
	.w2(32'hbcbc27a8),
	.w3(32'hbc821246),
	.w4(32'hbc93b2d7),
	.w5(32'hbc82e533),
	.w6(32'hbc4aad54),
	.w7(32'hbbefb6d2),
	.w8(32'hbc6ca36c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda18b6),
	.w1(32'h3b9245b1),
	.w2(32'h3bf35977),
	.w3(32'h3b8abb26),
	.w4(32'h3b2e66be),
	.w5(32'h3bb5f5ae),
	.w6(32'hba89842c),
	.w7(32'hb8ef9a2b),
	.w8(32'h3a9c7149),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7efee9),
	.w1(32'h3c1ecead),
	.w2(32'h3c30e081),
	.w3(32'h3bf8caec),
	.w4(32'h3b807938),
	.w5(32'h3c1fe1bb),
	.w6(32'h3b3bdba7),
	.w7(32'h3b28b999),
	.w8(32'h3bdc6942),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7bfb1d),
	.w1(32'hbb4d3256),
	.w2(32'hbaa32571),
	.w3(32'hbba29f39),
	.w4(32'hba46f5dc),
	.w5(32'hb8e6e716),
	.w6(32'hbba49ec9),
	.w7(32'h3b95d654),
	.w8(32'h3bd64057),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24a883),
	.w1(32'hbad827d8),
	.w2(32'h3aadfb16),
	.w3(32'hbb87db4f),
	.w4(32'h3b28b5eb),
	.w5(32'h3bb27cda),
	.w6(32'h3bdfd6df),
	.w7(32'h3b8a1f36),
	.w8(32'hbb4a2a06),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96320b),
	.w1(32'h3a569574),
	.w2(32'h3aec0043),
	.w3(32'h3c2e0846),
	.w4(32'h3a86ae89),
	.w5(32'h3b7efa33),
	.w6(32'hba6516a5),
	.w7(32'h3b1211fb),
	.w8(32'h3acb3100),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10de4f),
	.w1(32'h3aaa6bcd),
	.w2(32'h3a199cb9),
	.w3(32'h3bb037a5),
	.w4(32'h3b60b524),
	.w5(32'hbb938614),
	.w6(32'h3a370887),
	.w7(32'h3a451812),
	.w8(32'hbb407a3a),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2501a),
	.w1(32'h3aff7c20),
	.w2(32'h3ba08216),
	.w3(32'h3b52d871),
	.w4(32'h3b93c650),
	.w5(32'h3ba58110),
	.w6(32'h3b99e6f9),
	.w7(32'h3b0ae88f),
	.w8(32'h3b33e064),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b764894),
	.w1(32'hbb11c76b),
	.w2(32'h3924f89d),
	.w3(32'hbab542f8),
	.w4(32'hbb819b9c),
	.w5(32'hbba5a935),
	.w6(32'hba6aed53),
	.w7(32'hbb8574d2),
	.w8(32'hbb7c46e4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f97a6e),
	.w1(32'hbb7e03e7),
	.w2(32'hb802c1df),
	.w3(32'hbb538e59),
	.w4(32'h382ba5a9),
	.w5(32'hbb519695),
	.w6(32'hba9a6d4d),
	.w7(32'h3ad33662),
	.w8(32'hbb167cdc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891ff9),
	.w1(32'hb9aea245),
	.w2(32'h39020b2a),
	.w3(32'hba3d8f04),
	.w4(32'hbb96889c),
	.w5(32'h3c13ce79),
	.w6(32'hbae7852b),
	.w7(32'h3c5f6766),
	.w8(32'h3c690f95),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae96ce5),
	.w1(32'h3b0955b7),
	.w2(32'h3a25936e),
	.w3(32'h3c50d971),
	.w4(32'hbc09648f),
	.w5(32'hb92469cb),
	.w6(32'h3a19f702),
	.w7(32'h3bf426bf),
	.w8(32'h3bfd955d),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d4be7),
	.w1(32'hbad43edf),
	.w2(32'hbb8b445b),
	.w3(32'h3c35f307),
	.w4(32'hbb48a7b2),
	.w5(32'hbba84f2a),
	.w6(32'hbb99dc77),
	.w7(32'hbbd3d8ab),
	.w8(32'h3834a1f6),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ace1f),
	.w1(32'hba81bd34),
	.w2(32'h39e03c5e),
	.w3(32'hbbd3e620),
	.w4(32'hba2ff527),
	.w5(32'hbb8d5eca),
	.w6(32'hbb058654),
	.w7(32'h38e34b95),
	.w8(32'h3aa7b084),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b710c80),
	.w1(32'hba85d38a),
	.w2(32'hbb845a5f),
	.w3(32'hbc023fd4),
	.w4(32'h3a23bf29),
	.w5(32'h3b8bec9c),
	.w6(32'hba9c65a9),
	.w7(32'h3c0bbc18),
	.w8(32'h3b56c0ef),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c8b48),
	.w1(32'h3c239c63),
	.w2(32'h3bcf507f),
	.w3(32'h3cc928bf),
	.w4(32'h3bbb02a4),
	.w5(32'h3b1f8f40),
	.w6(32'h3be643b1),
	.w7(32'h3b43e0da),
	.w8(32'h3b86795d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48bd7c),
	.w1(32'h3c608b32),
	.w2(32'h3be8dc75),
	.w3(32'h3b2217be),
	.w4(32'hbac81c86),
	.w5(32'hbc0aea31),
	.w6(32'h3c4899b4),
	.w7(32'hba90da03),
	.w8(32'hb960211c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a366e),
	.w1(32'hbbaced07),
	.w2(32'hbaa1c496),
	.w3(32'hbb087ada),
	.w4(32'hbad9bffd),
	.w5(32'h3a9a31ae),
	.w6(32'hbb7a575d),
	.w7(32'hbb71bc29),
	.w8(32'hbb3c10d1),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fe353),
	.w1(32'hbbc63bed),
	.w2(32'hbbba53ff),
	.w3(32'hbab34ef5),
	.w4(32'h3b8ca9da),
	.w5(32'hbbab7cd4),
	.w6(32'h3b73e4cb),
	.w7(32'h3a7a5a1d),
	.w8(32'h3bd0e254),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988188b),
	.w1(32'hba96b4ae),
	.w2(32'hbbb22fd3),
	.w3(32'hbba4c622),
	.w4(32'hbab529d4),
	.w5(32'hbb2ae5a3),
	.w6(32'h3ac13c26),
	.w7(32'h3b2c4b58),
	.w8(32'hbaf91866),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2724da),
	.w1(32'hbc1ccdad),
	.w2(32'hbbcf3fa3),
	.w3(32'h3bb48ec6),
	.w4(32'h3b1d7469),
	.w5(32'hbb3bda0c),
	.w6(32'hbb37fff0),
	.w7(32'hbb05f041),
	.w8(32'h3b85031b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb339f1),
	.w1(32'hbb6113c3),
	.w2(32'h3b81f320),
	.w3(32'hbc1f1324),
	.w4(32'hbbcd108f),
	.w5(32'hbb8984e9),
	.w6(32'hba74fb8e),
	.w7(32'hbbd06e91),
	.w8(32'h38e8887b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf6a00),
	.w1(32'h3a3c2247),
	.w2(32'hb8bff183),
	.w3(32'hb90b8734),
	.w4(32'h3b5167f3),
	.w5(32'h3c79adc9),
	.w6(32'h3b17a09b),
	.w7(32'h3be67925),
	.w8(32'h3bb70ab8),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1adb6d),
	.w1(32'h3b6b013e),
	.w2(32'h3c0199aa),
	.w3(32'h3c5eb95c),
	.w4(32'hba17b27e),
	.w5(32'h3b7ae5b0),
	.w6(32'h3a92d49c),
	.w7(32'h3801ddaa),
	.w8(32'hbac5e346),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b188e69),
	.w1(32'h3b106c58),
	.w2(32'h3c22627c),
	.w3(32'hb892c482),
	.w4(32'hbb70083d),
	.w5(32'h3a2f39d2),
	.w6(32'hb9f6698b),
	.w7(32'hbbb49079),
	.w8(32'h3b47005d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36115e),
	.w1(32'hbc511312),
	.w2(32'hbc5bd2f6),
	.w3(32'hbca4d589),
	.w4(32'hbc6e4f92),
	.w5(32'hbc68ad27),
	.w6(32'hbc217f70),
	.w7(32'hbbcfc54b),
	.w8(32'hbc0650b5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6531a7),
	.w1(32'h3af54d5a),
	.w2(32'h3ab50648),
	.w3(32'hba11794d),
	.w4(32'hb9cd9754),
	.w5(32'h3b973345),
	.w6(32'h3ab21aa5),
	.w7(32'hbb1f9fee),
	.w8(32'hbadf2e01),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f7c2b),
	.w1(32'h3b5e40c3),
	.w2(32'h3b294697),
	.w3(32'h3b2164f2),
	.w4(32'h3b572881),
	.w5(32'h3b6b53c1),
	.w6(32'h3a1f969a),
	.w7(32'h3b8022d3),
	.w8(32'h39a93968),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcc168),
	.w1(32'hbb00ce72),
	.w2(32'hbb6476da),
	.w3(32'hbbb00ef0),
	.w4(32'hbad7a81e),
	.w5(32'hbb4cc25d),
	.w6(32'h3b27183a),
	.w7(32'hbb950964),
	.w8(32'hbb8443b6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc035986),
	.w1(32'hbac13650),
	.w2(32'hb79ca0de),
	.w3(32'hbb635ba1),
	.w4(32'hbb98871d),
	.w5(32'hbb7afb17),
	.w6(32'hba96855b),
	.w7(32'hb913c3d6),
	.w8(32'hbb80f3ba),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae23101),
	.w1(32'hbb90465f),
	.w2(32'hbc0add26),
	.w3(32'hb9bf2d90),
	.w4(32'hbab1c8df),
	.w5(32'h3ab9a15c),
	.w6(32'hbb5b66d2),
	.w7(32'h3b356d25),
	.w8(32'h3a7f1697),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d36a1),
	.w1(32'hbc04b973),
	.w2(32'hbc29a5dd),
	.w3(32'hb9fe37d2),
	.w4(32'hbbaadbfa),
	.w5(32'h399bcca4),
	.w6(32'hbb9d374b),
	.w7(32'hbac5820c),
	.w8(32'hbae5a268),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183a64),
	.w1(32'hbbbb12bc),
	.w2(32'hbb88af5a),
	.w3(32'h39b6d2cc),
	.w4(32'hbb37a7a8),
	.w5(32'hbba081d3),
	.w6(32'h3b13c0a9),
	.w7(32'hbb89dca3),
	.w8(32'hbb665787),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72ec5a),
	.w1(32'hbc0a7f61),
	.w2(32'hbc00d30e),
	.w3(32'hbbf12cc9),
	.w4(32'h3bdd98ba),
	.w5(32'hbb1da31d),
	.w6(32'hbb8e6796),
	.w7(32'hbaedb9d4),
	.w8(32'hbbed18a9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f131c),
	.w1(32'hbb1aa2ad),
	.w2(32'hbb965db1),
	.w3(32'hbbf25ef4),
	.w4(32'hbb4f696d),
	.w5(32'hbb83cfff),
	.w6(32'hbb8172e8),
	.w7(32'hba95ed08),
	.w8(32'hbb82482c),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79ab95),
	.w1(32'h3b83a30a),
	.w2(32'h3b920eca),
	.w3(32'h3ab3493d),
	.w4(32'h3ba7f7fc),
	.w5(32'h3b5225fd),
	.w6(32'hba9c6010),
	.w7(32'h3aa6b453),
	.w8(32'h3b6bff5e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63cdd5),
	.w1(32'hbb7884fa),
	.w2(32'hbb9583dc),
	.w3(32'h3aea52c9),
	.w4(32'hbad974ae),
	.w5(32'hbb82343f),
	.w6(32'h3ba48579),
	.w7(32'hbbb16f2c),
	.w8(32'h37d79a6e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c0474),
	.w1(32'h3b572545),
	.w2(32'h3c021b4a),
	.w3(32'hbb415116),
	.w4(32'h3ab14edf),
	.w5(32'h3acfbb72),
	.w6(32'h3aef450f),
	.w7(32'hbb5e2111),
	.w8(32'h3a7b1a7e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b631e),
	.w1(32'hbb4d7b56),
	.w2(32'hbab62b69),
	.w3(32'hbb57c2eb),
	.w4(32'hbb547348),
	.w5(32'hbac957fc),
	.w6(32'h3990e570),
	.w7(32'hbb62cb19),
	.w8(32'hbb285a21),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5740a6),
	.w1(32'hbb1baf42),
	.w2(32'hbb462878),
	.w3(32'hbbec2e1e),
	.w4(32'hbba5fcc3),
	.w5(32'hbc1e04f4),
	.w6(32'hb8c3b370),
	.w7(32'hbb9479ac),
	.w8(32'hbc0f72c0),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d950f5),
	.w1(32'hbbec77e9),
	.w2(32'h3a8ecfb2),
	.w3(32'h3b6c8ec0),
	.w4(32'h3b152a1a),
	.w5(32'hba889639),
	.w6(32'hbba0ed6b),
	.w7(32'hb9ebdaf9),
	.w8(32'h3b915607),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb965323e),
	.w1(32'h3a6501d5),
	.w2(32'hba028249),
	.w3(32'hbbd8f1d3),
	.w4(32'h3ae55ee5),
	.w5(32'h3adb18a7),
	.w6(32'hbb23bf0e),
	.w7(32'h39d508d1),
	.w8(32'hba6e312d),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b1bdd9),
	.w1(32'hbaf90cb6),
	.w2(32'h3a863c14),
	.w3(32'h3b0985d2),
	.w4(32'h3b19eccc),
	.w5(32'h3b85a4a9),
	.w6(32'hbac2f94c),
	.w7(32'hbb83d802),
	.w8(32'hbb135b01),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5bf15d),
	.w1(32'h3b0887ba),
	.w2(32'hbb568236),
	.w3(32'hb885b0d6),
	.w4(32'h3ab0bf95),
	.w5(32'h3b9095da),
	.w6(32'h3acbcf69),
	.w7(32'h3ba044ab),
	.w8(32'hb89e25e3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc122f30),
	.w1(32'hbb833792),
	.w2(32'h3a16b60d),
	.w3(32'h3be58fc3),
	.w4(32'hbc0689b2),
	.w5(32'hba0f82f7),
	.w6(32'hbb802d6f),
	.w7(32'hbaedb905),
	.w8(32'hb9f30729),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaca96),
	.w1(32'h39cf1cc9),
	.w2(32'h3ae4a91b),
	.w3(32'hba6cabcd),
	.w4(32'h39a60b2a),
	.w5(32'h3a889b9a),
	.w6(32'h3ac39114),
	.w7(32'h3b019baf),
	.w8(32'h397f45cb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5cb0d),
	.w1(32'hbbb81b3d),
	.w2(32'hbbef5f0a),
	.w3(32'hbbaea24f),
	.w4(32'hbbf7180d),
	.w5(32'hbc47772e),
	.w6(32'hbb9e1b45),
	.w7(32'hbbdb4893),
	.w8(32'hbb65f359),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b834124),
	.w1(32'h3c0ce493),
	.w2(32'h3c38775d),
	.w3(32'h3c125a9f),
	.w4(32'h3bc49af4),
	.w5(32'h3c28bc27),
	.w6(32'h3b9c38b4),
	.w7(32'h3b795e5f),
	.w8(32'h3c021454),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b2f09),
	.w1(32'hba5e5e98),
	.w2(32'hb9ded07d),
	.w3(32'h3aa6944b),
	.w4(32'hba97ae5b),
	.w5(32'hbb16e6ff),
	.w6(32'h3a10e03e),
	.w7(32'hb8bf5f80),
	.w8(32'h390adfaa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7944fe),
	.w1(32'h3a75ccd5),
	.w2(32'h3a194e62),
	.w3(32'hba888f13),
	.w4(32'h38f13833),
	.w5(32'hbae65f21),
	.w6(32'hb97f890c),
	.w7(32'hba66a282),
	.w8(32'hbac739a9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e67e72),
	.w1(32'hb848aa78),
	.w2(32'hb9c0df56),
	.w3(32'h39f02372),
	.w4(32'h3ac5d290),
	.w5(32'h397b7080),
	.w6(32'hb919887f),
	.w7(32'h3ad5661e),
	.w8(32'h3a387422),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ad3a8),
	.w1(32'hbb0087c5),
	.w2(32'hbaeeae9c),
	.w3(32'hba7c3f94),
	.w4(32'hba847856),
	.w5(32'hbac10a10),
	.w6(32'hba5ea704),
	.w7(32'hbadf6ae8),
	.w8(32'hbb0506e6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3bc1c52),
	.w1(32'hb9f8c8eb),
	.w2(32'hba21f5c3),
	.w3(32'hb945dc0e),
	.w4(32'hba97eace),
	.w5(32'hbad90a22),
	.w6(32'hba93c2a2),
	.w7(32'h3931e411),
	.w8(32'h3a9745ea),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92bd0b),
	.w1(32'hbbe1052a),
	.w2(32'hbb80b7a3),
	.w3(32'hbbef1990),
	.w4(32'hbc05a965),
	.w5(32'hbb9fc13b),
	.w6(32'hbbd91f7f),
	.w7(32'hbb42f54e),
	.w8(32'hbab84ecf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9539e3),
	.w1(32'hbc3a71e2),
	.w2(32'hbc4d849c),
	.w3(32'hbc118dd5),
	.w4(32'hbc5f4a7c),
	.w5(32'hbc27a97c),
	.w6(32'hbc4241ff),
	.w7(32'hbc08172e),
	.w8(32'hbc10d690),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1d35d),
	.w1(32'h3b6f678b),
	.w2(32'h3b32c337),
	.w3(32'h3a4932d9),
	.w4(32'h3b4a31aa),
	.w5(32'h3b87b2da),
	.w6(32'h3b0b41cd),
	.w7(32'h3b3b97c7),
	.w8(32'h3b5343d0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb354f30),
	.w1(32'hbafea368),
	.w2(32'hba807c93),
	.w3(32'hbb25846e),
	.w4(32'hba778bb8),
	.w5(32'hba22b046),
	.w6(32'hbb61a499),
	.w7(32'hba9cd3cf),
	.w8(32'h39ab9d20),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabd352),
	.w1(32'hbb128cd1),
	.w2(32'hba3fd5d0),
	.w3(32'hb994aea9),
	.w4(32'hbb067346),
	.w5(32'h3a9ce0f4),
	.w6(32'hbacbfaf6),
	.w7(32'hbafa0aba),
	.w8(32'hbb43b923),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba228bd6),
	.w1(32'h3b46291f),
	.w2(32'h3b2d2179),
	.w3(32'hba848db6),
	.w4(32'h3af2a36f),
	.w5(32'h3af69e3d),
	.w6(32'hb9e4f379),
	.w7(32'h3ab6bdff),
	.w8(32'h3af97c2a),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c197),
	.w1(32'hbbaab160),
	.w2(32'hbb84f0c5),
	.w3(32'hbb3af734),
	.w4(32'hbb4836d3),
	.w5(32'hbb3a0a22),
	.w6(32'hbb22730f),
	.w7(32'hbaebbefd),
	.w8(32'hbab5a3bc),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6746e1),
	.w1(32'h3a609892),
	.w2(32'h3a315370),
	.w3(32'h39bee9c1),
	.w4(32'h396e2cf2),
	.w5(32'hb9ba22c4),
	.w6(32'h3a6f15cd),
	.w7(32'h3a151d3e),
	.w8(32'h3a7f39d0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c380f6),
	.w1(32'hba75958b),
	.w2(32'hbb02bf17),
	.w3(32'hb98ab0c8),
	.w4(32'hba62a263),
	.w5(32'hba27d88c),
	.w6(32'h3a41420e),
	.w7(32'hbb002ac7),
	.w8(32'hbafba1e1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381d0063),
	.w1(32'hba0991a2),
	.w2(32'h39887153),
	.w3(32'h3a9df512),
	.w4(32'h399de13b),
	.w5(32'h3a3a27f4),
	.w6(32'hba464fe4),
	.w7(32'h38ba076c),
	.w8(32'h3a01cdf4),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3117b),
	.w1(32'hbab7b32e),
	.w2(32'h39efbd98),
	.w3(32'hba52915b),
	.w4(32'hba760dd2),
	.w5(32'h3b3159c7),
	.w6(32'h3930ef42),
	.w7(32'hba615265),
	.w8(32'hba7c17ce),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d2523),
	.w1(32'h3b702c7d),
	.w2(32'h3b805fff),
	.w3(32'h3a8c82e4),
	.w4(32'h3b20396a),
	.w5(32'h3baa7350),
	.w6(32'h3a3e1a52),
	.w7(32'h3b39fab4),
	.w8(32'h3b710629),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c480d2),
	.w1(32'hb90e72cf),
	.w2(32'hb8a0b3fe),
	.w3(32'h3aad98fe),
	.w4(32'h3a473959),
	.w5(32'h39aea5d7),
	.w6(32'h3a8d88a5),
	.w7(32'h3aee6e1b),
	.w8(32'hba0d2b23),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16c895),
	.w1(32'hbb41e08e),
	.w2(32'hbaec41a4),
	.w3(32'h39b0cf06),
	.w4(32'hbb52d001),
	.w5(32'hbb2a349a),
	.w6(32'hb9d345ac),
	.w7(32'hbb47acdd),
	.w8(32'hba8e38cf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc448d04),
	.w1(32'hbc39c1f1),
	.w2(32'hbc16af8c),
	.w3(32'hbc784fb4),
	.w4(32'hbc329f93),
	.w5(32'hbc282f52),
	.w6(32'hbc73bb08),
	.w7(32'hbbba0eec),
	.w8(32'hbbd39d55),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f946f),
	.w1(32'h3a9677d0),
	.w2(32'hb9378586),
	.w3(32'h3b7b6f5f),
	.w4(32'h3a2cff39),
	.w5(32'h3a95f08b),
	.w6(32'h3b297814),
	.w7(32'h39d28efd),
	.w8(32'hba393acd),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9ff96),
	.w1(32'hba6bae9e),
	.w2(32'h3af07928),
	.w3(32'hbaf1d6c2),
	.w4(32'h3a239a5d),
	.w5(32'h3b5d2996),
	.w6(32'hba1958c7),
	.w7(32'h3b2e1c6d),
	.w8(32'h3a8ed34e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f6ef0),
	.w1(32'h3b5e0650),
	.w2(32'h3b4c7514),
	.w3(32'h3b1ea688),
	.w4(32'h3abfed98),
	.w5(32'h3ab8437c),
	.w6(32'h3b4b10ec),
	.w7(32'h3a11f375),
	.w8(32'h39115597),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb888b17),
	.w1(32'hbac5ebad),
	.w2(32'h3b0cab83),
	.w3(32'hbb614ef7),
	.w4(32'hbada2478),
	.w5(32'h3b04b7eb),
	.w6(32'hbb3b2b5b),
	.w7(32'hbb39ee4e),
	.w8(32'hbaaf8692),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba011771),
	.w1(32'hb9b00568),
	.w2(32'h3abfd37a),
	.w3(32'hb9bda07e),
	.w4(32'hbb189553),
	.w5(32'hba76a32d),
	.w6(32'hbb043f0d),
	.w7(32'hba74be0a),
	.w8(32'hba5290f5),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae28fef),
	.w1(32'h3b59f7fe),
	.w2(32'h3b2d0588),
	.w3(32'h3a7707be),
	.w4(32'h3a9b9d74),
	.w5(32'h3a14c99b),
	.w6(32'h3af750f4),
	.w7(32'hba32dd51),
	.w8(32'hba26bb97),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c8602),
	.w1(32'hb9e6bfc2),
	.w2(32'h3b02c3cd),
	.w3(32'hbae38f2b),
	.w4(32'h3a1a38c1),
	.w5(32'h39f26a61),
	.w6(32'hbaa4fb4c),
	.w7(32'h398d7c46),
	.w8(32'hba984fa6),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43fff0),
	.w1(32'hba4d7409),
	.w2(32'h3ae03876),
	.w3(32'hbb80f949),
	.w4(32'hba75355d),
	.w5(32'h3ad66d98),
	.w6(32'hbad79c3e),
	.w7(32'hb86aabeb),
	.w8(32'h3ad9b4aa),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41c00),
	.w1(32'hbaa877fc),
	.w2(32'hba5b319a),
	.w3(32'h3a021455),
	.w4(32'hb9c6100a),
	.w5(32'hbaca3f96),
	.w6(32'h3b0a2721),
	.w7(32'h3a1bdd04),
	.w8(32'hbb122f1c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd21f5),
	.w1(32'hbc52a2cf),
	.w2(32'hbc201e86),
	.w3(32'hbc4e06d6),
	.w4(32'hbc3fc1eb),
	.w5(32'hbc24dd96),
	.w6(32'hbc86f4ea),
	.w7(32'hbbccf25a),
	.w8(32'hbb9e95a8),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9c1c2),
	.w1(32'h3bec0bc4),
	.w2(32'h3b9e80c5),
	.w3(32'h3c07314f),
	.w4(32'h3b8b762a),
	.w5(32'h3af19db1),
	.w6(32'h3c09bd20),
	.w7(32'h3bb539ed),
	.w8(32'h3ad87220),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a60e0c),
	.w1(32'h3ba4b5ad),
	.w2(32'h3bf1294c),
	.w3(32'h3b54240c),
	.w4(32'h3b863c6d),
	.w5(32'h3bfb19d5),
	.w6(32'h3b44d61b),
	.w7(32'h3b5390ec),
	.w8(32'h3bc6f558),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb20bb7),
	.w1(32'hbbf49623),
	.w2(32'hbba3954c),
	.w3(32'hbb94be3d),
	.w4(32'hbb8d2b34),
	.w5(32'hbbb1914f),
	.w6(32'hbb70ab1c),
	.w7(32'hba977b4a),
	.w8(32'hbb9025c3),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24376e),
	.w1(32'hb8b3f08c),
	.w2(32'hba625ee3),
	.w3(32'h3843a214),
	.w4(32'h38bb6290),
	.w5(32'hbae32fc8),
	.w6(32'h3ab2229e),
	.w7(32'hb995e031),
	.w8(32'hb92af94e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc242da2),
	.w1(32'hbc9291aa),
	.w2(32'hbc862802),
	.w3(32'hbc5cf43b),
	.w4(32'hbc7b053b),
	.w5(32'hbc455395),
	.w6(32'hbc81faee),
	.w7(32'hbc0afc1a),
	.w8(32'hbb8d4cbb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef7c49),
	.w1(32'h3a4297b3),
	.w2(32'h3b086530),
	.w3(32'h3b168b4e),
	.w4(32'hb88c3799),
	.w5(32'h3aefe430),
	.w6(32'h3b3f84b9),
	.w7(32'h3b13a32e),
	.w8(32'h3b30d4ec),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7c708),
	.w1(32'hba5c0342),
	.w2(32'hb95e2149),
	.w3(32'h39b6c106),
	.w4(32'hba69c16f),
	.w5(32'hba8080d8),
	.w6(32'h3a10f2ae),
	.w7(32'hb9c48976),
	.w8(32'hb8cb8c42),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0523f3),
	.w1(32'hb8d91652),
	.w2(32'h39ee9089),
	.w3(32'hb81d269c),
	.w4(32'hba6c4544),
	.w5(32'h3a5ccbe1),
	.w6(32'hba03d1cc),
	.w7(32'hbab79c0d),
	.w8(32'h3951d8b8),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadfcb00),
	.w1(32'h3b29a6dd),
	.w2(32'h3b75db9b),
	.w3(32'h3a6606fa),
	.w4(32'h3a2d21c4),
	.w5(32'h3b20a9c0),
	.w6(32'h3a03ee3b),
	.w7(32'h3b00823f),
	.w8(32'h3b69ded2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a11d8cb),
	.w1(32'h3b6507ac),
	.w2(32'h3b79fb03),
	.w3(32'h3b77c6df),
	.w4(32'h3ad642dc),
	.w5(32'h3ba0875c),
	.w6(32'h3b91ad0f),
	.w7(32'h3a8cc358),
	.w8(32'h3b4b3418),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b03f9),
	.w1(32'hbae3617c),
	.w2(32'hbb5e3733),
	.w3(32'hbaea1050),
	.w4(32'hb967fca8),
	.w5(32'hbb4a6d19),
	.w6(32'hbab05613),
	.w7(32'hba0d1573),
	.w8(32'hbb02c3ab),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1229d),
	.w1(32'h3a9999c4),
	.w2(32'h3b0a2c7a),
	.w3(32'h3ad79590),
	.w4(32'h3a21c0b5),
	.w5(32'h3a87ff3a),
	.w6(32'h3a6a7fc3),
	.w7(32'hb822cd88),
	.w8(32'h393980fb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3de283),
	.w1(32'hba1d3efc),
	.w2(32'h3ae6c4ed),
	.w3(32'hbb12f8ef),
	.w4(32'h3ad5765e),
	.w5(32'h3b24ac05),
	.w6(32'hbb327fdc),
	.w7(32'h3b48845a),
	.w8(32'h3af76447),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbc59f),
	.w1(32'hbb6ec768),
	.w2(32'h397fe251),
	.w3(32'hbafac931),
	.w4(32'hbb64af95),
	.w5(32'hba93d574),
	.w6(32'hba3573e1),
	.w7(32'hbb888d91),
	.w8(32'hbb12a133),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a195396),
	.w1(32'h3a55f7bc),
	.w2(32'h3ae61ced),
	.w3(32'h39ad0ee3),
	.w4(32'h3aa2b6b0),
	.w5(32'h3b114811),
	.w6(32'hba0c95fc),
	.w7(32'h3aaea0ea),
	.w8(32'h3b15e97c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cdae49),
	.w1(32'hb9af6179),
	.w2(32'hb929810a),
	.w3(32'hba1241e1),
	.w4(32'hba0f07a9),
	.w5(32'hba2fbb82),
	.w6(32'h3a06535c),
	.w7(32'h3900682d),
	.w8(32'hb8b74d63),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c2701),
	.w1(32'h3a80ec6e),
	.w2(32'hb98649a3),
	.w3(32'h39b949c9),
	.w4(32'h39400f76),
	.w5(32'h38ff272f),
	.w6(32'h3a691b76),
	.w7(32'hb8e8472c),
	.w8(32'hba96ded0),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4808b3),
	.w1(32'h3a5299a8),
	.w2(32'h3a334ed4),
	.w3(32'h380d234a),
	.w4(32'h39dc9a84),
	.w5(32'h396f2734),
	.w6(32'h3a0eb81c),
	.w7(32'hba29281e),
	.w8(32'hba2164c6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba299c3e),
	.w1(32'h3b141b81),
	.w2(32'h3b09fabe),
	.w3(32'hbb01bcf3),
	.w4(32'h3b2437be),
	.w5(32'h3ab46db8),
	.w6(32'hbb15035e),
	.w7(32'h3af3a84a),
	.w8(32'h3ab55db2),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac05aaf),
	.w1(32'h3afbb88d),
	.w2(32'h3b4b14e3),
	.w3(32'h3b675c33),
	.w4(32'h3abce870),
	.w5(32'h3b30c85c),
	.w6(32'h3b3086c8),
	.w7(32'h3ab5512d),
	.w8(32'h3b11dc67),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39537b74),
	.w1(32'hba6bcbc0),
	.w2(32'hbadb956a),
	.w3(32'h39b7d372),
	.w4(32'hb9d7620b),
	.w5(32'hbaa3c41f),
	.w6(32'h3a6bba49),
	.w7(32'hba2917ac),
	.w8(32'hba8db395),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b4d14),
	.w1(32'hbb5e906e),
	.w2(32'hbb765f10),
	.w3(32'hbaff93d3),
	.w4(32'hbb705c37),
	.w5(32'hbb68118d),
	.w6(32'hbb1fd144),
	.w7(32'hbb604b57),
	.w8(32'hbb034077),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f009),
	.w1(32'h3bb4a139),
	.w2(32'h3ba67a1b),
	.w3(32'h3b9c4d95),
	.w4(32'h3b4f4970),
	.w5(32'h3a6f51f2),
	.w6(32'h3babc1d8),
	.w7(32'h3aea4035),
	.w8(32'hb91c2523),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a3990),
	.w1(32'h38d8e9c1),
	.w2(32'h3a855bb4),
	.w3(32'hba5d68a2),
	.w4(32'hb968071f),
	.w5(32'h3a87394a),
	.w6(32'h3a6e75a9),
	.w7(32'h3800b2c6),
	.w8(32'h39934ad4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f5e32),
	.w1(32'h3aaebb6e),
	.w2(32'h3a40c5ac),
	.w3(32'h3937b5b2),
	.w4(32'h38fe6ae9),
	.w5(32'hb967e3cd),
	.w6(32'h3962a3c5),
	.w7(32'h384bea9f),
	.w8(32'h3a5ae284),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38161bdc),
	.w1(32'h380df935),
	.w2(32'h3ac306ad),
	.w3(32'h3a0481e3),
	.w4(32'h3964ae5e),
	.w5(32'hb97f6345),
	.w6(32'h3a7e6db4),
	.w7(32'hb92cda9c),
	.w8(32'hb96f9d0c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cdc09),
	.w1(32'hbac335b5),
	.w2(32'hbb0caea4),
	.w3(32'h3a38f046),
	.w4(32'hbabdcca0),
	.w5(32'h3a20063b),
	.w6(32'hba545729),
	.w7(32'h39bc0f1e),
	.w8(32'h3b19abce),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ec171),
	.w1(32'hbb88a635),
	.w2(32'hbaa0aa88),
	.w3(32'hbac5d45a),
	.w4(32'hba331de9),
	.w5(32'hbaebbc50),
	.w6(32'hbb19cbbd),
	.w7(32'hbafbd49e),
	.w8(32'hbb0a447e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb403920),
	.w1(32'hb93aea91),
	.w2(32'h3b304a62),
	.w3(32'hbae5c84a),
	.w4(32'hbaa7a160),
	.w5(32'h3aba69f3),
	.w6(32'hb9be995e),
	.w7(32'h3a2d3753),
	.w8(32'h3ae9b979),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4e231),
	.w1(32'hbb1f58d7),
	.w2(32'hbaa135dd),
	.w3(32'hbab845ad),
	.w4(32'hbaf0b8e5),
	.w5(32'hb9d57403),
	.w6(32'hbaa36fde),
	.w7(32'hbb210d97),
	.w8(32'hbacd34ad),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46aa10),
	.w1(32'hba4e3c12),
	.w2(32'hbadaa610),
	.w3(32'hbb19cfaa),
	.w4(32'hb98709fb),
	.w5(32'hba150b4c),
	.w6(32'hbb0be596),
	.w7(32'hba194d6a),
	.w8(32'hbb2b22fe),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac92b57),
	.w1(32'h3a437581),
	.w2(32'h3a9fefb8),
	.w3(32'h3acb0fce),
	.w4(32'h39e2e154),
	.w5(32'hba78691f),
	.w6(32'h3a45a72c),
	.w7(32'hba33d314),
	.w8(32'hb9c4af4f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bc433c),
	.w1(32'hba26f5f1),
	.w2(32'h3a054651),
	.w3(32'hba595a44),
	.w4(32'hb9e30da5),
	.w5(32'h39ddbb01),
	.w6(32'hba39dcdd),
	.w7(32'hb857a36d),
	.w8(32'h3a0c2fc8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114a3c),
	.w1(32'h3b4a4be0),
	.w2(32'h3b86d6cf),
	.w3(32'h3907dd08),
	.w4(32'h3afbc185),
	.w5(32'h3b8a57e7),
	.w6(32'h3a162719),
	.w7(32'h3acaf000),
	.w8(32'h3b1cfed0),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6cc16),
	.w1(32'hbbdafcb3),
	.w2(32'hbb856c08),
	.w3(32'hbc2207aa),
	.w4(32'hbbb5c0f2),
	.w5(32'hbbb2d94b),
	.w6(32'hbbe7fc12),
	.w7(32'hbb438a1f),
	.w8(32'hbba2a228),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e111b),
	.w1(32'h3b41e6bb),
	.w2(32'h3b50e7eb),
	.w3(32'h3b44e2f2),
	.w4(32'h3b270bde),
	.w5(32'h3b5d7ae5),
	.w6(32'h3b0dd984),
	.w7(32'hb9c5e9c3),
	.w8(32'h3a536ca6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2c09da),
	.w1(32'hbb471deb),
	.w2(32'hbab4ae4b),
	.w3(32'hba5f2a01),
	.w4(32'hbaeb411e),
	.w5(32'hbb189212),
	.w6(32'hbb00c60f),
	.w7(32'hbb0e1165),
	.w8(32'hbb6522b0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb782c3),
	.w1(32'hbb902546),
	.w2(32'hbad6ef34),
	.w3(32'hbc0abb4d),
	.w4(32'hbb3166d7),
	.w5(32'hbb83cbd5),
	.w6(32'hbbd6219a),
	.w7(32'h39822206),
	.w8(32'hbaac97dc),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd6de8),
	.w1(32'h3a816978),
	.w2(32'h3afdd3ed),
	.w3(32'h3a51d198),
	.w4(32'h39c90228),
	.w5(32'h3b0e8eba),
	.w6(32'h3a0ba652),
	.w7(32'h3a845c26),
	.w8(32'h3b29a279),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f872d),
	.w1(32'hbb098728),
	.w2(32'h39c19771),
	.w3(32'hbb3ff19c),
	.w4(32'hbb132104),
	.w5(32'h3943445b),
	.w6(32'hba8ce09f),
	.w7(32'hba1ef0b1),
	.w8(32'hba4e9388),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1a607),
	.w1(32'hba10a7ff),
	.w2(32'h3b113f96),
	.w3(32'hba4f0e3a),
	.w4(32'h38c471d0),
	.w5(32'h3a1b4141),
	.w6(32'hb8e79eae),
	.w7(32'h39ff2087),
	.w8(32'h3906b146),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0f3ca),
	.w1(32'h3bdbced1),
	.w2(32'h3bc614ab),
	.w3(32'h3c014776),
	.w4(32'h3b991401),
	.w5(32'h3b823f36),
	.w6(32'h3bbdaca9),
	.w7(32'h3b50dbb2),
	.w8(32'h3b9d5199),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e4961),
	.w1(32'hbb530c34),
	.w2(32'hbb21247c),
	.w3(32'hbb1efb9d),
	.w4(32'hbb3bf9a9),
	.w5(32'hba580576),
	.w6(32'hbb0e2efd),
	.w7(32'hbb206ad0),
	.w8(32'hbab9e297),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef6a68),
	.w1(32'hb906e366),
	.w2(32'h392e702a),
	.w3(32'h393c9d46),
	.w4(32'hb933637e),
	.w5(32'h3741ec75),
	.w6(32'h3a676eb2),
	.w7(32'h399114da),
	.w8(32'h3a73295e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e1da),
	.w1(32'hb9c1ee5f),
	.w2(32'hb989206a),
	.w3(32'h3ad933c4),
	.w4(32'h36ce2eff),
	.w5(32'h3a2f8c85),
	.w6(32'h3ac91145),
	.w7(32'hbaa1c452),
	.w8(32'hbaa00cdb),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c9b6c8),
	.w1(32'h3a57a639),
	.w2(32'h3a8e5e2d),
	.w3(32'h3a752b47),
	.w4(32'hb96d34f9),
	.w5(32'h3accba81),
	.w6(32'h398cceb3),
	.w7(32'h3a93fb09),
	.w8(32'h3aae4f6d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad087b1),
	.w1(32'hb8a29781),
	.w2(32'hba75beb3),
	.w3(32'h3ab2e8d9),
	.w4(32'hba329bbe),
	.w5(32'h3a5b916a),
	.w6(32'hb98d9fdb),
	.w7(32'h38aba19c),
	.w8(32'h39bfd6b0),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad364de),
	.w1(32'hba2e042c),
	.w2(32'h3b39961c),
	.w3(32'hb842ab48),
	.w4(32'h38d15ade),
	.w5(32'h3abc7d6e),
	.w6(32'h3ad235a1),
	.w7(32'h3a9815b6),
	.w8(32'h3aa1333c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04be0d),
	.w1(32'hb82d5174),
	.w2(32'h3a0822cb),
	.w3(32'hbb04ab95),
	.w4(32'hb9efe60e),
	.w5(32'h3a59ca6d),
	.w6(32'hbaf64bea),
	.w7(32'hb9ff1c48),
	.w8(32'hb8997ac5),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaabc524),
	.w1(32'h39230337),
	.w2(32'h3b5b98a5),
	.w3(32'hba66330d),
	.w4(32'hbac387c2),
	.w5(32'h3b78c155),
	.w6(32'hb952439c),
	.w7(32'hba2a7120),
	.w8(32'h3b08e44d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33c6bb),
	.w1(32'h3a04da48),
	.w2(32'h3b1c7826),
	.w3(32'h3adeaabd),
	.w4(32'hba8746ce),
	.w5(32'h3b032cc5),
	.w6(32'h3b1566d7),
	.w7(32'hba053a85),
	.w8(32'h3aede09a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9185fb),
	.w1(32'hbbaab0ac),
	.w2(32'hbbd4745d),
	.w3(32'hbb8e4b90),
	.w4(32'hbb88c219),
	.w5(32'hbb8008ac),
	.w6(32'hbb0dee38),
	.w7(32'hba2503e6),
	.w8(32'hbb1343eb),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacae449),
	.w1(32'h3a3f5531),
	.w2(32'h3a4b3482),
	.w3(32'h3a1436c3),
	.w4(32'h3a639a0e),
	.w5(32'h3acefcde),
	.w6(32'h3b4c1656),
	.w7(32'h39dff570),
	.w8(32'h3aa267ec),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3845a115),
	.w1(32'h3914858b),
	.w2(32'hba89d4b6),
	.w3(32'h3aebb028),
	.w4(32'hba87d568),
	.w5(32'hba96f4fe),
	.w6(32'h3b022689),
	.w7(32'hbae02ee8),
	.w8(32'hb9e004d1),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e0226),
	.w1(32'hba9a9dcb),
	.w2(32'h379e8b0a),
	.w3(32'hba2f2a44),
	.w4(32'hba4fe700),
	.w5(32'hb9b8c623),
	.w6(32'hb98d90c9),
	.w7(32'h39a715ec),
	.w8(32'h39ac7bab),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8da9a28),
	.w1(32'h3a89e9b8),
	.w2(32'h3a8adc69),
	.w3(32'h3b3fa299),
	.w4(32'h3afccb14),
	.w5(32'h3aa98979),
	.w6(32'h3b47c5dc),
	.w7(32'h3b0378f5),
	.w8(32'h3ad800a9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2b9c4),
	.w1(32'h39f1c3c8),
	.w2(32'h37253404),
	.w3(32'h3a5a7336),
	.w4(32'hbaf9fe99),
	.w5(32'hbaa42e22),
	.w6(32'h3ab8f3ca),
	.w7(32'hbb4d15d3),
	.w8(32'h35926e09),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a0e5c),
	.w1(32'h3a8eb266),
	.w2(32'h39919ff1),
	.w3(32'h3af5f689),
	.w4(32'h3a93d26a),
	.w5(32'h3a830a67),
	.w6(32'h3a22e8f7),
	.w7(32'h3a61174c),
	.w8(32'h3a40771e),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f0d44),
	.w1(32'hbb3bed05),
	.w2(32'hbb1359ac),
	.w3(32'hbada45d3),
	.w4(32'hbb12e957),
	.w5(32'hbafaaf0d),
	.w6(32'hbaee8884),
	.w7(32'hbafbf649),
	.w8(32'hba9b97b0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7a140),
	.w1(32'hb9d18f5e),
	.w2(32'h38676852),
	.w3(32'h3a4f26a4),
	.w4(32'h39a7d7d8),
	.w5(32'hb90d3ae3),
	.w6(32'hb9ec1387),
	.w7(32'h384ede97),
	.w8(32'hba5e2cbb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bdea0),
	.w1(32'hba5bda4b),
	.w2(32'h3a56f32c),
	.w3(32'hba9651ab),
	.w4(32'hb95b1dd0),
	.w5(32'h3953849d),
	.w6(32'hbac3df9c),
	.w7(32'h398963a7),
	.w8(32'h38ad1616),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812dd6a),
	.w1(32'h387ebe7e),
	.w2(32'h37a0020e),
	.w3(32'h3a00c301),
	.w4(32'hba1c1f1b),
	.w5(32'hba68e149),
	.w6(32'h3a6adc48),
	.w7(32'h398dc2f9),
	.w8(32'hba8ac9ee),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac001d6),
	.w1(32'h3b096f13),
	.w2(32'h3b19cc2f),
	.w3(32'h3a4d8ae3),
	.w4(32'h3a13a80e),
	.w5(32'h3a74c1ca),
	.w6(32'h3a4f3d1c),
	.w7(32'hb8f4729b),
	.w8(32'h39a9142d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a782f36),
	.w1(32'h395c4468),
	.w2(32'hb9d7df1f),
	.w3(32'hb90086b2),
	.w4(32'h39143d0b),
	.w5(32'hb921c733),
	.w6(32'h399687bf),
	.w7(32'hb98e4ba6),
	.w8(32'hb8478d2b),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2c31b),
	.w1(32'h3acb79cd),
	.w2(32'h3a767009),
	.w3(32'h3adb8eb5),
	.w4(32'h3b0f6d11),
	.w5(32'h3aa1c2ff),
	.w6(32'h39a56cb5),
	.w7(32'h3ade8988),
	.w8(32'hb8b47731),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b76ce0),
	.w1(32'h3971a116),
	.w2(32'h380e14cb),
	.w3(32'hb9295528),
	.w4(32'h3a8bc304),
	.w5(32'h38cd0f35),
	.w6(32'h3915b853),
	.w7(32'h3a2dc1fe),
	.w8(32'hb92e0cc7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f8f79e),
	.w1(32'h395d820e),
	.w2(32'hb99e4b26),
	.w3(32'h3981f443),
	.w4(32'hb9f5aeb0),
	.w5(32'h39c8a129),
	.w6(32'hb96b8656),
	.w7(32'hb853bd60),
	.w8(32'hb9b4724f),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf3c6f),
	.w1(32'h39df1b3e),
	.w2(32'hba57eecd),
	.w3(32'hba42a6f7),
	.w4(32'h3998d0cf),
	.w5(32'h39985172),
	.w6(32'h3ae54587),
	.w7(32'hb954c78b),
	.w8(32'h3a104876),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6309ad),
	.w1(32'hbb9eec48),
	.w2(32'hbb9cc7a7),
	.w3(32'hbb8c17a0),
	.w4(32'hbba7d0c0),
	.w5(32'hbb2d9632),
	.w6(32'hbbab67ea),
	.w7(32'hbb517950),
	.w8(32'hbb3161e1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a279953),
	.w1(32'h37bd2742),
	.w2(32'h3a87d99d),
	.w3(32'h3abee49f),
	.w4(32'h383eaa9b),
	.w5(32'h3a176030),
	.w6(32'h399ab668),
	.w7(32'hb9c51f8b),
	.w8(32'hba204afa),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba2c6a),
	.w1(32'hb978e4f4),
	.w2(32'h39eb0f5f),
	.w3(32'h3b1dd264),
	.w4(32'h3a6d4cff),
	.w5(32'h3898e0ac),
	.w6(32'h3b5b0c95),
	.w7(32'hb8df59b1),
	.w8(32'h3946b936),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9880002),
	.w1(32'h3a84283a),
	.w2(32'h3a9197e6),
	.w3(32'hba2dc07c),
	.w4(32'h3a01f74d),
	.w5(32'h3aa48cec),
	.w6(32'hba5f6989),
	.w7(32'hb84b8e96),
	.w8(32'hb99e832e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c67a5),
	.w1(32'h3905ba45),
	.w2(32'h3a05c76a),
	.w3(32'h3ae3a144),
	.w4(32'h39d5df8c),
	.w5(32'hba29cad6),
	.w6(32'h3b3bbabd),
	.w7(32'h3a81c62a),
	.w8(32'h3ad5bcb6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f3630),
	.w1(32'hbacea74f),
	.w2(32'hbaaf59c2),
	.w3(32'hbadda988),
	.w4(32'hbae99634),
	.w5(32'hba134512),
	.w6(32'hba237010),
	.w7(32'hba82d1a2),
	.w8(32'hb921947b),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3a085),
	.w1(32'hbb9f2574),
	.w2(32'hbad59fcf),
	.w3(32'hbbc56108),
	.w4(32'hbba78ff3),
	.w5(32'hbb32cb6c),
	.w6(32'hbba50a81),
	.w7(32'hbb95950f),
	.w8(32'hbb309169),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04f7ae),
	.w1(32'h39a904fb),
	.w2(32'h3986920f),
	.w3(32'hba95f253),
	.w4(32'hb95118d2),
	.w5(32'h39adefce),
	.w6(32'hbabea300),
	.w7(32'hb9bbb4d4),
	.w8(32'hba75075b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad32055),
	.w1(32'hba2e9259),
	.w2(32'h39c8b55f),
	.w3(32'hbad04a71),
	.w4(32'hbac16b7f),
	.w5(32'h39cd4254),
	.w6(32'hb926830b),
	.w7(32'hbaaf6dd9),
	.w8(32'hb971cd0d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5efb1),
	.w1(32'h38a85dd3),
	.w2(32'hb7918b0c),
	.w3(32'hba5b3ef2),
	.w4(32'hb9190422),
	.w5(32'h3a040bc6),
	.w6(32'hbacc3649),
	.w7(32'h3946b491),
	.w8(32'h3a0ea58d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4be75d),
	.w1(32'h398174a4),
	.w2(32'h3ad45e13),
	.w3(32'h3aac8044),
	.w4(32'h39e56811),
	.w5(32'h3aa9b646),
	.w6(32'hb91f35b7),
	.w7(32'h39a2406e),
	.w8(32'h3a76b92f),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98e84af),
	.w1(32'h3a3e3fcc),
	.w2(32'hb809474c),
	.w3(32'hba2a7e0b),
	.w4(32'hb9b5ee6e),
	.w5(32'h3a368d81),
	.w6(32'hb9a4c204),
	.w7(32'hba65d73e),
	.w8(32'hbaa82c8f),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf40a96),
	.w1(32'h3a1760d8),
	.w2(32'h39700a40),
	.w3(32'hbab58e41),
	.w4(32'h3a4e7c08),
	.w5(32'h3af5e0ce),
	.w6(32'h39d7e696),
	.w7(32'hb9899313),
	.w8(32'h38c4eedf),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8455ba3),
	.w1(32'h3abdd727),
	.w2(32'h3a641f2d),
	.w3(32'h385f19aa),
	.w4(32'h3b02e0ac),
	.w5(32'h3a217d04),
	.w6(32'hb94c9029),
	.w7(32'h3a42678f),
	.w8(32'hb9bfff71),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb957dc22),
	.w1(32'hb9b1947d),
	.w2(32'hbaa45c76),
	.w3(32'hb9dc0c27),
	.w4(32'h3a0b2962),
	.w5(32'h39c1de40),
	.w6(32'h39a4ac61),
	.w7(32'h3a5ffaf6),
	.w8(32'hb9dd183f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c1e01),
	.w1(32'hba380d76),
	.w2(32'hba07f080),
	.w3(32'h3b2d289c),
	.w4(32'h3a1bc451),
	.w5(32'h3a79e73c),
	.w6(32'h3a869cd5),
	.w7(32'h399afa69),
	.w8(32'h3a0b40f5),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f3bac),
	.w1(32'hba3c0a54),
	.w2(32'h3aee6fe2),
	.w3(32'h3ad568da),
	.w4(32'h3aa31ed3),
	.w5(32'h3b04c67e),
	.w6(32'h3a1f2d6c),
	.w7(32'h3b7b6601),
	.w8(32'h3b36de30),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba918865),
	.w1(32'hbacee516),
	.w2(32'hbabfe328),
	.w3(32'hbb0d4313),
	.w4(32'hbad1a7de),
	.w5(32'h39aca14c),
	.w6(32'hba7bda0f),
	.w7(32'hba3e8b50),
	.w8(32'h394d10ce),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36ab30),
	.w1(32'hba8bb02a),
	.w2(32'hbb1cf3e5),
	.w3(32'hbb251a7a),
	.w4(32'hba5f7095),
	.w5(32'hbb6eae21),
	.w6(32'hbafc8ba5),
	.w7(32'hba375060),
	.w8(32'hbb3779ea),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9403),
	.w1(32'hbbab046f),
	.w2(32'hba4bc75b),
	.w3(32'hbb80efca),
	.w4(32'hbb247ea0),
	.w5(32'h3a182b37),
	.w6(32'hba221953),
	.w7(32'h3a00a82d),
	.w8(32'h3b31fb3d),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a976578),
	.w1(32'h3b9126bf),
	.w2(32'h3bce831b),
	.w3(32'h3b4def0c),
	.w4(32'h3aeb7ce1),
	.w5(32'h3b5e40a4),
	.w6(32'h3b92b62a),
	.w7(32'h39d4f519),
	.w8(32'h39d53614),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af67187),
	.w1(32'h385152d7),
	.w2(32'h3a00f238),
	.w3(32'h38d5ead1),
	.w4(32'hb918aa29),
	.w5(32'h3a7722ba),
	.w6(32'hba0389ee),
	.w7(32'h3852d5a3),
	.w8(32'hb9fb53a9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37e14d),
	.w1(32'hb9d077cc),
	.w2(32'hba9d4607),
	.w3(32'h39c6d512),
	.w4(32'hb8c3a27f),
	.w5(32'hbaedcab2),
	.w6(32'h3a326b0b),
	.w7(32'hba75fbd8),
	.w8(32'hba7dc991),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02749b),
	.w1(32'hba540f6e),
	.w2(32'hba410f9d),
	.w3(32'hba1513ff),
	.w4(32'hba216eb7),
	.w5(32'hba85188b),
	.w6(32'hba370667),
	.w7(32'h39ab8baa),
	.w8(32'h39f2cb27),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5cb30),
	.w1(32'h3b069d5e),
	.w2(32'h3a91ee96),
	.w3(32'hba726793),
	.w4(32'h3a9ff529),
	.w5(32'hb98c24b0),
	.w6(32'h3a66a4e7),
	.w7(32'h3aed3c88),
	.w8(32'h3aac5bb2),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba0e60),
	.w1(32'hb951d187),
	.w2(32'h3a910317),
	.w3(32'h3a8d4808),
	.w4(32'h3a0dd384),
	.w5(32'h3afa14a6),
	.w6(32'h3a37d0ed),
	.w7(32'h3acb2db1),
	.w8(32'h3aad0983),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1f02b),
	.w1(32'hbb1b7a0a),
	.w2(32'hbb061ecb),
	.w3(32'hba31baa0),
	.w4(32'hba46ad52),
	.w5(32'hba96d704),
	.w6(32'hba2de219),
	.w7(32'hbaca65f8),
	.w8(32'hbb05d6cd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f84c),
	.w1(32'h3bb11ae6),
	.w2(32'h3be9a7d9),
	.w3(32'h3b252ba2),
	.w4(32'h3b8d989b),
	.w5(32'h3bcbbcdc),
	.w6(32'h3a96e7a2),
	.w7(32'h3b7e0161),
	.w8(32'h3b8b1958),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43dc14),
	.w1(32'h3ae02ff1),
	.w2(32'h3a63f9ce),
	.w3(32'h3a8ec5c8),
	.w4(32'h3ab4e997),
	.w5(32'h3af209b2),
	.w6(32'hba1b95eb),
	.w7(32'hba857854),
	.w8(32'h39e9103a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f3869),
	.w1(32'h3ab1b530),
	.w2(32'hba6327fa),
	.w3(32'h3875ecd4),
	.w4(32'hbbca6bd8),
	.w5(32'hbbef5830),
	.w6(32'h3b11ef11),
	.w7(32'hba627feb),
	.w8(32'hbb14f50c),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950f142),
	.w1(32'hbb1262be),
	.w2(32'h3a0229e3),
	.w3(32'hbb33d7a6),
	.w4(32'hbb9ac0a0),
	.w5(32'hbbafab40),
	.w6(32'h3a468af0),
	.w7(32'hbac3c7ba),
	.w8(32'h3b95ff53),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9d416),
	.w1(32'hbba2f160),
	.w2(32'hb9cdcc31),
	.w3(32'hbb9b57da),
	.w4(32'h3a41c0b7),
	.w5(32'h3b751997),
	.w6(32'h39d17a5a),
	.w7(32'hbb0acf2b),
	.w8(32'h3b898b07),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73c73f),
	.w1(32'h3aa1b984),
	.w2(32'h39d040b5),
	.w3(32'h3af2bd59),
	.w4(32'hbb4c18a3),
	.w5(32'hbb7f3599),
	.w6(32'hb8643485),
	.w7(32'h3adfa1d6),
	.w8(32'hbaf259bb),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d2a6f),
	.w1(32'h3bb37e39),
	.w2(32'h39863fe6),
	.w3(32'h395cd94d),
	.w4(32'h3b7951c3),
	.w5(32'h3ba752c0),
	.w6(32'hbb9ad63d),
	.w7(32'hb751faa9),
	.w8(32'h39aff89f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b6e3),
	.w1(32'hbc5a7417),
	.w2(32'hbb9ee228),
	.w3(32'h3addd211),
	.w4(32'hbbca9a17),
	.w5(32'h3ad8ebb6),
	.w6(32'h3a8ee672),
	.w7(32'h3bc6c7b0),
	.w8(32'h3b81f52f),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd43d2b),
	.w1(32'h3c0a18c4),
	.w2(32'h3c338280),
	.w3(32'h3ab5cba3),
	.w4(32'h3a22af44),
	.w5(32'h3c8de5bd),
	.w6(32'h3a10ff1c),
	.w7(32'hbba1c322),
	.w8(32'hba26acf0),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9462920),
	.w1(32'h3b047db6),
	.w2(32'h3b0c62f7),
	.w3(32'h3c194b36),
	.w4(32'h3a5d9292),
	.w5(32'hbbf60727),
	.w6(32'h3b5f599b),
	.w7(32'h3b8339ed),
	.w8(32'hbab53cd4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51c42b),
	.w1(32'hbb9f778e),
	.w2(32'h3b5235e3),
	.w3(32'h3b3a39c5),
	.w4(32'h3bc40fba),
	.w5(32'h3c99e9d4),
	.w6(32'h3a50cd52),
	.w7(32'hbac4337e),
	.w8(32'h3b86550d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb128026),
	.w1(32'h3b958857),
	.w2(32'h3b47b0b6),
	.w3(32'h3c94573f),
	.w4(32'h3b2e3ad4),
	.w5(32'h3b1fc472),
	.w6(32'h3bf5362e),
	.w7(32'h3a949dbe),
	.w8(32'h3aa49010),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fb62e),
	.w1(32'hbb9ad51f),
	.w2(32'h39cdf327),
	.w3(32'h3b67b7d8),
	.w4(32'h3bd4886b),
	.w5(32'hbb4ec1a4),
	.w6(32'hbad5dcb0),
	.w7(32'h3c3b9b4e),
	.w8(32'h3b87bbb7),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5aea5),
	.w1(32'h3bd4d87a),
	.w2(32'h3a9f9f57),
	.w3(32'h3c00637e),
	.w4(32'hba26afa4),
	.w5(32'hba767b4b),
	.w6(32'h3b6c9c17),
	.w7(32'hba40cce4),
	.w8(32'h3b897cce),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba830652),
	.w1(32'hbaf52d5f),
	.w2(32'hbb8a1776),
	.w3(32'hba935d39),
	.w4(32'hb9b8202c),
	.w5(32'hb8a4c883),
	.w6(32'hbab31cd5),
	.w7(32'h3af7e80a),
	.w8(32'h3bca9620),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f85bd6),
	.w1(32'h3aecd5b0),
	.w2(32'h3b11026c),
	.w3(32'h3bb342a1),
	.w4(32'h3a725510),
	.w5(32'h3a8418ff),
	.w6(32'h3bc263df),
	.w7(32'hbadef613),
	.w8(32'h3b9bfc4a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ca9f8),
	.w1(32'h3bc7ee74),
	.w2(32'hb9805981),
	.w3(32'h3c23051d),
	.w4(32'hb996ea61),
	.w5(32'h3adf2918),
	.w6(32'h3bb94d79),
	.w7(32'h3b244b1a),
	.w8(32'h3bfe2f72),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec545f),
	.w1(32'hbc175c7b),
	.w2(32'h3b12f5fb),
	.w3(32'hbbab8fd7),
	.w4(32'hbc0058d2),
	.w5(32'h3ba1f2e8),
	.w6(32'hbbdc8a4c),
	.w7(32'hbbbfb51f),
	.w8(32'hbb9ab5c1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34cc0),
	.w1(32'hbb889db9),
	.w2(32'h3c16ef68),
	.w3(32'h3c1c4c3c),
	.w4(32'hb8bf18b0),
	.w5(32'hbc5323e5),
	.w6(32'h3c323583),
	.w7(32'hbb85a816),
	.w8(32'hbb315a1d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8569b1),
	.w1(32'hbb58162c),
	.w2(32'h37d746d1),
	.w3(32'hbc5d40ea),
	.w4(32'h3bb7fb80),
	.w5(32'h39ccee3d),
	.w6(32'hbbbb93c6),
	.w7(32'h3a9730fc),
	.w8(32'h3b97944d),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939bf6e),
	.w1(32'hbbc083c2),
	.w2(32'hba4b3e9e),
	.w3(32'hbbafa55a),
	.w4(32'h3b7bab3d),
	.w5(32'hbaed4eb2),
	.w6(32'hbb47a068),
	.w7(32'h3bccd496),
	.w8(32'h3bd229aa),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01c806),
	.w1(32'hbb3054a8),
	.w2(32'hba1e0442),
	.w3(32'hbbe6006b),
	.w4(32'hbb85291c),
	.w5(32'hbbc97c15),
	.w6(32'hbaa82836),
	.w7(32'h3b8d6e35),
	.w8(32'hb98fd9e0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbedcf6),
	.w1(32'hbb017375),
	.w2(32'hbaddd0e3),
	.w3(32'hbc288235),
	.w4(32'h3c0c41bc),
	.w5(32'h3beee883),
	.w6(32'hbbd169b5),
	.w7(32'h3aaafa08),
	.w8(32'h3c72d391),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8acf6f),
	.w1(32'hbc065c3a),
	.w2(32'hbc0bd5c6),
	.w3(32'hbbc91039),
	.w4(32'hbbfdb8ae),
	.w5(32'hbbbfb25c),
	.w6(32'h3baaf4d4),
	.w7(32'hbba1957b),
	.w8(32'hba338d2c),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ede71),
	.w1(32'hbbbcc99e),
	.w2(32'hbc1529af),
	.w3(32'hbc3afa7b),
	.w4(32'hbc267583),
	.w5(32'hbbe65632),
	.w6(32'hbc241d83),
	.w7(32'hbba2ee13),
	.w8(32'hbb87fa62),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32055c),
	.w1(32'hba4961a0),
	.w2(32'hbb38e521),
	.w3(32'h3b859f91),
	.w4(32'hbbc62b78),
	.w5(32'hbb24fadc),
	.w6(32'h3b84f395),
	.w7(32'h395a27c2),
	.w8(32'hb9874ae2),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8a568),
	.w1(32'h3b3d46ba),
	.w2(32'h38f7f600),
	.w3(32'h3b840659),
	.w4(32'h390a40dd),
	.w5(32'h3b187747),
	.w6(32'h3a4f2f0a),
	.w7(32'hba735c55),
	.w8(32'h39e0da9c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20de1d),
	.w1(32'hbaa7bf87),
	.w2(32'h3b9bdf1e),
	.w3(32'hba2b062a),
	.w4(32'h3b340b41),
	.w5(32'h3b02c971),
	.w6(32'h3ae91eb0),
	.w7(32'h3c96e4fb),
	.w8(32'h3b4daf08),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3776bec7),
	.w1(32'h3b7ed4ed),
	.w2(32'hbb85a575),
	.w3(32'h3ac848c5),
	.w4(32'h38a4b709),
	.w5(32'hbc06e4b6),
	.w6(32'h3ad2c684),
	.w7(32'hbb8d0546),
	.w8(32'hbc14bbd8),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adfb9c9),
	.w1(32'hbbcd104b),
	.w2(32'hbb19f3c4),
	.w3(32'hbc27b605),
	.w4(32'hbbe48d0b),
	.w5(32'hbb62819d),
	.w6(32'hbc5420fd),
	.w7(32'hb99d7618),
	.w8(32'hbb8174c6),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaf19c),
	.w1(32'h3abea609),
	.w2(32'hbaac2df2),
	.w3(32'hbb41e06e),
	.w4(32'h3b952d0f),
	.w5(32'h3ba655a1),
	.w6(32'h3b2a7a50),
	.w7(32'hbac6eb43),
	.w8(32'h3b845334),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f0b0d),
	.w1(32'h3aacd164),
	.w2(32'hb94ff1ca),
	.w3(32'hba9ea092),
	.w4(32'h3ba49dbe),
	.w5(32'hbbd3a68b),
	.w6(32'hbb2457b0),
	.w7(32'h3c0540bc),
	.w8(32'h3b4f4263),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698da8),
	.w1(32'h3c12c3f3),
	.w2(32'hbb35b97f),
	.w3(32'hbbde5800),
	.w4(32'h3c3a9dde),
	.w5(32'h3d153278),
	.w6(32'hba02386f),
	.w7(32'hbacaf177),
	.w8(32'hbb9ff99f),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34782a),
	.w1(32'hbab8102e),
	.w2(32'hbb32e7da),
	.w3(32'h3c8e0e5c),
	.w4(32'hbab020d3),
	.w5(32'hb817f0bf),
	.w6(32'hba989137),
	.w7(32'h3bc1baf0),
	.w8(32'h3a7bedf6),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88259e),
	.w1(32'h39589e43),
	.w2(32'h3a182e21),
	.w3(32'hbb8ae4f2),
	.w4(32'hbbc9e120),
	.w5(32'h3c1aca3d),
	.w6(32'hb9de2add),
	.w7(32'hbba968c5),
	.w8(32'hbbbde8fd),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc46cd29),
	.w1(32'hbc0b4ea3),
	.w2(32'hbc01f6d4),
	.w3(32'hbbc636c2),
	.w4(32'hbaa95ce3),
	.w5(32'hb9be84b8),
	.w6(32'hbc33790e),
	.w7(32'hbb2f6294),
	.w8(32'hbb18e908),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd98c52),
	.w1(32'hba9f0ee6),
	.w2(32'hbb2951ef),
	.w3(32'hbc057e5b),
	.w4(32'hbaa608e7),
	.w5(32'h3bcb8b5b),
	.w6(32'hbbb57da0),
	.w7(32'h3b086e75),
	.w8(32'h3acb306e),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7b52a),
	.w1(32'hbb7902bf),
	.w2(32'hbb74d39d),
	.w3(32'h3c2396d6),
	.w4(32'hbb57ab85),
	.w5(32'hbb534cf7),
	.w6(32'h3b95aa8b),
	.w7(32'hbac820d8),
	.w8(32'h3a6a2904),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e02c9),
	.w1(32'hbbd2cbb5),
	.w2(32'hbba97c9c),
	.w3(32'hbc172af4),
	.w4(32'hbbb066cb),
	.w5(32'hbb62f625),
	.w6(32'hbb9dfa9d),
	.w7(32'hba91e27e),
	.w8(32'h3b19eac7),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56f2d1),
	.w1(32'hb98c141a),
	.w2(32'hbb80e204),
	.w3(32'h3a1e3899),
	.w4(32'h3b871aab),
	.w5(32'hba01e912),
	.w6(32'h3b825243),
	.w7(32'h3b51bed2),
	.w8(32'h3b7b2a1c),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdc0b2),
	.w1(32'h3bb8697d),
	.w2(32'h3be22bf4),
	.w3(32'h3a41db3f),
	.w4(32'h3a2c5fb3),
	.w5(32'h3bfaf84d),
	.w6(32'hbb6d4997),
	.w7(32'h3b482c7d),
	.w8(32'hbafab92d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2c3c6),
	.w1(32'hba81da29),
	.w2(32'hbb2e8a21),
	.w3(32'hba8f2c93),
	.w4(32'hbb9de63c),
	.w5(32'h3be9f6b4),
	.w6(32'hbba7292c),
	.w7(32'hbc0c72cd),
	.w8(32'hbb1ce128),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b41b2),
	.w1(32'h3ba28e73),
	.w2(32'h3b8e3f12),
	.w3(32'h3b0961eb),
	.w4(32'hbae3f400),
	.w5(32'h3bd74bba),
	.w6(32'hba228853),
	.w7(32'h3b8e4076),
	.w8(32'h3a2842f6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea5314),
	.w1(32'h3b472557),
	.w2(32'h37f74cd4),
	.w3(32'h3a7f22b9),
	.w4(32'h3a0c0064),
	.w5(32'hba6413b7),
	.w6(32'hbb60a712),
	.w7(32'h3be2daa4),
	.w8(32'h3c10ba9b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a376864),
	.w1(32'h3b3a50d7),
	.w2(32'h3bef1530),
	.w3(32'hb86697ed),
	.w4(32'h3b32d2ab),
	.w5(32'h3c1ce3d9),
	.w6(32'hbb0f26d5),
	.w7(32'hbbc7af2c),
	.w8(32'h3a5451a2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285fb6),
	.w1(32'hb945bb2c),
	.w2(32'h3b22bf5e),
	.w3(32'hbb0b044c),
	.w4(32'hbc2bdd58),
	.w5(32'hbb476be2),
	.w6(32'h3c06e0d7),
	.w7(32'hbaad3528),
	.w8(32'hbb259629),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8420cc),
	.w1(32'h3a4d3139),
	.w2(32'h3b28349d),
	.w3(32'hbac601dd),
	.w4(32'hba0f05b6),
	.w5(32'h3b4f39a6),
	.w6(32'hbb1d167c),
	.w7(32'h3a15874d),
	.w8(32'hba4b2425),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8c44),
	.w1(32'hbb0504b5),
	.w2(32'h3aebacd3),
	.w3(32'hba33feac),
	.w4(32'h3b909245),
	.w5(32'hbb2a1739),
	.w6(32'h3b0e66ac),
	.w7(32'h3bc13b67),
	.w8(32'h3bff38a1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c410646),
	.w1(32'h3b3c3a41),
	.w2(32'h3ad9711e),
	.w3(32'h39bb9b7b),
	.w4(32'hb92c8373),
	.w5(32'hb8e732a1),
	.w6(32'h3c292e0f),
	.w7(32'h3ab93734),
	.w8(32'h3ad604fc),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f8cfd),
	.w1(32'hb8ebcd0b),
	.w2(32'h3bb05f06),
	.w3(32'h3bc37608),
	.w4(32'hbb43ad53),
	.w5(32'hbacbf629),
	.w6(32'h3bddd27a),
	.w7(32'h3b8d57fe),
	.w8(32'h3b6f32e6),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b9f43),
	.w1(32'h3ba4d849),
	.w2(32'hbaa02d61),
	.w3(32'h3be8b094),
	.w4(32'hbb065f8c),
	.w5(32'hba8075af),
	.w6(32'h3adb236e),
	.w7(32'h3b961488),
	.w8(32'h3b35a451),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37baf4),
	.w1(32'hbbe5ffa5),
	.w2(32'hb908025c),
	.w3(32'hb9743a82),
	.w4(32'hbb811082),
	.w5(32'hbb647134),
	.w6(32'h3b8d22d6),
	.w7(32'hbbf575f1),
	.w8(32'hbb8287ca),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f29db),
	.w1(32'h3a3b5fa7),
	.w2(32'hbb4386e0),
	.w3(32'hb99117e0),
	.w4(32'hba904512),
	.w5(32'hb80663fd),
	.w6(32'hbbb99955),
	.w7(32'hbaa3d6ca),
	.w8(32'h3a997f94),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32241b),
	.w1(32'hba8122b9),
	.w2(32'hbb310ccb),
	.w3(32'h3b73bed6),
	.w4(32'hbbe1346e),
	.w5(32'hbc086245),
	.w6(32'h3b797a36),
	.w7(32'h3b0b6e2d),
	.w8(32'hbbbad33b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be73311),
	.w1(32'hb90a97a5),
	.w2(32'hbbc64614),
	.w3(32'hbbabbce1),
	.w4(32'hbc1891d2),
	.w5(32'hbc0ec99c),
	.w6(32'hbbe4f8ba),
	.w7(32'hbb880355),
	.w8(32'h3a28a527),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeae764),
	.w1(32'hbbead914),
	.w2(32'h3b37ed77),
	.w3(32'hbb35d079),
	.w4(32'hbc012d6d),
	.w5(32'hbbbd91c2),
	.w6(32'hbb1e3fc7),
	.w7(32'h3a55ed13),
	.w8(32'h3aa0c29d),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd896),
	.w1(32'h3af81b69),
	.w2(32'h3ba660d6),
	.w3(32'hb9f0d608),
	.w4(32'hba77ae38),
	.w5(32'h3c80cb4b),
	.w6(32'h3b9f52bc),
	.w7(32'hba4acedd),
	.w8(32'h3a83db1e),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8d004),
	.w1(32'hba24c7e1),
	.w2(32'h3bb3bc81),
	.w3(32'h3c0d58cf),
	.w4(32'h38875f1b),
	.w5(32'h3ca7a17a),
	.w6(32'h3bef20f7),
	.w7(32'hbba39474),
	.w8(32'hb92b112c),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba652b2),
	.w1(32'hbbc6f3a7),
	.w2(32'hbbbc20d1),
	.w3(32'h3ab9e177),
	.w4(32'hbc1538da),
	.w5(32'hbc3016bb),
	.w6(32'h3a8cc4b2),
	.w7(32'hbb9ec9b1),
	.w8(32'hbbc9e3cb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34dd93),
	.w1(32'hbaf0b3a0),
	.w2(32'h3c07262d),
	.w3(32'hbc21cab1),
	.w4(32'hba25e5ec),
	.w5(32'hbabefbfd),
	.w6(32'hbab53fb1),
	.w7(32'h3b82253c),
	.w8(32'hbb950895),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55dc7d),
	.w1(32'hbb5a19ca),
	.w2(32'hbb7f30ce),
	.w3(32'h3b180fba),
	.w4(32'hbb109ae1),
	.w5(32'hbaf5bb93),
	.w6(32'hbafa3f7d),
	.w7(32'hbaadf8f1),
	.w8(32'h3b644061),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule