module layer_8_featuremap_41(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32b4af),
	.w1(32'h3ad69081),
	.w2(32'h3b146811),
	.w3(32'hbb8cb81c),
	.w4(32'h392acc3c),
	.w5(32'h3ae869b8),
	.w6(32'hb9c2c902),
	.w7(32'h39055227),
	.w8(32'hbb0102cd),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09bfde),
	.w1(32'hbb10a681),
	.w2(32'hbab53b65),
	.w3(32'hbb0be4f6),
	.w4(32'hbb070e0f),
	.w5(32'hba26d56b),
	.w6(32'hbb1d19d9),
	.w7(32'hbad698e5),
	.w8(32'hb8edc5ff),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d1dc9b),
	.w1(32'hba1e9838),
	.w2(32'hb8b828ed),
	.w3(32'hba0c6ba0),
	.w4(32'hb9c6fa80),
	.w5(32'h3a37739e),
	.w6(32'hb9a87a92),
	.w7(32'hb61ca77d),
	.w8(32'h395c02e3),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb493fa4),
	.w1(32'hbbaa7f07),
	.w2(32'hbac1274d),
	.w3(32'h3b393376),
	.w4(32'h3a17dd85),
	.w5(32'h3b3d024e),
	.w6(32'hba74f0be),
	.w7(32'h3b2828f9),
	.w8(32'h3b75e255),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b445471),
	.w1(32'h3a99b86b),
	.w2(32'h3a3b20ae),
	.w3(32'h3adc8e9f),
	.w4(32'h3a958edf),
	.w5(32'h3af2b429),
	.w6(32'h3af38d71),
	.w7(32'h3a367e84),
	.w8(32'hb91ded80),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ba6bf),
	.w1(32'hbc90a25e),
	.w2(32'hbc913820),
	.w3(32'hbc1d7053),
	.w4(32'hbc8ec648),
	.w5(32'hbc743c85),
	.w6(32'hbc44446a),
	.w7(32'hbc5780c1),
	.w8(32'hb8ebcd12),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba08c71a),
	.w1(32'hb9c726cd),
	.w2(32'h3a245924),
	.w3(32'hbad896fa),
	.w4(32'hba1b858e),
	.w5(32'h3ac34f26),
	.w6(32'h38590b61),
	.w7(32'h3a58444b),
	.w8(32'h3af61ec1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a34dd0e),
	.w1(32'hbacf5c18),
	.w2(32'hba84d17d),
	.w3(32'h398970ac),
	.w4(32'hba82d5f8),
	.w5(32'h38b06823),
	.w6(32'h3841f11c),
	.w7(32'hb95f4143),
	.w8(32'h3a13cbac),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3919335c),
	.w1(32'hba4297af),
	.w2(32'h3a2c9b3c),
	.w3(32'hba45b7fc),
	.w4(32'hb9b67d77),
	.w5(32'h3b113804),
	.w6(32'hb9be90f7),
	.w7(32'h3a5bac99),
	.w8(32'h3a385eca),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa00511),
	.w1(32'hbb6656f2),
	.w2(32'hbb821485),
	.w3(32'h3baf1c15),
	.w4(32'h3a87bae1),
	.w5(32'hbb854111),
	.w6(32'h3a7960d2),
	.w7(32'hbb58517f),
	.w8(32'h3b230467),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f3220),
	.w1(32'hba9f76a9),
	.w2(32'h3a4893bb),
	.w3(32'h3ab7e642),
	.w4(32'h39c6ace6),
	.w5(32'h3b152a54),
	.w6(32'h3ad0e7c3),
	.w7(32'h3b5d36b3),
	.w8(32'hbb0628d4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5331f),
	.w1(32'hba92c56e),
	.w2(32'hba957571),
	.w3(32'hbb2dfd14),
	.w4(32'hbaaf4466),
	.w5(32'hb9342021),
	.w6(32'hbade2197),
	.w7(32'hbaec0ff8),
	.w8(32'hba82f9e9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08839f),
	.w1(32'hbb4ff74b),
	.w2(32'hba5150bc),
	.w3(32'hba87c958),
	.w4(32'hbaa218ff),
	.w5(32'h3a8a31c9),
	.w6(32'hbad7555f),
	.w7(32'h3a361deb),
	.w8(32'h3b3a1bf1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1824fe),
	.w1(32'hbca318ff),
	.w2(32'hbc9fd264),
	.w3(32'hbc11eff9),
	.w4(32'hbc9e1d33),
	.w5(32'hbc84c9ea),
	.w6(32'hbc49320a),
	.w7(32'hbc579fae),
	.w8(32'hbb77441b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc018133),
	.w1(32'hbc4750ad),
	.w2(32'hbc36cf95),
	.w3(32'hbc098c9b),
	.w4(32'hbc3c4d21),
	.w5(32'hbc12a77a),
	.w6(32'hbc11507e),
	.w7(32'hbc1acae2),
	.w8(32'hbb9bdba8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb44425),
	.w1(32'hbb9adebd),
	.w2(32'hbb19dfe0),
	.w3(32'hbb8fdbbd),
	.w4(32'hbb9460be),
	.w5(32'hbab01f57),
	.w6(32'hbb91c768),
	.w7(32'hbb21f3c5),
	.w8(32'hbad2254a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b571fa1),
	.w1(32'h3bb370c8),
	.w2(32'h3bc7380a),
	.w3(32'hb997d757),
	.w4(32'hbb6794dd),
	.w5(32'hbb992729),
	.w6(32'hbb5035b3),
	.w7(32'hbb7461be),
	.w8(32'hbaab3f11),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2ae86),
	.w1(32'hbb156126),
	.w2(32'hb9f0ae43),
	.w3(32'hb9d9e347),
	.w4(32'hba1fbb0e),
	.w5(32'h396464a8),
	.w6(32'hbad933f0),
	.w7(32'h3a4ab713),
	.w8(32'h396223a5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2aad25),
	.w1(32'hbbe17210),
	.w2(32'hbb827009),
	.w3(32'h3a43fe0a),
	.w4(32'hbb8ffa19),
	.w5(32'hbac4320b),
	.w6(32'hbb8a7dd9),
	.w7(32'hbaee23ae),
	.w8(32'hbb9f1aad),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0769bb),
	.w1(32'h3b8d8156),
	.w2(32'h3b15f305),
	.w3(32'hba5bdb17),
	.w4(32'h39aefadf),
	.w5(32'hbbedb728),
	.w6(32'hbbb5c6fd),
	.w7(32'hbb0c68bf),
	.w8(32'h3bdee459),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3abc3),
	.w1(32'h3b9ad6a9),
	.w2(32'h3c01cfd0),
	.w3(32'h3c0ff626),
	.w4(32'h3bec6f4d),
	.w5(32'h3be8b573),
	.w6(32'h3bbc8702),
	.w7(32'h3c0b5396),
	.w8(32'h3c025702),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be811b9),
	.w1(32'h3b9be551),
	.w2(32'h3b545c09),
	.w3(32'h3ba263ba),
	.w4(32'h3b77d3e5),
	.w5(32'h3b8b9bbd),
	.w6(32'h3bb08fe8),
	.w7(32'h3b7478b8),
	.w8(32'h3cddf3b9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9956e3),
	.w1(32'h3c5df020),
	.w2(32'h3c9eda7c),
	.w3(32'h3cbe28ef),
	.w4(32'h3c87bac8),
	.w5(32'h3c992054),
	.w6(32'h3c95e627),
	.w7(32'h3ccbba33),
	.w8(32'hb884079a),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7c82e),
	.w1(32'hbb80d452),
	.w2(32'hba8d36e6),
	.w3(32'hb88dbe86),
	.w4(32'hbb264da5),
	.w5(32'hb7a2c2f3),
	.w6(32'hbb233e40),
	.w7(32'hb9276a97),
	.w8(32'hbb81fda8),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb3873),
	.w1(32'hbc197cad),
	.w2(32'hbb5e80e7),
	.w3(32'hba9470fc),
	.w4(32'hbbf5e240),
	.w5(32'hbba85ceb),
	.w6(32'hbc281fba),
	.w7(32'hbb2bf11c),
	.w8(32'h3cd224e9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c909d87),
	.w1(32'h3c4ecfa3),
	.w2(32'h3c92e0eb),
	.w3(32'h3cb36551),
	.w4(32'h3c7c127a),
	.w5(32'h3c8d2826),
	.w6(32'h3c8eee6e),
	.w7(32'h3cbedf3c),
	.w8(32'h3cb108e2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c1144),
	.w1(32'h3c350b9e),
	.w2(32'h3c807a88),
	.w3(32'h3c9b0860),
	.w4(32'h3c5aacb8),
	.w5(32'h3c75e58f),
	.w6(32'h3c775b7a),
	.w7(32'h3ca3e926),
	.w8(32'h3c3f41fe),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3598a3),
	.w1(32'h3c6a6aa7),
	.w2(32'h3c87cfc1),
	.w3(32'h3c76b0ac),
	.w4(32'h3c82ddfe),
	.w5(32'h3c713881),
	.w6(32'h3c6a6100),
	.w7(32'h3c8faa4b),
	.w8(32'hbb851426),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f5c05),
	.w1(32'hbbc7b6a4),
	.w2(32'hbb4e2c15),
	.w3(32'h3b336bdb),
	.w4(32'hbab489da),
	.w5(32'h3b83e610),
	.w6(32'hbbca7e36),
	.w7(32'h3ad17732),
	.w8(32'hba8c6b51),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba540c98),
	.w1(32'hba3e21f8),
	.w2(32'hba84bf0e),
	.w3(32'hba6daf4b),
	.w4(32'hba1e5874),
	.w5(32'hba031ac9),
	.w6(32'hba35bc9e),
	.w7(32'hba99dbea),
	.w8(32'hbb2087a8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96596f),
	.w1(32'hbb49d09d),
	.w2(32'h3ab6fa98),
	.w3(32'hba6c1a45),
	.w4(32'hbb25a447),
	.w5(32'h3b129a38),
	.w6(32'hbbc88ea8),
	.w7(32'hba6a7fd7),
	.w8(32'h37893978),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5ee7d),
	.w1(32'hbbd5173f),
	.w2(32'h3a726aff),
	.w3(32'h3b8a86bd),
	.w4(32'hbaf693c3),
	.w5(32'hb9f42462),
	.w6(32'hbbc306c3),
	.w7(32'h39bafb2c),
	.w8(32'hbb28647c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd3401),
	.w1(32'hbb5a5966),
	.w2(32'hba2e7bc6),
	.w3(32'hbbad7950),
	.w4(32'hbb260811),
	.w5(32'h3a5de7a6),
	.w6(32'h3ad73729),
	.w7(32'h3afbb237),
	.w8(32'hbb82f680),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f0b08),
	.w1(32'h3a1fe255),
	.w2(32'h39ecb408),
	.w3(32'h3b5e64ab),
	.w4(32'hba076049),
	.w5(32'hbae8cf62),
	.w6(32'hbbc02921),
	.w7(32'hba87c6e7),
	.w8(32'h3b209ead),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04ee2a),
	.w1(32'hbc8e1944),
	.w2(32'hbc8b6040),
	.w3(32'hbbfcb543),
	.w4(32'hbc891618),
	.w5(32'hbc66dba3),
	.w6(32'hbc2f3329),
	.w7(32'hbc3a8da7),
	.w8(32'hbaa99d5c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5871e7),
	.w1(32'hbb646435),
	.w2(32'h3938d3ea),
	.w3(32'hbb437dca),
	.w4(32'hbb27bdb6),
	.w5(32'h3a90b60c),
	.w6(32'hbb2d5d70),
	.w7(32'h388949ac),
	.w8(32'h3bf1fa09),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c35cc38),
	.w1(32'h3c7018b8),
	.w2(32'h3c517e9b),
	.w3(32'h3c3f30e2),
	.w4(32'h3c51c719),
	.w5(32'h3c21c8a9),
	.w6(32'h3c1e6d68),
	.w7(32'h3c40c8e8),
	.w8(32'hb8ff843c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95594c2),
	.w1(32'hba804c85),
	.w2(32'hba640f9e),
	.w3(32'hb97e211e),
	.w4(32'hb9b9e216),
	.w5(32'h388d32c1),
	.w6(32'hba183b37),
	.w7(32'hba38a093),
	.w8(32'hbc00052a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5bcd8d),
	.w1(32'hbc9af573),
	.w2(32'hbc885380),
	.w3(32'hbc7408c0),
	.w4(32'hbc931221),
	.w5(32'hbc5aab24),
	.w6(32'hbc679e52),
	.w7(32'hbc796777),
	.w8(32'h3b6573e1),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6aa91),
	.w1(32'h3bfeb162),
	.w2(32'h3c26f0fa),
	.w3(32'h3c19fd20),
	.w4(32'h3c225b2f),
	.w5(32'h3c1614c5),
	.w6(32'h3bc14147),
	.w7(32'h3c1a60e1),
	.w8(32'h3c1f4612),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcfcc8),
	.w1(32'h3bb00590),
	.w2(32'h3bf2ddc5),
	.w3(32'h3c096783),
	.w4(32'h3bd3b57a),
	.w5(32'h3be85d0e),
	.w6(32'h3bddec0e),
	.w7(32'h3c183c74),
	.w8(32'hba2f987a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09257e),
	.w1(32'hb9ee1151),
	.w2(32'hb9abffd9),
	.w3(32'hb9a36894),
	.w4(32'hb89ca924),
	.w5(32'hb95dda5f),
	.w6(32'hb9f2f2e4),
	.w7(32'hb7a86ba5),
	.w8(32'h3a6b6679),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399ab462),
	.w1(32'h3706b96b),
	.w2(32'hba045612),
	.w3(32'h3a1c8436),
	.w4(32'hbaa33538),
	.w5(32'h39a6fa94),
	.w6(32'hb9c0caf8),
	.w7(32'hbab267a6),
	.w8(32'hb9f21845),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e315d4),
	.w1(32'hba130625),
	.w2(32'hb88c9016),
	.w3(32'hb8a38893),
	.w4(32'hb996f7a0),
	.w5(32'hb92b8631),
	.w6(32'hba1c8685),
	.w7(32'h37a1919f),
	.w8(32'h386c6a23),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396fb55b),
	.w1(32'h39afd4b4),
	.w2(32'h39226738),
	.w3(32'h3a1f11e6),
	.w4(32'h39fae056),
	.w5(32'h3913443e),
	.w6(32'h3a2e246c),
	.w7(32'h3a217337),
	.w8(32'hba33a176),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba797359),
	.w1(32'hb9ca8eb3),
	.w2(32'hba06ab3d),
	.w3(32'hb9e286ee),
	.w4(32'hb94d78ec),
	.w5(32'h38b2d867),
	.w6(32'hba0aa089),
	.w7(32'hb8d5cd39),
	.w8(32'hbb09288e),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e1866),
	.w1(32'hba1c8859),
	.w2(32'hb9aee18d),
	.w3(32'hbaff3b00),
	.w4(32'hbb4627c8),
	.w5(32'h3aa098c6),
	.w6(32'hbb285c70),
	.w7(32'hbad28ea5),
	.w8(32'hba2f8211),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d4d1),
	.w1(32'hbad4421d),
	.w2(32'hb9c43f94),
	.w3(32'hba9a9c2d),
	.w4(32'hba86ab54),
	.w5(32'hba2f2441),
	.w6(32'hb9c188be),
	.w7(32'h38ea4d78),
	.w8(32'h3a9b5fa9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26bee2),
	.w1(32'hba1fd617),
	.w2(32'hba55cb0c),
	.w3(32'h3a9bd968),
	.w4(32'h3988b379),
	.w5(32'h38bf890d),
	.w6(32'hb9de7260),
	.w7(32'hba2669a6),
	.w8(32'hb866796d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d88c11),
	.w1(32'h38ef855b),
	.w2(32'h3998b5ae),
	.w3(32'h39ef05f5),
	.w4(32'h3a08fe0f),
	.w5(32'h3a0b5b9d),
	.w6(32'h39ce65e2),
	.w7(32'h3a3e05b1),
	.w8(32'hb84df56b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba134475),
	.w1(32'hb9cce93b),
	.w2(32'hb99e3c5b),
	.w3(32'hb9b0b688),
	.w4(32'hb92dbdac),
	.w5(32'hb9b8873a),
	.w6(32'hb9b2deca),
	.w7(32'hb97fa089),
	.w8(32'hba6f38be),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfc0ec),
	.w1(32'hba04829c),
	.w2(32'hba6c216f),
	.w3(32'h389ed7fd),
	.w4(32'hb92731ec),
	.w5(32'hba818b14),
	.w6(32'hb94ce844),
	.w7(32'hb9a46bbb),
	.w8(32'hb9e19293),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a159da0),
	.w1(32'h37931ba5),
	.w2(32'hb9c0ff23),
	.w3(32'hba28340c),
	.w4(32'hb92396fc),
	.w5(32'hba6a3607),
	.w6(32'h3a926599),
	.w7(32'hba06c970),
	.w8(32'hb97ac57e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d4f84a),
	.w1(32'hba1f823c),
	.w2(32'hb9e2f58f),
	.w3(32'h3929ee5b),
	.w4(32'hb80f86ba),
	.w5(32'h39520a6f),
	.w6(32'hb9fb433e),
	.w7(32'hb9d9b214),
	.w8(32'hba7b1cbe),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2bd615),
	.w1(32'h3b1f77c6),
	.w2(32'h3ac001ec),
	.w3(32'hbaba47ae),
	.w4(32'h3a826614),
	.w5(32'h3a9be70a),
	.w6(32'h398953ed),
	.w7(32'h39649a4e),
	.w8(32'hbaa21bb6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245c2e),
	.w1(32'hbb3ab5d0),
	.w2(32'hba8f659a),
	.w3(32'hbb0c231c),
	.w4(32'hbb2fdcb2),
	.w5(32'hba963e89),
	.w6(32'hbb2156c8),
	.w7(32'hba669301),
	.w8(32'hba7a3106),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8536ea),
	.w1(32'hbabb11aa),
	.w2(32'h3a1ccc76),
	.w3(32'hba8d1b18),
	.w4(32'hbb198cab),
	.w5(32'h39dce565),
	.w6(32'hbb160d80),
	.w7(32'hba0419e5),
	.w8(32'h3a1914b6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b89b8),
	.w1(32'hbb19630a),
	.w2(32'hbad02d1e),
	.w3(32'hbae4023d),
	.w4(32'hb9e90863),
	.w5(32'hba95b604),
	.w6(32'hbacbadbc),
	.w7(32'hbaf06f73),
	.w8(32'h3b0e4293),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb627f),
	.w1(32'hb8f9724f),
	.w2(32'hb7095e66),
	.w3(32'h3b065913),
	.w4(32'h39dcd252),
	.w5(32'h39349489),
	.w6(32'h3955b35a),
	.w7(32'h39a581aa),
	.w8(32'hba70b900),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48471b),
	.w1(32'h3a3a55f9),
	.w2(32'hba9d2285),
	.w3(32'hbaafb5c9),
	.w4(32'hb9db0a61),
	.w5(32'hba2870f0),
	.w6(32'hba6c93c1),
	.w7(32'hbad141ea),
	.w8(32'h3a0ae972),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0a66a),
	.w1(32'h3a76d33f),
	.w2(32'h399d517b),
	.w3(32'hbae0bf13),
	.w4(32'hbacb5e25),
	.w5(32'h3a3125cf),
	.w6(32'hbb175650),
	.w7(32'h3765cc7e),
	.w8(32'hba54dfd8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9407c2),
	.w1(32'hba6c79db),
	.w2(32'hb9ab72f5),
	.w3(32'hba66532f),
	.w4(32'hba2635ff),
	.w5(32'hb962c493),
	.w6(32'hba168816),
	.w7(32'hb9f727e8),
	.w8(32'h39c18d04),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f70952),
	.w1(32'hb9bd2f0b),
	.w2(32'hb917f06e),
	.w3(32'h39f33719),
	.w4(32'h383cff58),
	.w5(32'hb984a835),
	.w6(32'h38dc4809),
	.w7(32'h3a0c2738),
	.w8(32'hbafa42e5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58fe66),
	.w1(32'hbb80b37f),
	.w2(32'hbb05d677),
	.w3(32'hbb434417),
	.w4(32'hbb88a981),
	.w5(32'hbb255e68),
	.w6(32'hba3337c4),
	.w7(32'hbaffcaf6),
	.w8(32'hb90d3be0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb57cd3d5),
	.w1(32'hb9a6a3fd),
	.w2(32'h3928b7c3),
	.w3(32'h39c201b4),
	.w4(32'hb93182a7),
	.w5(32'h38faa824),
	.w6(32'hb931d0ab),
	.w7(32'h39d93f7c),
	.w8(32'hb9e6e1cc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd21e9),
	.w1(32'hb9c3005f),
	.w2(32'hb94df0ab),
	.w3(32'hb9ced875),
	.w4(32'hb9d2ad4a),
	.w5(32'hb9b3b493),
	.w6(32'hb9f3f664),
	.w7(32'hb97655bc),
	.w8(32'hb962276c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0f8b4b),
	.w1(32'hba05d188),
	.w2(32'hba1a6ded),
	.w3(32'hb9fe7996),
	.w4(32'hb9ce1586),
	.w5(32'hba275d1e),
	.w6(32'hba11b25b),
	.w7(32'hb9b5e981),
	.w8(32'hba4d7832),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e74e6),
	.w1(32'hba670aca),
	.w2(32'hb8aa5d01),
	.w3(32'hba3917fc),
	.w4(32'hba4da27f),
	.w5(32'hb8f1d7bd),
	.w6(32'hba164648),
	.w7(32'hb9b21282),
	.w8(32'h390c8991),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a89be),
	.w1(32'hb85d9e50),
	.w2(32'h398b8029),
	.w3(32'h383fd974),
	.w4(32'h3930aaa7),
	.w5(32'h399b1205),
	.w6(32'hb891da85),
	.w7(32'h3925962c),
	.w8(32'h3b0bc6d1),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af0baa5),
	.w1(32'h3a3a2f0d),
	.w2(32'h3a9f21c6),
	.w3(32'h3b015513),
	.w4(32'h3a38344d),
	.w5(32'h3a36c6b6),
	.w6(32'h3a82e482),
	.w7(32'h3ac51a8d),
	.w8(32'hb904f47c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab7352),
	.w1(32'hb991566f),
	.w2(32'hb8c348de),
	.w3(32'h3778a166),
	.w4(32'h387b5014),
	.w5(32'hb93ca84e),
	.w6(32'hb988aa0d),
	.w7(32'h3937c52c),
	.w8(32'hb92a3efd),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d11a7),
	.w1(32'hb90a8ce6),
	.w2(32'h38663a69),
	.w3(32'hb88f91be),
	.w4(32'h39b58bd6),
	.w5(32'h39cdd0de),
	.w6(32'hb76ab95a),
	.w7(32'h39db29b3),
	.w8(32'hb9ff3641),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c0e11e),
	.w1(32'h38f67f0d),
	.w2(32'h38eceba8),
	.w3(32'h399a773f),
	.w4(32'h39bfc002),
	.w5(32'hb8585fe2),
	.w6(32'hb7b7de1e),
	.w7(32'h3949a4eb),
	.w8(32'hba9a9ac0),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c681c),
	.w1(32'hbb447f53),
	.w2(32'hbab59fe9),
	.w3(32'hbb5e473c),
	.w4(32'hbb37a2eb),
	.w5(32'hbb013431),
	.w6(32'h39a4d073),
	.w7(32'hb959c9ea),
	.w8(32'hba3540f3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2be5cb),
	.w1(32'hb9015b4f),
	.w2(32'hb98b419e),
	.w3(32'hb9b26c4e),
	.w4(32'h3931ec66),
	.w5(32'hb8b7bd81),
	.w6(32'h38a06ff6),
	.w7(32'hb883b8d7),
	.w8(32'hb9ba4411),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a78a3),
	.w1(32'hb9c98e20),
	.w2(32'hb84a3003),
	.w3(32'hb9b745ab),
	.w4(32'hb924f6b3),
	.w5(32'hb970f9a2),
	.w6(32'hba2805cd),
	.w7(32'hb8dc0101),
	.w8(32'hb9bbb715),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb960dada),
	.w1(32'hb9523a4c),
	.w2(32'hb910b0b3),
	.w3(32'h387250b5),
	.w4(32'h392636ce),
	.w5(32'hb64976ff),
	.w6(32'hb831ea96),
	.w7(32'h379e8935),
	.w8(32'h3b3701f8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b241c46),
	.w1(32'h3a2d4479),
	.w2(32'h3a886883),
	.w3(32'h3b2fe336),
	.w4(32'h3a42bfc8),
	.w5(32'h39e9e252),
	.w6(32'h3a896e6b),
	.w7(32'h3ac9cfe9),
	.w8(32'h3a86f998),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84a725),
	.w1(32'h398d2366),
	.w2(32'h3a2712ab),
	.w3(32'h3a5c3d80),
	.w4(32'h384a927c),
	.w5(32'h382a1b05),
	.w6(32'h3a2efa05),
	.w7(32'h3a97bbd5),
	.w8(32'hb927f4b2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9435cee),
	.w1(32'hba5f497c),
	.w2(32'hb8fe3cd3),
	.w3(32'h3811f663),
	.w4(32'hba24130b),
	.w5(32'hb88e906f),
	.w6(32'hba42da1b),
	.w7(32'hb9405848),
	.w8(32'hbaa39d25),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d47f3),
	.w1(32'hbb0f7a31),
	.w2(32'hbab66610),
	.w3(32'hba6142e8),
	.w4(32'hba832786),
	.w5(32'hba40539f),
	.w6(32'hbb051c41),
	.w7(32'hbaec4419),
	.w8(32'hba101d7d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39352d),
	.w1(32'hb9b65f09),
	.w2(32'hb9b5d4ff),
	.w3(32'hb987c9bc),
	.w4(32'hb7336dbb),
	.w5(32'hb92be8f4),
	.w6(32'hb9586d37),
	.w7(32'hb95526fa),
	.w8(32'hb9780864),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988a260),
	.w1(32'hb8c6a8fc),
	.w2(32'h37b40be8),
	.w3(32'h39f366c2),
	.w4(32'h39ddc439),
	.w5(32'h39dc5d6a),
	.w6(32'hb92b788b),
	.w7(32'h39d9071b),
	.w8(32'h39c83aba),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a1e67),
	.w1(32'h3aef7765),
	.w2(32'h3a7b9621),
	.w3(32'hb7c33228),
	.w4(32'hb9853df7),
	.w5(32'h39d6c8cf),
	.w6(32'hba04d037),
	.w7(32'hb9ff8624),
	.w8(32'h3900f846),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2a8f),
	.w1(32'hb95b9510),
	.w2(32'h39bcc647),
	.w3(32'hb94ec3b0),
	.w4(32'h38eac87a),
	.w5(32'h39e713cc),
	.w6(32'hb9aa46b4),
	.w7(32'h39ae931d),
	.w8(32'hb895d880),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9521e3d),
	.w1(32'hb9862149),
	.w2(32'h389feb69),
	.w3(32'h38e9f13c),
	.w4(32'h392d0e3f),
	.w5(32'h391d03cc),
	.w6(32'h39701a6d),
	.w7(32'h39aac695),
	.w8(32'h3aa38930),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a759fbb),
	.w1(32'hba5c834d),
	.w2(32'hba99b377),
	.w3(32'h3adad609),
	.w4(32'h39987022),
	.w5(32'hb731d134),
	.w6(32'hba034460),
	.w7(32'hba6f1496),
	.w8(32'hb8e6f9cd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38cc6c66),
	.w1(32'h399a3948),
	.w2(32'h39ba06d4),
	.w3(32'h3775250e),
	.w4(32'h399cb9c3),
	.w5(32'h39b8d807),
	.w6(32'h3817d025),
	.w7(32'h399eae02),
	.w8(32'hbab1ac28),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70ad2f),
	.w1(32'hba6b6030),
	.w2(32'hbaaddc3a),
	.w3(32'hbad481cc),
	.w4(32'hbac0caef),
	.w5(32'hbab3ffcf),
	.w6(32'hbaeaba56),
	.w7(32'hbb093c3b),
	.w8(32'h3ab5b73f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a554e89),
	.w1(32'hba51ca27),
	.w2(32'hba8a5f25),
	.w3(32'h3ac633c5),
	.w4(32'h39a44a55),
	.w5(32'h383f95dc),
	.w6(32'hba009359),
	.w7(32'hba5c8fd5),
	.w8(32'h3a88573c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2bd8c9),
	.w1(32'hba3061ea),
	.w2(32'hba79818b),
	.w3(32'h3aa87931),
	.w4(32'h39688abe),
	.w5(32'h33ff9a90),
	.w6(32'hb9ccbed7),
	.w7(32'hba2fa2ee),
	.w8(32'hba25ba51),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba108b76),
	.w1(32'hba4122df),
	.w2(32'hb9de04b7),
	.w3(32'hb9fa08d3),
	.w4(32'hba66d093),
	.w5(32'hb98b4893),
	.w6(32'hba81a051),
	.w7(32'hba5f1c51),
	.w8(32'hb952ce82),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba135478),
	.w1(32'hbb644f15),
	.w2(32'h3adbb03d),
	.w3(32'hb9fac0db),
	.w4(32'hbb930524),
	.w5(32'h3a8c1321),
	.w6(32'hbb25acae),
	.w7(32'h39e9836d),
	.w8(32'hb94049a2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c67455),
	.w1(32'h39b12d39),
	.w2(32'h39a2f7a2),
	.w3(32'h391f93c4),
	.w4(32'h397da3b9),
	.w5(32'hb7a8cc3c),
	.w6(32'h39c18477),
	.w7(32'h3a0ad446),
	.w8(32'hbb1c461c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba854aa2),
	.w1(32'hbabab214),
	.w2(32'hbab78971),
	.w3(32'hbb150bf5),
	.w4(32'hbaf46b26),
	.w5(32'hbb15c888),
	.w6(32'hbb115e4d),
	.w7(32'hbb21850a),
	.w8(32'hba72ab87),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabba31b),
	.w1(32'hbab16e63),
	.w2(32'hba5b34b3),
	.w3(32'hba80c1ee),
	.w4(32'hba8c92ec),
	.w5(32'hba2a92a4),
	.w6(32'hba84adff),
	.w7(32'hb9e551e2),
	.w8(32'h3912d8d6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba862a76),
	.w1(32'hbadabeed),
	.w2(32'hba6ecb30),
	.w3(32'hbaaa5dc3),
	.w4(32'hba1930f9),
	.w5(32'hb9bb18cb),
	.w6(32'hba8fcfe5),
	.w7(32'hba8fd6a1),
	.w8(32'hb98bfb7d),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26b171),
	.w1(32'h3978e7cd),
	.w2(32'h3a8c9db3),
	.w3(32'hbab7451d),
	.w4(32'hbaec8a72),
	.w5(32'h3a152f23),
	.w6(32'h37a78fe3),
	.w7(32'hbaab8c0d),
	.w8(32'h3b1d499f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15190c),
	.w1(32'h39f2577a),
	.w2(32'h3a552387),
	.w3(32'h3b195c23),
	.w4(32'h3a08c7c0),
	.w5(32'h399fb227),
	.w6(32'h3a718569),
	.w7(32'h3aa26580),
	.w8(32'h37fe089b),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39982e5a),
	.w1(32'h39dd661b),
	.w2(32'h3a25faab),
	.w3(32'h3a08a305),
	.w4(32'h39c228df),
	.w5(32'h3a171647),
	.w6(32'h38bf48b3),
	.w7(32'h39ea30bc),
	.w8(32'hbab9ec6c),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959933),
	.w1(32'hb9b1f2c9),
	.w2(32'hba67ec5d),
	.w3(32'hbab5454a),
	.w4(32'hba6e8f85),
	.w5(32'hb9217015),
	.w6(32'hbad37512),
	.w7(32'hbaa39569),
	.w8(32'hb98c3f0e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07d5c6),
	.w1(32'hba2620a2),
	.w2(32'hba719ce4),
	.w3(32'hb7b1f736),
	.w4(32'hb911af09),
	.w5(32'hba0f6f68),
	.w6(32'hb9d52da9),
	.w7(32'hb9610137),
	.w8(32'h3a814aed),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a50699a),
	.w1(32'hb98ef60c),
	.w2(32'h3a988e3a),
	.w3(32'h3a9c0188),
	.w4(32'h393599f9),
	.w5(32'h3a04d978),
	.w6(32'h39ec4a99),
	.w7(32'h3ac8254f),
	.w8(32'hba42124b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dfadf7),
	.w1(32'hb99d442e),
	.w2(32'hb9b34c29),
	.w3(32'hb95052de),
	.w4(32'hb9e70be0),
	.w5(32'hb943294d),
	.w6(32'hba617ddd),
	.w7(32'hba108e26),
	.w8(32'h39b60dcd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399643b0),
	.w1(32'hb98bd1f1),
	.w2(32'hb9c3f86c),
	.w3(32'h3a141859),
	.w4(32'h38f4f377),
	.w5(32'h3846ea58),
	.w6(32'hb94a0ec8),
	.w7(32'hb9afcd81),
	.w8(32'h38a5935e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95358b5),
	.w1(32'h3778d428),
	.w2(32'h39a555a5),
	.w3(32'h3934f3d5),
	.w4(32'h386c558d),
	.w5(32'h39a187df),
	.w6(32'h398a8db7),
	.w7(32'h39285e76),
	.w8(32'h3a1f774c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ae55f),
	.w1(32'hb95e3e29),
	.w2(32'hba14b341),
	.w3(32'h39ac2d10),
	.w4(32'h38109f02),
	.w5(32'hb983a1a8),
	.w6(32'h39179e6e),
	.w7(32'hb6c12c6a),
	.w8(32'hb8fdfc3c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86fd765),
	.w1(32'hb92ca9b3),
	.w2(32'hb98882b5),
	.w3(32'h3818e823),
	.w4(32'hb8d4046c),
	.w5(32'hb92f608b),
	.w6(32'hb61ca9b1),
	.w7(32'h389a5d5b),
	.w8(32'h35e217e4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc0e89),
	.w1(32'h399c51cb),
	.w2(32'h39b6bef4),
	.w3(32'h39308748),
	.w4(32'h399f37df),
	.w5(32'h39a3e163),
	.w6(32'h386408a8),
	.w7(32'h39889fed),
	.w8(32'h39929f6e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926a319),
	.w1(32'hb9ef88ad),
	.w2(32'hba0b5ced),
	.w3(32'hb8c8703b),
	.w4(32'hb99dbc22),
	.w5(32'hb9ea1b9f),
	.w6(32'hb921c9a4),
	.w7(32'hb98bdc8e),
	.w8(32'hb9a4c9d6),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942917f),
	.w1(32'hb8c20a12),
	.w2(32'hb9286ca5),
	.w3(32'hb896dbad),
	.w4(32'h38739ece),
	.w5(32'h3824d06c),
	.w6(32'hb97e9c65),
	.w7(32'hb868d557),
	.w8(32'h379fd86d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99e3ff1),
	.w1(32'hb716d31f),
	.w2(32'h39089893),
	.w3(32'hb95c3db6),
	.w4(32'h36bef994),
	.w5(32'h38e70e40),
	.w6(32'hb9367163),
	.w7(32'h38dd22be),
	.w8(32'h3932366c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3860ce46),
	.w1(32'h36b13ac9),
	.w2(32'h372ba5fe),
	.w3(32'h3856a383),
	.w4(32'h383c75f6),
	.w5(32'h388539a1),
	.w6(32'h37efab99),
	.w7(32'h38877e59),
	.w8(32'h3906ed6c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3839a84b),
	.w1(32'hb6f77456),
	.w2(32'h36b93780),
	.w3(32'h3847efe8),
	.w4(32'hb6897333),
	.w5(32'h36944403),
	.w6(32'h37f1f646),
	.w7(32'hb79ef11b),
	.w8(32'hb7ddda43),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376939ab),
	.w1(32'hb4aaab24),
	.w2(32'hb7a36359),
	.w3(32'h37cd5c0e),
	.w4(32'hb6263c36),
	.w5(32'hb7c1f92a),
	.w6(32'h38218168),
	.w7(32'hb70ce883),
	.w8(32'hb82a1130),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9674343),
	.w1(32'hb95cc554),
	.w2(32'hb8e7df2b),
	.w3(32'hb9725b06),
	.w4(32'hb9441801),
	.w5(32'hb9023795),
	.w6(32'hb9754fdf),
	.w7(32'hb9248514),
	.w8(32'hb801e93d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb875ae88),
	.w1(32'h390a896c),
	.w2(32'h3974de66),
	.w3(32'hb87c0d74),
	.w4(32'h3904088c),
	.w5(32'h39460ce6),
	.w6(32'h368dc01c),
	.w7(32'h3903a1a5),
	.w8(32'h3944dc73),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f112f5),
	.w1(32'h384e2c2a),
	.w2(32'h38b62d84),
	.w3(32'hb8e5c0d6),
	.w4(32'h37e933f5),
	.w5(32'h389a1a8b),
	.w6(32'hb8d325c2),
	.w7(32'h3827076e),
	.w8(32'h38af4e86),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3648431f),
	.w1(32'h34d49127),
	.w2(32'hb5291a0f),
	.w3(32'h365db641),
	.w4(32'h353dd344),
	.w5(32'hb44d0c90),
	.w6(32'h368c4df4),
	.w7(32'hb5305485),
	.w8(32'hb49af963),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7190c06),
	.w1(32'h36cae212),
	.w2(32'hb610e6b8),
	.w3(32'hb6ccf37c),
	.w4(32'h360d5406),
	.w5(32'hb6e04e60),
	.w6(32'h37538b78),
	.w7(32'h35aaed59),
	.w8(32'hb6bf1a63),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ac64e),
	.w1(32'hb919e9ef),
	.w2(32'hb8db1f5e),
	.w3(32'hb8aeffb7),
	.w4(32'h38698e3b),
	.w5(32'h38370cbf),
	.w6(32'hb945a55b),
	.w7(32'hb8f34a8c),
	.w8(32'hb86e3ace),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b113b2),
	.w1(32'hb971efa9),
	.w2(32'hb966d37e),
	.w3(32'h397762d6),
	.w4(32'hb8d1cf83),
	.w5(32'hb9209a5e),
	.w6(32'h39382617),
	.w7(32'hb8b859b0),
	.w8(32'hb87e25a9),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83002f8),
	.w1(32'hb85bc89d),
	.w2(32'hb70c36fd),
	.w3(32'hb849a7a4),
	.w4(32'hb7f94a81),
	.w5(32'hb8209a93),
	.w6(32'hb8a2e37b),
	.w7(32'hb8b24059),
	.w8(32'hb78c0652),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb896589b),
	.w1(32'hb83f7172),
	.w2(32'h38b510ae),
	.w3(32'hb9402cfa),
	.w4(32'hb8bace56),
	.w5(32'h38db9fa6),
	.w6(32'hb94880cd),
	.w7(32'hb89c817d),
	.w8(32'h38f448eb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e4a92b),
	.w1(32'hb97329b1),
	.w2(32'hba05e0b0),
	.w3(32'hb94b45b7),
	.w4(32'hb9d0eeef),
	.w5(32'hb9feb3dc),
	.w6(32'hb9b077e3),
	.w7(32'hb9dcf2f5),
	.w8(32'hb9e40c13),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93275c3),
	.w1(32'hb8e02183),
	.w2(32'hb8da1837),
	.w3(32'hb9368f31),
	.w4(32'hb8d418da),
	.w5(32'hb8a8741d),
	.w6(32'hb92e46cf),
	.w7(32'hb9046e19),
	.w8(32'hb8ac9739),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c5e77),
	.w1(32'hb9b7df06),
	.w2(32'hb9737689),
	.w3(32'hb90fb7da),
	.w4(32'hb94c4cb0),
	.w5(32'hb8a6a232),
	.w6(32'hb97e0359),
	.w7(32'hb930ee0c),
	.w8(32'h36cd1326),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6681ccc),
	.w1(32'h38a043bc),
	.w2(32'h38e86beb),
	.w3(32'h3912c458),
	.w4(32'h3791c84b),
	.w5(32'h3896d239),
	.w6(32'h392f8441),
	.w7(32'h375d70de),
	.w8(32'h391b00ab),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule