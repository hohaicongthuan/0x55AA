module layer_10_featuremap_310(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c480f),
	.w1(32'hbb29f461),
	.w2(32'h3b6373df),
	.w3(32'hb9d6bc50),
	.w4(32'h3b0fa18d),
	.w5(32'hba14829d),
	.w6(32'h3aa00018),
	.w7(32'h3bb93079),
	.w8(32'h3adcf2c0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0a10a),
	.w1(32'h3af8e7af),
	.w2(32'h3b306c32),
	.w3(32'h3a275470),
	.w4(32'h39d37234),
	.w5(32'h3b212580),
	.w6(32'h3c09c0d5),
	.w7(32'h3b230a35),
	.w8(32'hbb01f2c5),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9806aa),
	.w1(32'h3a621cfa),
	.w2(32'h3b3fe30f),
	.w3(32'hba718de7),
	.w4(32'hba44be0d),
	.w5(32'hba9916cd),
	.w6(32'hbaef171c),
	.w7(32'hb7e01c77),
	.w8(32'hbb6fc078),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e6d15),
	.w1(32'hbb7ab077),
	.w2(32'hbb809790),
	.w3(32'hbb266c92),
	.w4(32'hbb7287a1),
	.w5(32'hbb5fdbdb),
	.w6(32'hbbcbd211),
	.w7(32'hbbc7ab22),
	.w8(32'hbbec2319),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8218b0),
	.w1(32'hbb8e1804),
	.w2(32'hbb73193f),
	.w3(32'hbb42ad51),
	.w4(32'hbb6669df),
	.w5(32'h3a7aa421),
	.w6(32'hbc09652d),
	.w7(32'hbbbff36d),
	.w8(32'h3a73de16),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d12ef4),
	.w1(32'h3a96dd1e),
	.w2(32'h3ba2c17b),
	.w3(32'h3a203a77),
	.w4(32'h3b81ea21),
	.w5(32'hb9723224),
	.w6(32'h3a93de73),
	.w7(32'h3bb4e552),
	.w8(32'hba4216d2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a2a17),
	.w1(32'h39e7b9e2),
	.w2(32'h3b174d1b),
	.w3(32'h3aadc54d),
	.w4(32'h3b259b4e),
	.w5(32'hbaa00e72),
	.w6(32'h3a0eb1fc),
	.w7(32'h392d8c5c),
	.w8(32'hbb9df13a),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9842a2),
	.w1(32'hbb6f2073),
	.w2(32'hbb03409f),
	.w3(32'hbadc9e34),
	.w4(32'hbb036a97),
	.w5(32'hb9b29dd9),
	.w6(32'hbbbcdd5b),
	.w7(32'hbbd054c3),
	.w8(32'h39fdc3c0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398dac92),
	.w1(32'h3abb4cf9),
	.w2(32'h3b35f515),
	.w3(32'h39d62c82),
	.w4(32'h3b198137),
	.w5(32'hb97c9a43),
	.w6(32'h3a881a99),
	.w7(32'h3b5a6907),
	.w8(32'hba5758c2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb5f23),
	.w1(32'hba5599b1),
	.w2(32'h3b62a503),
	.w3(32'hb5d98e53),
	.w4(32'h3b40da87),
	.w5(32'h39623d1d),
	.w6(32'hba591775),
	.w7(32'h3b8e9d92),
	.w8(32'h3a145774),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9797e),
	.w1(32'hb8a67c49),
	.w2(32'h3b4eb4e0),
	.w3(32'hba8fba42),
	.w4(32'h39865bde),
	.w5(32'h3b9d669f),
	.w6(32'h394e4d70),
	.w7(32'h3b1ef57f),
	.w8(32'h3afe473b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aee57),
	.w1(32'h3bc85810),
	.w2(32'h3bae9d6c),
	.w3(32'h3b3cdec2),
	.w4(32'h3aa70f52),
	.w5(32'hbaf4ec78),
	.w6(32'h3b8e92fa),
	.w7(32'h3b5e887d),
	.w8(32'hb9c60b39),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53a3bb),
	.w1(32'h3846cceb),
	.w2(32'h37c8e09d),
	.w3(32'hbaf7b01c),
	.w4(32'h3a1cda85),
	.w5(32'hba99be7b),
	.w6(32'h3ae82910),
	.w7(32'hb9b20d24),
	.w8(32'hbaa9060b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74d40e),
	.w1(32'h39960a31),
	.w2(32'hbaa491ec),
	.w3(32'hba881b8f),
	.w4(32'h3936a28f),
	.w5(32'h3bcac52c),
	.w6(32'hba835c15),
	.w7(32'hbaa1c7bb),
	.w8(32'h3b9d91bf),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a0efe),
	.w1(32'h3aa5546c),
	.w2(32'h3a646c6a),
	.w3(32'h3ba23396),
	.w4(32'h3b5a532b),
	.w5(32'hbbd3aec9),
	.w6(32'h3b41c272),
	.w7(32'h3ac9de9f),
	.w8(32'hbbd294f4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d91b7),
	.w1(32'hbb9c0e43),
	.w2(32'hba374c8f),
	.w3(32'hbba3fce6),
	.w4(32'hbb37c7ff),
	.w5(32'h3bffa1e2),
	.w6(32'hbb01351d),
	.w7(32'h3aacec1e),
	.w8(32'h3ba74579),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bed99),
	.w1(32'h3bfe377f),
	.w2(32'h3c3d3d4a),
	.w3(32'h3b9767ad),
	.w4(32'h3c1f7185),
	.w5(32'hba598bcb),
	.w6(32'h3bd8e513),
	.w7(32'h3c1119fe),
	.w8(32'hbab50230),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad04287),
	.w1(32'hbb0ba37a),
	.w2(32'hbb162ba0),
	.w3(32'hbb1bf5b4),
	.w4(32'hbb0a8b99),
	.w5(32'hbb261fe0),
	.w6(32'hbb0c0a25),
	.w7(32'hbb3a6ee3),
	.w8(32'hb9aa730a),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1ad07),
	.w1(32'hbb65bbdd),
	.w2(32'hba0281c3),
	.w3(32'hbae28083),
	.w4(32'hbab4ce8c),
	.w5(32'hbbd1b6d5),
	.w6(32'hbae03e37),
	.w7(32'hbaa07209),
	.w8(32'hbb9c7dc9),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79ca93),
	.w1(32'hbb5324d4),
	.w2(32'hbbe2008d),
	.w3(32'hbbaf90f4),
	.w4(32'hbaec71d6),
	.w5(32'hbb4111bc),
	.w6(32'hbb9f305a),
	.w7(32'hbb992687),
	.w8(32'hbb2ea22a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e2414),
	.w1(32'hbb13c7b8),
	.w2(32'hbb2ed093),
	.w3(32'hbafb2c04),
	.w4(32'hbb45edcc),
	.w5(32'h3ba87c9f),
	.w6(32'hbb36990b),
	.w7(32'hbac57d8d),
	.w8(32'h3b17f8dd),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35e1de),
	.w1(32'h3aa6809d),
	.w2(32'h3a6be304),
	.w3(32'h3b91c5b9),
	.w4(32'h3b683083),
	.w5(32'hbb502f6c),
	.w6(32'hb9cd15cb),
	.w7(32'hba7056f3),
	.w8(32'hbb41ed7b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6198),
	.w1(32'hbb17ac0d),
	.w2(32'hbb1b094e),
	.w3(32'hbb5c39b1),
	.w4(32'hbb66c196),
	.w5(32'hbb5764de),
	.w6(32'hbb04e4d5),
	.w7(32'hbb1c8f25),
	.w8(32'hbb326956),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833365),
	.w1(32'hb9ad1081),
	.w2(32'h39a20852),
	.w3(32'hbb23c8d2),
	.w4(32'hbba013fa),
	.w5(32'h3aee3805),
	.w6(32'hbb239eec),
	.w7(32'hb9591fe2),
	.w8(32'hbab66990),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1528d1),
	.w1(32'h3a8ce7a0),
	.w2(32'h3b13d720),
	.w3(32'h3ad606bd),
	.w4(32'h3a55e332),
	.w5(32'h3b8f35dc),
	.w6(32'hb86a9601),
	.w7(32'h39eab76b),
	.w8(32'h3b2e1c6d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a33f5c4),
	.w1(32'hba6f4655),
	.w2(32'h3b0bf0d1),
	.w3(32'h3b88eafa),
	.w4(32'h3bc853a5),
	.w5(32'h3b910973),
	.w6(32'h3a7e06c7),
	.w7(32'h3b8014dc),
	.w8(32'h3b435ba1),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816578),
	.w1(32'h3b3188d4),
	.w2(32'h3bd6c791),
	.w3(32'h3b660e8a),
	.w4(32'h3c059b26),
	.w5(32'hbaa9dddd),
	.w6(32'h3a91fa31),
	.w7(32'h3bbb4f91),
	.w8(32'hba4e3fad),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a0b24),
	.w1(32'h3b514aea),
	.w2(32'h3c0980ee),
	.w3(32'h3aecfc08),
	.w4(32'h3bcc7a83),
	.w5(32'hb9ca1908),
	.w6(32'h3bb8d762),
	.w7(32'h3c3fba0e),
	.w8(32'hbab62949),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ce8ed),
	.w1(32'hba7abf86),
	.w2(32'hbb75ca5e),
	.w3(32'hb922f729),
	.w4(32'h3a9d6a67),
	.w5(32'h395db93f),
	.w6(32'hbb354803),
	.w7(32'hba67d73d),
	.w8(32'h3a57dd69),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1d3ae),
	.w1(32'h3ac60230),
	.w2(32'hbb1cc718),
	.w3(32'h3a11d127),
	.w4(32'h3ae90c59),
	.w5(32'hbadb3057),
	.w6(32'hba99952f),
	.w7(32'hba84cccc),
	.w8(32'h3b5ff123),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0f449),
	.w1(32'h3a7ad332),
	.w2(32'hbaa326df),
	.w3(32'h3ac8da4b),
	.w4(32'hbaf397e2),
	.w5(32'h3adb92df),
	.w6(32'h3bc08051),
	.w7(32'h3b75798a),
	.w8(32'h3b08c07e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc38afd),
	.w1(32'h3c40ce2d),
	.w2(32'h3c09d2e4),
	.w3(32'h3bcff64a),
	.w4(32'h3bc73e87),
	.w5(32'h3a6cf4f7),
	.w6(32'h3b213b07),
	.w7(32'hb9bea5e6),
	.w8(32'h3b8a1455),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba320086),
	.w1(32'h3aa254d7),
	.w2(32'h3a565f1f),
	.w3(32'h3bd10df7),
	.w4(32'h3b7b6006),
	.w5(32'hbaec3246),
	.w6(32'h3ba943b2),
	.w7(32'h3b9dd603),
	.w8(32'hbb92aa35),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65f1ef),
	.w1(32'hbb81b8de),
	.w2(32'hbb252e68),
	.w3(32'hbb5ec543),
	.w4(32'hbb5bc944),
	.w5(32'hbb1d0948),
	.w6(32'hbb4d0ec1),
	.w7(32'hbb7b45e4),
	.w8(32'hbb57841e),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cf1f70),
	.w1(32'hb9f7cc35),
	.w2(32'hba1e8f26),
	.w3(32'hba8df05a),
	.w4(32'h3aac75d5),
	.w5(32'hbb2e9e4f),
	.w6(32'hbafefc02),
	.w7(32'hba7fb2d4),
	.w8(32'hbaff9c74),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1bee1a),
	.w1(32'hbb296d89),
	.w2(32'h3a89afef),
	.w3(32'hbb85c8de),
	.w4(32'hbb828c2e),
	.w5(32'h3976e6a8),
	.w6(32'hba951aeb),
	.w7(32'hb969c3f1),
	.w8(32'h3bd9cec4),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b554f8c),
	.w1(32'h3b25207a),
	.w2(32'h3a5d090c),
	.w3(32'h3b97c104),
	.w4(32'h3b8e6c5d),
	.w5(32'h3b4b4b90),
	.w6(32'h3c3e181e),
	.w7(32'h3c0c33c6),
	.w8(32'h3b911cc7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a1df2),
	.w1(32'h3b4bf8d5),
	.w2(32'h3c1ce20a),
	.w3(32'h3b0103c0),
	.w4(32'h3bf8b10c),
	.w5(32'hbbb29714),
	.w6(32'h3aaa3101),
	.w7(32'h3c126f1d),
	.w8(32'hbac87dde),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40f190),
	.w1(32'hbb6b19e0),
	.w2(32'hbaabf9b1),
	.w3(32'hbbbc2258),
	.w4(32'hbbc4ef1c),
	.w5(32'h3c1bc16a),
	.w6(32'hbaab822d),
	.w7(32'h378a6b33),
	.w8(32'h3b9b6d79),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3b080),
	.w1(32'h3b95e9df),
	.w2(32'h3ade48f1),
	.w3(32'h3c0aec07),
	.w4(32'h3ba1fb99),
	.w5(32'hbad7d71e),
	.w6(32'h3b0746da),
	.w7(32'h3abed19e),
	.w8(32'hbad5c309),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4835d0),
	.w1(32'hbb7c4708),
	.w2(32'hbb4ba577),
	.w3(32'hbb203164),
	.w4(32'hbb3402ea),
	.w5(32'h3ad34681),
	.w6(32'hbb43d79c),
	.w7(32'hba8920ee),
	.w8(32'hbb07bd23),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd5fc3),
	.w1(32'hbb2b6b98),
	.w2(32'h3a97df2b),
	.w3(32'h39908551),
	.w4(32'h3b75364e),
	.w5(32'hbb5487ce),
	.w6(32'hbbe6b33a),
	.w7(32'hbaa99932),
	.w8(32'hbac70308),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b724),
	.w1(32'hbbcc7bcf),
	.w2(32'hbb5092f4),
	.w3(32'hbb48b8f1),
	.w4(32'hba85b50a),
	.w5(32'hba6dd2bc),
	.w6(32'hbbb546a9),
	.w7(32'hbaa1c684),
	.w8(32'hba3fca60),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12ac16),
	.w1(32'h3ac3a1e5),
	.w2(32'h3baff808),
	.w3(32'hbb526617),
	.w4(32'h3b0a2f40),
	.w5(32'hbb2f07d5),
	.w6(32'h3b39c8f1),
	.w7(32'h3b7920cd),
	.w8(32'hbb80db2e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf2e976),
	.w1(32'hbc095604),
	.w2(32'hbbfb4a4d),
	.w3(32'hbafb6ded),
	.w4(32'hbafd9c24),
	.w5(32'h3b328b77),
	.w6(32'hbbb572d5),
	.w7(32'hbb6c4bc5),
	.w8(32'h3a89c4f2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b218d1f),
	.w1(32'h3a8151bb),
	.w2(32'h3a9fed44),
	.w3(32'h3b1c3695),
	.w4(32'h3b5b3b59),
	.w5(32'h394a35f1),
	.w6(32'h3ac2fbcd),
	.w7(32'h3b3f043b),
	.w8(32'hbb894b34),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb374e01),
	.w1(32'hbbad008f),
	.w2(32'hbb0a57a1),
	.w3(32'hbae070af),
	.w4(32'h39c39c50),
	.w5(32'h3b46fa16),
	.w6(32'hbba3eeb1),
	.w7(32'hba9a96fc),
	.w8(32'h3af24486),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5621a2),
	.w1(32'h3b1c128c),
	.w2(32'h3af33aaa),
	.w3(32'h3b0ec2e5),
	.w4(32'h3b31d5c5),
	.w5(32'hb8fbda9b),
	.w6(32'hb8831bf2),
	.w7(32'h3b1be373),
	.w8(32'h3b501422),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa98541),
	.w1(32'h3b04eaac),
	.w2(32'h3ac8756a),
	.w3(32'h39053187),
	.w4(32'h3b09c01a),
	.w5(32'h3a81229c),
	.w6(32'h3b95bec5),
	.w7(32'h3bb1300a),
	.w8(32'hbacc4f3d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09465c),
	.w1(32'hb9f7f3fb),
	.w2(32'h3a1668fa),
	.w3(32'h3a96658d),
	.w4(32'h3af2407a),
	.w5(32'hbb1f3356),
	.w6(32'hbb6f23ca),
	.w7(32'hbb33db4e),
	.w8(32'hbb65a22b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd38532),
	.w1(32'hba14f425),
	.w2(32'hbb045567),
	.w3(32'hb948b4a5),
	.w4(32'hba8341ab),
	.w5(32'h39b1fbba),
	.w6(32'h3abb669e),
	.w7(32'hbb1f9465),
	.w8(32'hba891b9c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc6694),
	.w1(32'h3a74f056),
	.w2(32'hb8bbc860),
	.w3(32'hbadc7909),
	.w4(32'hbaa980b5),
	.w5(32'h39bbcbd7),
	.w6(32'hba93f080),
	.w7(32'hbb836c74),
	.w8(32'hb9cb234f),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3788d),
	.w1(32'hbbdb5c1d),
	.w2(32'hb83abaea),
	.w3(32'hbadb316b),
	.w4(32'hbb11dc9c),
	.w5(32'h3c301239),
	.w6(32'hbb57d1b4),
	.w7(32'hb9b89a58),
	.w8(32'h3bd8eb31),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c062504),
	.w1(32'h3b921ee2),
	.w2(32'hba11ba1f),
	.w3(32'h3bd86a2a),
	.w4(32'h3b90726e),
	.w5(32'hbb94c027),
	.w6(32'h3b24aab6),
	.w7(32'h3b2a39a5),
	.w8(32'hba745b0f),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68200e),
	.w1(32'hb99ea405),
	.w2(32'hbb125357),
	.w3(32'hbb757f36),
	.w4(32'hba38e3ec),
	.w5(32'hbb76b7ae),
	.w6(32'hbacad823),
	.w7(32'hbb072c1a),
	.w8(32'hbb8b5038),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb434e80),
	.w1(32'hb8f6b5bf),
	.w2(32'hb931168f),
	.w3(32'hba72380c),
	.w4(32'h3aa84830),
	.w5(32'hba17d9ec),
	.w6(32'hbab2c3be),
	.w7(32'h3a90dcc2),
	.w8(32'hba571ae4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f7a5c),
	.w1(32'h3abf6b57),
	.w2(32'hb9f96317),
	.w3(32'h39a5b91c),
	.w4(32'hba12bd7f),
	.w5(32'hb9bf4f55),
	.w6(32'h3938fdf3),
	.w7(32'h3a861247),
	.w8(32'hbae9ee60),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f5206),
	.w1(32'hbb6f2b7b),
	.w2(32'hbb8fcbfa),
	.w3(32'hb98d7cc2),
	.w4(32'hbadad043),
	.w5(32'h3a78c01d),
	.w6(32'hbad152fb),
	.w7(32'hba9d88da),
	.w8(32'hba96b26b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a48f822),
	.w1(32'h3a3de6e5),
	.w2(32'h3af21f3f),
	.w3(32'h3aeda043),
	.w4(32'h3b431b23),
	.w5(32'h3a678b61),
	.w6(32'hbb1f3e01),
	.w7(32'hba643e80),
	.w8(32'hba49f679),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d63de),
	.w1(32'hb67e38d6),
	.w2(32'h3a78905e),
	.w3(32'hba3eb854),
	.w4(32'hb98b7fac),
	.w5(32'hbb44cfff),
	.w6(32'hba5e5a82),
	.w7(32'hba8f3eb8),
	.w8(32'hbb02afc8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac73798),
	.w1(32'hbaa7a04e),
	.w2(32'hba9a38b8),
	.w3(32'hbaf0aa8e),
	.w4(32'hba914129),
	.w5(32'hbb8ec3f2),
	.w6(32'hba54e867),
	.w7(32'hb8fde20c),
	.w8(32'hbb2e6629),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbace39e),
	.w1(32'hbb8acd71),
	.w2(32'hbb3af772),
	.w3(32'hbb58c8c0),
	.w4(32'hba98b88e),
	.w5(32'h3a1a0871),
	.w6(32'h3b26ffa1),
	.w7(32'h39f3428a),
	.w8(32'hbac183e7),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c9c9c),
	.w1(32'hb918b62d),
	.w2(32'h3b15d298),
	.w3(32'h3a63c1b7),
	.w4(32'h3ae961bb),
	.w5(32'hbb1cd591),
	.w6(32'hbb14c212),
	.w7(32'hb92dc932),
	.w8(32'hbb25debc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5cb556),
	.w1(32'hbab4e076),
	.w2(32'h3992fd42),
	.w3(32'hb911b54e),
	.w4(32'h3b1603f6),
	.w5(32'hbbfa7077),
	.w6(32'hbab2e96b),
	.w7(32'h3a8ce196),
	.w8(32'hbba34988),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05cadd),
	.w1(32'hba87aa86),
	.w2(32'hbb60351f),
	.w3(32'hbb38c284),
	.w4(32'h3a94acbf),
	.w5(32'hbbcde1cc),
	.w6(32'hbb5c6606),
	.w7(32'hb9bd3f09),
	.w8(32'hbb4fbd24),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73e3c5),
	.w1(32'hbb301cc2),
	.w2(32'h3a5bea04),
	.w3(32'hbb9b5872),
	.w4(32'hbb8e5da4),
	.w5(32'hba0a59fb),
	.w6(32'hbb270eb1),
	.w7(32'h39fa0973),
	.w8(32'hbaef7c97),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810da9),
	.w1(32'hbbc0ede6),
	.w2(32'hbbb5d112),
	.w3(32'hbb000134),
	.w4(32'hbaac9172),
	.w5(32'hba4ec63f),
	.w6(32'hba909d5e),
	.w7(32'hbafa2ec2),
	.w8(32'h3b664e60),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f6566),
	.w1(32'hba7a8784),
	.w2(32'hb98eb5e0),
	.w3(32'hbae515cc),
	.w4(32'h3b49c57a),
	.w5(32'hbbaa54fb),
	.w6(32'h3ab58486),
	.w7(32'h3ae402fc),
	.w8(32'hbb873880),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb843190),
	.w1(32'hb9d8dae6),
	.w2(32'hbb6cafb6),
	.w3(32'hb9cf6ac6),
	.w4(32'h38af67c6),
	.w5(32'hba8c6cd9),
	.w6(32'hbb348a59),
	.w7(32'hbb7767bc),
	.w8(32'hbb8f821a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb408cd4),
	.w1(32'hbbcd2170),
	.w2(32'hba91068a),
	.w3(32'hbbbf6136),
	.w4(32'hbb068912),
	.w5(32'h3a34c6a9),
	.w6(32'hbb986940),
	.w7(32'hbb9e3d09),
	.w8(32'h3a7b99ae),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb073236),
	.w1(32'hbb98891b),
	.w2(32'hbaed1c87),
	.w3(32'h3a7152c9),
	.w4(32'h3a8616fe),
	.w5(32'h3b6b1efd),
	.w6(32'hba812fa3),
	.w7(32'h3a3e7d7e),
	.w8(32'h3ba2cd55),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b532ab4),
	.w1(32'h3a9695dc),
	.w2(32'h3bbbee1a),
	.w3(32'h3b9ff90e),
	.w4(32'h3afec71b),
	.w5(32'hbb4ff509),
	.w6(32'h3bf1ec5a),
	.w7(32'h3b899751),
	.w8(32'h3b732fba),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6b8ea),
	.w1(32'hba28577a),
	.w2(32'h3b94b107),
	.w3(32'hbbb04d4a),
	.w4(32'hbb1d3db7),
	.w5(32'h39ba45a1),
	.w6(32'h3be3bde8),
	.w7(32'h3b986d89),
	.w8(32'h3a2eb3af),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06df61),
	.w1(32'h39af38c1),
	.w2(32'hb9d13b55),
	.w3(32'h3a1f48ed),
	.w4(32'hb9c4caab),
	.w5(32'h3b2a0ecd),
	.w6(32'h3b41092a),
	.w7(32'h3a3a9d2c),
	.w8(32'h3b7812d8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bf64c),
	.w1(32'hba69b94f),
	.w2(32'h3b0cf97d),
	.w3(32'h38d7b864),
	.w4(32'h3a8a80a3),
	.w5(32'h3aca05b3),
	.w6(32'h3b91ac96),
	.w7(32'h3bd7b535),
	.w8(32'h3a643eba),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac45a15),
	.w1(32'h3b1b9796),
	.w2(32'h3b0bd8d1),
	.w3(32'h3a20c86a),
	.w4(32'h39c96786),
	.w5(32'hbb8951d6),
	.w6(32'h3aa2ae31),
	.w7(32'h3a37c264),
	.w8(32'hbb0cc9b0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f4e5),
	.w1(32'hbb713252),
	.w2(32'hb9e2e984),
	.w3(32'hbb113073),
	.w4(32'hbabb0b11),
	.w5(32'hbb65e362),
	.w6(32'hba244e04),
	.w7(32'h39e5e812),
	.w8(32'hbbba2657),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8fb9ce),
	.w1(32'hbb872c0d),
	.w2(32'hbad95ee1),
	.w3(32'hbba0f68c),
	.w4(32'hbb4d4695),
	.w5(32'h3a9fa350),
	.w6(32'hbbbb8fcf),
	.w7(32'hbb866a1c),
	.w8(32'h3aed811c),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a369688),
	.w1(32'hb9c18f2b),
	.w2(32'h3a0b8e1b),
	.w3(32'h3a3220fc),
	.w4(32'hba986412),
	.w5(32'h3a7df81c),
	.w6(32'h3b08999d),
	.w7(32'h38ac2b0e),
	.w8(32'h3a687883),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a938d55),
	.w1(32'hb9bddfbd),
	.w2(32'h3ab0efc5),
	.w3(32'h3a5542e9),
	.w4(32'h3b654fb1),
	.w5(32'h3b848895),
	.w6(32'h3b4df99d),
	.w7(32'h3b98b6f7),
	.w8(32'hba6a82a4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe24e5),
	.w1(32'hba534d2d),
	.w2(32'hbb3cd577),
	.w3(32'h3bb6f455),
	.w4(32'h3a1af5ef),
	.w5(32'hbab4404c),
	.w6(32'hbb0c8fec),
	.w7(32'hbb8b1e52),
	.w8(32'hba4a0cf1),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3269a),
	.w1(32'hbb0bba7f),
	.w2(32'hbac1bd45),
	.w3(32'hbb3910a2),
	.w4(32'hbb6dd9cd),
	.w5(32'hbb9f8cf9),
	.w6(32'hbb0915e5),
	.w7(32'hbaed17b2),
	.w8(32'hbbab5521),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c7d4),
	.w1(32'hbae71e8d),
	.w2(32'hbae0418a),
	.w3(32'hba990063),
	.w4(32'hbb074646),
	.w5(32'h3bddbf29),
	.w6(32'hbab010c8),
	.w7(32'hbb12c6dd),
	.w8(32'h3c2d251e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d7186),
	.w1(32'h3bc9d9a6),
	.w2(32'h3b9d8695),
	.w3(32'h3b57df00),
	.w4(32'h3b7a85b3),
	.w5(32'hbb439cd5),
	.w6(32'h3b59235f),
	.w7(32'h3b9b4176),
	.w8(32'hbb4cb21b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c71bf),
	.w1(32'hbad5b3ce),
	.w2(32'hbae2304f),
	.w3(32'hbb5881a4),
	.w4(32'hbb0d86b2),
	.w5(32'hbbcb9f7b),
	.w6(32'hbab38826),
	.w7(32'hbaa6f2e9),
	.w8(32'hbb642796),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb465f),
	.w1(32'hbb289263),
	.w2(32'hbafaa29e),
	.w3(32'hbb8c4c2f),
	.w4(32'hbba04bd8),
	.w5(32'h3b759a3b),
	.w6(32'h3a6baf75),
	.w7(32'hb946643d),
	.w8(32'hb9a1a20a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a2864),
	.w1(32'h3b3c8a63),
	.w2(32'h3b846a17),
	.w3(32'h398b5ad0),
	.w4(32'h3b28f299),
	.w5(32'hbb91ad9d),
	.w6(32'hb99047b4),
	.w7(32'h3b6c6db5),
	.w8(32'hbb2dd26e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39a132),
	.w1(32'hbb2c2e19),
	.w2(32'hbb4812a1),
	.w3(32'hbb80f737),
	.w4(32'hbacec737),
	.w5(32'h3b4c811d),
	.w6(32'hbb46f5f7),
	.w7(32'hbab4c9cf),
	.w8(32'h3b17752f),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4431f6),
	.w1(32'h3b440b4d),
	.w2(32'h3bb51c4b),
	.w3(32'h3b917782),
	.w4(32'h3be49f61),
	.w5(32'hbb8986cd),
	.w6(32'h3b5ca87f),
	.w7(32'h3b94a52c),
	.w8(32'hbb1d2daa),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb399075),
	.w1(32'hb9b0515e),
	.w2(32'hbb688124),
	.w3(32'hbb12a218),
	.w4(32'hba52aaa3),
	.w5(32'h3ad31d77),
	.w6(32'hb9960020),
	.w7(32'hba96c690),
	.w8(32'h3b3637d4),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a965c),
	.w1(32'h3b152f71),
	.w2(32'h39c2ffc6),
	.w3(32'h3aabee6c),
	.w4(32'h3a193a18),
	.w5(32'hb999d8be),
	.w6(32'h3b592e3a),
	.w7(32'h3a8a4c1f),
	.w8(32'hb9139b29),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0bab9),
	.w1(32'h3a06ad87),
	.w2(32'hbb0ad298),
	.w3(32'h3b2549f4),
	.w4(32'h3a611c6c),
	.w5(32'hbb03d8b1),
	.w6(32'hba207944),
	.w7(32'hbb01f75b),
	.w8(32'h3b1a984f),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf789e),
	.w1(32'h3c0acab9),
	.w2(32'h3c0ad4fb),
	.w3(32'h3aae47d5),
	.w4(32'h3bb73fb9),
	.w5(32'hbb6d3ce9),
	.w6(32'h3b8886bb),
	.w7(32'h3b03df8f),
	.w8(32'hbb7e22ec),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973ba0),
	.w1(32'hba76bfff),
	.w2(32'h3934ea47),
	.w3(32'hbaca5d3e),
	.w4(32'hb98a97da),
	.w5(32'hba4c18a5),
	.w6(32'hbae6dba9),
	.w7(32'hba87fa7a),
	.w8(32'h3a89b0cd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac294d0),
	.w1(32'hbab4709c),
	.w2(32'h3b1671b1),
	.w3(32'hba097f55),
	.w4(32'h39a93d38),
	.w5(32'hbb033e92),
	.w6(32'hba8858eb),
	.w7(32'h3b5ab0c6),
	.w8(32'hba96c06a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526413),
	.w1(32'h3b704a46),
	.w2(32'h3bd431dc),
	.w3(32'hbb103e61),
	.w4(32'h3a747c62),
	.w5(32'hb9e0410b),
	.w6(32'hbb7a6ba7),
	.w7(32'h39ab6e71),
	.w8(32'h3aa143ec),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a8e958),
	.w1(32'h3ad6947a),
	.w2(32'hbb3d2793),
	.w3(32'h3a40981d),
	.w4(32'hbba51b44),
	.w5(32'h3ac9e546),
	.w6(32'h3b04c5de),
	.w7(32'hbb6454eb),
	.w8(32'h3acc5dec),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97cf49),
	.w1(32'h3bb1d79f),
	.w2(32'h3bcd3741),
	.w3(32'h3bfd2204),
	.w4(32'h3bfd28a2),
	.w5(32'h3b8c017f),
	.w6(32'h3b7e62c2),
	.w7(32'h3c288bea),
	.w8(32'h3b9ea927),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1db915),
	.w1(32'h3ae1771b),
	.w2(32'h3aa11d64),
	.w3(32'h3ad14070),
	.w4(32'h3a6967d6),
	.w5(32'hba4bbec3),
	.w6(32'h3b807512),
	.w7(32'h3b0b87f2),
	.w8(32'hbb8e7c0a),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8bbbd),
	.w1(32'hbb3e3046),
	.w2(32'hbb33710b),
	.w3(32'hbb4e2dca),
	.w4(32'hbb058a82),
	.w5(32'hbb6d698b),
	.w6(32'h38ae2e2b),
	.w7(32'hbba1beff),
	.w8(32'hbb1bc696),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1a0e2),
	.w1(32'hbb92d585),
	.w2(32'hbb032694),
	.w3(32'hbbab2a58),
	.w4(32'hbafcdd26),
	.w5(32'h3a31b559),
	.w6(32'h381eb087),
	.w7(32'h37a07e10),
	.w8(32'hbaa736c5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba137c6b),
	.w1(32'h398b2ab2),
	.w2(32'hbab97294),
	.w3(32'h3a3ca6c6),
	.w4(32'hba7d1d1d),
	.w5(32'h3b98d55f),
	.w6(32'hb89a6d2d),
	.w7(32'hbb33393a),
	.w8(32'h3b4f14ff),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b336453),
	.w1(32'h3b07c75c),
	.w2(32'h3943b447),
	.w3(32'h394ece24),
	.w4(32'hbb00d59c),
	.w5(32'hbb8f1b3d),
	.w6(32'hba704073),
	.w7(32'hba929b22),
	.w8(32'hbbb6fbdf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeaf33c),
	.w1(32'hbbb47d13),
	.w2(32'hbb469ddb),
	.w3(32'hbbcbd6bc),
	.w4(32'hbbc542b9),
	.w5(32'hbb03e7be),
	.w6(32'hbbc76672),
	.w7(32'hbb991c64),
	.w8(32'h3aab562f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ba91e),
	.w1(32'h392e932f),
	.w2(32'hba522482),
	.w3(32'hba82028a),
	.w4(32'hbaa4198b),
	.w5(32'hb92f7ae4),
	.w6(32'h3aecb688),
	.w7(32'hbb7e3f26),
	.w8(32'h3a4fdbac),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6fd61),
	.w1(32'hba2da451),
	.w2(32'hbb0133d7),
	.w3(32'h39e0b18e),
	.w4(32'h39ae50e5),
	.w5(32'h3ba9abdb),
	.w6(32'hba38a669),
	.w7(32'hba26ea19),
	.w8(32'h3b3e684c),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393def07),
	.w1(32'h3abc9780),
	.w2(32'h3ad08616),
	.w3(32'h3b580efc),
	.w4(32'h3a36ae05),
	.w5(32'hbaa23b3c),
	.w6(32'h3b82d7ff),
	.w7(32'h3ac7eeef),
	.w8(32'hba6b9a80),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00a1fd),
	.w1(32'h3b0f5546),
	.w2(32'hbafbfac2),
	.w3(32'h3b20a9fa),
	.w4(32'hb9d8f012),
	.w5(32'h3b934bbc),
	.w6(32'h3be7703a),
	.w7(32'h36d536fb),
	.w8(32'h3bca9b03),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5de4eb),
	.w1(32'hb8efeb46),
	.w2(32'h3ab6f298),
	.w3(32'hb79d84c1),
	.w4(32'h3a68e59c),
	.w5(32'hba9011bd),
	.w6(32'h3b5e992d),
	.w7(32'h3b5c00d2),
	.w8(32'hba12caaa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4035ce),
	.w1(32'h3b81881f),
	.w2(32'h3a953863),
	.w3(32'h3b52418b),
	.w4(32'hba362dd5),
	.w5(32'h3bab6c78),
	.w6(32'h3bd2709c),
	.w7(32'h3ae7cfce),
	.w8(32'h3b948793),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3905d8),
	.w1(32'h3bbb490e),
	.w2(32'h3bb46463),
	.w3(32'h3ba82a8a),
	.w4(32'h3aface0f),
	.w5(32'h3a7cfde0),
	.w6(32'h3c568eed),
	.w7(32'h3bb0d8a4),
	.w8(32'hba61e918),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976f004),
	.w1(32'h3b83ec60),
	.w2(32'h3af39e89),
	.w3(32'h3b2eaf7b),
	.w4(32'h3b85d65c),
	.w5(32'hbac6ca30),
	.w6(32'h3b56c310),
	.w7(32'h3bace89a),
	.w8(32'hba03db28),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f6e00),
	.w1(32'h3b0a6cd1),
	.w2(32'hbb0c0893),
	.w3(32'h3a68fd0e),
	.w4(32'hbb0daf62),
	.w5(32'h3ad18dd8),
	.w6(32'h3a959c1d),
	.w7(32'hbaca5dd2),
	.w8(32'hbaf2e016),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01a6f1),
	.w1(32'hba9b0ad6),
	.w2(32'h39644ac3),
	.w3(32'h3a432eb1),
	.w4(32'h3a187d49),
	.w5(32'h38c11148),
	.w6(32'hbb1b7d80),
	.w7(32'h3a8da916),
	.w8(32'hbb8566e1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41abd2),
	.w1(32'hbbd8dd88),
	.w2(32'hbb8fe319),
	.w3(32'hba944b85),
	.w4(32'h3a81029f),
	.w5(32'h3b408f8f),
	.w6(32'hbb2bee05),
	.w7(32'hbaf5d81f),
	.w8(32'h3b43d85f),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3233a1),
	.w1(32'h3ad5607c),
	.w2(32'hbaf8e778),
	.w3(32'h3b1679b7),
	.w4(32'h3ad0e498),
	.w5(32'hbac4a5a0),
	.w6(32'h3a461bd3),
	.w7(32'hb95b802d),
	.w8(32'hbb3f5602),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d45b1),
	.w1(32'hbb3d74e8),
	.w2(32'hb97fcf95),
	.w3(32'hbaf9ded7),
	.w4(32'hbb186fc6),
	.w5(32'hbb8dde5b),
	.w6(32'hbb4d6e2f),
	.w7(32'hbb02eaf4),
	.w8(32'hba660065),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b0ffb),
	.w1(32'hb980aa8a),
	.w2(32'hba105385),
	.w3(32'hbb8f35dc),
	.w4(32'hbac59012),
	.w5(32'hbafac5ea),
	.w6(32'hbbad741c),
	.w7(32'hbb47b029),
	.w8(32'hbb68adcf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9e9a9),
	.w1(32'h3baf214e),
	.w2(32'h39f5dbd3),
	.w3(32'h3b8234f0),
	.w4(32'hb800db46),
	.w5(32'h3b891aa7),
	.w6(32'h3b8d0684),
	.w7(32'hb8283c90),
	.w8(32'h3ba1a40b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a773d45),
	.w1(32'hba800812),
	.w2(32'h3b9c4f97),
	.w3(32'hbafec9b2),
	.w4(32'h39a80f8e),
	.w5(32'hbb058066),
	.w6(32'hbaf6bb23),
	.w7(32'h3b59f2b2),
	.w8(32'hbb35f865),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba970c3b),
	.w1(32'h3b65c243),
	.w2(32'h39e9e525),
	.w3(32'hbb446292),
	.w4(32'h3a6448f2),
	.w5(32'hbaf373a6),
	.w6(32'hbb035dda),
	.w7(32'h3b4b47e0),
	.w8(32'hbb0ffa93),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac80ba7),
	.w1(32'h398ac811),
	.w2(32'hb9c07316),
	.w3(32'hbaafc392),
	.w4(32'h3a8f8995),
	.w5(32'hbb29a88b),
	.w6(32'hbb2f2d62),
	.w7(32'h3b2a8fab),
	.w8(32'h398db8eb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a8ffc),
	.w1(32'h39cf4c88),
	.w2(32'hbb82d647),
	.w3(32'hbb8519c8),
	.w4(32'hbb31e95d),
	.w5(32'hba50b348),
	.w6(32'hba4422ac),
	.w7(32'hbb3f3cf5),
	.w8(32'hbb2a1003),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0befaa),
	.w1(32'hbb127bc7),
	.w2(32'hbb2ef2e0),
	.w3(32'hbb2f8d41),
	.w4(32'hbae1b3f0),
	.w5(32'hbb0ffebb),
	.w6(32'hbaae30e2),
	.w7(32'hba3e3773),
	.w8(32'hba40b790),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb0f62),
	.w1(32'h3a8efd1a),
	.w2(32'hbb7d2917),
	.w3(32'hbb681fe9),
	.w4(32'hbad1c5b3),
	.w5(32'h39d11c41),
	.w6(32'hba8ab0b7),
	.w7(32'hb98ac1f7),
	.w8(32'hbb4f1c46),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb724583),
	.w1(32'hba37c659),
	.w2(32'h3b0c0d2a),
	.w3(32'h3b6d69fa),
	.w4(32'h3b9a6984),
	.w5(32'hbb2753a4),
	.w6(32'hb9cb383a),
	.w7(32'h3ac1eb25),
	.w8(32'hba5cb536),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c1d6c),
	.w1(32'hbb29f31b),
	.w2(32'hba1c406f),
	.w3(32'hbb3df16b),
	.w4(32'hbb26f30b),
	.w5(32'hb90b0f9a),
	.w6(32'hbaa080b5),
	.w7(32'hbb20b456),
	.w8(32'hba52353d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75080f),
	.w1(32'hb97eacfb),
	.w2(32'hba25786a),
	.w3(32'h3b1e0f9f),
	.w4(32'h3a9fc3a2),
	.w5(32'hbac97f18),
	.w6(32'h3a25dc2b),
	.w7(32'hb9d80db0),
	.w8(32'h3b431485),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d6f7d),
	.w1(32'h3bbe421f),
	.w2(32'h3b5d118a),
	.w3(32'h3ba1e10d),
	.w4(32'h3b07b36e),
	.w5(32'hbb2fb0b5),
	.w6(32'h3baeea8d),
	.w7(32'h3b42e77f),
	.w8(32'hbae4cd91),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82b3f51),
	.w1(32'hbb1e9dac),
	.w2(32'hbb4fd431),
	.w3(32'hbb97b6f0),
	.w4(32'hbb2ce01c),
	.w5(32'h38b3f898),
	.w6(32'hbbe85e6a),
	.w7(32'hbb90f7d5),
	.w8(32'hba9c0205),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46793c),
	.w1(32'h3b914ad0),
	.w2(32'h3ab24f34),
	.w3(32'h3b6162f0),
	.w4(32'h3a16a122),
	.w5(32'hba2edd2d),
	.w6(32'h3b772444),
	.w7(32'h3b4d103d),
	.w8(32'h3a85d0a4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52036d),
	.w1(32'hba50f7fc),
	.w2(32'h3aea23dc),
	.w3(32'hb9970c1a),
	.w4(32'h3aa194df),
	.w5(32'h3b1a5d4f),
	.w6(32'h3b289430),
	.w7(32'h3b1b2e5e),
	.w8(32'h3ad82bdf),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71073d),
	.w1(32'hbb6c5f72),
	.w2(32'hbb0612e8),
	.w3(32'h3904c473),
	.w4(32'h3af9a3fe),
	.w5(32'hba72f94b),
	.w6(32'hba83f43b),
	.w7(32'h3a9fe9db),
	.w8(32'h37aa232e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0e38a),
	.w1(32'h39eacd1b),
	.w2(32'hb9bc590a),
	.w3(32'hb9e9af4c),
	.w4(32'hb8718b16),
	.w5(32'hbb790f72),
	.w6(32'h3b779d03),
	.w7(32'h3aabd795),
	.w8(32'hbb36d992),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb122a55),
	.w1(32'hbb6139e3),
	.w2(32'hbaf35aef),
	.w3(32'hbbb4781f),
	.w4(32'hbaf94841),
	.w5(32'h3b241bae),
	.w6(32'hbb6c24f1),
	.w7(32'hbabfc8ef),
	.w8(32'h3b971490),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19abb2),
	.w1(32'h3bf7fd4d),
	.w2(32'h3b3863b1),
	.w3(32'h3bf31656),
	.w4(32'h3b5a1a48),
	.w5(32'hbb05ee9f),
	.w6(32'h3c464bde),
	.w7(32'h3b8e7997),
	.w8(32'hbb2d3f19),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae66ac),
	.w1(32'hba012c20),
	.w2(32'hbb0df704),
	.w3(32'hba15cc30),
	.w4(32'hba871b5e),
	.w5(32'h39813d15),
	.w6(32'h3a632010),
	.w7(32'hba2599a5),
	.w8(32'h3a9902b2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00db04),
	.w1(32'h39967931),
	.w2(32'h3b0118cf),
	.w3(32'h3a104a8e),
	.w4(32'h3a12657d),
	.w5(32'h3a143c9d),
	.w6(32'h3b775126),
	.w7(32'h3b3559f6),
	.w8(32'h3b0c824c),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acee057),
	.w1(32'h378ab3a7),
	.w2(32'hb89d030c),
	.w3(32'hb770588b),
	.w4(32'h3a61e015),
	.w5(32'h3b1ee855),
	.w6(32'h3b609167),
	.w7(32'h3b009560),
	.w8(32'h3a2f1237),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab9d424),
	.w1(32'h3b9442f7),
	.w2(32'h3aef722d),
	.w3(32'h3ad9d386),
	.w4(32'h3b7d3d28),
	.w5(32'h3b804ba2),
	.w6(32'h3bbfce3b),
	.w7(32'h3bce75b6),
	.w8(32'h3b9206dc),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ba2e2),
	.w1(32'h3b29612c),
	.w2(32'h3ac3f0df),
	.w3(32'h3b861128),
	.w4(32'h3b171403),
	.w5(32'hb9f30fc2),
	.w6(32'h3b721a1f),
	.w7(32'h3af3b12d),
	.w8(32'h39ec3b68),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c068c),
	.w1(32'h3ad523d0),
	.w2(32'h3b34b6d2),
	.w3(32'h3a42e446),
	.w4(32'h3b4950e1),
	.w5(32'h3ae5138f),
	.w6(32'h3af00c5d),
	.w7(32'h3b8d6ff8),
	.w8(32'h3b6ce6ff),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c8279),
	.w1(32'h3b63c978),
	.w2(32'h3b904b51),
	.w3(32'h3b090b6f),
	.w4(32'h3b164459),
	.w5(32'hba47a335),
	.w6(32'h3c263911),
	.w7(32'h3bb31375),
	.w8(32'h3b68115e),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40cac1),
	.w1(32'h39db861d),
	.w2(32'hbac4b673),
	.w3(32'h3a034062),
	.w4(32'hbabf46b9),
	.w5(32'hbb29bebe),
	.w6(32'h3a0637b5),
	.w7(32'hbb200874),
	.w8(32'h3a5ec328),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaccf06a),
	.w1(32'h3aef5a5d),
	.w2(32'hbb910210),
	.w3(32'h3abc2e28),
	.w4(32'hbae75bc6),
	.w5(32'hba0cd24c),
	.w6(32'h3bd4a991),
	.w7(32'hba47737c),
	.w8(32'hba946b43),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e175e4),
	.w1(32'hb88b6656),
	.w2(32'hbb2e267b),
	.w3(32'h3a85c36f),
	.w4(32'hba006a9b),
	.w5(32'hbb41349d),
	.w6(32'h39ad4b9d),
	.w7(32'hbaf749ab),
	.w8(32'hbb89f24a),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9129c3),
	.w1(32'hbb0a6ef0),
	.w2(32'hbad5bcb7),
	.w3(32'hbb7b7b35),
	.w4(32'hbb2d0f08),
	.w5(32'hbb07cf40),
	.w6(32'h3a53f432),
	.w7(32'hbb6e638e),
	.w8(32'hbb4687ec),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55b54d),
	.w1(32'hbad0ae23),
	.w2(32'h3a1b2d5e),
	.w3(32'h3ac9b2d5),
	.w4(32'h3ad25ab7),
	.w5(32'hbb290019),
	.w6(32'hb7ade4a3),
	.w7(32'h3b404b95),
	.w8(32'h39c3baa3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e8538),
	.w1(32'hbaf52c81),
	.w2(32'hba8db790),
	.w3(32'hb9f291da),
	.w4(32'hba857f1d),
	.w5(32'hba9b4992),
	.w6(32'hbad4aaf5),
	.w7(32'hbab6f7c8),
	.w8(32'hbacb3568),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb202469),
	.w1(32'hba35c747),
	.w2(32'h3ac93823),
	.w3(32'hbb20e11e),
	.w4(32'hbb257e00),
	.w5(32'h3b8f0cd0),
	.w6(32'hbabb0412),
	.w7(32'hbaa70ec8),
	.w8(32'h3a4d455c),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c18314),
	.w1(32'h38d7d680),
	.w2(32'h3a4ed792),
	.w3(32'h39cebbf0),
	.w4(32'hbac0af15),
	.w5(32'h3b50f077),
	.w6(32'hbb30a3bb),
	.w7(32'hb8847f80),
	.w8(32'h3bc6dc2a),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b630a5d),
	.w1(32'hbb0ccbe5),
	.w2(32'h3b4606a8),
	.w3(32'h3b4fa034),
	.w4(32'hba7e4989),
	.w5(32'hb95d0d26),
	.w6(32'hbb0c82c3),
	.w7(32'h3b420dcf),
	.w8(32'h3b181ec0),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3fafef),
	.w1(32'h3aa609d2),
	.w2(32'h398aad3d),
	.w3(32'hbaa04c6b),
	.w4(32'hba5d244b),
	.w5(32'hb9ea2d87),
	.w6(32'h3a773fba),
	.w7(32'hba34bdca),
	.w8(32'h3b57ab51),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a82f414),
	.w1(32'h3b1dc8cf),
	.w2(32'h3a1bd35d),
	.w3(32'h3acb4d51),
	.w4(32'hb9cc4f33),
	.w5(32'hba6ff653),
	.w6(32'h3c163580),
	.w7(32'h3a38f11f),
	.w8(32'h3a3ba6ba),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7da779),
	.w1(32'hbae04c43),
	.w2(32'h3a001058),
	.w3(32'hbb7bab88),
	.w4(32'h39cfdf99),
	.w5(32'hba3008be),
	.w6(32'hb9d7b29e),
	.w7(32'h3a816c6d),
	.w8(32'hb9918dc7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13f17b),
	.w1(32'h3b0693aa),
	.w2(32'hb964d4c2),
	.w3(32'h3b277c46),
	.w4(32'hbb0f697c),
	.w5(32'hbb21ea07),
	.w6(32'h3b7cf959),
	.w7(32'hb8c70aea),
	.w8(32'hbb177b63),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb081419),
	.w1(32'hbb1b064b),
	.w2(32'h39b7d5f9),
	.w3(32'hbb8cf51d),
	.w4(32'hb9c72244),
	.w5(32'hbadf2867),
	.w6(32'hbb5fd6c5),
	.w7(32'hba79b335),
	.w8(32'hbaefafef),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafeeb6d),
	.w1(32'hba9c00d0),
	.w2(32'hba4db7fc),
	.w3(32'hbafdb2f5),
	.w4(32'h39d23af2),
	.w5(32'h3b298a3a),
	.w6(32'hbb1f53fe),
	.w7(32'h397c2a92),
	.w8(32'hbaaa1376),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad88b53),
	.w1(32'h39e31412),
	.w2(32'h3b2dbc10),
	.w3(32'hbb43dc66),
	.w4(32'h3931ca01),
	.w5(32'hbac64456),
	.w6(32'hbb63da78),
	.w7(32'h39fb9d6f),
	.w8(32'hbbadc902),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba29782),
	.w1(32'hbb5b4874),
	.w2(32'hbb030c3c),
	.w3(32'hbb277f7c),
	.w4(32'hba91a3b4),
	.w5(32'hba3de7fe),
	.w6(32'hbb8424ff),
	.w7(32'h39d32956),
	.w8(32'hbae48dc8),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ab1ae9),
	.w1(32'hb92a0fc6),
	.w2(32'hbb5da19e),
	.w3(32'h3a5ac39d),
	.w4(32'h3923b18d),
	.w5(32'hb98a1bdd),
	.w6(32'h3b1a4a39),
	.w7(32'hbb3bc1a9),
	.w8(32'h381546ea),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad54bfc),
	.w1(32'h3a8ee561),
	.w2(32'hbabaf7d3),
	.w3(32'h3a3e0e90),
	.w4(32'hb9a847b5),
	.w5(32'hbab746c7),
	.w6(32'h3a8102fa),
	.w7(32'hba0c129c),
	.w8(32'h3afd1365),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaa59f),
	.w1(32'h3a96931b),
	.w2(32'h3a5209d2),
	.w3(32'hba8d2983),
	.w4(32'hba722251),
	.w5(32'h3b501f06),
	.w6(32'h3a8d0aa6),
	.w7(32'h396fa44f),
	.w8(32'h3b1b1355),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a7bd1),
	.w1(32'hba827233),
	.w2(32'hbac3fdb2),
	.w3(32'h3a9ff3d4),
	.w4(32'hba2c6837),
	.w5(32'hbb05ba54),
	.w6(32'hba620e66),
	.w7(32'hb92085f3),
	.w8(32'h3a865969),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b2373),
	.w1(32'h3a547315),
	.w2(32'hbb1c2cc7),
	.w3(32'hbb257660),
	.w4(32'hbb4f1c2e),
	.w5(32'hbb500400),
	.w6(32'hbb2c0552),
	.w7(32'hbb7e7075),
	.w8(32'hbb2acffa),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6efc8f),
	.w1(32'hbad2088f),
	.w2(32'hba2f75ae),
	.w3(32'hbbb1cfdc),
	.w4(32'hb98fc5f2),
	.w5(32'hba6a0682),
	.w6(32'hbb3990df),
	.w7(32'hba70406f),
	.w8(32'hbb450a0e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad951d),
	.w1(32'hbb243582),
	.w2(32'hbb1e1bfe),
	.w3(32'h3a6d98e9),
	.w4(32'hbb60aa42),
	.w5(32'hba3de770),
	.w6(32'hbb5278cd),
	.w7(32'hbade427f),
	.w8(32'hb9631596),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacfa84f),
	.w1(32'h3b0b02e2),
	.w2(32'h3b6ff6df),
	.w3(32'hba2ec274),
	.w4(32'h390a2dda),
	.w5(32'h3a1d1426),
	.w6(32'h3a1f23b3),
	.w7(32'h3a23d0de),
	.w8(32'h39e78604),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88a728),
	.w1(32'h3abeab6d),
	.w2(32'hba3f0b8b),
	.w3(32'hba01e8bd),
	.w4(32'h3a0201f6),
	.w5(32'hbb08b3cb),
	.w6(32'hba8f242e),
	.w7(32'h39805ce1),
	.w8(32'h39b12566),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26c43b),
	.w1(32'hbac8345a),
	.w2(32'hb932dc77),
	.w3(32'hbb0d14fa),
	.w4(32'hba9ccaa0),
	.w5(32'h393c86e8),
	.w6(32'h3b4d4e23),
	.w7(32'h3a3e313e),
	.w8(32'hbb2b5487),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3964dea3),
	.w1(32'hbb239ed9),
	.w2(32'hbb849789),
	.w3(32'hbb2b818f),
	.w4(32'hba99c58d),
	.w5(32'h3b1fc951),
	.w6(32'hbb5a8eab),
	.w7(32'hbb5042b3),
	.w8(32'h3b48ae8c),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b459802),
	.w1(32'hb989c3e4),
	.w2(32'hbb8915f6),
	.w3(32'hbafa9784),
	.w4(32'hbb8e75bf),
	.w5(32'hbb765a3e),
	.w6(32'h3b97310b),
	.w7(32'hbb8f65d9),
	.w8(32'hbb4e6926),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba09c44),
	.w1(32'hbb5559ed),
	.w2(32'hba49e480),
	.w3(32'hbba263ad),
	.w4(32'hbb654607),
	.w5(32'h3975fd91),
	.w6(32'hbad89d36),
	.w7(32'hbb0c2df0),
	.w8(32'h3aaa53c8),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22004c),
	.w1(32'hb95ea46a),
	.w2(32'h3a038d7e),
	.w3(32'h3b34e6bf),
	.w4(32'hb94154cc),
	.w5(32'hbb65feda),
	.w6(32'h3baa7ff3),
	.w7(32'h3ac597da),
	.w8(32'hba9c2b39),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba62c1a),
	.w1(32'hbb2b1443),
	.w2(32'hbab812b1),
	.w3(32'hbb8a6670),
	.w4(32'hbb86a16a),
	.w5(32'hbac8a6c6),
	.w6(32'hba8843f7),
	.w7(32'hbae95755),
	.w8(32'hba8066d4),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f25b3),
	.w1(32'hba9e48a9),
	.w2(32'hba95871e),
	.w3(32'hbac30d19),
	.w4(32'hbb44b700),
	.w5(32'h3afcfd7c),
	.w6(32'hbb166a64),
	.w7(32'hbad495ba),
	.w8(32'h3b6c814b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90384d),
	.w1(32'h3b767077),
	.w2(32'h3a175e97),
	.w3(32'h3b67c77d),
	.w4(32'h3b1849bc),
	.w5(32'hb9e2999c),
	.w6(32'h3b46eb97),
	.w7(32'h3b152982),
	.w8(32'h3a80214b),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadff8ca),
	.w1(32'h39e8122d),
	.w2(32'h3b103a57),
	.w3(32'hbb171312),
	.w4(32'hbb0b0557),
	.w5(32'h3bddf3c4),
	.w6(32'h39f1cfd2),
	.w7(32'h3a9234b6),
	.w8(32'h3b8e62ce),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce40cd),
	.w1(32'hba122cca),
	.w2(32'hb9eebd3e),
	.w3(32'hba479f7d),
	.w4(32'h3b3c8d4d),
	.w5(32'hbae3f62f),
	.w6(32'hba48ec36),
	.w7(32'h3b14f161),
	.w8(32'hbb275ac0),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394f1ee2),
	.w1(32'hbb4d55df),
	.w2(32'hbb40cb94),
	.w3(32'hbb06e586),
	.w4(32'h39e92674),
	.w5(32'hbb133861),
	.w6(32'hbada8ac8),
	.w7(32'hbacb0006),
	.w8(32'hbad7d2f6),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8724c0f),
	.w1(32'h3b36c5b8),
	.w2(32'hba24bcf0),
	.w3(32'h39b830ef),
	.w4(32'h39de6499),
	.w5(32'hba10c2ef),
	.w6(32'h3ae401e8),
	.w7(32'h37925c68),
	.w8(32'h39a2f424),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb540c),
	.w1(32'h3b99680f),
	.w2(32'h3b65d62f),
	.w3(32'h39dc5498),
	.w4(32'h3bb08223),
	.w5(32'hbb0e4a48),
	.w6(32'h3aafc5c7),
	.w7(32'h3bbc84c2),
	.w8(32'hbb3ca326),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc02e3),
	.w1(32'hbb339224),
	.w2(32'hbb19b517),
	.w3(32'hba16e381),
	.w4(32'hba8999b8),
	.w5(32'hba77bfda),
	.w6(32'hbb00eac9),
	.w7(32'hbabceb90),
	.w8(32'h3a9c4e4d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca2257),
	.w1(32'hbb324282),
	.w2(32'hbb31dd22),
	.w3(32'hbb83bdf1),
	.w4(32'hbb2741c1),
	.w5(32'h377d3d86),
	.w6(32'hbab1b66b),
	.w7(32'hbb235f07),
	.w8(32'h39ab8de3),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93c98e8),
	.w1(32'h3a4304f0),
	.w2(32'h36eaa01c),
	.w3(32'hbb0528d6),
	.w4(32'hba82ba0b),
	.w5(32'hb9b2e9db),
	.w6(32'hb990533f),
	.w7(32'h389a50d4),
	.w8(32'hb9f03b18),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394c5eda),
	.w1(32'h3b9f399b),
	.w2(32'h3a45ba0d),
	.w3(32'h3b55044a),
	.w4(32'h39bd7cbf),
	.w5(32'hb9dce1fe),
	.w6(32'h3b846e7b),
	.w7(32'h3a79ef3b),
	.w8(32'h3a2c819d),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39093331),
	.w1(32'h38f17f46),
	.w2(32'h3a9d9947),
	.w3(32'hbb143333),
	.w4(32'hbab2de10),
	.w5(32'hbb3ae2a9),
	.w6(32'h3a9f4249),
	.w7(32'h3b050fc9),
	.w8(32'hbb5b860e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb799e32),
	.w1(32'hba3fbfc2),
	.w2(32'hbabe503c),
	.w3(32'hbb7d8235),
	.w4(32'hbbb2f622),
	.w5(32'h3a2ec9be),
	.w6(32'hba95afae),
	.w7(32'hbb422848),
	.w8(32'hb9767bc3),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3850f),
	.w1(32'h3ab1c736),
	.w2(32'h3b002a5b),
	.w3(32'h3ba63b6c),
	.w4(32'h3a7ff529),
	.w5(32'hbb0da3b8),
	.w6(32'h3b942dc9),
	.w7(32'h3b38ba6d),
	.w8(32'h3b5280a4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1eb78),
	.w1(32'hbab07537),
	.w2(32'hba558cb5),
	.w3(32'hbacf735c),
	.w4(32'hbb52b9e7),
	.w5(32'hba430588),
	.w6(32'h3b8a499f),
	.w7(32'hbaaaa7f5),
	.w8(32'h3aba484d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa769de),
	.w1(32'hb86f2fba),
	.w2(32'hba79e30b),
	.w3(32'hbaa1c0cf),
	.w4(32'h3a633b2f),
	.w5(32'h3aa5e3bc),
	.w6(32'hb98991e8),
	.w7(32'h3a692a2e),
	.w8(32'h3b3bffa9),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fa316),
	.w1(32'hb9f0209c),
	.w2(32'hba429e1d),
	.w3(32'hbb4055ad),
	.w4(32'hbb28c7a4),
	.w5(32'hb8b07a6f),
	.w6(32'hba8d2f2d),
	.w7(32'hbafb86d4),
	.w8(32'h3ac4ebc5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bf8e9),
	.w1(32'hbac733b3),
	.w2(32'h37bf8188),
	.w3(32'hbaa1276b),
	.w4(32'hb8e9733e),
	.w5(32'hbabc5123),
	.w6(32'hb9b7ac9a),
	.w7(32'h3829d575),
	.w8(32'hbb3d0d86),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5569e),
	.w1(32'hbb1a41b0),
	.w2(32'hbb193fbe),
	.w3(32'hbaed862e),
	.w4(32'h3a3f0d54),
	.w5(32'hb92c3383),
	.w6(32'hbb071cb6),
	.w7(32'hbac5cdf1),
	.w8(32'h3b097268),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d56493),
	.w1(32'h3bfb8e7b),
	.w2(32'h3b2f683b),
	.w3(32'h3b81e751),
	.w4(32'h3b7ebeed),
	.w5(32'h3bbd0d22),
	.w6(32'h3c3dde61),
	.w7(32'h3bbd3e2f),
	.w8(32'h3bdc3f4a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bebb19d),
	.w1(32'hba691f8a),
	.w2(32'hba86bd4f),
	.w3(32'hbaae90fa),
	.w4(32'h3b1fcdf1),
	.w5(32'h3b8f4bbf),
	.w6(32'h3a366229),
	.w7(32'h3aa28b10),
	.w8(32'h3b91f675),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6aca13),
	.w1(32'h3b2d9f52),
	.w2(32'hbafceb48),
	.w3(32'h3b80cc92),
	.w4(32'h3a95b710),
	.w5(32'h3bb8113e),
	.w6(32'h3b8ea2b4),
	.w7(32'hb983ae3c),
	.w8(32'h3b9aff27),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14a316),
	.w1(32'h3b370aba),
	.w2(32'h3a200f3d),
	.w3(32'h3b02d7d0),
	.w4(32'h3abf87dc),
	.w5(32'h38867e9c),
	.w6(32'h3be7edcd),
	.w7(32'h3b219edf),
	.w8(32'h3a9b599f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3915ccad),
	.w1(32'hb8ec9e13),
	.w2(32'h39837e36),
	.w3(32'hbaa03e8f),
	.w4(32'h3a49d33b),
	.w5(32'hbb1b1a8b),
	.w6(32'h3a2eb4af),
	.w7(32'h398e50d7),
	.w8(32'h3b9381ee),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8bedc),
	.w1(32'h3b53a219),
	.w2(32'hb8ca8f94),
	.w3(32'h3c0d6bf7),
	.w4(32'h3b4f810d),
	.w5(32'hb8dbf6b2),
	.w6(32'h3bc0c5dc),
	.w7(32'h379fc56f),
	.w8(32'h3a37866f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacaedc1),
	.w1(32'hbafd2bec),
	.w2(32'hbb5da46f),
	.w3(32'h3abd9eb2),
	.w4(32'hb99ac762),
	.w5(32'hbafbb6c9),
	.w6(32'hbb1f7383),
	.w7(32'hbb1975a0),
	.w8(32'hbabd3640),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac11a84),
	.w1(32'hba310433),
	.w2(32'hbac7db70),
	.w3(32'hbb206e2e),
	.w4(32'hbb263ca2),
	.w5(32'hbac689ca),
	.w6(32'hbb2d059b),
	.w7(32'hbb2e58e4),
	.w8(32'h3a796ebc),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b18a56),
	.w1(32'h3bccda86),
	.w2(32'hb7f5811f),
	.w3(32'h3b1f810b),
	.w4(32'h3a36db2a),
	.w5(32'h397046d9),
	.w6(32'h3c076281),
	.w7(32'h3b0c0eb4),
	.w8(32'hba6fdcea),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39023a11),
	.w1(32'hb9f7a81b),
	.w2(32'hbb00d92f),
	.w3(32'h3a4c34a8),
	.w4(32'hba0ac1bb),
	.w5(32'h3b37377b),
	.w6(32'hba8b4bc4),
	.w7(32'hbb0db56f),
	.w8(32'h39c97c15),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da3505),
	.w1(32'hb93c33cd),
	.w2(32'h39ce6507),
	.w3(32'h39e61f0c),
	.w4(32'h39737fac),
	.w5(32'hbaa2729d),
	.w6(32'hbb3f21a2),
	.w7(32'hba4be6ca),
	.w8(32'hbaffdb52),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb422c7c),
	.w1(32'hbb6c1f09),
	.w2(32'hbb14d77a),
	.w3(32'hbb270a7a),
	.w4(32'hba424e3e),
	.w5(32'h3bf6d147),
	.w6(32'hba1b3709),
	.w7(32'hb89367f5),
	.w8(32'h3be9517e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13089),
	.w1(32'h3be8197a),
	.w2(32'h3bd9c03a),
	.w3(32'h3bff6a93),
	.w4(32'h3be73f2a),
	.w5(32'hba565c36),
	.w6(32'h3c2b8142),
	.w7(32'h3c07eaf8),
	.w8(32'h3b038495),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6b097d),
	.w1(32'h3b0ba89a),
	.w2(32'hbb2e24ab),
	.w3(32'h3b0c59eb),
	.w4(32'hba38b1b5),
	.w5(32'h3b638cb8),
	.w6(32'h3bcf7410),
	.w7(32'hb90812dd),
	.w8(32'h3b228f71),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58f852),
	.w1(32'h3b6b90d6),
	.w2(32'h3ba60b0b),
	.w3(32'h3b1bd8d4),
	.w4(32'h3aad52ef),
	.w5(32'h3a6363c6),
	.w6(32'h3b5a9667),
	.w7(32'h3aeb678e),
	.w8(32'h38ac3c84),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3905e671),
	.w1(32'h3991f94e),
	.w2(32'h39106e4f),
	.w3(32'h3a275179),
	.w4(32'h3aa098da),
	.w5(32'h3bc2e73e),
	.w6(32'h39dd3497),
	.w7(32'h39ad9dfb),
	.w8(32'h3b7b8e36),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f0727),
	.w1(32'hb99d5235),
	.w2(32'h39a5de29),
	.w3(32'hb9cd1fd4),
	.w4(32'hba9fa876),
	.w5(32'hbb2cefb4),
	.w6(32'hbb558b41),
	.w7(32'hb91562dd),
	.w8(32'h39c26929),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a926258),
	.w1(32'hbb7afbc6),
	.w2(32'hbb413fe1),
	.w3(32'hbb75574b),
	.w4(32'hb7dc51fd),
	.w5(32'h3b8a1cc2),
	.w6(32'hba9f149d),
	.w7(32'hba5cc743),
	.w8(32'h3afeb0b3),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7cbd90),
	.w1(32'hb99b39b1),
	.w2(32'h3a67cf60),
	.w3(32'h3b068ca1),
	.w4(32'h3a8ea046),
	.w5(32'h39c66ccd),
	.w6(32'hbad1553e),
	.w7(32'h3a6bc3e6),
	.w8(32'hba050966),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1c0e),
	.w1(32'hbb2bc6d2),
	.w2(32'hbb662a98),
	.w3(32'hbad5b688),
	.w4(32'hbb1808c9),
	.w5(32'h3b36a815),
	.w6(32'h3af834c8),
	.w7(32'hba9e8967),
	.w8(32'h3b25f7ef),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f4e5a),
	.w1(32'h3c1b472d),
	.w2(32'h3b935213),
	.w3(32'h3b94833b),
	.w4(32'h3b56d1b4),
	.w5(32'hba829a44),
	.w6(32'h3c3d74ff),
	.w7(32'h3c0aac9d),
	.w8(32'hbb72a11c),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf37ed7),
	.w1(32'hbb059dc8),
	.w2(32'hb9f24888),
	.w3(32'h39436515),
	.w4(32'h3addbdcc),
	.w5(32'hbb3a8b63),
	.w6(32'hbb6eb0af),
	.w7(32'hbaba151d),
	.w8(32'hbadf8c82),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17b15c),
	.w1(32'hba51d226),
	.w2(32'hbad5e507),
	.w3(32'hbb470cef),
	.w4(32'hbb251130),
	.w5(32'hbaa4795c),
	.w6(32'h3a57df59),
	.w7(32'hba833471),
	.w8(32'hb945692f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae88ae1),
	.w1(32'h3a4164b6),
	.w2(32'hbb425a1b),
	.w3(32'hbb5d5c26),
	.w4(32'h3b00d7ff),
	.w5(32'hbab9a423),
	.w6(32'h3a60cbdf),
	.w7(32'h3a3cbdf0),
	.w8(32'hb942205b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8634ee),
	.w1(32'h3a037889),
	.w2(32'hb8dc3a7f),
	.w3(32'h3b0eb68a),
	.w4(32'hba29bc81),
	.w5(32'hbb4e81bd),
	.w6(32'hb858b238),
	.w7(32'h3a7af62f),
	.w8(32'hb843a1f9),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944a96d),
	.w1(32'hbb283804),
	.w2(32'hbb5e30cf),
	.w3(32'h3a8aad5f),
	.w4(32'h3a2be334),
	.w5(32'hba3a4506),
	.w6(32'h3b173580),
	.w7(32'hbb3d0fd7),
	.w8(32'hb95f4faf),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed3774),
	.w1(32'hbaf6d8ed),
	.w2(32'hbb6a8f40),
	.w3(32'hbacfc1d6),
	.w4(32'hba8639e6),
	.w5(32'hbbc73eeb),
	.w6(32'h39b8eb1c),
	.w7(32'h3935756a),
	.w8(32'hbba16b8a),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856def),
	.w1(32'h3c26d916),
	.w2(32'h3a312518),
	.w3(32'h3bc955f1),
	.w4(32'hba7aa95c),
	.w5(32'hba30ed06),
	.w6(32'h3c1f96ec),
	.w7(32'hba34acc7),
	.w8(32'h3b113386),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b454f9a),
	.w1(32'h3b546c0c),
	.w2(32'h3ab2032b),
	.w3(32'h3b4c86cb),
	.w4(32'h3b46e612),
	.w5(32'hba25323e),
	.w6(32'h3b78c690),
	.w7(32'h3a668d4d),
	.w8(32'hbb60251e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb072a9e),
	.w1(32'hbb4d4a02),
	.w2(32'hbba4e40f),
	.w3(32'h38cc1f5c),
	.w4(32'hbad6715e),
	.w5(32'h3ad78e32),
	.w6(32'hba61dfa7),
	.w7(32'hbb0d67db),
	.w8(32'hba3cfe11),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb245671),
	.w1(32'hb9c93086),
	.w2(32'h3a53693b),
	.w3(32'hba7aac69),
	.w4(32'hb9cea5c4),
	.w5(32'hba1d59f6),
	.w6(32'hb9f7a5f2),
	.w7(32'hb9bbb7f9),
	.w8(32'hbb036424),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb0a31),
	.w1(32'hb9f190df),
	.w2(32'hba5767c3),
	.w3(32'h3a1f7bf5),
	.w4(32'hba8525bd),
	.w5(32'h35eafb33),
	.w6(32'h37424ca7),
	.w7(32'hbafe8957),
	.w8(32'h35975b7f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h359c43a4),
	.w1(32'h3794d6b7),
	.w2(32'h37662ad0),
	.w3(32'h37a7e870),
	.w4(32'h36a4507e),
	.w5(32'hb66b58dd),
	.w6(32'h380dbb60),
	.w7(32'h378d84b7),
	.w8(32'h3760ddc3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38598af4),
	.w1(32'h38719a7d),
	.w2(32'h385185a0),
	.w3(32'h37cb8379),
	.w4(32'h3838f132),
	.w5(32'hb548c3d9),
	.w6(32'h384d9166),
	.w7(32'h388083a8),
	.w8(32'h3868cfb6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371e0c90),
	.w1(32'h37300417),
	.w2(32'h37238cbd),
	.w3(32'h3669dcad),
	.w4(32'h3707ae3b),
	.w5(32'h37768637),
	.w6(32'h37a84a88),
	.w7(32'h37e24d43),
	.w8(32'h3731df7f),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3674a95e),
	.w1(32'h35933f5f),
	.w2(32'h34eb9824),
	.w3(32'h37445893),
	.w4(32'h36fcb34e),
	.w5(32'h346e853d),
	.w6(32'hb751dda6),
	.w7(32'hb76f8e2b),
	.w8(32'hb52ddf1e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380dd2f1),
	.w1(32'h356e5711),
	.w2(32'h379ba851),
	.w3(32'h37d71b8b),
	.w4(32'hb63cc6de),
	.w5(32'hb8763c29),
	.w6(32'h390a9532),
	.w7(32'h38de97a2),
	.w8(32'h3880a810),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e6803a),
	.w1(32'h350a15c5),
	.w2(32'h3779ea1e),
	.w3(32'hb7001ba1),
	.w4(32'hb6dd6909),
	.w5(32'h364894e1),
	.w6(32'h38217259),
	.w7(32'h3806e963),
	.w8(32'h37af93b6),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b72181),
	.w1(32'h368f8e0c),
	.w2(32'h365ebbf9),
	.w3(32'h3753b4e2),
	.w4(32'h37630945),
	.w5(32'h362221ad),
	.w6(32'hb70e34b1),
	.w7(32'hb6e4dc3b),
	.w8(32'hb6270e06),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6acd67b),
	.w1(32'hb6a0e888),
	.w2(32'h34cba926),
	.w3(32'h33c42052),
	.w4(32'hb76b9ec9),
	.w5(32'hb74d451f),
	.w6(32'h37e2274a),
	.w7(32'h37ec34ac),
	.w8(32'h37ae2201),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d9edff),
	.w1(32'h3675b3e1),
	.w2(32'hb6b3a809),
	.w3(32'h36daeddb),
	.w4(32'h363ecead),
	.w5(32'hb7197ece),
	.w6(32'h36a1e929),
	.w7(32'hb6bd673e),
	.w8(32'hb71600cb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h355a5aae),
	.w1(32'h36975200),
	.w2(32'h36261be8),
	.w3(32'h35799210),
	.w4(32'hb5c05aa0),
	.w5(32'h359a9345),
	.w6(32'h368a6d6e),
	.w7(32'h35744567),
	.w8(32'h36929142),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36387288),
	.w1(32'h36c531d2),
	.w2(32'h36112c6c),
	.w3(32'h363f6cf6),
	.w4(32'hb563bb41),
	.w5(32'h364d6573),
	.w6(32'h35f5dca0),
	.w7(32'hb624efe5),
	.w8(32'h3546a536),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a32a39),
	.w1(32'h369eaece),
	.w2(32'h36a28ee8),
	.w3(32'h363d82de),
	.w4(32'h36c42349),
	.w5(32'hb50f9b21),
	.w6(32'h353e9c21),
	.w7(32'h36803f8d),
	.w8(32'hb4e383b5),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68ea139),
	.w1(32'h36829dd4),
	.w2(32'hb780d319),
	.w3(32'h3631cda4),
	.w4(32'h36ced2f2),
	.w5(32'hb71ef0cd),
	.w6(32'h36675823),
	.w7(32'h36b6ed7b),
	.w8(32'h36124cfa),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38534663),
	.w1(32'h38a426b6),
	.w2(32'h38e422a1),
	.w3(32'hb7746683),
	.w4(32'h382b4e4c),
	.w5(32'h37cf1190),
	.w6(32'h38910a3d),
	.w7(32'h3818b7c2),
	.w8(32'h3886896b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36acad6f),
	.w1(32'h376802d7),
	.w2(32'h3809059e),
	.w3(32'hb77b19ba),
	.w4(32'hb69f08c5),
	.w5(32'h371e4502),
	.w6(32'h37fc9441),
	.w7(32'h380ecf5f),
	.w8(32'h3837a357),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37607c97),
	.w1(32'h3841ecb1),
	.w2(32'h38b06547),
	.w3(32'hb801de93),
	.w4(32'h36573dca),
	.w5(32'h37edc45f),
	.w6(32'h38a3d651),
	.w7(32'h388477a9),
	.w8(32'h38b51e57),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69954cf),
	.w1(32'hb64dcb59),
	.w2(32'h34e4ed04),
	.w3(32'h35b0fb55),
	.w4(32'hb50f5e2a),
	.w5(32'h33c0ab45),
	.w6(32'h36924a1d),
	.w7(32'h36b86b13),
	.w8(32'hb5ba6b82),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362f8131),
	.w1(32'h35ea1927),
	.w2(32'h370cb04d),
	.w3(32'hb647caad),
	.w4(32'hb6c44dfe),
	.w5(32'h363e0abe),
	.w6(32'h36583a32),
	.w7(32'hb70a33ff),
	.w8(32'hb665bed0),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ae2172),
	.w1(32'h357c284f),
	.w2(32'h3510ccd5),
	.w3(32'hb6a316b1),
	.w4(32'hb3849639),
	.w5(32'h37902f24),
	.w6(32'hb66783b8),
	.w7(32'h3565fc74),
	.w8(32'hb592578c),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370009db),
	.w1(32'h36595504),
	.w2(32'h35fee8f1),
	.w3(32'h375465b5),
	.w4(32'h3749ad45),
	.w5(32'h356aaeaa),
	.w6(32'hb6c5a5a3),
	.w7(32'hb60c6729),
	.w8(32'hb6970a62),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37328416),
	.w1(32'h3801db44),
	.w2(32'h384c47bc),
	.w3(32'hb7c8e494),
	.w4(32'hb7218a50),
	.w5(32'h37e5a036),
	.w6(32'h383c86b0),
	.w7(32'h38091ee1),
	.w8(32'h384a451d),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f4ef70),
	.w1(32'h3729b7d3),
	.w2(32'hb5b67524),
	.w3(32'h36fd8c87),
	.w4(32'h36b4f186),
	.w5(32'h358b02cd),
	.w6(32'h37853ee2),
	.w7(32'h3731927e),
	.w8(32'h36575eec),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h351364ef),
	.w1(32'hb67574fe),
	.w2(32'hb6dd673d),
	.w3(32'h369d6d1a),
	.w4(32'hb5fca79b),
	.w5(32'hb7022559),
	.w6(32'h372b9d70),
	.w7(32'h370c1694),
	.w8(32'hb59be372),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h361bb37f),
	.w1(32'h3757c0e8),
	.w2(32'h372f644f),
	.w3(32'h343e4cd3),
	.w4(32'h36999857),
	.w5(32'h3712f466),
	.w6(32'hb61c9c48),
	.w7(32'hb609ebce),
	.w8(32'h36e11158),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7355b03),
	.w1(32'hb6f6c21e),
	.w2(32'hb6677785),
	.w3(32'h36740f22),
	.w4(32'hb4a83147),
	.w5(32'h363b988c),
	.w6(32'h349eadd7),
	.w7(32'hb5d9084f),
	.w8(32'h34f73c0a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36702ce4),
	.w1(32'h36cd9805),
	.w2(32'h37b6d810),
	.w3(32'hb5515392),
	.w4(32'h3711ca4d),
	.w5(32'h3757f1ae),
	.w6(32'h37b0df00),
	.w7(32'h379208f2),
	.w8(32'h37f780ab),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d5bb5f),
	.w1(32'hb6091b57),
	.w2(32'hb4d91ace),
	.w3(32'h3631ba8a),
	.w4(32'h35e9969c),
	.w5(32'h37030b6b),
	.w6(32'h360024af),
	.w7(32'h362a2ca5),
	.w8(32'hb5a2488b),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6df6449),
	.w1(32'h384e5d40),
	.w2(32'h38d44844),
	.w3(32'h3419c76f),
	.w4(32'h3808d5e4),
	.w5(32'h37df9779),
	.w6(32'h3829a3ac),
	.w7(32'h365bf78f),
	.w8(32'h38c0d74f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36293eca),
	.w1(32'h36a885e5),
	.w2(32'h36ca4282),
	.w3(32'h36253aef),
	.w4(32'h365358b0),
	.w5(32'hb69df2ed),
	.w6(32'h36b3a6fd),
	.w7(32'h36b6615a),
	.w8(32'hb5b204a6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88185b0),
	.w1(32'hb7d6c2cf),
	.w2(32'hb73297ec),
	.w3(32'h378f58ec),
	.w4(32'h3681f619),
	.w5(32'h37f89d00),
	.w6(32'h37e55a89),
	.w7(32'h37ea2612),
	.w8(32'h3808dfba),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule