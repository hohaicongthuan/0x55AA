module layer_10_featuremap_177(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a31972),
	.w1(32'h3a0bcf5a),
	.w2(32'hb57bcd83),
	.w3(32'h39d30a19),
	.w4(32'hb7cfbf9c),
	.w5(32'hb8ebf3ce),
	.w6(32'h39cb0aa2),
	.w7(32'h391a4db0),
	.w8(32'h38a23974),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0db727),
	.w1(32'h39dcdab1),
	.w2(32'h3acc5a4b),
	.w3(32'hb9864261),
	.w4(32'hb9b33bb4),
	.w5(32'h3aba8496),
	.w6(32'hb9a0ac97),
	.w7(32'hba18be7e),
	.w8(32'h3ad2ce87),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980d19f),
	.w1(32'h39338189),
	.w2(32'h394d3bbb),
	.w3(32'h39bd8361),
	.w4(32'h39b95418),
	.w5(32'h39cdafea),
	.w6(32'h3980fda6),
	.w7(32'h39492664),
	.w8(32'h397d6fbd),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5c11b),
	.w1(32'hba039bd2),
	.w2(32'hba1368e1),
	.w3(32'h39f958e9),
	.w4(32'hb86c4fd3),
	.w5(32'hb9ae8bc6),
	.w6(32'hb96d7afd),
	.w7(32'hba2114a1),
	.w8(32'hba1fafbf),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a6ccd7),
	.w1(32'hb933fd53),
	.w2(32'h383d2582),
	.w3(32'hb919c230),
	.w4(32'hb9f128c7),
	.w5(32'hb71c3f73),
	.w6(32'h38c9c3f3),
	.w7(32'h399dec06),
	.w8(32'hb58bf864),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb855361f),
	.w1(32'h3996dbe4),
	.w2(32'hb7fc6708),
	.w3(32'h3999f081),
	.w4(32'h399d6880),
	.w5(32'h38e9eaab),
	.w6(32'h39939edd),
	.w7(32'h38be6f95),
	.w8(32'h392309fb),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb8a2e),
	.w1(32'h3afc2325),
	.w2(32'h3b246735),
	.w3(32'h3abd98b3),
	.w4(32'h3b072370),
	.w5(32'h3b1051ac),
	.w6(32'h392c6880),
	.w7(32'h3a789613),
	.w8(32'hb9205d67),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba591c),
	.w1(32'h3b82f0b1),
	.w2(32'h3b413767),
	.w3(32'h3bffcc7a),
	.w4(32'h3bd0af82),
	.w5(32'h3b22ffad),
	.w6(32'h3bbfb72b),
	.w7(32'h3b91bc33),
	.w8(32'h3b197742),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a668505),
	.w1(32'hb618d6fd),
	.w2(32'h3915cd6e),
	.w3(32'h3a1de069),
	.w4(32'hb9297b55),
	.w5(32'h399b57a5),
	.w6(32'h388236b3),
	.w7(32'h39873c7b),
	.w8(32'h3a1572ff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b912ed9),
	.w1(32'h3a1e6cab),
	.w2(32'h3bc4527d),
	.w3(32'h3b492288),
	.w4(32'hba07f57b),
	.w5(32'h3b50662f),
	.w6(32'h3af031e0),
	.w7(32'hbb08136c),
	.w8(32'h3b032fa8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c6768),
	.w1(32'h3a2ebf57),
	.w2(32'h39e6e090),
	.w3(32'hba3b6ae3),
	.w4(32'h3a173fde),
	.w5(32'h379cf2ff),
	.w6(32'h39799c34),
	.w7(32'h38d1f6c2),
	.w8(32'hb92eb3ad),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1a48c),
	.w1(32'h3ac91b38),
	.w2(32'h3913ac1d),
	.w3(32'h3b76289e),
	.w4(32'h39c4c781),
	.w5(32'hba397b02),
	.w6(32'h3afb8463),
	.w7(32'hb9fb4bd4),
	.w8(32'hbae69f46),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78897e),
	.w1(32'h3b01d91a),
	.w2(32'h3bd57d17),
	.w3(32'h3b5e4762),
	.w4(32'h3aa86ec1),
	.w5(32'h3b9bc42b),
	.w6(32'h3b20ead6),
	.w7(32'hb93afee1),
	.w8(32'h3b1fce28),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90009e3),
	.w1(32'h3ab9a854),
	.w2(32'h3b536652),
	.w3(32'hb93ff3d6),
	.w4(32'h3ac74d9c),
	.w5(32'h3b25aff4),
	.w6(32'h3a2a54c1),
	.w7(32'h3a6ebcb2),
	.w8(32'h3b2376be),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b1201),
	.w1(32'h39002ae3),
	.w2(32'h3af540e4),
	.w3(32'h3b02f302),
	.w4(32'hbb0adf3d),
	.w5(32'hb92db20d),
	.w6(32'hb9b8763d),
	.w7(32'hbb21d192),
	.w8(32'h3950fd69),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b585e1b),
	.w1(32'h3b35617c),
	.w2(32'h3bc2a223),
	.w3(32'h3adeaa4c),
	.w4(32'hb9fc62e6),
	.w5(32'h3b7006fc),
	.w6(32'h3ad89eab),
	.w7(32'hb9c71f08),
	.w8(32'h3b48f24c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f33336),
	.w1(32'hb6f0f98c),
	.w2(32'hb625e291),
	.w3(32'h398f10ed),
	.w4(32'h37f87bb6),
	.w5(32'hb93105b1),
	.w6(32'h38e5f35f),
	.w7(32'h3a056c83),
	.w8(32'hb8412158),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0bcbd),
	.w1(32'h3b55ffea),
	.w2(32'h3bb3156a),
	.w3(32'h3b90aeec),
	.w4(32'h3acb6b8e),
	.w5(32'h3b48defa),
	.w6(32'h3b4a24c5),
	.w7(32'hb9c90b76),
	.w8(32'hba3c07c0),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22efe4),
	.w1(32'h3b2fee26),
	.w2(32'h3b98f069),
	.w3(32'h3b064b48),
	.w4(32'h3afc8f35),
	.w5(32'h3b5111be),
	.w6(32'h3aadfa1a),
	.w7(32'h3933476c),
	.w8(32'h3a867f78),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39909e7d),
	.w1(32'h39371770),
	.w2(32'h39750a7f),
	.w3(32'h396cac4e),
	.w4(32'h38c22fd3),
	.w5(32'h39aa164e),
	.w6(32'h3972424e),
	.w7(32'h39890f98),
	.w8(32'h39aaf5ed),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397dd4ee),
	.w1(32'hb9c88a9e),
	.w2(32'hb9c7465d),
	.w3(32'h39a1f858),
	.w4(32'hb9a9722e),
	.w5(32'hb99e2b51),
	.w6(32'hba05c5e2),
	.w7(32'hb9fc8674),
	.w8(32'hba1a2c3f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86d632),
	.w1(32'hb98aed3a),
	.w2(32'h3a573aa1),
	.w3(32'hba58c03b),
	.w4(32'hba185378),
	.w5(32'h38875658),
	.w6(32'hb9ecdf60),
	.w7(32'hba5a6e58),
	.w8(32'h39a2cacc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec8a7d),
	.w1(32'h398dc431),
	.w2(32'h3b084d3c),
	.w3(32'h3b80f415),
	.w4(32'hbab1beb4),
	.w5(32'h3a8d5c69),
	.w6(32'h3b278487),
	.w7(32'hbb306964),
	.w8(32'hbad246b6),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9de293),
	.w1(32'h3a4e7f40),
	.w2(32'h3bae6755),
	.w3(32'h3937a17e),
	.w4(32'hba670bc3),
	.w5(32'h3b46ccc2),
	.w6(32'h3a588ba5),
	.w7(32'hbb22a5bb),
	.w8(32'h3ac1fda0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ade7530),
	.w1(32'hbb04aff4),
	.w2(32'h3b041781),
	.w3(32'h3b1101ab),
	.w4(32'hbb211c70),
	.w5(32'h3aa9f0d5),
	.w6(32'h3a51dead),
	.w7(32'hbb732ba3),
	.w8(32'h3a44940a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ff685),
	.w1(32'h3974f022),
	.w2(32'h3a128b45),
	.w3(32'hb90a119c),
	.w4(32'hb679a921),
	.w5(32'h3a0e85b0),
	.w6(32'h3a01d270),
	.w7(32'h39e539ca),
	.w8(32'h3a43a80a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b9fb4),
	.w1(32'h39987be1),
	.w2(32'h39579eea),
	.w3(32'h37ccc03c),
	.w4(32'h399d40aa),
	.w5(32'h39c528ae),
	.w6(32'h399e8b02),
	.w7(32'h39b9962c),
	.w8(32'h39553d41),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbbcb4),
	.w1(32'hbb0ead52),
	.w2(32'h3aea1600),
	.w3(32'hbb3d5d6f),
	.w4(32'h39d6199b),
	.w5(32'h3b5d0114),
	.w6(32'hbb6677a3),
	.w7(32'hba07cc26),
	.w8(32'h3af195aa),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa76ed7),
	.w1(32'hba7905fd),
	.w2(32'hbad75072),
	.w3(32'h3ac0dbd6),
	.w4(32'hb98ab4c5),
	.w5(32'hba811989),
	.w6(32'h3a8110d6),
	.w7(32'hb82b3644),
	.w8(32'hba58f7e9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2f294),
	.w1(32'hbb8a8ae4),
	.w2(32'h3b0ae987),
	.w3(32'hbad73991),
	.w4(32'hbad74022),
	.w5(32'h3b81dac8),
	.w6(32'hbab9d67b),
	.w7(32'hbb28796e),
	.w8(32'h3b82dfef),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cfd78),
	.w1(32'hb861e1a5),
	.w2(32'hb95d69fd),
	.w3(32'hb9c83aaa),
	.w4(32'h37f581f1),
	.w5(32'hb8a78f1b),
	.w6(32'hb8b6e4fe),
	.w7(32'hb91ce0c9),
	.w8(32'hb9768337),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb932496e),
	.w1(32'h3914f03d),
	.w2(32'h38e3f07a),
	.w3(32'hb7d323c8),
	.w4(32'h39382496),
	.w5(32'h391f89e6),
	.w6(32'h38f83206),
	.w7(32'h39184a68),
	.w8(32'hb7f63437),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9479e7),
	.w1(32'h38d707bb),
	.w2(32'h3b138e54),
	.w3(32'h39540475),
	.w4(32'hba2ab955),
	.w5(32'h3aa9ac44),
	.w6(32'hb8a0ae3c),
	.w7(32'hba57925c),
	.w8(32'h3a3afd8b),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd8371),
	.w1(32'h39c63330),
	.w2(32'h3a00f37b),
	.w3(32'h3abf24da),
	.w4(32'hb9791474),
	.w5(32'h3a304cd9),
	.w6(32'h3a982a63),
	.w7(32'hb95baa91),
	.w8(32'h3a082c08),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10000c),
	.w1(32'h39095e70),
	.w2(32'hba0d931e),
	.w3(32'h3a3fe85a),
	.w4(32'h39e8cfa6),
	.w5(32'hb8d37973),
	.w6(32'h39dfafe0),
	.w7(32'h38d8e03e),
	.w8(32'hb9fd5aca),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a28dcd7),
	.w1(32'h3aa9ac4f),
	.w2(32'h3b02e7d8),
	.w3(32'h39f9fbac),
	.w4(32'h3a9b2793),
	.w5(32'h3af1f2da),
	.w6(32'h37e5e38d),
	.w7(32'h390f13bb),
	.w8(32'hb98a4b8f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b5249),
	.w1(32'h3aa03e82),
	.w2(32'h3b4fccdf),
	.w3(32'h3b9aedd5),
	.w4(32'hbb9ab836),
	.w5(32'hba830435),
	.w6(32'h3b13cdb6),
	.w7(32'hbbcc99ef),
	.w8(32'hb996a74d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad38376),
	.w1(32'hbb43adc1),
	.w2(32'h3a575109),
	.w3(32'h3a861e21),
	.w4(32'hbbab2c63),
	.w5(32'hb9c064f2),
	.w6(32'hb986bd05),
	.w7(32'hbbb2d735),
	.w8(32'h3a16f45d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19951a),
	.w1(32'hbb942020),
	.w2(32'hbb0211a5),
	.w3(32'h3b060354),
	.w4(32'hbad9d8a0),
	.w5(32'h3b03d8e1),
	.w6(32'h3a381987),
	.w7(32'hbab69b5a),
	.w8(32'h3b479c7c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24e341),
	.w1(32'hb9ea93ae),
	.w2(32'h3a243369),
	.w3(32'h3a0515d8),
	.w4(32'hba47530d),
	.w5(32'h39cfc637),
	.w6(32'hb722e4e7),
	.w7(32'hba486cb4),
	.w8(32'h394441cc),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f636d1),
	.w1(32'hb898ae50),
	.w2(32'hb983881d),
	.w3(32'h39a70669),
	.w4(32'hb8e4163d),
	.w5(32'hb97792a1),
	.w6(32'hb8f242bf),
	.w7(32'hb8f9196c),
	.w8(32'h38a1c334),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8073507),
	.w1(32'h39c7aea2),
	.w2(32'h393cc14b),
	.w3(32'hb94aae08),
	.w4(32'h39babe78),
	.w5(32'h397c2826),
	.w6(32'h38677796),
	.w7(32'hb90d1d80),
	.w8(32'hb937455c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a621ee2),
	.w1(32'hba0cb260),
	.w2(32'hb9337b06),
	.w3(32'h3a586b7f),
	.w4(32'h390d208f),
	.w5(32'h3a1b9d28),
	.w6(32'h3a37a1ad),
	.w7(32'hb8a0e3ef),
	.w8(32'h3a6ea2e3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b844d97),
	.w1(32'h3ad5f009),
	.w2(32'h3bbd89cc),
	.w3(32'h3b726039),
	.w4(32'h38b5d367),
	.w5(32'h3b36fa35),
	.w6(32'h3b29c649),
	.w7(32'hba6c93d0),
	.w8(32'h3a66d55c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b1926),
	.w1(32'hbaa60c7f),
	.w2(32'h3b4e175e),
	.w3(32'h39273af1),
	.w4(32'hbb04b1d2),
	.w5(32'h3af93f68),
	.w6(32'hb9e52d36),
	.w7(32'hbb83bc26),
	.w8(32'h3a2e0010),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fc095),
	.w1(32'hb97a647f),
	.w2(32'h3b83d814),
	.w3(32'h3b02b1e9),
	.w4(32'hbabaa43f),
	.w5(32'h3b1b40db),
	.w6(32'h39bab6f9),
	.w7(32'hbb8c51f2),
	.w8(32'h39bdac68),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a69c2),
	.w1(32'h3908908e),
	.w2(32'h3b4724f5),
	.w3(32'h3afc307c),
	.w4(32'hbaf3f5a7),
	.w5(32'h3aa54be6),
	.w6(32'hb96d93f7),
	.w7(32'hbb4dc4e8),
	.w8(32'hb8b373e3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bf6c4),
	.w1(32'h3b8d604a),
	.w2(32'h3bf518a5),
	.w3(32'h3b6012fd),
	.w4(32'h3b66e07b),
	.w5(32'h3b9ad08a),
	.w6(32'h3ab14070),
	.w7(32'h3a648708),
	.w8(32'h3ac317f4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a486e9),
	.w1(32'hb774241e),
	.w2(32'hb8baa1ab),
	.w3(32'hb9474027),
	.w4(32'hb90a380c),
	.w5(32'hb8a29fc6),
	.w6(32'h3886b368),
	.w7(32'hb806d5c0),
	.w8(32'hb97888e0),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385f0a69),
	.w1(32'h3a364cb1),
	.w2(32'h3a24fddc),
	.w3(32'hb9227a98),
	.w4(32'h3a33b023),
	.w5(32'h3a496c02),
	.w6(32'h3a163686),
	.w7(32'h3a42cb4f),
	.w8(32'h3a655fdb),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a688610),
	.w1(32'hb947a7f9),
	.w2(32'hb9c8d446),
	.w3(32'h3a4ff6b2),
	.w4(32'hb9625867),
	.w5(32'hb99deb2f),
	.w6(32'hba165b85),
	.w7(32'hb9b82f18),
	.w8(32'hb9b91988),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af39520),
	.w1(32'h390cbe78),
	.w2(32'h3b08d515),
	.w3(32'h3a80fac2),
	.w4(32'h39b75cb4),
	.w5(32'h3ab9d160),
	.w6(32'h38d410a5),
	.w7(32'hbad49e85),
	.w8(32'h39150eed),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3872175c),
	.w1(32'hb9ed5fdd),
	.w2(32'hb7aad6a7),
	.w3(32'h3775e70e),
	.w4(32'hb9b54d97),
	.w5(32'h39700170),
	.w6(32'hb8e1ee3f),
	.w7(32'hba3a6ec5),
	.w8(32'hb8327f5f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7cbbf),
	.w1(32'h3b4e63cf),
	.w2(32'h3bf6e4f6),
	.w3(32'h3b643a48),
	.w4(32'h3a9a1a2a),
	.w5(32'h3b85a183),
	.w6(32'h3ac5e92b),
	.w7(32'hba5a22f4),
	.w8(32'h3a25e0c0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d60a46),
	.w1(32'hb96fdd71),
	.w2(32'h3876b324),
	.w3(32'h3a57e0d0),
	.w4(32'h3889e33f),
	.w5(32'hb8fc3dd2),
	.w6(32'h39576101),
	.w7(32'hba15c338),
	.w8(32'hb9f2bf8d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb980343d),
	.w1(32'hb91fb057),
	.w2(32'h36e1ed10),
	.w3(32'hb9cd83f6),
	.w4(32'h390e4803),
	.w5(32'h38d3b0c2),
	.w6(32'hb883919e),
	.w7(32'hb94fe0db),
	.w8(32'h3988205a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395805c4),
	.w1(32'h39594414),
	.w2(32'hb85fdec1),
	.w3(32'h399aa166),
	.w4(32'h39d9a8c5),
	.w5(32'h399a8aa5),
	.w6(32'h39944339),
	.w7(32'h39a3a30b),
	.w8(32'h39a53bd2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99dd45f),
	.w1(32'h39158b65),
	.w2(32'h39b2baf7),
	.w3(32'h39310cc1),
	.w4(32'h376796f5),
	.w5(32'h3a1aa1b1),
	.w6(32'h396e5ec3),
	.w7(32'h39ec1edb),
	.w8(32'h37d25e45),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939a703),
	.w1(32'hb910bf3c),
	.w2(32'hba6971e3),
	.w3(32'h39567468),
	.w4(32'h3955d229),
	.w5(32'hb9b020ec),
	.w6(32'h39a97d31),
	.w7(32'hb975dd78),
	.w8(32'hb9720488),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c81fc6),
	.w1(32'h3a57bc7d),
	.w2(32'h3a51720a),
	.w3(32'h39d63939),
	.w4(32'h3a48a6eb),
	.w5(32'h3a57e6f0),
	.w6(32'h3a42ad29),
	.w7(32'h3a406fd3),
	.w8(32'h3a410ec8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b872118),
	.w1(32'h3b0b74cf),
	.w2(32'h3b2469b2),
	.w3(32'h3b5cae6c),
	.w4(32'h3a9c9224),
	.w5(32'h3b0ef9d0),
	.w6(32'h3b104d08),
	.w7(32'hb77357c4),
	.w8(32'h3a187da5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b9e1e),
	.w1(32'h3a8740da),
	.w2(32'h3b567049),
	.w3(32'h3af7eeed),
	.w4(32'h3a191e5b),
	.w5(32'h3aca47f8),
	.w6(32'h3b28d534),
	.w7(32'h3979570f),
	.w8(32'h3a4eab8a),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a584027),
	.w1(32'hb90e5c83),
	.w2(32'hb98a05c9),
	.w3(32'h3a6a121c),
	.w4(32'hb9c5e5e0),
	.w5(32'hb9401664),
	.w6(32'h382fc440),
	.w7(32'hb73b9693),
	.w8(32'h3946317a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c809ee),
	.w1(32'hba01490b),
	.w2(32'hba5a0e70),
	.w3(32'h3a27a571),
	.w4(32'hb9d05b4f),
	.w5(32'hba34298e),
	.w6(32'hb9c7aaaa),
	.w7(32'hba29cfcc),
	.w8(32'hb9f7613f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48ca77),
	.w1(32'h37e6c8fc),
	.w2(32'hb83f7895),
	.w3(32'hba2dd61b),
	.w4(32'h38e79016),
	.w5(32'h3890865f),
	.w6(32'h36fe8d1d),
	.w7(32'h368b7b5b),
	.w8(32'h3926f4fc),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394b20b4),
	.w1(32'h380bdd6d),
	.w2(32'hb817f098),
	.w3(32'h399f5c35),
	.w4(32'h37d8f6c2),
	.w5(32'hb82f37f5),
	.w6(32'hb923a7a0),
	.w7(32'h399d63ac),
	.w8(32'h386ecdea),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd67d63),
	.w1(32'h3ba3c6ba),
	.w2(32'h3c00fb25),
	.w3(32'h3b604a21),
	.w4(32'h3a81588f),
	.w5(32'h3af940be),
	.w6(32'h3b4bd0c2),
	.w7(32'h3a8a7dcd),
	.w8(32'hb9b0e7da),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e5c18),
	.w1(32'hba4a93cc),
	.w2(32'h3ad46c2f),
	.w3(32'h3b520ffc),
	.w4(32'hb8ec93b4),
	.w5(32'h3b27af7a),
	.w6(32'hba7c051f),
	.w7(32'hbb9f7e02),
	.w8(32'hba19c513),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b265c),
	.w1(32'hbaa7ed13),
	.w2(32'h3a23f210),
	.w3(32'h3b1cf3c0),
	.w4(32'hbb1be9e4),
	.w5(32'hbaa66c97),
	.w6(32'h3afdeb69),
	.w7(32'hbb859a4f),
	.w8(32'hbb797e0d),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a16b6),
	.w1(32'hbb07b1fc),
	.w2(32'h3bb25062),
	.w3(32'h3a2055d9),
	.w4(32'hbb3cbce6),
	.w5(32'h3b1bf955),
	.w6(32'hb8b4dfc6),
	.w7(32'hbba88229),
	.w8(32'h3b0dd69e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17ab7a),
	.w1(32'h38d2adc5),
	.w2(32'hb9137c81),
	.w3(32'h3a115742),
	.w4(32'h39a574e3),
	.w5(32'h390e9edc),
	.w6(32'h3867b0aa),
	.w7(32'hb87c6a45),
	.w8(32'hb907088b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a6af5e),
	.w1(32'h39c9c4df),
	.w2(32'h39833aaf),
	.w3(32'hb9108b4e),
	.w4(32'h3a0f265a),
	.w5(32'h39dfa8aa),
	.w6(32'h39ab55e3),
	.w7(32'h399afe4a),
	.w8(32'h39af4930),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fb68e),
	.w1(32'h3a11b929),
	.w2(32'h39f7f21c),
	.w3(32'h39f5b841),
	.w4(32'h3a263cfb),
	.w5(32'h3a131eca),
	.w6(32'h39faf902),
	.w7(32'h3a08ae7d),
	.w8(32'h3a031f67),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b028b41),
	.w1(32'h39f7db9d),
	.w2(32'h3a409ca9),
	.w3(32'h3aacce40),
	.w4(32'h398e9a9c),
	.w5(32'h3a436d1c),
	.w6(32'h3a00e469),
	.w7(32'hb98c7832),
	.w8(32'hb953e893),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6fd90),
	.w1(32'h39ccf631),
	.w2(32'h39386a20),
	.w3(32'h384f5137),
	.w4(32'h3a04e6c5),
	.w5(32'h39da2454),
	.w6(32'h39ae9f4f),
	.w7(32'h394361c1),
	.w8(32'h39478aaf),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b729f60),
	.w1(32'h3b0149d3),
	.w2(32'h3aed3b36),
	.w3(32'h3b3af90e),
	.w4(32'h3a5eea4d),
	.w5(32'h39c9a3bf),
	.w6(32'hb9775af2),
	.w7(32'hba672a71),
	.w8(32'hbac0d7d0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8049b),
	.w1(32'h3ba3fd58),
	.w2(32'h3b93e4d8),
	.w3(32'h3bac9e51),
	.w4(32'h3b594da8),
	.w5(32'h3b3761ae),
	.w6(32'h3b456bd8),
	.w7(32'h39f29e53),
	.w8(32'h3abfb952),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19bced),
	.w1(32'h3ab26154),
	.w2(32'h3b882c5f),
	.w3(32'h3b506744),
	.w4(32'h3a8f02c9),
	.w5(32'h3b5e6574),
	.w6(32'h3abc917f),
	.w7(32'hba011b2c),
	.w8(32'h3b0600d1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5d4c5),
	.w1(32'hb98dad7c),
	.w2(32'h3b01b0fd),
	.w3(32'h3a81c9f6),
	.w4(32'hbaa067fa),
	.w5(32'h38851aef),
	.w6(32'h3a3482cd),
	.w7(32'hbaa084b6),
	.w8(32'hba681760),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1220f),
	.w1(32'h3ac32333),
	.w2(32'h3b3ae236),
	.w3(32'h3a52c415),
	.w4(32'h3a792d34),
	.w5(32'h3b07d6d7),
	.w6(32'h39b53400),
	.w7(32'h391dfc71),
	.w8(32'h39ef57f0),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397387ca),
	.w1(32'hba9d9688),
	.w2(32'h39fd8ce5),
	.w3(32'h393f181e),
	.w4(32'hba90df6c),
	.w5(32'h373ef2ca),
	.w6(32'hba3bc06b),
	.w7(32'hbafba050),
	.w8(32'hba04e38f),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a881d64),
	.w1(32'h3a804534),
	.w2(32'h3b186e11),
	.w3(32'h3a7e93f5),
	.w4(32'h3ab4ac11),
	.w5(32'h3b066d5e),
	.w6(32'h3a61d04c),
	.w7(32'hb9261fb1),
	.w8(32'h388728cf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37be7a88),
	.w1(32'hb9bbb3b8),
	.w2(32'hb9b8ac99),
	.w3(32'h395c039a),
	.w4(32'hb960fc7f),
	.w5(32'hb94d05fb),
	.w6(32'hb9817508),
	.w7(32'hb9c86bd7),
	.w8(32'hb93384ea),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb900c211),
	.w1(32'h3988e1ef),
	.w2(32'h386c474c),
	.w3(32'hb91af963),
	.w4(32'h39c12d78),
	.w5(32'h397dbb63),
	.w6(32'h3993a5b7),
	.w7(32'h392cc732),
	.w8(32'h3933b237),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e318e6),
	.w1(32'hb8e8e1a1),
	.w2(32'h361eab76),
	.w3(32'h39a1c913),
	.w4(32'h3944b591),
	.w5(32'hb7e050ca),
	.w6(32'hb9805d5c),
	.w7(32'hb9883283),
	.w8(32'hb8611277),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b8420),
	.w1(32'hb92fd276),
	.w2(32'hb96b172f),
	.w3(32'hb91d384f),
	.w4(32'h38583a32),
	.w5(32'h38675510),
	.w6(32'hb90555ad),
	.w7(32'hb8a699b9),
	.w8(32'h3857ac38),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7310),
	.w1(32'hbac752fd),
	.w2(32'h39ee7b47),
	.w3(32'h3a930802),
	.w4(32'hbb2f9ae0),
	.w5(32'hb99afac1),
	.w6(32'h38666a56),
	.w7(32'hbb619c21),
	.w8(32'h3975d763),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854a479),
	.w1(32'hb9c69676),
	.w2(32'hba07ff85),
	.w3(32'h39920113),
	.w4(32'h38ff1acb),
	.w5(32'hb944a5d3),
	.w6(32'h3a08a0c2),
	.w7(32'hb8582922),
	.w8(32'hb95e3ccd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25e178),
	.w1(32'hba83b868),
	.w2(32'h3a60a946),
	.w3(32'hb9e4646d),
	.w4(32'hbaa8aec3),
	.w5(32'h3a1958a6),
	.w6(32'hba6f3aa8),
	.w7(32'hbb3cdada),
	.w8(32'hb97b8474),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb84083),
	.w1(32'h3adbfda7),
	.w2(32'h3b02fa5d),
	.w3(32'h3b683aea),
	.w4(32'h3984c621),
	.w5(32'h39ed3a97),
	.w6(32'h3b3167da),
	.w7(32'hba282acb),
	.w8(32'hba9e76ed),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb049fea),
	.w1(32'hbb34227e),
	.w2(32'hba9116f1),
	.w3(32'hb76ece45),
	.w4(32'hba1d420c),
	.w5(32'h3adfbead),
	.w6(32'hba8af5d6),
	.w7(32'hbae23c25),
	.w8(32'h3a524687),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c005b88),
	.w1(32'h3bb18c33),
	.w2(32'h3b7edcff),
	.w3(32'h3bb2df6c),
	.w4(32'h3ad62bbe),
	.w5(32'h3b03cc33),
	.w6(32'h3b34a3dc),
	.w7(32'h3a5f08b3),
	.w8(32'h3ace1cd1),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb13877c),
	.w1(32'hbb02b9e8),
	.w2(32'hba17ddee),
	.w3(32'hba383810),
	.w4(32'hba6c51dd),
	.w5(32'h39ba48be),
	.w6(32'hbae5ce54),
	.w7(32'hbb1eeeb8),
	.w8(32'hbae8b9f4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63b34d),
	.w1(32'hb93504c3),
	.w2(32'h3b6d30e6),
	.w3(32'h3adc4033),
	.w4(32'hbb1ea81b),
	.w5(32'h38193362),
	.w6(32'h38616f4e),
	.w7(32'hbb539f8b),
	.w8(32'hbac385fa),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5b9f96),
	.w1(32'hba9d49a8),
	.w2(32'h3a297441),
	.w3(32'hbae86417),
	.w4(32'hbb4fd3a8),
	.w5(32'hb91cff02),
	.w6(32'hbaf2bfd7),
	.w7(32'hbb710326),
	.w8(32'hba5d59c7),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad7407),
	.w1(32'hba843e9e),
	.w2(32'h3b1c3f45),
	.w3(32'h39b93db5),
	.w4(32'hbada993b),
	.w5(32'h3b23f7ef),
	.w6(32'hba023811),
	.w7(32'hbb3606d4),
	.w8(32'h3adf7913),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb977da61),
	.w1(32'hba1dcbca),
	.w2(32'hba398469),
	.w3(32'hba6ebe92),
	.w4(32'hba69b787),
	.w5(32'hba4876bb),
	.w6(32'hba2b0ad9),
	.w7(32'hba4ab127),
	.w8(32'hb9cec7b8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ea934),
	.w1(32'h3aaa41d4),
	.w2(32'h3b9b90c6),
	.w3(32'h3a73bcce),
	.w4(32'hba0abdaf),
	.w5(32'h3b092c54),
	.w6(32'h3a52ce26),
	.w7(32'hbafffb2b),
	.w8(32'h3a55cf30),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9edc60),
	.w1(32'h3ad2b4dd),
	.w2(32'h3b07bcd5),
	.w3(32'h3b04c790),
	.w4(32'hbac0deaa),
	.w5(32'hba82abbe),
	.w6(32'hbaaa24a2),
	.w7(32'hbb80736c),
	.w8(32'hbb6404d0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd53c55),
	.w1(32'hba348258),
	.w2(32'h39a5d0d2),
	.w3(32'h3bc91594),
	.w4(32'hbb30480c),
	.w5(32'h39cbc604),
	.w6(32'h3b1eaf9b),
	.w7(32'hbbc2e88f),
	.w8(32'hbadd31df),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b9406),
	.w1(32'hbbe001b2),
	.w2(32'hbb9f48df),
	.w3(32'h3a6aaf71),
	.w4(32'hbbe3a4bc),
	.w5(32'hbb849350),
	.w6(32'hba1a511b),
	.w7(32'hbbd8d3b8),
	.w8(32'hbb456d6a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb7020),
	.w1(32'hba8ded55),
	.w2(32'h3ba3d9ed),
	.w3(32'hba37ed59),
	.w4(32'hba94f53a),
	.w5(32'h3b76aaf5),
	.w6(32'h3a17e965),
	.w7(32'hbb070ec0),
	.w8(32'h3b532896),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc6b67),
	.w1(32'h3b0af586),
	.w2(32'h3b0bec83),
	.w3(32'h3b8fd17f),
	.w4(32'hb9a1d687),
	.w5(32'hba235418),
	.w6(32'h3b1232cb),
	.w7(32'hbb40d2db),
	.w8(32'hbb101cd8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad12925),
	.w1(32'h38329b5f),
	.w2(32'hba40d4a4),
	.w3(32'h3aa8d5c8),
	.w4(32'h37b1aab1),
	.w5(32'hba143555),
	.w6(32'hb98f0590),
	.w7(32'hb9d5ed2b),
	.w8(32'hba08f2b1),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17fd90),
	.w1(32'h3b5dc783),
	.w2(32'h3bb05f85),
	.w3(32'h3bb31562),
	.w4(32'hba2b48b9),
	.w5(32'h3b89dd2f),
	.w6(32'h3b0520e5),
	.w7(32'hbb881954),
	.w8(32'h3a8bbdde),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b77a3a6),
	.w1(32'h3ad42d18),
	.w2(32'h3b3d3647),
	.w3(32'h3b6c27d6),
	.w4(32'h3b01ae8c),
	.w5(32'h3b2f3bdd),
	.w6(32'h3b15202c),
	.w7(32'h3a9eba2d),
	.w8(32'h3ac48754),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913a688),
	.w1(32'h359c0be7),
	.w2(32'h38c6e9d6),
	.w3(32'h392bdddf),
	.w4(32'h389acc54),
	.w5(32'h392a7932),
	.w6(32'hb97eaf78),
	.w7(32'hb96c95ca),
	.w8(32'hb86c1e7d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa56a4f),
	.w1(32'h3a74b23b),
	.w2(32'h3a477386),
	.w3(32'h3a513754),
	.w4(32'h392856f2),
	.w5(32'h39c73f1b),
	.w6(32'hb6b23131),
	.w7(32'hba259fcd),
	.w8(32'hb9810ed4),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39710e39),
	.w1(32'h3b00a0b0),
	.w2(32'h3bbb3e78),
	.w3(32'h39a64378),
	.w4(32'h3a988318),
	.w5(32'h3b875ee8),
	.w6(32'h3af3364d),
	.w7(32'h3a97729c),
	.w8(32'h3b837466),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05a499),
	.w1(32'hbae5ffa0),
	.w2(32'h3afafea0),
	.w3(32'h3a32a71b),
	.w4(32'hba95fdf8),
	.w5(32'h3b0bb276),
	.w6(32'hba0cf6a7),
	.w7(32'hbafac271),
	.w8(32'h3ab94bfa),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23df7b),
	.w1(32'hba0f5f64),
	.w2(32'h3aa489b7),
	.w3(32'hb9d5e586),
	.w4(32'hba9de665),
	.w5(32'h3a8cddc2),
	.w6(32'h3991f084),
	.w7(32'hbacbe5f7),
	.w8(32'h3a9431b7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ca1b98),
	.w1(32'hbafbe159),
	.w2(32'h391cf30d),
	.w3(32'hb829a8fb),
	.w4(32'hbb10df09),
	.w5(32'h3958f207),
	.w6(32'hb9ef1b64),
	.w7(32'hbacfb8dc),
	.w8(32'h39f340d3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa64337),
	.w1(32'hba01d11d),
	.w2(32'h39f1889b),
	.w3(32'h3adce919),
	.w4(32'hb8cd8bc6),
	.w5(32'h3a8b92a4),
	.w6(32'h39ef29a9),
	.w7(32'hbad7d856),
	.w8(32'hbaaca9ee),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33da85),
	.w1(32'h3af240ff),
	.w2(32'h3b654ca6),
	.w3(32'h3a8eee6c),
	.w4(32'hb946d604),
	.w5(32'h3ab9d112),
	.w6(32'h3b08cbdd),
	.w7(32'h39de866b),
	.w8(32'h3aa73be1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399d7a9e),
	.w1(32'hb968b7bd),
	.w2(32'h3ae1480c),
	.w3(32'h3a04b857),
	.w4(32'hb957211d),
	.w5(32'h3acb7ad6),
	.w6(32'h3a32e57a),
	.w7(32'hba57e039),
	.w8(32'h3a8793ea),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f7901),
	.w1(32'h3a7d9db4),
	.w2(32'h3a664d4e),
	.w3(32'h3a52c095),
	.w4(32'h3a8232b7),
	.w5(32'h3a655a2a),
	.w6(32'h3a8502f5),
	.w7(32'h3a7deb00),
	.w8(32'h3a895306),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abff2a2),
	.w1(32'h3a61bfee),
	.w2(32'h3a50a054),
	.w3(32'h3ab52a41),
	.w4(32'h3a51d228),
	.w5(32'h3a3293fd),
	.w6(32'h3a7100f2),
	.w7(32'h3a635500),
	.w8(32'h3a5fceaf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd3b6e),
	.w1(32'h39e8dfcd),
	.w2(32'h39ef8df9),
	.w3(32'h3a388650),
	.w4(32'h3a1415f5),
	.w5(32'h3a155f32),
	.w6(32'h3a196a28),
	.w7(32'h39e4055f),
	.w8(32'h3a0b28d4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a125d7a),
	.w1(32'h3914f40f),
	.w2(32'h399982d5),
	.w3(32'h3a3962df),
	.w4(32'h3982a556),
	.w5(32'h38c7493d),
	.w6(32'h388fee59),
	.w7(32'h394a3413),
	.w8(32'h38c880c5),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b91a4),
	.w1(32'hba5c00aa),
	.w2(32'h3af68a14),
	.w3(32'h3a51f905),
	.w4(32'hbaaaecc6),
	.w5(32'h3a8eff89),
	.w6(32'hb6446f4d),
	.w7(32'hbaf9f6d0),
	.w8(32'h39cd4a07),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4781d),
	.w1(32'h39e9c43b),
	.w2(32'h39b4c0d5),
	.w3(32'h3947476a),
	.w4(32'h390992a5),
	.w5(32'h3933da5f),
	.w6(32'h393a87fc),
	.w7(32'h37d8c256),
	.w8(32'hb8823420),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae239dd),
	.w1(32'h3aa7aedf),
	.w2(32'h3b03f0ad),
	.w3(32'h3ac089a0),
	.w4(32'h3a421d5b),
	.w5(32'h3aa2ec0a),
	.w6(32'h3a45cabc),
	.w7(32'h38ff6800),
	.w8(32'hb98051e6),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5be04),
	.w1(32'hba50b95b),
	.w2(32'h3b2a6fed),
	.w3(32'h38f8925e),
	.w4(32'hb8d8d6ec),
	.w5(32'h3b4041b8),
	.w6(32'h39d7a0c7),
	.w7(32'hba0ec14b),
	.w8(32'h3b911462),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4800ea),
	.w1(32'h37eec3bd),
	.w2(32'h39b2e0a4),
	.w3(32'h3a5abc84),
	.w4(32'hb934207b),
	.w5(32'hb988d6c8),
	.w6(32'hb9dc104c),
	.w7(32'hb936b990),
	.w8(32'hb89f5573),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787c2f2),
	.w1(32'hb991b82b),
	.w2(32'hba4715ea),
	.w3(32'hb9c2beed),
	.w4(32'hb9dfc925),
	.w5(32'hba441ebf),
	.w6(32'hb9baef18),
	.w7(32'hba14248b),
	.w8(32'hb9a4052c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f7b029),
	.w1(32'hb92ebf69),
	.w2(32'hb986ce70),
	.w3(32'hb9bbd8d2),
	.w4(32'hb86ff08e),
	.w5(32'hb8ea13bf),
	.w6(32'hb9428aff),
	.w7(32'hb9555e68),
	.w8(32'hb993bc64),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb648b),
	.w1(32'hba29f19c),
	.w2(32'hb9d20588),
	.w3(32'hb987a1fc),
	.w4(32'hbac9a295),
	.w5(32'hbb5d3896),
	.w6(32'hbab92cf8),
	.w7(32'hbaf389d9),
	.w8(32'hb9f5b89d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3494c),
	.w1(32'h3b33f34c),
	.w2(32'h3a78e480),
	.w3(32'h3b155aeb),
	.w4(32'h3b82ef72),
	.w5(32'h3ae8ca8b),
	.w6(32'hb92c7278),
	.w7(32'hba840e3c),
	.w8(32'hba9811bb),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3da26c),
	.w1(32'h3b265405),
	.w2(32'h3bc4a6d9),
	.w3(32'h3b4f0da7),
	.w4(32'hba62497e),
	.w5(32'h3b357a2c),
	.w6(32'h3ad91265),
	.w7(32'h3a75ff5a),
	.w8(32'h3b4616d6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaba9e7),
	.w1(32'h39e4f2ef),
	.w2(32'h3a828cae),
	.w3(32'h3b2b5dd7),
	.w4(32'h3aa50987),
	.w5(32'h3b1c63c8),
	.w6(32'hb7fb37fa),
	.w7(32'h3a0da0d2),
	.w8(32'h39eee158),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44bf26),
	.w1(32'hb8c93700),
	.w2(32'h3934c452),
	.w3(32'h3b71b515),
	.w4(32'h3a95197c),
	.w5(32'h3afac6d9),
	.w6(32'h3a3021ae),
	.w7(32'h383d7f77),
	.w8(32'h39811dd4),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ce1ed0),
	.w1(32'h39d582cd),
	.w2(32'h3bb5f339),
	.w3(32'h3a9e35ca),
	.w4(32'hbb2c4409),
	.w5(32'hbb34052b),
	.w6(32'hba96fbff),
	.w7(32'hbaff6176),
	.w8(32'h3b034790),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9731af),
	.w1(32'h3b0b66a6),
	.w2(32'h3b46a1af),
	.w3(32'h39bc2f08),
	.w4(32'h3aec47a7),
	.w5(32'h3b5d1044),
	.w6(32'h3a8b94af),
	.w7(32'hba1b602e),
	.w8(32'h387050d0),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a855b68),
	.w1(32'h3a0a087b),
	.w2(32'h3b243d68),
	.w3(32'h3a6c174a),
	.w4(32'h3a730388),
	.w5(32'h3b246bdb),
	.w6(32'hba980645),
	.w7(32'hbaffbece),
	.w8(32'hb91e31ed),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbcbb9),
	.w1(32'h3b89d784),
	.w2(32'h3bcca10c),
	.w3(32'h3bd2f629),
	.w4(32'h3b718f92),
	.w5(32'h3bb6237a),
	.w6(32'h3ad0526c),
	.w7(32'h39d1d667),
	.w8(32'h3ae9d95b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad07e24),
	.w1(32'h3959186d),
	.w2(32'h3aed97f3),
	.w3(32'h3b69e441),
	.w4(32'h3a327258),
	.w5(32'h3b0872a3),
	.w6(32'h3ab12daa),
	.w7(32'hba5c2cb2),
	.w8(32'h3b3a56f4),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48ca19),
	.w1(32'h3a5b829a),
	.w2(32'hb904033a),
	.w3(32'h3b0e4944),
	.w4(32'hba755e04),
	.w5(32'hbb0bff4f),
	.w6(32'hba1c13f2),
	.w7(32'hbb5071c9),
	.w8(32'hba83f52a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b758313),
	.w1(32'hba5e8a3e),
	.w2(32'h3a7a9f5c),
	.w3(32'h3b5f5dcd),
	.w4(32'h39c6c38e),
	.w5(32'h3ad7a198),
	.w6(32'hba03bcf0),
	.w7(32'hbb887e0b),
	.w8(32'hbb22d506),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3c0983),
	.w1(32'h3aef873d),
	.w2(32'h3ab1b34c),
	.w3(32'h3a1f5c4e),
	.w4(32'h3b165865),
	.w5(32'hba4c2fee),
	.w6(32'h39b2fd20),
	.w7(32'hb9c4ae4f),
	.w8(32'hba7f3945),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d2d3d),
	.w1(32'hbadfb2da),
	.w2(32'h3a867361),
	.w3(32'h3bee5ffc),
	.w4(32'hbafe4ea8),
	.w5(32'h3981a726),
	.w6(32'hbacda646),
	.w7(32'hb9f6351d),
	.w8(32'h3b509294),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97953ab),
	.w1(32'hba2b509c),
	.w2(32'h39a67f21),
	.w3(32'h392363ca),
	.w4(32'hba79167e),
	.w5(32'hbad97b7d),
	.w6(32'hb9c2cada),
	.w7(32'hba765694),
	.w8(32'hb9e80d0f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7b562),
	.w1(32'hbb62dcd3),
	.w2(32'h3ab89471),
	.w3(32'hbb57d371),
	.w4(32'h39d411d2),
	.w5(32'h3b6d6af4),
	.w6(32'hba91b934),
	.w7(32'hbad63b5e),
	.w8(32'h3b85e590),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983e8c1),
	.w1(32'hbab6e98f),
	.w2(32'hbadefce3),
	.w3(32'hb966026f),
	.w4(32'hbb87fcc6),
	.w5(32'hbb827a71),
	.w6(32'hba321ed9),
	.w7(32'hbb344b92),
	.w8(32'hba717d01),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad39e38),
	.w1(32'h3a0ea7c9),
	.w2(32'hbaf13356),
	.w3(32'hbaa88dd3),
	.w4(32'h3a8b4887),
	.w5(32'hba47fcf9),
	.w6(32'h3a250beb),
	.w7(32'hba70e735),
	.w8(32'hba0516ae),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3901be19),
	.w1(32'h3a88f6ec),
	.w2(32'h3bca1f04),
	.w3(32'h3a47fbe1),
	.w4(32'h3b618831),
	.w5(32'h3c0f0e6c),
	.w6(32'hbb4baf9a),
	.w7(32'h3b0e08db),
	.w8(32'hbb5a86e0),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32ab73),
	.w1(32'h3a429155),
	.w2(32'hba8c3417),
	.w3(32'hbaa8c7c3),
	.w4(32'h3adde620),
	.w5(32'hb7cb8b8d),
	.w6(32'h3a67bb57),
	.w7(32'hba3fb5c6),
	.w8(32'hb96b9074),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a57461),
	.w1(32'hba85bff5),
	.w2(32'hba2662cb),
	.w3(32'h3a34c847),
	.w4(32'hbad9c857),
	.w5(32'hb6bb1a76),
	.w6(32'hba13dbda),
	.w7(32'hbb8b256a),
	.w8(32'hb84b55a9),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3c616),
	.w1(32'hb8c65f41),
	.w2(32'h3a547dd8),
	.w3(32'h3b68500c),
	.w4(32'h3a56268f),
	.w5(32'h3a312620),
	.w6(32'h3ac8379c),
	.w7(32'hbb0d0c68),
	.w8(32'h3a72f852),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ac2cc),
	.w1(32'h3a89abe9),
	.w2(32'h3b946f09),
	.w3(32'hb97e3849),
	.w4(32'hbaadc65d),
	.w5(32'h39e83ee5),
	.w6(32'hba4dfaec),
	.w7(32'h3aa3497b),
	.w8(32'hb982b775),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5deae6),
	.w1(32'hb8a0fa3f),
	.w2(32'h3b34698e),
	.w3(32'h3abe15f0),
	.w4(32'hbaf93413),
	.w5(32'h38e25cea),
	.w6(32'h39a6ee7a),
	.w7(32'hb9b5bc2b),
	.w8(32'h3b20df27),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed60af),
	.w1(32'h3aa23e67),
	.w2(32'h3c44bb0f),
	.w3(32'hbb3848c4),
	.w4(32'hbb889766),
	.w5(32'h3bbb247c),
	.w6(32'hbbf44483),
	.w7(32'h3941fce4),
	.w8(32'hbb1a9236),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c673c4b),
	.w1(32'h3bb7b828),
	.w2(32'h3ba4fecc),
	.w3(32'h3b8625f6),
	.w4(32'h3b6088db),
	.w5(32'h3b3746eb),
	.w6(32'h3b60f7cc),
	.w7(32'h3aa059ad),
	.w8(32'hb927516f),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d314a),
	.w1(32'hbb880ade),
	.w2(32'h3ba16279),
	.w3(32'hb98ab6fc),
	.w4(32'hbae97592),
	.w5(32'h3ba01d26),
	.w6(32'hbbcd711d),
	.w7(32'hbb9c6552),
	.w8(32'h3a8a34d5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71ddc2),
	.w1(32'hbb98f83d),
	.w2(32'hbae079e5),
	.w3(32'hba4a9e53),
	.w4(32'hba77c8a4),
	.w5(32'h3a892731),
	.w6(32'hbbd811b5),
	.w7(32'hbbe2d4fc),
	.w8(32'hba78a62e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80276ec),
	.w1(32'hbb10227f),
	.w2(32'hbb45ff37),
	.w3(32'hbb4cdac3),
	.w4(32'hbaa4187d),
	.w5(32'hbb2bdb0d),
	.w6(32'hbb1973f6),
	.w7(32'hbb2a2693),
	.w8(32'hbac0b3ef),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93fa8f),
	.w1(32'hbae5106b),
	.w2(32'h38b11ffc),
	.w3(32'h3906bb87),
	.w4(32'hbb27ebd7),
	.w5(32'hb9ec8267),
	.w6(32'hbadec934),
	.w7(32'hbb640118),
	.w8(32'hbaa0833c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba801525),
	.w1(32'hbb89e1f6),
	.w2(32'h3baf86dc),
	.w3(32'hbb070ff2),
	.w4(32'hbb10d9a3),
	.w5(32'h3baeed77),
	.w6(32'hbbcd5f6c),
	.w7(32'hba4180b7),
	.w8(32'hbb511c90),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad31941),
	.w1(32'hba1e9ce8),
	.w2(32'h3c55803d),
	.w3(32'h3b87e65c),
	.w4(32'h3896d4fa),
	.w5(32'h3c6a047c),
	.w6(32'h3a472ba4),
	.w7(32'h3c28e0fa),
	.w8(32'hbbc00eb5),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20300d),
	.w1(32'h3a8f2170),
	.w2(32'h3ac36ea7),
	.w3(32'hbbd29fbe),
	.w4(32'h39f99ef1),
	.w5(32'h39914e88),
	.w6(32'hb84b84e0),
	.w7(32'h3a1d96f9),
	.w8(32'h396b2e7a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842a438),
	.w1(32'hb9e1fb28),
	.w2(32'hb9c07311),
	.w3(32'h3829b6da),
	.w4(32'h37735517),
	.w5(32'hba61d810),
	.w6(32'hba9e9334),
	.w7(32'hba925856),
	.w8(32'hba04bbef),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c8cca),
	.w1(32'hba07a635),
	.w2(32'h3acc70a9),
	.w3(32'h3ade8d20),
	.w4(32'hb985ec20),
	.w5(32'h3aa125f6),
	.w6(32'hb9de88d7),
	.w7(32'hbaae974f),
	.w8(32'hbaaa2209),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1eed8b),
	.w1(32'h3ab5e4f8),
	.w2(32'hbb9dac61),
	.w3(32'hbaf83de9),
	.w4(32'hbaebd8a9),
	.w5(32'hbb36de00),
	.w6(32'h3b106bb5),
	.w7(32'hbaaff433),
	.w8(32'hbb29722e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a825c),
	.w1(32'hbb393771),
	.w2(32'hbb10b6de),
	.w3(32'h39ada77b),
	.w4(32'hb88901ff),
	.w5(32'hb7d998c3),
	.w6(32'hbaafada0),
	.w7(32'hbb52f143),
	.w8(32'hb922a7fd),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd359d),
	.w1(32'hba409b7f),
	.w2(32'hb83e526c),
	.w3(32'h3a0be7ff),
	.w4(32'hb9ebcda0),
	.w5(32'hbabf31ce),
	.w6(32'hbac02406),
	.w7(32'hb9b7027c),
	.w8(32'h38614a4e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8be416),
	.w1(32'hb9a8fc2c),
	.w2(32'hba9eca1a),
	.w3(32'h3af8e49a),
	.w4(32'h3a8ef129),
	.w5(32'h3a30aa5f),
	.w6(32'hb9bc9b2b),
	.w7(32'hb90ad9cb),
	.w8(32'hba850b2e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4ce39),
	.w1(32'h3a1772cc),
	.w2(32'h3a1f9568),
	.w3(32'hba088f8b),
	.w4(32'h3ab8bfe3),
	.w5(32'h3b2c1d7b),
	.w6(32'h3a20e225),
	.w7(32'h3ac1c471),
	.w8(32'h3a7f2b09),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefa5e1),
	.w1(32'h3a6dd443),
	.w2(32'h370652ba),
	.w3(32'h3ae3897e),
	.w4(32'h3abf8ccd),
	.w5(32'h39c50f4b),
	.w6(32'h3a391960),
	.w7(32'hb8fed2f0),
	.w8(32'h383e2886),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb0a7),
	.w1(32'hba3fc85c),
	.w2(32'h3ac3a274),
	.w3(32'h3a1246b2),
	.w4(32'hba58ada3),
	.w5(32'h3b1440e5),
	.w6(32'hb95e25d1),
	.w7(32'hbab488b8),
	.w8(32'hb7adbc54),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5829b9),
	.w1(32'h3b74f90c),
	.w2(32'h3ccd9c20),
	.w3(32'h3b8193bc),
	.w4(32'hbade2aca),
	.w5(32'h3cb375de),
	.w6(32'h3bb1b045),
	.w7(32'h3c72d185),
	.w8(32'hbb156dcb),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f29ad7),
	.w1(32'hba22c438),
	.w2(32'hbb1560cd),
	.w3(32'hbc07b382),
	.w4(32'h3ab410ab),
	.w5(32'h3a048547),
	.w6(32'h3ad4fc0b),
	.w7(32'h3a069c76),
	.w8(32'h3a0f1606),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecac4e),
	.w1(32'hbb68f9c7),
	.w2(32'h3aab3980),
	.w3(32'h3a8c668c),
	.w4(32'hbb3423f5),
	.w5(32'h3a12d36a),
	.w6(32'hbb187c5f),
	.w7(32'hbb2b45ee),
	.w8(32'h39ff3a15),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3b76),
	.w1(32'h38828c53),
	.w2(32'h3ab99259),
	.w3(32'hba987fb7),
	.w4(32'h3b5f3de7),
	.w5(32'h3b8652bb),
	.w6(32'h38d38666),
	.w7(32'hbab34ce0),
	.w8(32'hb903c81f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc75c45),
	.w1(32'h3b59bd49),
	.w2(32'h3bbccca0),
	.w3(32'h3bacf702),
	.w4(32'h3b184560),
	.w5(32'h3ba54e91),
	.w6(32'h3b3f0608),
	.w7(32'hbb0a5d0f),
	.w8(32'h39c9f237),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b64ed),
	.w1(32'hba609264),
	.w2(32'h3a8035c9),
	.w3(32'h3b2dc7fe),
	.w4(32'hba1cebb6),
	.w5(32'h395558e8),
	.w6(32'hb9ff6900),
	.w7(32'hbb36aa41),
	.w8(32'hba3368c9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28fb42),
	.w1(32'h3b3eb0a7),
	.w2(32'h3bf2a84c),
	.w3(32'h3b56bec5),
	.w4(32'h3ab8b72e),
	.w5(32'h3b86c4fa),
	.w6(32'h3b02d37b),
	.w7(32'h3ad31c9b),
	.w8(32'h3b453f14),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1807),
	.w1(32'h39c7c3e8),
	.w2(32'h3b3c44f9),
	.w3(32'h3acb261e),
	.w4(32'h3b85d8c7),
	.w5(32'h3bc1080c),
	.w6(32'hba87010d),
	.w7(32'h3aadb97a),
	.w8(32'hbb2f3737),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5c4a8),
	.w1(32'hbb36d79b),
	.w2(32'h39d6294e),
	.w3(32'h3bb482a2),
	.w4(32'hbb32be83),
	.w5(32'hbab968a4),
	.w6(32'hbb84149c),
	.w7(32'hbb6a1c23),
	.w8(32'hbb11fc1d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc9171),
	.w1(32'h3ad73285),
	.w2(32'h3a29f98a),
	.w3(32'hb8a4cd39),
	.w4(32'h3afe45d8),
	.w5(32'h3a929210),
	.w6(32'h3b113c86),
	.w7(32'h3aaf7715),
	.w8(32'h3a8e4cd7),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad78a0),
	.w1(32'h39892e73),
	.w2(32'h3b274817),
	.w3(32'h3af6de8a),
	.w4(32'h3a222cc9),
	.w5(32'h3b2d733c),
	.w6(32'h3a58fa7d),
	.w7(32'h3b179fae),
	.w8(32'h3aee4efe),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110a4a),
	.w1(32'hbaf9a3cc),
	.w2(32'hba5402c9),
	.w3(32'h3ad0fb48),
	.w4(32'h3a50ab29),
	.w5(32'h3b569ed2),
	.w6(32'hba9fba2d),
	.w7(32'hbad44109),
	.w8(32'h3b13af7e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce5e5c),
	.w1(32'h3b759f45),
	.w2(32'h3c03803a),
	.w3(32'h3b8d0d91),
	.w4(32'h3af8ca65),
	.w5(32'h3bd52a05),
	.w6(32'h3b35ab73),
	.w7(32'h3b719bae),
	.w8(32'h3b500c7e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8655cf),
	.w1(32'h3aa6f049),
	.w2(32'h3a5ab59c),
	.w3(32'h3b377f4a),
	.w4(32'h3ae57c12),
	.w5(32'h3b0dfe45),
	.w6(32'hbac24c55),
	.w7(32'hba321669),
	.w8(32'hba2c5193),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae52c92),
	.w1(32'hb9ea115a),
	.w2(32'h3b4d11fb),
	.w3(32'hb964b81d),
	.w4(32'h3995cb51),
	.w5(32'h3b353abf),
	.w6(32'hbaa41f40),
	.w7(32'h3aca9643),
	.w8(32'hbaa67a80),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7a98a),
	.w1(32'h3b22706a),
	.w2(32'h3c8e6470),
	.w3(32'hbb24463e),
	.w4(32'hbb9ae6be),
	.w5(32'h3bfdad67),
	.w6(32'h3be69b42),
	.w7(32'h3ca90b8b),
	.w8(32'h3b8d9ea6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91f37c),
	.w1(32'hba449234),
	.w2(32'h3b6eaa5b),
	.w3(32'hbc01e142),
	.w4(32'hbb980524),
	.w5(32'h3ac3c8b1),
	.w6(32'h3b2ef441),
	.w7(32'h3b510678),
	.w8(32'hbb4c1709),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fae057),
	.w1(32'h3a8ccc52),
	.w2(32'hba7ecb3a),
	.w3(32'hbb6a39d7),
	.w4(32'h3a2cfa7d),
	.w5(32'hba367d11),
	.w6(32'hba0fe283),
	.w7(32'hbbb0f476),
	.w8(32'h3afcd0bd),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa73d15),
	.w1(32'h3a5cb45e),
	.w2(32'h3a50483b),
	.w3(32'h3b52661c),
	.w4(32'h3ae12fdf),
	.w5(32'h3b20439b),
	.w6(32'h3a1afa04),
	.w7(32'h385dc2c9),
	.w8(32'h3a1dab31),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ac2d4),
	.w1(32'h3be62189),
	.w2(32'h3c2e1a85),
	.w3(32'h3c255753),
	.w4(32'h3bb7adf1),
	.w5(32'h3bef89ac),
	.w6(32'h3bad71be),
	.w7(32'h39beb4ec),
	.w8(32'h3ad395f2),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ca51),
	.w1(32'hba87decc),
	.w2(32'h3b62daff),
	.w3(32'h395b850e),
	.w4(32'hbb7ece06),
	.w5(32'h3b6503c1),
	.w6(32'hbba05f61),
	.w7(32'hbbdfae54),
	.w8(32'h39bd473c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7041b9),
	.w1(32'h3a670897),
	.w2(32'h3a1a7aa6),
	.w3(32'h3ad1e769),
	.w4(32'h3abd7231),
	.w5(32'h3a7beed5),
	.w6(32'h39303d28),
	.w7(32'h39f823e8),
	.w8(32'hb73dbea7),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba661773),
	.w1(32'hb939e904),
	.w2(32'hba698811),
	.w3(32'h398060c3),
	.w4(32'hbb00b606),
	.w5(32'hb90c4b6e),
	.w6(32'hba5080bd),
	.w7(32'hba7381e8),
	.w8(32'h388e3244),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2f7a),
	.w1(32'h39043994),
	.w2(32'hb8cae368),
	.w3(32'h3a4ebcbd),
	.w4(32'h3b2e58d9),
	.w5(32'h3b07552d),
	.w6(32'h399bd56b),
	.w7(32'hba2dc71d),
	.w8(32'hb97aeaca),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936af06),
	.w1(32'hbb0bb436),
	.w2(32'hbab439d6),
	.w3(32'h39fc27ad),
	.w4(32'hba8559c9),
	.w5(32'hbad4a7d9),
	.w6(32'hbadc67fa),
	.w7(32'hbaad27c5),
	.w8(32'hba8df558),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73e4d1),
	.w1(32'h38d8dd50),
	.w2(32'h3a47fc57),
	.w3(32'hb8daa71b),
	.w4(32'hba258f25),
	.w5(32'hbab19949),
	.w6(32'hbaac9f2d),
	.w7(32'hbab98ac2),
	.w8(32'h3a810048),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86a46b),
	.w1(32'h3bc46518),
	.w2(32'h3c75f62d),
	.w3(32'hb988f3cc),
	.w4(32'hba42dbff),
	.w5(32'h3c204323),
	.w6(32'h3beb0d85),
	.w7(32'h3c3b6674),
	.w8(32'h3bb7098e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c186159),
	.w1(32'h3baec253),
	.w2(32'h3cdd785b),
	.w3(32'h3a3835f2),
	.w4(32'hbb289237),
	.w5(32'h3ca5f009),
	.w6(32'hbb1f6daf),
	.w7(32'h3c206f09),
	.w8(32'h39fe9219),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c27dbee),
	.w1(32'h3a38c286),
	.w2(32'hb9d29298),
	.w3(32'h3aa2d07b),
	.w4(32'h3a91293c),
	.w5(32'h3a68be4f),
	.w6(32'h3aa0a5a0),
	.w7(32'h3932b2ae),
	.w8(32'hba23297f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bf960),
	.w1(32'hb8e98ab1),
	.w2(32'h3bad8ca0),
	.w3(32'h3b0cab93),
	.w4(32'hb937e9f4),
	.w5(32'h3b181c79),
	.w6(32'h3a4ce9fe),
	.w7(32'hba7bfa21),
	.w8(32'h3ba1ac9e),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86e4f9),
	.w1(32'h39efb0bd),
	.w2(32'hba1f8767),
	.w3(32'h3b9bcf04),
	.w4(32'h3af1d954),
	.w5(32'h3a973114),
	.w6(32'h3a639845),
	.w7(32'hb8e6f2a3),
	.w8(32'hba31de54),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7e4412),
	.w1(32'h3a29627c),
	.w2(32'h392ef1e8),
	.w3(32'h3a17d3ed),
	.w4(32'h399f6774),
	.w5(32'hb81a8cc0),
	.w6(32'hb7566bf4),
	.w7(32'h38bd991f),
	.w8(32'hb95f66f8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa82273),
	.w1(32'h3aa4ae46),
	.w2(32'h3a57574c),
	.w3(32'h3a80ab41),
	.w4(32'h3aa2173d),
	.w5(32'h3a5c496b),
	.w6(32'h3a838c61),
	.w7(32'h395b413a),
	.w8(32'h3a818497),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a070b96),
	.w1(32'hba565e56),
	.w2(32'hb8c99c69),
	.w3(32'h3aa84d58),
	.w4(32'hb9891bc2),
	.w5(32'hba50123e),
	.w6(32'hba8d025a),
	.w7(32'hb9216b69),
	.w8(32'h39a063ee),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62d0e1),
	.w1(32'hb8ac64fa),
	.w2(32'h3a9a01b9),
	.w3(32'h3ab99c85),
	.w4(32'h3a925985),
	.w5(32'h3b4fbfac),
	.w6(32'hba1a0636),
	.w7(32'hba8aa010),
	.w8(32'h3a1bfca9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b427b30),
	.w1(32'hbb90c72c),
	.w2(32'hba9cb6f1),
	.w3(32'h3b16d5ae),
	.w4(32'hbb9a4b05),
	.w5(32'hbb218740),
	.w6(32'hbb91ad0d),
	.w7(32'hbba887f2),
	.w8(32'h3a2a826b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad52a17),
	.w1(32'h384404b6),
	.w2(32'h3b1b9fd5),
	.w3(32'hbb35c63f),
	.w4(32'h3a0abd30),
	.w5(32'h3a92c179),
	.w6(32'h3a319c64),
	.w7(32'hbb06ae71),
	.w8(32'h3a788bcf),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a40f210),
	.w1(32'hb935619d),
	.w2(32'hbb50e02a),
	.w3(32'h3a9257d3),
	.w4(32'h3a0f10a5),
	.w5(32'hb9adeae8),
	.w6(32'h3954390c),
	.w7(32'hbaafde4d),
	.w8(32'hb8e4cb8a),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba350ab4),
	.w1(32'hbba3323e),
	.w2(32'h3ba7e4ae),
	.w3(32'h3a25e2cd),
	.w4(32'hba27a49f),
	.w5(32'h3bb6978a),
	.w6(32'hbbca8ac4),
	.w7(32'hba3fd989),
	.w8(32'h3b104fc8),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63afb2),
	.w1(32'h3a00b0fc),
	.w2(32'h3b2eba27),
	.w3(32'hba179fde),
	.w4(32'hba1f3347),
	.w5(32'hb99f4983),
	.w6(32'h39b4cadb),
	.w7(32'hb92b91dd),
	.w8(32'h3acaa6c9),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e2167),
	.w1(32'h3ba6e6ec),
	.w2(32'h3cafe34b),
	.w3(32'h3b907722),
	.w4(32'hbb9eba8d),
	.w5(32'h3c68b7d9),
	.w6(32'h3b4c1df9),
	.w7(32'h3c3843bd),
	.w8(32'h3b1bd8ae),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f45dd),
	.w1(32'h3ae2bee4),
	.w2(32'h3a1138a5),
	.w3(32'hb98c50d5),
	.w4(32'h3b32c65c),
	.w5(32'h3b333e3b),
	.w6(32'h3a025c76),
	.w7(32'h3a1f6351),
	.w8(32'h3a4f30f0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa91519),
	.w1(32'h39907313),
	.w2(32'h3b93fe30),
	.w3(32'h3b062bf9),
	.w4(32'h389d7094),
	.w5(32'h3b7a4ba4),
	.w6(32'hb9c7a56d),
	.w7(32'h3b2d00c8),
	.w8(32'hbac7dfa2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9696d1),
	.w1(32'h3af08395),
	.w2(32'h3b087eb5),
	.w3(32'h3a0139c6),
	.w4(32'h3a2d401f),
	.w5(32'h3b29a082),
	.w6(32'h386a18ae),
	.w7(32'hbb56dcea),
	.w8(32'hba3d78a6),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a3508),
	.w1(32'h3bd7e9f4),
	.w2(32'h3c2b327f),
	.w3(32'h3b863a6c),
	.w4(32'h3bd52c86),
	.w5(32'h3c498307),
	.w6(32'hbb209fd4),
	.w7(32'h38a582ea),
	.w8(32'hbad9c0d2),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34f1bc),
	.w1(32'h3a1fe4d0),
	.w2(32'h3bc42929),
	.w3(32'h3ca47b32),
	.w4(32'hbab965cb),
	.w5(32'h3b988cea),
	.w6(32'h3a3577aa),
	.w7(32'h3a7defa1),
	.w8(32'h3acf97be),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8450b1),
	.w1(32'h3ba81d79),
	.w2(32'h3aa380f2),
	.w3(32'h3ab251f9),
	.w4(32'h3b555201),
	.w5(32'h391e270a),
	.w6(32'h3ad830b3),
	.w7(32'h3a97c8e9),
	.w8(32'h393c9201),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c8f66),
	.w1(32'h39c68c48),
	.w2(32'h3aba2f57),
	.w3(32'h38b25870),
	.w4(32'hba260047),
	.w5(32'hb84e392d),
	.w6(32'h389f0c2c),
	.w7(32'h3a875584),
	.w8(32'h3a285608),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6b321),
	.w1(32'h3a3a96e2),
	.w2(32'h3b668061),
	.w3(32'h38b965d3),
	.w4(32'h3aae1f38),
	.w5(32'h3b8dd3ae),
	.w6(32'hb925ad86),
	.w7(32'h3b159abd),
	.w8(32'hba64125d),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b971cb1),
	.w1(32'h3a218fb3),
	.w2(32'h3b0b3683),
	.w3(32'h3b7a9f76),
	.w4(32'h3a82cc05),
	.w5(32'h3b334c3d),
	.w6(32'h39b0dd08),
	.w7(32'hba48512d),
	.w8(32'h3a477d43),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ab24e),
	.w1(32'h3ba852e7),
	.w2(32'h3bccbef0),
	.w3(32'h3bc9b089),
	.w4(32'h3b8d9cf9),
	.w5(32'h3b71988d),
	.w6(32'h3bb6f286),
	.w7(32'h3aed5e93),
	.w8(32'hba92c9c8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b638a25),
	.w1(32'h3af2e0cb),
	.w2(32'h3b55dd51),
	.w3(32'h3b533fc3),
	.w4(32'h3abb390b),
	.w5(32'h3b715e0d),
	.w6(32'hb7d8fb76),
	.w7(32'hb9939296),
	.w8(32'h3a3ec374),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a894dd),
	.w1(32'hbaf399de),
	.w2(32'h3a3db034),
	.w3(32'h3a089647),
	.w4(32'hba8aea3d),
	.w5(32'h3b087132),
	.w6(32'h3980112e),
	.w7(32'hba32d822),
	.w8(32'hba43ae20),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af78ab8),
	.w1(32'h3afc3709),
	.w2(32'h3cc0e515),
	.w3(32'h3aa55fd2),
	.w4(32'hbc046c66),
	.w5(32'h3c6d9c1a),
	.w6(32'hbb5855c2),
	.w7(32'h3c371ad9),
	.w8(32'h3ab4b2e9),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29ad7c),
	.w1(32'hba30a17b),
	.w2(32'hba28361b),
	.w3(32'hbb0aa8a3),
	.w4(32'hba801bca),
	.w5(32'h395a2c0e),
	.w6(32'hbaa4d6f2),
	.w7(32'hb9dddda4),
	.w8(32'hba5c35ce),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b0e97),
	.w1(32'h3a71ba81),
	.w2(32'h3a782023),
	.w3(32'hba3ba4fe),
	.w4(32'h3a3628d9),
	.w5(32'hbae1311f),
	.w6(32'hb9bbd835),
	.w7(32'h39a6a9e0),
	.w8(32'h38994ba4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4ca593),
	.w1(32'hbb59af21),
	.w2(32'h3ada7317),
	.w3(32'hba98da0a),
	.w4(32'hbbdaf865),
	.w5(32'h3a562615),
	.w6(32'hbbb5a450),
	.w7(32'hba5ae4ce),
	.w8(32'hbba8ff0f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c0a14b),
	.w1(32'hb9b08367),
	.w2(32'h391eada0),
	.w3(32'hbb806ea1),
	.w4(32'hba3f468a),
	.w5(32'hb95c541e),
	.w6(32'h389f9d51),
	.w7(32'hbaac0455),
	.w8(32'h39995970),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37b745),
	.w1(32'h3a86e707),
	.w2(32'h39d89108),
	.w3(32'h3b70f048),
	.w4(32'h3b2b7f2e),
	.w5(32'h3b59358f),
	.w6(32'h39f2604a),
	.w7(32'h3a3825a8),
	.w8(32'hba3e9e5c),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec8797),
	.w1(32'h39cd9ab0),
	.w2(32'h3bb235a3),
	.w3(32'h3b5e45f7),
	.w4(32'h39e25f1a),
	.w5(32'h3bbe15da),
	.w6(32'hb9c15637),
	.w7(32'h3a8620cb),
	.w8(32'h3a7298f8),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10eef5),
	.w1(32'hbba03c32),
	.w2(32'h3aa4ddb3),
	.w3(32'h3b0704fe),
	.w4(32'hbb1d8e59),
	.w5(32'h3b57a803),
	.w6(32'hbb392f05),
	.w7(32'h38a04046),
	.w8(32'hbb037784),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dbd5d),
	.w1(32'h3aae8075),
	.w2(32'h3b71dcf4),
	.w3(32'hba28b25f),
	.w4(32'h39e298c4),
	.w5(32'h3ae50a8c),
	.w6(32'hb9d74f5a),
	.w7(32'hb915a236),
	.w8(32'h3a9dc899),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205135),
	.w1(32'h3b8c7424),
	.w2(32'h3b900968),
	.w3(32'h3b70137b),
	.w4(32'h3b80c21a),
	.w5(32'h3ae99fd3),
	.w6(32'h3b914517),
	.w7(32'hba55314a),
	.w8(32'h39642a73),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2395a4),
	.w1(32'h3ad67495),
	.w2(32'h3b37ccf2),
	.w3(32'h3b08291a),
	.w4(32'h39c425aa),
	.w5(32'h3a9cd752),
	.w6(32'hb9a164b3),
	.w7(32'hb9bb6167),
	.w8(32'h3908ba6f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa1348),
	.w1(32'h3a022ddb),
	.w2(32'h39a58146),
	.w3(32'h3a089d5d),
	.w4(32'h3ac3e5a6),
	.w5(32'h387afe3d),
	.w6(32'h3a664a14),
	.w7(32'h38d51ae6),
	.w8(32'h39b1ea5f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3baac4),
	.w1(32'hb9a34387),
	.w2(32'hba6991f4),
	.w3(32'h3b17007f),
	.w4(32'h398fddb4),
	.w5(32'hbafd2262),
	.w6(32'hb9a3b374),
	.w7(32'hbad20e27),
	.w8(32'hba4dc23e),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7672a5),
	.w1(32'h3a352d12),
	.w2(32'h3a68d032),
	.w3(32'hb9340ae1),
	.w4(32'h3a631b68),
	.w5(32'h3ae1188b),
	.w6(32'hba831cc9),
	.w7(32'hb9a10b92),
	.w8(32'h38c365b1),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aafcdc8),
	.w1(32'h3b178b56),
	.w2(32'h3b6e6c37),
	.w3(32'h3b03f1fc),
	.w4(32'h38819299),
	.w5(32'h3a9a7bd3),
	.w6(32'h394b82dc),
	.w7(32'h3ad4bd00),
	.w8(32'hb90739d6),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a638f6c),
	.w1(32'h3a0126b7),
	.w2(32'h39af326f),
	.w3(32'h398bcb3d),
	.w4(32'h3aad9317),
	.w5(32'hb8cff0b9),
	.w6(32'h3a58940f),
	.w7(32'h370477d3),
	.w8(32'h39791cf2),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394466ca),
	.w1(32'h39c78131),
	.w2(32'h3ac451f7),
	.w3(32'h39e39ec8),
	.w4(32'h3adbd909),
	.w5(32'h3b51b16e),
	.w6(32'hbad6da7d),
	.w7(32'h3a409628),
	.w8(32'h3a781699),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7db9e4),
	.w1(32'hbaccfa01),
	.w2(32'hbb4cbdb6),
	.w3(32'h3b2a45ab),
	.w4(32'h38385927),
	.w5(32'hbaa14fca),
	.w6(32'h3ad810f9),
	.w7(32'hbace8d9e),
	.w8(32'h3a33ec9b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b983f5a),
	.w1(32'h3b6317cc),
	.w2(32'h3b9b989f),
	.w3(32'h3b85cff9),
	.w4(32'h3aaa60f7),
	.w5(32'h3b65dcaa),
	.w6(32'h3b066473),
	.w7(32'hbade0853),
	.w8(32'hba29b047),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7de37),
	.w1(32'h3ac2014e),
	.w2(32'h3a90d422),
	.w3(32'h3aa8e48c),
	.w4(32'h3a84618b),
	.w5(32'h3a11a879),
	.w6(32'h3add590d),
	.w7(32'hbaf66a6c),
	.w8(32'h39b2acde),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2d6c1),
	.w1(32'h3b46b782),
	.w2(32'h3b8912ee),
	.w3(32'h3b8dd7b3),
	.w4(32'h3b02c24a),
	.w5(32'h3b6e816e),
	.w6(32'h3b10a9ac),
	.w7(32'h39d2bd39),
	.w8(32'h3b1f3d91),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7ffa4),
	.w1(32'hbb0f0158),
	.w2(32'hbb41bb16),
	.w3(32'h3af9280c),
	.w4(32'hbb6dbf65),
	.w5(32'hbb810807),
	.w6(32'hba952892),
	.w7(32'hba960b33),
	.w8(32'hba7d43d9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39cf19),
	.w1(32'h3a393c0e),
	.w2(32'h3a007b67),
	.w3(32'hbb77319f),
	.w4(32'h3b087541),
	.w5(32'hb810733f),
	.w6(32'h3a9d412d),
	.w7(32'h391ea313),
	.w8(32'h3a187bf5),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c60eb4),
	.w1(32'h3a02a594),
	.w2(32'h378b334c),
	.w3(32'h3a4df82b),
	.w4(32'h3ace3eab),
	.w5(32'h39ae4f9a),
	.w6(32'h3a4a1ab0),
	.w7(32'h396a2817),
	.w8(32'h39f34029),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d6de37),
	.w1(32'h3a1efef7),
	.w2(32'hb6e6e9d5),
	.w3(32'h3ae28773),
	.w4(32'h3b1105f2),
	.w5(32'h39f3b87b),
	.w6(32'h3a9888a4),
	.w7(32'h393b3b97),
	.w8(32'h3a0b90de),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cda41),
	.w1(32'hba9fac96),
	.w2(32'h3b2bd4ba),
	.w3(32'h3b2d8f48),
	.w4(32'hbae2d9df),
	.w5(32'h398ad837),
	.w6(32'hba12c2fe),
	.w7(32'hbb5f231b),
	.w8(32'hba832458),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecddbc),
	.w1(32'hbb486ee2),
	.w2(32'hbaf0fba2),
	.w3(32'hb9394364),
	.w4(32'hbb22e283),
	.w5(32'hba9e782e),
	.w6(32'hbb29a3ac),
	.w7(32'hbac85647),
	.w8(32'hbb14c80c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d942f),
	.w1(32'h396b4903),
	.w2(32'hbadb69af),
	.w3(32'hbaad7c60),
	.w4(32'hba910004),
	.w5(32'hbb14ebcb),
	.w6(32'hba9c73fb),
	.w7(32'hbb196258),
	.w8(32'hbab2f6de),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383f1a4e),
	.w1(32'h3a30d315),
	.w2(32'hbb0bbaae),
	.w3(32'h3a9adb7d),
	.w4(32'h3951a8d2),
	.w5(32'hbadbada0),
	.w6(32'h3a0cb161),
	.w7(32'hbb2fc256),
	.w8(32'hbb40f13b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06067b),
	.w1(32'h3a8aafa2),
	.w2(32'h3a17f718),
	.w3(32'hb9d5d03d),
	.w4(32'h3add4c05),
	.w5(32'h3a77c5a1),
	.w6(32'h3a8520a2),
	.w7(32'h3a166647),
	.w8(32'h3a368423),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b2b2),
	.w1(32'hba963207),
	.w2(32'h3a41af99),
	.w3(32'h3b30bf81),
	.w4(32'hbb1cb422),
	.w5(32'hb9831c62),
	.w6(32'hba96e941),
	.w7(32'hbb4a8931),
	.w8(32'h3ace3156),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57afed),
	.w1(32'h3b2e5349),
	.w2(32'h3b8e86cc),
	.w3(32'h38b81f6c),
	.w4(32'h3b03fa99),
	.w5(32'h3b859372),
	.w6(32'h3a7f73bd),
	.w7(32'h3b520db7),
	.w8(32'h38af3094),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be57f5a),
	.w1(32'h3b8ccb5d),
	.w2(32'h3bee9c77),
	.w3(32'h3b494a39),
	.w4(32'hbad4a2bd),
	.w5(32'hba9c20dd),
	.w6(32'h3afa85a9),
	.w7(32'hba861361),
	.w8(32'hbaf1a9b9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8fe9236),
	.w1(32'hb940705a),
	.w2(32'hb95e963a),
	.w3(32'h37954a54),
	.w4(32'hb8e070b9),
	.w5(32'hb90a2952),
	.w6(32'hb97bf86a),
	.w7(32'hb980f604),
	.w8(32'hba0c7710),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9781911),
	.w1(32'hbada5115),
	.w2(32'hbb2d9416),
	.w3(32'h39ccf43d),
	.w4(32'hbafd363d),
	.w5(32'hbb1b8cdf),
	.w6(32'h3addd72e),
	.w7(32'hbad33182),
	.w8(32'hbb314fad),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule