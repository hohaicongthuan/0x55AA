module layer_5 (
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 512;
	parameter IMG_SIZE = 104;

	wire	valid_out_0,
		valid_out_1,
		valid_out_2,
		valid_out_3,
		valid_out_4,
		valid_out_5,
		valid_out_6,
		valid_out_7,
		valid_out_8,
		valid_out_9,
		valid_out_10,
		valid_out_11,
		valid_out_12,
		valid_out_13,
		valid_out_14,
		valid_out_15,
		valid_out_16,
		valid_out_17,
		valid_out_18,
		valid_out_19,
		valid_out_20,
		valid_out_21,
		valid_out_22,
		valid_out_23,
		valid_out_24,
		valid_out_25,
		valid_out_26,
		valid_out_27,
		valid_out_28,
		valid_out_29,
		valid_out_30,
		valid_out_31,
		valid_out_32,
		valid_out_33,
		valid_out_34,
		valid_out_35,
		valid_out_36,
		valid_out_37,
		valid_out_38,
		valid_out_39,
		valid_out_40,
		valid_out_41,
		valid_out_42,
		valid_out_43,
		valid_out_44,
		valid_out_45,
		valid_out_46,
		valid_out_47,
		valid_out_48,
		valid_out_49,
		valid_out_50,
		valid_out_51,
		valid_out_52,
		valid_out_53,
		valid_out_54,
		valid_out_55,
		valid_out_56,
		valid_out_57,
		valid_out_58,
		valid_out_59,
		valid_out_60,
		valid_out_61,
		valid_out_62,
		valid_out_63;
Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7:0]),
	.valid_in(valid_in),
	.data_out(data_out[7:0]),
	.valid_out(valid_out_0)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[15:8]),
	.valid_in(valid_in),
	.data_out(data_out[15:8]),
	.valid_out(valid_out_1)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[23:16]),
	.valid_in(valid_in),
	.data_out(data_out[23:16]),
	.valid_out(valid_out_2)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:24]),
	.valid_in(valid_in),
	.data_out(data_out[31:24]),
	.valid_out(valid_out_3)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[39:32]),
	.valid_in(valid_in),
	.data_out(data_out[39:32]),
	.valid_out(valid_out_4)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[47:40]),
	.valid_in(valid_in),
	.data_out(data_out[47:40]),
	.valid_out(valid_out_5)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[55:48]),
	.valid_in(valid_in),
	.data_out(data_out[55:48]),
	.valid_out(valid_out_6)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:56]),
	.valid_in(valid_in),
	.data_out(data_out[63:56]),
	.valid_out(valid_out_7)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[71:64]),
	.valid_in(valid_in),
	.data_out(data_out[71:64]),
	.valid_out(valid_out_8)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[79:72]),
	.valid_in(valid_in),
	.data_out(data_out[79:72]),
	.valid_out(valid_out_9)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[87:80]),
	.valid_in(valid_in),
	.data_out(data_out[87:80]),
	.valid_out(valid_out_10)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:88]),
	.valid_in(valid_in),
	.data_out(data_out[95:88]),
	.valid_out(valid_out_11)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[103:96]),
	.valid_in(valid_in),
	.data_out(data_out[103:96]),
	.valid_out(valid_out_12)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[111:104]),
	.valid_in(valid_in),
	.data_out(data_out[111:104]),
	.valid_out(valid_out_13)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[119:112]),
	.valid_in(valid_in),
	.data_out(data_out[119:112]),
	.valid_out(valid_out_14)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:120]),
	.valid_in(valid_in),
	.data_out(data_out[127:120]),
	.valid_out(valid_out_15)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[135:128]),
	.valid_in(valid_in),
	.data_out(data_out[135:128]),
	.valid_out(valid_out_16)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[143:136]),
	.valid_in(valid_in),
	.data_out(data_out[143:136]),
	.valid_out(valid_out_17)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[151:144]),
	.valid_in(valid_in),
	.data_out(data_out[151:144]),
	.valid_out(valid_out_18)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:152]),
	.valid_in(valid_in),
	.data_out(data_out[159:152]),
	.valid_out(valid_out_19)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[167:160]),
	.valid_in(valid_in),
	.data_out(data_out[167:160]),
	.valid_out(valid_out_20)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[175:168]),
	.valid_in(valid_in),
	.data_out(data_out[175:168]),
	.valid_out(valid_out_21)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[183:176]),
	.valid_in(valid_in),
	.data_out(data_out[183:176]),
	.valid_out(valid_out_22)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:184]),
	.valid_in(valid_in),
	.data_out(data_out[191:184]),
	.valid_out(valid_out_23)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[199:192]),
	.valid_in(valid_in),
	.data_out(data_out[199:192]),
	.valid_out(valid_out_24)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[207:200]),
	.valid_in(valid_in),
	.data_out(data_out[207:200]),
	.valid_out(valid_out_25)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[215:208]),
	.valid_in(valid_in),
	.data_out(data_out[215:208]),
	.valid_out(valid_out_26)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:216]),
	.valid_in(valid_in),
	.data_out(data_out[223:216]),
	.valid_out(valid_out_27)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[231:224]),
	.valid_in(valid_in),
	.data_out(data_out[231:224]),
	.valid_out(valid_out_28)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[239:232]),
	.valid_in(valid_in),
	.data_out(data_out[239:232]),
	.valid_out(valid_out_29)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[247:240]),
	.valid_in(valid_in),
	.data_out(data_out[247:240]),
	.valid_out(valid_out_30)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:248]),
	.valid_in(valid_in),
	.data_out(data_out[255:248]),
	.valid_out(valid_out_31)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[263:256]),
	.valid_in(valid_in),
	.data_out(data_out[263:256]),
	.valid_out(valid_out_32)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[271:264]),
	.valid_in(valid_in),
	.data_out(data_out[271:264]),
	.valid_out(valid_out_33)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[279:272]),
	.valid_in(valid_in),
	.data_out(data_out[279:272]),
	.valid_out(valid_out_34)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:280]),
	.valid_in(valid_in),
	.data_out(data_out[287:280]),
	.valid_out(valid_out_35)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[295:288]),
	.valid_in(valid_in),
	.data_out(data_out[295:288]),
	.valid_out(valid_out_36)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[303:296]),
	.valid_in(valid_in),
	.data_out(data_out[303:296]),
	.valid_out(valid_out_37)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[311:304]),
	.valid_in(valid_in),
	.data_out(data_out[311:304]),
	.valid_out(valid_out_38)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:312]),
	.valid_in(valid_in),
	.data_out(data_out[319:312]),
	.valid_out(valid_out_39)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[327:320]),
	.valid_in(valid_in),
	.data_out(data_out[327:320]),
	.valid_out(valid_out_40)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[335:328]),
	.valid_in(valid_in),
	.data_out(data_out[335:328]),
	.valid_out(valid_out_41)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[343:336]),
	.valid_in(valid_in),
	.data_out(data_out[343:336]),
	.valid_out(valid_out_42)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:344]),
	.valid_in(valid_in),
	.data_out(data_out[351:344]),
	.valid_out(valid_out_43)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[359:352]),
	.valid_in(valid_in),
	.data_out(data_out[359:352]),
	.valid_out(valid_out_44)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[367:360]),
	.valid_in(valid_in),
	.data_out(data_out[367:360]),
	.valid_out(valid_out_45)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[375:368]),
	.valid_in(valid_in),
	.data_out(data_out[375:368]),
	.valid_out(valid_out_46)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:376]),
	.valid_in(valid_in),
	.data_out(data_out[383:376]),
	.valid_out(valid_out_47)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[391:384]),
	.valid_in(valid_in),
	.data_out(data_out[391:384]),
	.valid_out(valid_out_48)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[399:392]),
	.valid_in(valid_in),
	.data_out(data_out[399:392]),
	.valid_out(valid_out_49)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[407:400]),
	.valid_in(valid_in),
	.data_out(data_out[407:400]),
	.valid_out(valid_out_50)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:408]),
	.valid_in(valid_in),
	.data_out(data_out[415:408]),
	.valid_out(valid_out_51)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[423:416]),
	.valid_in(valid_in),
	.data_out(data_out[423:416]),
	.valid_out(valid_out_52)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[431:424]),
	.valid_in(valid_in),
	.data_out(data_out[431:424]),
	.valid_out(valid_out_53)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[439:432]),
	.valid_in(valid_in),
	.data_out(data_out[439:432]),
	.valid_out(valid_out_54)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:440]),
	.valid_in(valid_in),
	.data_out(data_out[447:440]),
	.valid_out(valid_out_55)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[455:448]),
	.valid_in(valid_in),
	.data_out(data_out[455:448]),
	.valid_out(valid_out_56)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[463:456]),
	.valid_in(valid_in),
	.data_out(data_out[463:456]),
	.valid_out(valid_out_57)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[471:464]),
	.valid_in(valid_in),
	.data_out(data_out[471:464]),
	.valid_out(valid_out_58)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:472]),
	.valid_in(valid_in),
	.data_out(data_out[479:472]),
	.valid_out(valid_out_59)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[487:480]),
	.valid_in(valid_in),
	.data_out(data_out[487:480]),
	.valid_out(valid_out_60)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[495:488]),
	.valid_in(valid_in),
	.data_out(data_out[495:488]),
	.valid_out(valid_out_61)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[503:496]),
	.valid_in(valid_in),
	.data_out(data_out[503:496]),
	.valid_out(valid_out_62)
);

Maxpool2D2x2s2 #(
	.IMG_SIZE(IMG_SIZE)
)
Maxpool2D2x2s2_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:504]),
	.valid_in(valid_in),
	.data_out(data_out[511:504]),
	.valid_out(valid_out_63)
);

	assign valid_out = valid_out_0 & valid_out_1 & valid_out_2 & valid_out_3 & valid_out_4 & valid_out_5 & valid_out_6 & valid_out_7 & valid_out_8 & valid_out_9 & valid_out_10 & valid_out_11 & valid_out_12 & valid_out_13 & valid_out_14 & valid_out_15 & valid_out_16 & valid_out_17 & valid_out_18 & valid_out_19 & valid_out_20 & valid_out_21 & valid_out_22 & valid_out_23 & valid_out_24 & valid_out_25 & valid_out_26 & valid_out_27 & valid_out_28 & valid_out_29 & valid_out_30 & valid_out_31 & valid_out_32 & valid_out_33 & valid_out_34 & valid_out_35 & valid_out_36 & valid_out_37 & valid_out_38 & valid_out_39 & valid_out_40 & valid_out_41 & valid_out_42 & valid_out_43 & valid_out_44 & valid_out_45 & valid_out_46 & valid_out_47 & valid_out_48 & valid_out_49 & valid_out_50 & valid_out_51 & valid_out_52 & valid_out_53 & valid_out_54 & valid_out_55 & valid_out_56 & valid_out_57 & valid_out_58 & valid_out_59 & valid_out_60 & valid_out_61 & valid_out_62 & valid_out_63;
endmodule