module layer_10_featuremap_312(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379b47e9),
	.w1(32'h362a3cdd),
	.w2(32'h3710b2dd),
	.w3(32'h371f4ce3),
	.w4(32'h35c5951f),
	.w5(32'h366d860b),
	.w6(32'h3757457d),
	.w7(32'h36b06161),
	.w8(32'h371fa397),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b337f),
	.w1(32'hb90376c6),
	.w2(32'h3a5d2bcf),
	.w3(32'h39aef686),
	.w4(32'h3a77010a),
	.w5(32'h3969bea2),
	.w6(32'h3ad679b5),
	.w7(32'h3a3ab76f),
	.w8(32'h38c86879),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h357e91d1),
	.w1(32'h36a8288d),
	.w2(32'hb514b29d),
	.w3(32'h362a720b),
	.w4(32'hb6e789c6),
	.w5(32'h36ac4c45),
	.w6(32'h377f1679),
	.w7(32'h369c8c5a),
	.w8(32'h3704202f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ac84ff),
	.w1(32'h3a302234),
	.w2(32'h3940da84),
	.w3(32'h39446df1),
	.w4(32'h399ae07b),
	.w5(32'hb8e43580),
	.w6(32'h382779a3),
	.w7(32'h38e66c95),
	.w8(32'h388b0596),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e2aae),
	.w1(32'h397135bc),
	.w2(32'h390ce626),
	.w3(32'h396ec139),
	.w4(32'h3981cc97),
	.w5(32'h391e45fd),
	.w6(32'h393e0dbe),
	.w7(32'h39506206),
	.w8(32'h392343ad),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3700c7ac),
	.w1(32'h361a1155),
	.w2(32'h376209fc),
	.w3(32'h3740a0c8),
	.w4(32'h36e8d090),
	.w5(32'h3711c472),
	.w6(32'h36fa6d44),
	.w7(32'h35396514),
	.w8(32'h36c8eae0),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76cad0),
	.w1(32'h3ad6a53e),
	.w2(32'h3a05ce3b),
	.w3(32'h3af3f0ca),
	.w4(32'h3a652c20),
	.w5(32'h38212a3c),
	.w6(32'h390dc05f),
	.w7(32'h38de8943),
	.w8(32'hb9a6092f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabae674),
	.w1(32'hbb386f3b),
	.w2(32'hbb36929f),
	.w3(32'hbbbb808f),
	.w4(32'hbb885609),
	.w5(32'h3a0d6d4c),
	.w6(32'hbba4e401),
	.w7(32'hbb9980bb),
	.w8(32'hbb728ea4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6918f0),
	.w1(32'hba6d8d2b),
	.w2(32'hba27f669),
	.w3(32'hba6fc42b),
	.w4(32'hba427394),
	.w5(32'hb9a6896c),
	.w6(32'hba050896),
	.w7(32'hb9abe4ba),
	.w8(32'hb8117ed9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bf63a7),
	.w1(32'hb9fd5c59),
	.w2(32'h3a498665),
	.w3(32'hb9198926),
	.w4(32'h3987c157),
	.w5(32'h3a75c8d0),
	.w6(32'hbaa262bf),
	.w7(32'hbaaf99d2),
	.w8(32'hb9007a54),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3918fe73),
	.w1(32'h38a7fbb6),
	.w2(32'h390f876f),
	.w3(32'h3980f7e7),
	.w4(32'h38d339b2),
	.w5(32'hb850bc55),
	.w6(32'h39cd3854),
	.w7(32'h39959329),
	.w8(32'h38eeca41),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399eb27d),
	.w1(32'h3af7018f),
	.w2(32'h3a031d45),
	.w3(32'h3b2d60dd),
	.w4(32'h3b25fe4d),
	.w5(32'h3a21768f),
	.w6(32'h3a445f5b),
	.w7(32'h3ae83003),
	.w8(32'h39df0590),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b839c),
	.w1(32'h3a94c50b),
	.w2(32'h3afe9f5e),
	.w3(32'h3a8bf4ec),
	.w4(32'h3ac0d26e),
	.w5(32'h3b0103b2),
	.w6(32'hba902d98),
	.w7(32'hba97dc77),
	.w8(32'h3a467abe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb9dd6),
	.w1(32'h3a1086b0),
	.w2(32'h3a2dacd8),
	.w3(32'h398bde10),
	.w4(32'h39a293d9),
	.w5(32'h3a7c57b8),
	.w6(32'h39ab2d45),
	.w7(32'h39b6e697),
	.w8(32'h3a29e803),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb910e2a9),
	.w1(32'hba5be060),
	.w2(32'h38f2961f),
	.w3(32'h3a29a4dc),
	.w4(32'h393d4599),
	.w5(32'h39363ef5),
	.w6(32'h3a8d3e0d),
	.w7(32'h376810db),
	.w8(32'h39c34b38),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f32b5),
	.w1(32'hb9b6eb00),
	.w2(32'hb992b085),
	.w3(32'hba6292f1),
	.w4(32'hba41b046),
	.w5(32'hba01609d),
	.w6(32'hbaf61c2c),
	.w7(32'hbb1fc905),
	.w8(32'hba66c840),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d97f10),
	.w1(32'h39063d28),
	.w2(32'h3989bd5e),
	.w3(32'h374fb00f),
	.w4(32'h3926b2fd),
	.w5(32'h39c9f0db),
	.w6(32'h3855cb7e),
	.w7(32'h3989427b),
	.w8(32'h39fe1463),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44640f),
	.w1(32'hbb0a72c5),
	.w2(32'hbb952414),
	.w3(32'hbadb3bdd),
	.w4(32'hbb86f940),
	.w5(32'hbb7e3b4c),
	.w6(32'hbc12fd79),
	.w7(32'hbbdc9d76),
	.w8(32'hbb99ba50),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38febb2e),
	.w1(32'hba2fa0f1),
	.w2(32'hba9177f2),
	.w3(32'hba64f7d4),
	.w4(32'hbacf1fd2),
	.w5(32'hba93d25f),
	.w6(32'hbb8249c2),
	.w7(32'hbb4b977a),
	.w8(32'hbad06346),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb744e909),
	.w1(32'hb560671b),
	.w2(32'h37d5e03a),
	.w3(32'h37852a45),
	.w4(32'h37d99873),
	.w5(32'h384d570f),
	.w6(32'h37ba0d44),
	.w7(32'h371f985b),
	.w8(32'hb7adf409),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69f6390),
	.w1(32'hb81d2b7c),
	.w2(32'h37c8c7d4),
	.w3(32'h362f9e34),
	.w4(32'hb88b66ab),
	.w5(32'hb65f0826),
	.w6(32'h371fe7dc),
	.w7(32'hb7407eb3),
	.w8(32'h382401c8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a50931),
	.w1(32'h386e82cc),
	.w2(32'hb90e4f03),
	.w3(32'h3a0f1184),
	.w4(32'h39cc1556),
	.w5(32'hb9292b4c),
	.w6(32'h3a30c753),
	.w7(32'h39f2f38b),
	.w8(32'hb687f8d4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9da598),
	.w1(32'hbb22d94f),
	.w2(32'hbc066e3c),
	.w3(32'hba930626),
	.w4(32'hbbea64f2),
	.w5(32'hbc107a99),
	.w6(32'hbc1f1c8b),
	.w7(32'hbc01efed),
	.w8(32'hbc0c2e88),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e1eae),
	.w1(32'h39b04938),
	.w2(32'h3afe80b5),
	.w3(32'h3a2ccee8),
	.w4(32'h3a8f7cfd),
	.w5(32'h3b03c139),
	.w6(32'h39d6aeea),
	.w7(32'h394f69db),
	.w8(32'h3a9180e2),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39df912a),
	.w1(32'hb675da7c),
	.w2(32'h3a82d48c),
	.w3(32'h3a5f89f3),
	.w4(32'h3af34513),
	.w5(32'h3a8e27b2),
	.w6(32'h3afed37b),
	.w7(32'h3a8b54f4),
	.w8(32'hba09e352),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8976803),
	.w1(32'hb7810f1a),
	.w2(32'hb7460c4d),
	.w3(32'hb9a8b782),
	.w4(32'hb930fcea),
	.w5(32'hb8a613b6),
	.w6(32'hb93ad508),
	.w7(32'hb7de340b),
	.w8(32'h391f87b6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3880490d),
	.w1(32'h388f2043),
	.w2(32'h3903f555),
	.w3(32'h387b6d4e),
	.w4(32'h389279bf),
	.w5(32'h38f3c2a3),
	.w6(32'h390c875f),
	.w7(32'h38e61f56),
	.w8(32'h3914951e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39918b68),
	.w1(32'hbaa54d93),
	.w2(32'h38d41783),
	.w3(32'h3a909a69),
	.w4(32'h3a46d93e),
	.w5(32'h3a3e3de1),
	.w6(32'h3b570afb),
	.w7(32'h3aa8fb55),
	.w8(32'h3aeef320),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb766),
	.w1(32'h3a851b14),
	.w2(32'h39b93418),
	.w3(32'h3a9d07ea),
	.w4(32'h3aae9413),
	.w5(32'h39fbd157),
	.w6(32'h3aae9c24),
	.w7(32'h3ac4a7b4),
	.w8(32'h3a8f0367),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985f1c8),
	.w1(32'hb9b71fb8),
	.w2(32'h3a85927d),
	.w3(32'h3a1636bf),
	.w4(32'h3a078d30),
	.w5(32'h3a237e22),
	.w6(32'h3b2e8c49),
	.w7(32'h3a9cf5ab),
	.w8(32'h3aa927cd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d52e91),
	.w1(32'h377ad032),
	.w2(32'h382deb74),
	.w3(32'h38072177),
	.w4(32'h37c89f59),
	.w5(32'h3809eea8),
	.w6(32'h3836c0cd),
	.w7(32'h3837d6ea),
	.w8(32'h3870c4fe),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364f5182),
	.w1(32'h3764b4d2),
	.w2(32'h3875be29),
	.w3(32'hb79f084e),
	.w4(32'h384fe562),
	.w5(32'h38c3ba42),
	.w6(32'hb7528111),
	.w7(32'h38cc3ace),
	.w8(32'h3902d752),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b4f50b),
	.w1(32'hb8cfb882),
	.w2(32'h3894fdda),
	.w3(32'hba041e07),
	.w4(32'hb997b6ea),
	.w5(32'h3958f429),
	.w6(32'hbacab6dd),
	.w7(32'hba8b61cb),
	.w8(32'hb94af74e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05184b),
	.w1(32'hb90c3226),
	.w2(32'h3a0f301a),
	.w3(32'hb9a1b6b7),
	.w4(32'h38fe8f60),
	.w5(32'h39f3e42b),
	.w6(32'h3a2346a3),
	.w7(32'h395b1df9),
	.w8(32'h39a500af),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88dfdbd),
	.w1(32'hb7201052),
	.w2(32'h37f700e0),
	.w3(32'h39394b33),
	.w4(32'h38ac01ae),
	.w5(32'hb8d8f58d),
	.w6(32'h392c0a04),
	.w7(32'h384b4928),
	.w8(32'h394a4064),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5bc30),
	.w1(32'h3a1588f1),
	.w2(32'h39aae3c4),
	.w3(32'h37389fef),
	.w4(32'h3941842f),
	.w5(32'h39afb628),
	.w6(32'hba57f139),
	.w7(32'hb89dd06d),
	.w8(32'hb9477074),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d6e8b),
	.w1(32'hb9f38c03),
	.w2(32'h3a174137),
	.w3(32'h3a3152f7),
	.w4(32'hba4d406a),
	.w5(32'hba613a1a),
	.w6(32'hb9e56784),
	.w7(32'hbb452ec4),
	.w8(32'hbb7a7ea6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2b56d),
	.w1(32'h3ab26605),
	.w2(32'h3b527e21),
	.w3(32'h3b5fe202),
	.w4(32'h3bb0c3d3),
	.w5(32'h3b38c035),
	.w6(32'h3bf0c675),
	.w7(32'h3bc2ff13),
	.w8(32'h3b712d14),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b102b29),
	.w1(32'h3af459c9),
	.w2(32'h3ad05b3d),
	.w3(32'h3bc0f644),
	.w4(32'h3bac1dcf),
	.w5(32'h3abc4cd7),
	.w6(32'h3c2009b5),
	.w7(32'h3bbe0e33),
	.w8(32'h3b323654),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ab22b),
	.w1(32'h3a27a3cb),
	.w2(32'h3a504093),
	.w3(32'h39f6648b),
	.w4(32'h3a3fbe81),
	.w5(32'h3a052728),
	.w6(32'h3a680ea0),
	.w7(32'h39cf4832),
	.w8(32'h39dc228e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb988a9f7),
	.w1(32'hb937bfea),
	.w2(32'hb8b40408),
	.w3(32'hb9a7430a),
	.w4(32'hb97c5ad3),
	.w5(32'hb8d2528d),
	.w6(32'hb8f92418),
	.w7(32'hb8c58e5c),
	.w8(32'hb863c4e7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f629e),
	.w1(32'h3788fda9),
	.w2(32'h38d74910),
	.w3(32'h38ee3b66),
	.w4(32'h384e4de7),
	.w5(32'h38caa67e),
	.w6(32'h396f1dd4),
	.w7(32'h39056637),
	.w8(32'h3908b8af),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9506bfd),
	.w1(32'h397b1e7d),
	.w2(32'h39faf878),
	.w3(32'h38ae9064),
	.w4(32'h3a11045c),
	.w5(32'h3a05c569),
	.w6(32'hb90984c5),
	.w7(32'h39830ed1),
	.w8(32'h397c9b2b),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d07b1f),
	.w1(32'hb981dd21),
	.w2(32'hb9bb122f),
	.w3(32'hbafb61f9),
	.w4(32'hbad5c9f7),
	.w5(32'hb8fd53dd),
	.w6(32'hbb91cedf),
	.w7(32'hbb3d0ee8),
	.w8(32'h38a28486),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22eb5d),
	.w1(32'hba0b40b0),
	.w2(32'h39bcdb19),
	.w3(32'hba02d3f5),
	.w4(32'h36673ed2),
	.w5(32'h39cc8d6c),
	.w6(32'h3a0ea688),
	.w7(32'h39a6866b),
	.w8(32'h39fb16d1),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a0a7e4),
	.w1(32'hb96adbc8),
	.w2(32'h3a905da0),
	.w3(32'h37a200f5),
	.w4(32'h3937a458),
	.w5(32'h3a8a6f01),
	.w6(32'hb9e2ac48),
	.w7(32'hba893a60),
	.w8(32'hb9e6dc5b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7c5f2),
	.w1(32'hba46300c),
	.w2(32'hba4fefd7),
	.w3(32'hba6687d8),
	.w4(32'hba12925a),
	.w5(32'hba4391e6),
	.w6(32'hbb1af570),
	.w7(32'hbaf1acfe),
	.w8(32'hbacc8dc8),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0d6a9),
	.w1(32'hbabbc69d),
	.w2(32'hbb9f253b),
	.w3(32'hbaeb14dc),
	.w4(32'hbb7a4f0b),
	.w5(32'hbb666b01),
	.w6(32'hbc24b300),
	.w7(32'hbbfde400),
	.w8(32'hbbabf4e3),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390101b7),
	.w1(32'h39423ed1),
	.w2(32'h372d8eb4),
	.w3(32'h39775445),
	.w4(32'h39896a70),
	.w5(32'h3853a1e3),
	.w6(32'h39622b55),
	.w7(32'h393e37d8),
	.w8(32'h385b495c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86757c6),
	.w1(32'hb960f722),
	.w2(32'hb9809f92),
	.w3(32'hb8e5a89f),
	.w4(32'hb9c82312),
	.w5(32'hb9c0538b),
	.w6(32'hb9b951bb),
	.w7(32'hba2739d7),
	.w8(32'hba4ef300),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0effe8),
	.w1(32'h399137d5),
	.w2(32'hb915cbe8),
	.w3(32'h3a31346c),
	.w4(32'h39b73ec0),
	.w5(32'hb8fa5699),
	.w6(32'h3a185824),
	.w7(32'h39be42ce),
	.w8(32'hb8f15f62),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3994c229),
	.w1(32'h399c863b),
	.w2(32'h392b201d),
	.w3(32'hb87acd39),
	.w4(32'hb9f92574),
	.w5(32'h38fce2cc),
	.w6(32'hb9b21c4e),
	.w7(32'hba38727c),
	.w8(32'hba320658),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3881c86a),
	.w1(32'hb9d1510c),
	.w2(32'hba2cdf33),
	.w3(32'hb9cc1fbd),
	.w4(32'hba2ce067),
	.w5(32'hba1d163f),
	.w6(32'hba683454),
	.w7(32'hba7b5ee1),
	.w8(32'hba57de35),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6cf1),
	.w1(32'hba6ca7e2),
	.w2(32'hba5e44a2),
	.w3(32'hb9982347),
	.w4(32'hb9db352e),
	.w5(32'h3a346226),
	.w6(32'hbbbbf28c),
	.w7(32'hbb8387e9),
	.w8(32'hba2188c7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394bbae4),
	.w1(32'hb982868a),
	.w2(32'hba29938a),
	.w3(32'hb999e099),
	.w4(32'hb9e5a4b7),
	.w5(32'hb969fd82),
	.w6(32'hb919398a),
	.w7(32'hb99a5ca5),
	.w8(32'hba16d2c2),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cbd0af),
	.w1(32'hb8217696),
	.w2(32'hb836c639),
	.w3(32'h3805befe),
	.w4(32'h37f1a233),
	.w5(32'hb7a0b46e),
	.w6(32'h386cd380),
	.w7(32'h389c6133),
	.w8(32'h381a88c6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c31ce3),
	.w1(32'hb7055fb9),
	.w2(32'h348f06fc),
	.w3(32'hb6a283d9),
	.w4(32'hb6c3973d),
	.w5(32'h3680cf75),
	.w6(32'h37b519a1),
	.w7(32'h378830ff),
	.w8(32'h379ef954),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed57f7),
	.w1(32'h37c1ac2f),
	.w2(32'h376471d8),
	.w3(32'h3897ce48),
	.w4(32'hb896b89a),
	.w5(32'hb819a829),
	.w6(32'h394d3c27),
	.w7(32'h38028b5e),
	.w8(32'h38553d6e),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ef9c0c),
	.w1(32'h38f56862),
	.w2(32'h390ae946),
	.w3(32'h3764e77e),
	.w4(32'h3953f034),
	.w5(32'h38dc9542),
	.w6(32'h37f21922),
	.w7(32'h39131b94),
	.w8(32'h38c49bab),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8bf4351),
	.w1(32'h38e423cb),
	.w2(32'h39b48d23),
	.w3(32'h38808c6a),
	.w4(32'h38eeafd9),
	.w5(32'h39d2b579),
	.w6(32'h369e1dae),
	.w7(32'hb61dcda1),
	.w8(32'h39851526),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39af7d1b),
	.w1(32'hb9ac0d6e),
	.w2(32'hbab20e9a),
	.w3(32'hba2d3934),
	.w4(32'hba4f219a),
	.w5(32'hba8667c8),
	.w6(32'hbb1dc81b),
	.w7(32'hbac9ba45),
	.w8(32'hbab7d6bc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21e94e),
	.w1(32'hbad08802),
	.w2(32'hbb0ae5b9),
	.w3(32'hbaf8c484),
	.w4(32'hbb19fecf),
	.w5(32'hbafa25b4),
	.w6(32'hbb03de45),
	.w7(32'hbab322ab),
	.w8(32'hba9f023b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35913902),
	.w1(32'h3811306c),
	.w2(32'h38461ecd),
	.w3(32'hb7b82ba6),
	.w4(32'h385e1651),
	.w5(32'h38882dfb),
	.w6(32'hb80e0329),
	.w7(32'h37dee77b),
	.w8(32'h38981fb8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb748e90a),
	.w1(32'hb7c62890),
	.w2(32'hb7163ea5),
	.w3(32'hb78cb0b7),
	.w4(32'hb7ef2152),
	.w5(32'h35dcae12),
	.w6(32'hb75ca08e),
	.w7(32'hb787d774),
	.w8(32'h37652061),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39063b06),
	.w1(32'h38c818da),
	.w2(32'h38e8bd4d),
	.w3(32'h38ba2126),
	.w4(32'h38731249),
	.w5(32'h386f374c),
	.w6(32'h38d6b576),
	.w7(32'h38b515cd),
	.w8(32'h38aa8b9a),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3649df13),
	.w1(32'h3716f069),
	.w2(32'h3841cc7f),
	.w3(32'h370724b8),
	.w4(32'h379993e0),
	.w5(32'h3843d8c7),
	.w6(32'h382c18b6),
	.w7(32'h382c11c2),
	.w8(32'h38962c85),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39deccf0),
	.w1(32'hb9f8a3ce),
	.w2(32'h3945b5ef),
	.w3(32'h3b1bde0b),
	.w4(32'h3ac7a831),
	.w5(32'h3a2d313e),
	.w6(32'hbab3aaf7),
	.w7(32'hbab6a4c6),
	.w8(32'h3a07e714),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd02df),
	.w1(32'h3a87028e),
	.w2(32'h3a596522),
	.w3(32'h392c3d42),
	.w4(32'hb9090857),
	.w5(32'h3a1bd1de),
	.w6(32'h39821099),
	.w7(32'hb9eb239a),
	.w8(32'hbac9c0f7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e92d44),
	.w1(32'hbacc31d4),
	.w2(32'hbb453390),
	.w3(32'hba7ed69f),
	.w4(32'hbae4020b),
	.w5(32'hbb25e4f8),
	.w6(32'hbb7ff6c4),
	.w7(32'hbb632153),
	.w8(32'hbb8833a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3814414a),
	.w1(32'h3abc1ec9),
	.w2(32'h3b642235),
	.w3(32'h3b0d7cd9),
	.w4(32'h3b7169d2),
	.w5(32'h3b615af9),
	.w6(32'h3b865855),
	.w7(32'h3b4a6298),
	.w8(32'h3b1b1467),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370c67b9),
	.w1(32'h3658508d),
	.w2(32'h378e73bb),
	.w3(32'h342cc07d),
	.w4(32'hb76afb8e),
	.w5(32'hb6dd4041),
	.w6(32'h3707a59f),
	.w7(32'hb71a4e69),
	.w8(32'hb64ae0e0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3577f19a),
	.w1(32'h349174e0),
	.w2(32'h38490ef0),
	.w3(32'hb7371bc8),
	.w4(32'hb70e631c),
	.w5(32'h38079d02),
	.w6(32'h37a6cf98),
	.w7(32'h37afa0fc),
	.w8(32'h384cdc09),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f57f62),
	.w1(32'hb7af951b),
	.w2(32'h37d8ddf2),
	.w3(32'hb7707c0e),
	.w4(32'hb82d7b8f),
	.w5(32'h376bbabc),
	.w6(32'h36366c33),
	.w7(32'hb75c522e),
	.w8(32'h37cf3d11),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3856620c),
	.w1(32'hb988081a),
	.w2(32'hb9d6efdb),
	.w3(32'hb832f188),
	.w4(32'hb96fa56a),
	.w5(32'hb88b06c2),
	.w6(32'hba25d891),
	.w7(32'hba69057e),
	.w8(32'hba2801b0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c45cb4),
	.w1(32'h355800c1),
	.w2(32'h3808acc5),
	.w3(32'h382dbdf4),
	.w4(32'h367df44e),
	.w5(32'h37df6702),
	.w6(32'h388b2ee4),
	.w7(32'h380aef94),
	.w8(32'h3840bf5d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caedb2),
	.w1(32'hbad2b21d),
	.w2(32'hbb14344c),
	.w3(32'hb99359db),
	.w4(32'hba9522d5),
	.w5(32'hbafd9e71),
	.w6(32'hbb7ad704),
	.w7(32'hbb6d69ec),
	.w8(32'hbb0a3784),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d39b14),
	.w1(32'hbb851f48),
	.w2(32'hbb7237d3),
	.w3(32'hbb31fecf),
	.w4(32'hbb8f771a),
	.w5(32'hbb81cfdf),
	.w6(32'hbbb56504),
	.w7(32'hbbf27774),
	.w8(32'hbbb1b83d),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9407609),
	.w1(32'h3a26d687),
	.w2(32'h3acc8339),
	.w3(32'h3aa77459),
	.w4(32'h3ae0e0f7),
	.w5(32'h3ab25191),
	.w6(32'h3b01960f),
	.w7(32'h3a8dd8d9),
	.w8(32'h3a857327),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3827e86c),
	.w1(32'hb9fcf100),
	.w2(32'hb997bfbe),
	.w3(32'hba142665),
	.w4(32'hb9cec905),
	.w5(32'h38b7ab3a),
	.w6(32'hba9495c2),
	.w7(32'hba96062f),
	.w8(32'hba053ede),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ca5a1),
	.w1(32'hb8c8dae8),
	.w2(32'h3a12cc9e),
	.w3(32'h3a5ce54c),
	.w4(32'h3a88b221),
	.w5(32'h3a4c61f3),
	.w6(32'hb997163d),
	.w7(32'hba1cc1cf),
	.w8(32'hb9834693),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d47745),
	.w1(32'hba4c54a4),
	.w2(32'hba015e0c),
	.w3(32'hb965d85f),
	.w4(32'hb98e32bf),
	.w5(32'hb984f28c),
	.w6(32'h39806681),
	.w7(32'hb74b23f8),
	.w8(32'h38713243),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95b713d),
	.w1(32'hba86e352),
	.w2(32'hbb146e50),
	.w3(32'hb99c8ee1),
	.w4(32'hbab0d177),
	.w5(32'hbaf2c2c3),
	.w6(32'hbb6b008b),
	.w7(32'hbb3ac61e),
	.w8(32'hbafa7961),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37189fb6),
	.w1(32'h36d87bf4),
	.w2(32'h37c98d07),
	.w3(32'h371eeef6),
	.w4(32'h373fa026),
	.w5(32'h37541391),
	.w6(32'h37428d9f),
	.w7(32'h373db80a),
	.w8(32'h37921786),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35760319),
	.w1(32'h36933963),
	.w2(32'h3789e184),
	.w3(32'h36b32fa2),
	.w4(32'hb560a735),
	.w5(32'h353adbc5),
	.w6(32'h37bb6996),
	.w7(32'h371ed35a),
	.w8(32'hb6d592ad),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39105b43),
	.w1(32'h38f59964),
	.w2(32'h3931f933),
	.w3(32'h39829ed1),
	.w4(32'h395ae8c3),
	.w5(32'h3981442f),
	.w6(32'h39c44b1c),
	.w7(32'h3965fbb3),
	.w8(32'h39800eec),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3771cd8f),
	.w1(32'hb8329f96),
	.w2(32'hb827ce28),
	.w3(32'h380e1914),
	.w4(32'hb665fbb8),
	.w5(32'h36167578),
	.w6(32'h388f018b),
	.w7(32'hb6cd0272),
	.w8(32'h37ab11a2),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d2ef41),
	.w1(32'h3a659272),
	.w2(32'h3b029c96),
	.w3(32'h3988f110),
	.w4(32'h3ab23750),
	.w5(32'h3ab06b44),
	.w6(32'h3ada5cc5),
	.w7(32'h38d2be06),
	.w8(32'h39f8c339),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92f78df),
	.w1(32'h38eed630),
	.w2(32'h396d2444),
	.w3(32'h390854f0),
	.w4(32'h39b9f620),
	.w5(32'h3993326e),
	.w6(32'h399ef31c),
	.w7(32'h39df59d9),
	.w8(32'h39a8a0a5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90af465),
	.w1(32'hba0a27b8),
	.w2(32'hb8c7eda9),
	.w3(32'hba055988),
	.w4(32'hb9ddba1c),
	.w5(32'h37256d09),
	.w6(32'hb9ca5ca8),
	.w7(32'hba21111f),
	.w8(32'hba2dd7c6),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374d8b9b),
	.w1(32'hbb4807c5),
	.w2(32'hbb8cb397),
	.w3(32'hbb8f2118),
	.w4(32'hbbbfed03),
	.w5(32'hbb8a29a0),
	.w6(32'hbc1b0e73),
	.w7(32'hbc0537c1),
	.w8(32'hbbad5d91),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5be3d),
	.w1(32'h3a7cc1fc),
	.w2(32'h3a03bf9e),
	.w3(32'h3b0a4a64),
	.w4(32'h3b222b98),
	.w5(32'h3a149dba),
	.w6(32'h3b32acdb),
	.w7(32'h3b0327f6),
	.w8(32'h3a82444b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba847831),
	.w1(32'h3b1e0c29),
	.w2(32'h3aab0502),
	.w3(32'h3b0564ca),
	.w4(32'h39e70dac),
	.w5(32'hb9b352b1),
	.w6(32'hb9ef7f97),
	.w7(32'hb97e638b),
	.w8(32'hb8b55017),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06a44a),
	.w1(32'h3a92a181),
	.w2(32'h3ab55c18),
	.w3(32'h3976e1ae),
	.w4(32'h3a9452cc),
	.w5(32'h3a964057),
	.w6(32'h3a05e68f),
	.w7(32'h3a918412),
	.w8(32'h3a496498),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b8f46),
	.w1(32'hba40089d),
	.w2(32'h3a4a17ae),
	.w3(32'h3804e820),
	.w4(32'h38c5115b),
	.w5(32'h3ac55c59),
	.w6(32'hba86c82e),
	.w7(32'hbaf380a9),
	.w8(32'hba27211f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba316bc6),
	.w1(32'hba786613),
	.w2(32'h3888b4d3),
	.w3(32'h39cfa771),
	.w4(32'h393302b4),
	.w5(32'h39245e23),
	.w6(32'hb9868336),
	.w7(32'hba8270bb),
	.w8(32'hba03977d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923c150),
	.w1(32'h3a6863a6),
	.w2(32'h3ade8af5),
	.w3(32'h3ab50a7c),
	.w4(32'h3ad3e61f),
	.w5(32'h3aca401a),
	.w6(32'h3b180a97),
	.w7(32'h3ad03fb5),
	.w8(32'h3b08e3c4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954203e),
	.w1(32'h3a318085),
	.w2(32'h39c0f438),
	.w3(32'h3960bc7e),
	.w4(32'h39987175),
	.w5(32'h39cd59b1),
	.w6(32'h39f50ba8),
	.w7(32'h399b3858),
	.w8(32'h3a1d39ed),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0c5052),
	.w1(32'hb9a71b02),
	.w2(32'hbaa7ef37),
	.w3(32'hb9c18437),
	.w4(32'hbaa58ed3),
	.w5(32'hbac7a7fd),
	.w6(32'hbb4e7a30),
	.w7(32'hbb578e01),
	.w8(32'hbb32279d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93d8f65),
	.w1(32'h3a09f66e),
	.w2(32'h3a725ea0),
	.w3(32'h3a9c999c),
	.w4(32'h3ad92ee3),
	.w5(32'h398a9284),
	.w6(32'hba309a83),
	.w7(32'hbabcfdbb),
	.w8(32'hbacb41a8),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad29b23),
	.w1(32'hbb0d39f5),
	.w2(32'hbb5750d1),
	.w3(32'hbb236247),
	.w4(32'hbbb22480),
	.w5(32'hbbae0556),
	.w6(32'hbbc66d02),
	.w7(32'hbbe20778),
	.w8(32'hbbe8a379),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabc913d),
	.w1(32'h3ac30976),
	.w2(32'h3b72ce95),
	.w3(32'h3b1867b8),
	.w4(32'h3bb1c2eb),
	.w5(32'h3b8d859f),
	.w6(32'h3b96146b),
	.w7(32'h3aca857a),
	.w8(32'h3ae65e1d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e89cc8),
	.w1(32'hb9d74532),
	.w2(32'h3a8af7b4),
	.w3(32'hb889159c),
	.w4(32'h3812250d),
	.w5(32'hb888afee),
	.w6(32'h3a160dfa),
	.w7(32'hb95c461e),
	.w8(32'hba0cba4a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398579cc),
	.w1(32'h3a88d237),
	.w2(32'hb93e03ca),
	.w3(32'h3add3e09),
	.w4(32'h3a177e26),
	.w5(32'h3a7debfa),
	.w6(32'hbb24e64b),
	.w7(32'hbb1e3487),
	.w8(32'hba5351f6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa157cb),
	.w1(32'h3aff2e2d),
	.w2(32'h3a88ae2f),
	.w3(32'h3a3bafc8),
	.w4(32'h3a17b578),
	.w5(32'h390e5fc5),
	.w6(32'hb98b809d),
	.w7(32'h3a55483a),
	.w8(32'hb9a8f97e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a1ff4),
	.w1(32'hbbb0c203),
	.w2(32'hbbe39fc9),
	.w3(32'hbb39421b),
	.w4(32'hbb7df60a),
	.w5(32'hbbb4fea5),
	.w6(32'hbbbcca54),
	.w7(32'hbc2d44a8),
	.w8(32'hbbfa8bec),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb845f728),
	.w1(32'hb93014de),
	.w2(32'h3889afd9),
	.w3(32'h3a9da982),
	.w4(32'h3a8f749b),
	.w5(32'hba1aa624),
	.w6(32'h3a806062),
	.w7(32'h39274b2a),
	.w8(32'hb9f9352b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3af60e),
	.w1(32'hba176def),
	.w2(32'hba4bb391),
	.w3(32'hb9dfafd8),
	.w4(32'hba02648c),
	.w5(32'h39ea5ba9),
	.w6(32'hba511797),
	.w7(32'hba235909),
	.w8(32'h38a24d9d),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9adf999),
	.w1(32'h39c6c145),
	.w2(32'hb926ad59),
	.w3(32'h39a0b919),
	.w4(32'hb6c41025),
	.w5(32'hba1ef108),
	.w6(32'h364cae1b),
	.w7(32'hb932ad4c),
	.w8(32'hba1e03a0),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77e852),
	.w1(32'h39ba3901),
	.w2(32'h3a4601fb),
	.w3(32'hba2735dd),
	.w4(32'hb96861f9),
	.w5(32'h39f138ea),
	.w6(32'hbb0fc0cf),
	.w7(32'hbb0ba66b),
	.w8(32'hba2e6839),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e7212),
	.w1(32'hba161934),
	.w2(32'h396538fc),
	.w3(32'h3a3e1b71),
	.w4(32'h39d00496),
	.w5(32'hba309a02),
	.w6(32'h3b064c0f),
	.w7(32'h3a4f9cc9),
	.w8(32'hb7984356),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba46351c),
	.w1(32'hba9d3f0a),
	.w2(32'hbaac50dc),
	.w3(32'h39f7b905),
	.w4(32'hba6ad2c3),
	.w5(32'hba536dbf),
	.w6(32'h3b10dae3),
	.w7(32'hba3501f7),
	.w8(32'hb9ad9122),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f41ce6),
	.w1(32'h389777ee),
	.w2(32'h3a5fa63f),
	.w3(32'h39baf6ad),
	.w4(32'h39e5bdcd),
	.w5(32'h397de60f),
	.w6(32'h39101046),
	.w7(32'hb9317971),
	.w8(32'hba9c4778),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2479),
	.w1(32'h396931d2),
	.w2(32'h3a3433ab),
	.w3(32'hba6d4337),
	.w4(32'h3a9fafe3),
	.w5(32'h3abbce0c),
	.w6(32'hba26e409),
	.w7(32'h3aaac43b),
	.w8(32'h3a85b83f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b24c),
	.w1(32'h396e2aa1),
	.w2(32'h38c125f4),
	.w3(32'h39d22434),
	.w4(32'h3812445b),
	.w5(32'hba4e4f3d),
	.w6(32'hbab8ef60),
	.w7(32'hbab78301),
	.w8(32'hba925063),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20e891),
	.w1(32'hb95617a0),
	.w2(32'h3a118eb5),
	.w3(32'hb8fb27f6),
	.w4(32'h39b67119),
	.w5(32'hb9a0c64b),
	.w6(32'h3a971413),
	.w7(32'h39a9de78),
	.w8(32'hb9ca81bf),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91200c5),
	.w1(32'h3873d43a),
	.w2(32'h39ab2c83),
	.w3(32'hb8e37741),
	.w4(32'h383784b3),
	.w5(32'h3a0cd54d),
	.w6(32'hb981954d),
	.w7(32'h3982238a),
	.w8(32'h39d925c5),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dc0e1d),
	.w1(32'h392c74a2),
	.w2(32'h38f9b480),
	.w3(32'h39a84406),
	.w4(32'h3910083b),
	.w5(32'hb9607d44),
	.w6(32'h393926b0),
	.w7(32'hb835980c),
	.w8(32'h38b729e2),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3666e7a1),
	.w1(32'hb9dce381),
	.w2(32'hb9ca963d),
	.w3(32'hba80467e),
	.w4(32'hba13adec),
	.w5(32'hb9de9015),
	.w6(32'hba01e30c),
	.w7(32'hb98c17b5),
	.w8(32'hba088a5a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5768e),
	.w1(32'hba38d4ec),
	.w2(32'hba0460f4),
	.w3(32'hba362e20),
	.w4(32'hba585f15),
	.w5(32'h38b69f39),
	.w6(32'hba83abeb),
	.w7(32'hba320e79),
	.w8(32'h37b00d3c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa2d36),
	.w1(32'hba1bde7a),
	.w2(32'h3a13b2a7),
	.w3(32'hb98cacfe),
	.w4(32'hb91aac3f),
	.w5(32'h3a885ea3),
	.w6(32'h376a97d4),
	.w7(32'hb9ddecfc),
	.w8(32'h3a653c6e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ed89a2),
	.w1(32'h3943709f),
	.w2(32'h3a58df95),
	.w3(32'h39fe6b20),
	.w4(32'h39c4ca4c),
	.w5(32'h3abd59cf),
	.w6(32'h395cf515),
	.w7(32'h3a518cea),
	.w8(32'h3a94be72),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a71823c),
	.w1(32'h398831ff),
	.w2(32'hb868cb9e),
	.w3(32'hba473b42),
	.w4(32'h3958c470),
	.w5(32'hba89bd03),
	.w6(32'hbb05f4d5),
	.w7(32'hbaa0185b),
	.w8(32'hba7bf2ab),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8055ba),
	.w1(32'hb888ade4),
	.w2(32'h3a4cc004),
	.w3(32'h39d9bec3),
	.w4(32'h3ac2f6b1),
	.w5(32'h3a8e5d63),
	.w6(32'h3b38baed),
	.w7(32'h3a736779),
	.w8(32'h3a06d150),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a216272),
	.w1(32'h39f2dcdf),
	.w2(32'h39466d91),
	.w3(32'h39d4afa8),
	.w4(32'h39283388),
	.w5(32'hba5b538b),
	.w6(32'h3a0a7fa7),
	.w7(32'h399168b4),
	.w8(32'hb9d92531),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c84d08),
	.w1(32'hb6364eb6),
	.w2(32'hb9cb430c),
	.w3(32'hb9121414),
	.w4(32'h38e00b78),
	.w5(32'h3a48d286),
	.w6(32'hb9c37bce),
	.w7(32'h39454061),
	.w8(32'h3a37760f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0cac3),
	.w1(32'h39e4a20e),
	.w2(32'h398c9a3b),
	.w3(32'h39d5ad7c),
	.w4(32'h3a349631),
	.w5(32'h395cf8f8),
	.w6(32'h3a617f1c),
	.w7(32'h3a376d18),
	.w8(32'h38a23019),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ebf77),
	.w1(32'h3a38d4a8),
	.w2(32'h3a62fbf4),
	.w3(32'h3a1dcc51),
	.w4(32'h3a9fb127),
	.w5(32'h3a44c971),
	.w6(32'h3982271c),
	.w7(32'h39be29b0),
	.w8(32'h3a27aa93),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac0f6fc),
	.w1(32'hb95dae70),
	.w2(32'hbaac257a),
	.w3(32'h39bbaeee),
	.w4(32'hbaf23048),
	.w5(32'hbaf007e9),
	.w6(32'hbae3c9be),
	.w7(32'hba8f6810),
	.w8(32'hbaf02bef),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fb07b),
	.w1(32'hbaad6bc2),
	.w2(32'hba8b19a5),
	.w3(32'hba938fbe),
	.w4(32'hba1a5bdd),
	.w5(32'h390fd603),
	.w6(32'hbb3bf1e6),
	.w7(32'hbb042fd8),
	.w8(32'hba161e3c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb876aba9),
	.w1(32'hba56b9d9),
	.w2(32'hba446ff3),
	.w3(32'hb93cbd83),
	.w4(32'hb8944844),
	.w5(32'hba7e7725),
	.w6(32'hba399f28),
	.w7(32'hba397b54),
	.w8(32'hba90422a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3dd41),
	.w1(32'hbabbbf2c),
	.w2(32'hb9ce58a7),
	.w3(32'hbb0d038a),
	.w4(32'hba6e2c29),
	.w5(32'hb99605e0),
	.w6(32'hbaed174a),
	.w7(32'hba38f0aa),
	.w8(32'hba3bcb7b),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90020bd),
	.w1(32'hb8850071),
	.w2(32'h39d1b2a6),
	.w3(32'h39a0c8fd),
	.w4(32'h3a0af97d),
	.w5(32'hb932bcae),
	.w6(32'h3a1625dc),
	.w7(32'h39c68444),
	.w8(32'hba81e29d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9a525),
	.w1(32'hb965393f),
	.w2(32'hb9cb1f29),
	.w3(32'hb9e7e0f9),
	.w4(32'hb85b2a52),
	.w5(32'h3932c168),
	.w6(32'hbaddaec6),
	.w7(32'hbaa6f686),
	.w8(32'hb94853ef),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb308193),
	.w1(32'hbb1a3af9),
	.w2(32'h39395731),
	.w3(32'hbb0d33af),
	.w4(32'hb9e3e947),
	.w5(32'h3a2124c5),
	.w6(32'hba855571),
	.w7(32'h399e3b56),
	.w8(32'h39fefe8d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398e0761),
	.w1(32'hba858433),
	.w2(32'hbb158810),
	.w3(32'h388fe9dc),
	.w4(32'hba83bc20),
	.w5(32'hbad5d590),
	.w6(32'hbbb4e174),
	.w7(32'hbb96f6aa),
	.w8(32'hbb40b6fa),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba376a10),
	.w1(32'hba0e198c),
	.w2(32'h3a062db2),
	.w3(32'h3a80cafa),
	.w4(32'h395a9ee5),
	.w5(32'h3a3733cd),
	.w6(32'h3ab7a9ac),
	.w7(32'h39ec7445),
	.w8(32'h3a83b491),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388faa13),
	.w1(32'hba2661b8),
	.w2(32'hba9277f6),
	.w3(32'h3a06ba84),
	.w4(32'h3a678165),
	.w5(32'h38cb8f23),
	.w6(32'hba6aa6fe),
	.w7(32'hba964e63),
	.w8(32'hba1b2aae),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a865a4d),
	.w1(32'hb93b1304),
	.w2(32'hba0a0efb),
	.w3(32'h385dc32e),
	.w4(32'hba8e7186),
	.w5(32'hb909942e),
	.w6(32'hbb8114cd),
	.w7(32'hbb161940),
	.w8(32'hba6b2005),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9843125),
	.w1(32'h395b8378),
	.w2(32'h3a389e30),
	.w3(32'hbaa60263),
	.w4(32'hba07a2fa),
	.w5(32'h3961a762),
	.w6(32'hba001676),
	.w7(32'hb9910288),
	.w8(32'h3910a0d2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38708635),
	.w1(32'hb9e1a6fd),
	.w2(32'h3a05bf19),
	.w3(32'h389cf40f),
	.w4(32'hb8e2a786),
	.w5(32'h3a6ad9d0),
	.w6(32'hbab8c312),
	.w7(32'hba85379c),
	.w8(32'hb962f3c1),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3866005c),
	.w1(32'h37ded312),
	.w2(32'hb809bfff),
	.w3(32'h3992aec2),
	.w4(32'h399e3955),
	.w5(32'hb7fd04c4),
	.w6(32'hb9bef704),
	.w7(32'hb96791eb),
	.w8(32'hb9f69031),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b0199),
	.w1(32'h3accaf6d),
	.w2(32'h3b131b93),
	.w3(32'h3b558194),
	.w4(32'h3afd4b70),
	.w5(32'h3ac821ff),
	.w6(32'h3b9aa3f5),
	.w7(32'h3ae8eb21),
	.w8(32'h3a343e91),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37e72d),
	.w1(32'hba8db5e9),
	.w2(32'hba9c7499),
	.w3(32'hba9d0216),
	.w4(32'hba86a548),
	.w5(32'hba38a6c8),
	.w6(32'hbab71cf9),
	.w7(32'hbaabbfb2),
	.w8(32'hba9faafb),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb809f0f8),
	.w1(32'h38d4dc4c),
	.w2(32'h3965ec16),
	.w3(32'h39718f12),
	.w4(32'h3a24da5c),
	.w5(32'h396d9511),
	.w6(32'h39eff580),
	.w7(32'h3a03ee65),
	.w8(32'hb9389fcf),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb944cb4d),
	.w1(32'hb9b78f55),
	.w2(32'h3826d994),
	.w3(32'h39738572),
	.w4(32'h390e2d75),
	.w5(32'hb94523b7),
	.w6(32'h395cecea),
	.w7(32'hb7878f0b),
	.w8(32'h385a25b8),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e21120),
	.w1(32'h392c6cd6),
	.w2(32'h3a11d912),
	.w3(32'h38ebf079),
	.w4(32'h3879ab41),
	.w5(32'hba3fb4f5),
	.w6(32'h39d77f15),
	.w7(32'hba0098d1),
	.w8(32'hba679ef6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3977678e),
	.w1(32'h3a069c86),
	.w2(32'h3a81add6),
	.w3(32'h3a1ebe23),
	.w4(32'h3a92cf11),
	.w5(32'h3ac94b28),
	.w6(32'h3a79bbba),
	.w7(32'hb94a5554),
	.w8(32'h3a66bdf6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f61969),
	.w1(32'h3ab34d17),
	.w2(32'h3b31a7a2),
	.w3(32'h39d6d380),
	.w4(32'h3adb1e7d),
	.w5(32'h3b35b17a),
	.w6(32'h3900077e),
	.w7(32'h3a02d472),
	.w8(32'h3ab25e98),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e56890),
	.w1(32'h39d9b843),
	.w2(32'h397c4e90),
	.w3(32'h38e38893),
	.w4(32'h3a3193d6),
	.w5(32'h3a42ecbc),
	.w6(32'h3a1f7323),
	.w7(32'h3a0e5475),
	.w8(32'h3a0b9ef0),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a166148),
	.w1(32'h39e8fd62),
	.w2(32'h3a67dcbe),
	.w3(32'h38c3b550),
	.w4(32'h3948256d),
	.w5(32'h3a2d979e),
	.w6(32'hba853cbe),
	.w7(32'hbab00e9c),
	.w8(32'hb9222902),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ad6d9),
	.w1(32'hb9128a0c),
	.w2(32'h3995b35a),
	.w3(32'h395029db),
	.w4(32'hba5083df),
	.w5(32'hb99a410c),
	.w6(32'hb8f6bfd6),
	.w7(32'hba8e393a),
	.w8(32'hb9e03f37),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3845dc52),
	.w1(32'hba272afe),
	.w2(32'hbadf3205),
	.w3(32'h3a46fe2f),
	.w4(32'hb992f220),
	.w5(32'hba800bf8),
	.w6(32'hbb305b2e),
	.w7(32'hbad5cb31),
	.w8(32'hbada7301),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6489514),
	.w1(32'hba16e766),
	.w2(32'hb86812fa),
	.w3(32'h3a9df087),
	.w4(32'h3ad696f5),
	.w5(32'h395f44f6),
	.w6(32'h3b064398),
	.w7(32'h3afb1ae7),
	.w8(32'h3a499382),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393af6d0),
	.w1(32'h39ccfc50),
	.w2(32'h3a2ca041),
	.w3(32'h3a638e0a),
	.w4(32'h3a2c0d1a),
	.w5(32'h39a9eb09),
	.w6(32'h3b1df07d),
	.w7(32'h3a67de9c),
	.w8(32'h384e6fe9),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e6c3a),
	.w1(32'h399d34f2),
	.w2(32'h39ed2b38),
	.w3(32'h3a8b78fa),
	.w4(32'h3ad41a16),
	.w5(32'h3aa8aac4),
	.w6(32'h3aa636f0),
	.w7(32'h3a94cc98),
	.w8(32'h3a4b31c6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e7712),
	.w1(32'hba36dc60),
	.w2(32'hb96cfbd6),
	.w3(32'hb9ca8913),
	.w4(32'hb9954f98),
	.w5(32'h3901294b),
	.w6(32'h37945930),
	.w7(32'hb7c9d23c),
	.w8(32'h3807bc91),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b5574),
	.w1(32'h3956807a),
	.w2(32'h3a945a40),
	.w3(32'h3a7f364c),
	.w4(32'h3acebbb4),
	.w5(32'h3b089598),
	.w6(32'h3b27dcd2),
	.w7(32'h3a7c88f5),
	.w8(32'h3a29c1a4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985ebd0),
	.w1(32'h3a187734),
	.w2(32'h3a0178b3),
	.w3(32'h3a77e13a),
	.w4(32'h3ab905ee),
	.w5(32'hba0a43b3),
	.w6(32'h3a9029ce),
	.w7(32'h3a99930d),
	.w8(32'hb984ef12),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba599748),
	.w1(32'hba9079ac),
	.w2(32'hbac2ac68),
	.w3(32'hb9d61f49),
	.w4(32'hb99a7bea),
	.w5(32'hba6c02f2),
	.w6(32'hbb0d547b),
	.w7(32'hba36b746),
	.w8(32'hb87c80b2),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15268e),
	.w1(32'h3a18a937),
	.w2(32'h3a46e01f),
	.w3(32'h3a0e0c7b),
	.w4(32'hb8e4d269),
	.w5(32'hb9d4ef77),
	.w6(32'h3a4959e2),
	.w7(32'h3a2326ab),
	.w8(32'hb7f08cb1),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6e0615),
	.w1(32'h39eec5bf),
	.w2(32'h3a8c9551),
	.w3(32'h3a8cdf34),
	.w4(32'h39c44c4d),
	.w5(32'h3a7290c4),
	.w6(32'hb9c9ead6),
	.w7(32'hba0e0227),
	.w8(32'h395bcded),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38350c08),
	.w1(32'h394217bc),
	.w2(32'hb9838b5b),
	.w3(32'h399e5b10),
	.w4(32'h38cbbaa4),
	.w5(32'h39ad32d9),
	.w6(32'hb8736984),
	.w7(32'hb7f3afa1),
	.w8(32'h3a031c80),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3813c2b0),
	.w1(32'hb82a3230),
	.w2(32'h3a3f768e),
	.w3(32'hb90872ae),
	.w4(32'h3a0d378e),
	.w5(32'h3a82d929),
	.w6(32'h3a21e288),
	.w7(32'h3a8345a5),
	.w8(32'h396d9145),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38848851),
	.w1(32'hb61772de),
	.w2(32'h3822aa72),
	.w3(32'hb89c2ac3),
	.w4(32'h39519a7a),
	.w5(32'h3974ca2a),
	.w6(32'hb9738e93),
	.w7(32'h38d4d66e),
	.w8(32'h38f67c37),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a85e11d),
	.w1(32'h39dbdab7),
	.w2(32'hb9ab83ae),
	.w3(32'h3ac2ef3c),
	.w4(32'h3a381669),
	.w5(32'hb92a95c8),
	.w6(32'h3a684a9b),
	.w7(32'hb90ae3ac),
	.w8(32'hba5d780d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b424f5),
	.w1(32'hb93357b2),
	.w2(32'hb898a2c7),
	.w3(32'h38a3ecc7),
	.w4(32'h3a018f70),
	.w5(32'h3934c246),
	.w6(32'h3a264cd1),
	.w7(32'h39c8d12d),
	.w8(32'h38302473),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990cf5b),
	.w1(32'h388413dd),
	.w2(32'hb99fbfc2),
	.w3(32'h3779c57f),
	.w4(32'hb9670d88),
	.w5(32'h3a84c723),
	.w6(32'h3944677d),
	.w7(32'h39af91d2),
	.w8(32'h39d54cf5),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7b59f),
	.w1(32'h39c5c823),
	.w2(32'h3af62735),
	.w3(32'h3a993e22),
	.w4(32'h3ac42417),
	.w5(32'h3ac9c38f),
	.w6(32'h3ae3332e),
	.w7(32'h3af63031),
	.w8(32'h3ae13f31),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ce44de),
	.w1(32'hbaba8092),
	.w2(32'hbb31e6a5),
	.w3(32'hbb053889),
	.w4(32'hbb729b08),
	.w5(32'hbb42dd5e),
	.w6(32'hbbbb56b5),
	.w7(32'hbbcd464f),
	.w8(32'hbb9970ca),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35ae09),
	.w1(32'h3a2aea4e),
	.w2(32'h398eb72a),
	.w3(32'h3a94d01f),
	.w4(32'h3a9f1b72),
	.w5(32'hba2f1c1b),
	.w6(32'h3aadca4e),
	.w7(32'h3a741323),
	.w8(32'h37aff477),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8be44ab),
	.w1(32'hb8f047fe),
	.w2(32'hb95db102),
	.w3(32'h39a4c5f8),
	.w4(32'hba069406),
	.w5(32'hbb195dd2),
	.w6(32'h3aef5aa7),
	.w7(32'hb988284f),
	.w8(32'hbb0d2a65),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca2759),
	.w1(32'hbaa16b66),
	.w2(32'hba8eec94),
	.w3(32'hba8d4f58),
	.w4(32'hba19974a),
	.w5(32'hba36a79f),
	.w6(32'hb74101cc),
	.w7(32'hba4d1a51),
	.w8(32'hb8eee319),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b798b5),
	.w1(32'h3a6e28cc),
	.w2(32'h3a57f021),
	.w3(32'hb9e842ed),
	.w4(32'hb97e0b38),
	.w5(32'h3a99e763),
	.w6(32'hbaeecd74),
	.w7(32'hbaaa31c3),
	.w8(32'h3a47cc5a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a6cffd),
	.w1(32'hb94f5972),
	.w2(32'hb961c394),
	.w3(32'h3935972e),
	.w4(32'h3a54d075),
	.w5(32'hb95569de),
	.w6(32'hbac6527f),
	.w7(32'hba3a8e01),
	.w8(32'hba41efcb),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9925320),
	.w1(32'hbb0185d6),
	.w2(32'hbb1582c6),
	.w3(32'hbb3514ec),
	.w4(32'hbb4212e2),
	.w5(32'hbaec54e4),
	.w6(32'hbbc05899),
	.w7(32'hbba49d5f),
	.w8(32'hbb377c19),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a24828d),
	.w1(32'hb752afcd),
	.w2(32'h39ac1242),
	.w3(32'h3a136f9d),
	.w4(32'h3a4991c4),
	.w5(32'h39f5c3d9),
	.w6(32'h39c21a47),
	.w7(32'h3a665e26),
	.w8(32'h3a2866f9),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918b1b2),
	.w1(32'hba3295bf),
	.w2(32'hb911923e),
	.w3(32'h3a3f3a79),
	.w4(32'h39f86614),
	.w5(32'h3ac2ce8d),
	.w6(32'hb9171e1a),
	.w7(32'hb90b57ad),
	.w8(32'h3a833c6e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e21ce),
	.w1(32'hb67262e5),
	.w2(32'h395f9b4c),
	.w3(32'h38a69f32),
	.w4(32'h39be68fd),
	.w5(32'hb9a3397b),
	.w6(32'hb9344f4a),
	.w7(32'hb78a104e),
	.w8(32'hb991491e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba093c5f),
	.w1(32'h3912a3fb),
	.w2(32'h3a321a57),
	.w3(32'h39e3399d),
	.w4(32'h3a200571),
	.w5(32'h38da6719),
	.w6(32'hb90b35d8),
	.w7(32'h392dcd6f),
	.w8(32'h3a243cf9),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ad8447),
	.w1(32'hba1c2361),
	.w2(32'h3872b2f5),
	.w3(32'hb9656800),
	.w4(32'h390679e7),
	.w5(32'hb7f0a355),
	.w6(32'hb8f8548c),
	.w7(32'h39e3c8ef),
	.w8(32'hb8fdaeda),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90728de),
	.w1(32'hb7ba3b60),
	.w2(32'hb4e26750),
	.w3(32'h38e62d0e),
	.w4(32'hb9a8f0e6),
	.w5(32'h3a5d9a18),
	.w6(32'hb9ba6322),
	.w7(32'hba7c5727),
	.w8(32'hb922255a),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb885b44e),
	.w1(32'hba8a2742),
	.w2(32'h3a1edda8),
	.w3(32'hba4bfa1d),
	.w4(32'h39f65453),
	.w5(32'h3881ce01),
	.w6(32'hba531ef9),
	.w7(32'h3a00b24b),
	.w8(32'h3833e319),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4578f),
	.w1(32'h39ebe5a1),
	.w2(32'h396bed2b),
	.w3(32'h39accc69),
	.w4(32'h3a368cfd),
	.w5(32'hb959316f),
	.w6(32'h39a37a30),
	.w7(32'h3a160972),
	.w8(32'hb8d79488),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6dfe0e),
	.w1(32'h3909a9eb),
	.w2(32'h37f102a3),
	.w3(32'h396a0efd),
	.w4(32'h38751f6a),
	.w5(32'h3a7ff858),
	.w6(32'h3a061519),
	.w7(32'h384fb7b3),
	.w8(32'h3a1a3bd8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4673cf),
	.w1(32'h3b255764),
	.w2(32'h3b02ee57),
	.w3(32'h3b5b806c),
	.w4(32'h3ab8f2e7),
	.w5(32'h3a959afa),
	.w6(32'h3b116948),
	.w7(32'h39aefd96),
	.w8(32'hba00ec7a),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade4685),
	.w1(32'hba09a82b),
	.w2(32'hb84682ff),
	.w3(32'hba4c3209),
	.w4(32'h394f6471),
	.w5(32'h3a80833d),
	.w6(32'hba989953),
	.w7(32'hba9273e8),
	.w8(32'hba7a6868),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ce8e6e),
	.w1(32'hba916376),
	.w2(32'hba998e3f),
	.w3(32'hba7bef06),
	.w4(32'hba6b8b69),
	.w5(32'hbab2f3b7),
	.w6(32'hbacfce2a),
	.w7(32'hba919d36),
	.w8(32'hbb09e398),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae50ee),
	.w1(32'hba91a3b5),
	.w2(32'hbabb62cf),
	.w3(32'h3a161649),
	.w4(32'hbae5b3cf),
	.w5(32'hb97247b8),
	.w6(32'hbb9558b0),
	.w7(32'hbb8ab045),
	.w8(32'hbab6a10f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba235ac3),
	.w1(32'hba9ca981),
	.w2(32'h38d84d62),
	.w3(32'h3b2a6f2f),
	.w4(32'h3b49a55d),
	.w5(32'h3aa86bf2),
	.w6(32'h3b81962a),
	.w7(32'h3b354173),
	.w8(32'h3b1aa027),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2398aa),
	.w1(32'h3983bba6),
	.w2(32'h39754238),
	.w3(32'h3a32c810),
	.w4(32'h3a98c34f),
	.w5(32'h3a11dbd6),
	.w6(32'h39ed8d53),
	.w7(32'h38b6c351),
	.w8(32'hb9ca4e77),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eae2b8),
	.w1(32'h390fbc05),
	.w2(32'h38de6542),
	.w3(32'h398b8124),
	.w4(32'h3a0f6809),
	.w5(32'h39cba5ea),
	.w6(32'hb938eb0c),
	.w7(32'h38c208af),
	.w8(32'h3988e7ce),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36856eea),
	.w1(32'h382b84d6),
	.w2(32'hb604f80c),
	.w3(32'h38a658b6),
	.w4(32'hb8673c1d),
	.w5(32'h39e1e493),
	.w6(32'h38e3e936),
	.w7(32'hb8de89e6),
	.w8(32'h3918973d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4f8f0),
	.w1(32'h39e08609),
	.w2(32'h3a3ea36e),
	.w3(32'h3a1f6703),
	.w4(32'h3a78ffcd),
	.w5(32'hb9ce1c25),
	.w6(32'h39e2314b),
	.w7(32'h3a87df74),
	.w8(32'hb9cb5dc5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e635e),
	.w1(32'h3a46a401),
	.w2(32'h39b4f32d),
	.w3(32'h3a887e48),
	.w4(32'h3a2c2792),
	.w5(32'h39958d94),
	.w6(32'hba15069e),
	.w7(32'h37535502),
	.w8(32'hb9846fec),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38518dd3),
	.w1(32'hb9039a03),
	.w2(32'hb8fd880e),
	.w3(32'h39dba59d),
	.w4(32'hb95915a4),
	.w5(32'hb99c205a),
	.w6(32'hbaaa67ce),
	.w7(32'hbb09fb49),
	.w8(32'hbb2c403c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c50672),
	.w1(32'hb901040a),
	.w2(32'h3b25f594),
	.w3(32'hb86ad09c),
	.w4(32'h3ade5545),
	.w5(32'h3b0d1ad4),
	.w6(32'h3aa35be3),
	.w7(32'h3ae611fd),
	.w8(32'h3b0141bb),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a63d6f),
	.w1(32'h3a198d55),
	.w2(32'h3a8e7f31),
	.w3(32'h398be63b),
	.w4(32'h3a2993e5),
	.w5(32'h368d170a),
	.w6(32'h3a12299f),
	.w7(32'h3a2a5f7b),
	.w8(32'hb9a81061),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154f97),
	.w1(32'h3a1e160b),
	.w2(32'h39c0d317),
	.w3(32'h3a9c276f),
	.w4(32'h3a574971),
	.w5(32'hba16ec23),
	.w6(32'hb9d33903),
	.w7(32'hbae88d79),
	.w8(32'hbac643de),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b372a2),
	.w1(32'h394a8c70),
	.w2(32'h399be1fa),
	.w3(32'hb85e66e8),
	.w4(32'hb8bc2a0e),
	.w5(32'h39bfd7b0),
	.w6(32'h3a5e5c27),
	.w7(32'h38cf8f36),
	.w8(32'h39141a4e),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8617498),
	.w1(32'hb8df6d17),
	.w2(32'hb980b69e),
	.w3(32'h3965366a),
	.w4(32'hb96df4cf),
	.w5(32'h3884d82e),
	.w6(32'hb73a53a2),
	.w7(32'h375f578e),
	.w8(32'hb95086be),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39916a98),
	.w1(32'hb966a9a8),
	.w2(32'hb9f8661b),
	.w3(32'hba8f1a17),
	.w4(32'hba810e5b),
	.w5(32'hb963c7f4),
	.w6(32'hba814f53),
	.w7(32'hb9e14025),
	.w8(32'hb8963c71),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b53fa),
	.w1(32'h399ec0f6),
	.w2(32'h38e6ecc5),
	.w3(32'hb8fcb16f),
	.w4(32'hb8f3445e),
	.w5(32'hb8020b15),
	.w6(32'h39af0ab6),
	.w7(32'hb8eda3f5),
	.w8(32'h39bea45a),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a35c97),
	.w1(32'hba1ec7c6),
	.w2(32'hb9b90911),
	.w3(32'hbab20605),
	.w4(32'hb9a3ec6c),
	.w5(32'hb9d37265),
	.w6(32'hbab67add),
	.w7(32'hba423334),
	.w8(32'hba4784f3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c3330),
	.w1(32'hb81093f5),
	.w2(32'h3a31bd05),
	.w3(32'h3a878f32),
	.w4(32'h3aa728e8),
	.w5(32'h3a834526),
	.w6(32'h3b307fd9),
	.w7(32'h3a9a0286),
	.w8(32'h3a163d9a),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380956fd),
	.w1(32'hb99f0fbc),
	.w2(32'h37710a32),
	.w3(32'h3a48dee8),
	.w4(32'h38d057b5),
	.w5(32'hba2460c8),
	.w6(32'h3a64580b),
	.w7(32'h396c5c7d),
	.w8(32'hb99d0a74),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb995db4c),
	.w1(32'hb8fac47e),
	.w2(32'hb989ef90),
	.w3(32'hb908f0b0),
	.w4(32'h38f5ca38),
	.w5(32'h3945c9e1),
	.w6(32'hb8af1833),
	.w7(32'h3949035d),
	.w8(32'h39c4242b),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c56f0),
	.w1(32'h3a683be9),
	.w2(32'h3b03a05b),
	.w3(32'h3ad2c4f3),
	.w4(32'h3aab7d85),
	.w5(32'h3a8a176c),
	.w6(32'h3b1bc37d),
	.w7(32'h3ae92b28),
	.w8(32'h3abd5d81),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba202664),
	.w1(32'hba9d8103),
	.w2(32'hb9f6f1a5),
	.w3(32'hba91982a),
	.w4(32'hba3e88fc),
	.w5(32'hb9833fba),
	.w6(32'hbabfd680),
	.w7(32'hba9fd6b8),
	.w8(32'hb9e97c29),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb962b96f),
	.w1(32'h39fbb76c),
	.w2(32'h3a9fdabe),
	.w3(32'h3aaa724a),
	.w4(32'h3a3abdb7),
	.w5(32'h3b20502e),
	.w6(32'hb8989eb4),
	.w7(32'hbaaa587b),
	.w8(32'h399f4c7b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ceebb8),
	.w1(32'hb80598fc),
	.w2(32'hb8db740c),
	.w3(32'h3397edf5),
	.w4(32'hb9267f1c),
	.w5(32'hb8d29244),
	.w6(32'h38ff26a1),
	.w7(32'hb98aeae5),
	.w8(32'hb8b6df1a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b93c49),
	.w1(32'hb9140a1f),
	.w2(32'h3968856d),
	.w3(32'hb90b5d43),
	.w4(32'h39375bf4),
	.w5(32'h39a0325d),
	.w6(32'hb88c9fa6),
	.w7(32'h39fb1111),
	.w8(32'h39967acf),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12054f),
	.w1(32'h3ac7f9dc),
	.w2(32'h3b093b5e),
	.w3(32'h3a959c00),
	.w4(32'h3b0318ce),
	.w5(32'h3a63db0c),
	.w6(32'h3b013c54),
	.w7(32'h3a0b060d),
	.w8(32'h3913e8b9),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abaa2a3),
	.w1(32'hba3208f4),
	.w2(32'hbb1c445c),
	.w3(32'hbadbb4fa),
	.w4(32'hbb4ca991),
	.w5(32'hbb22e6f8),
	.w6(32'hbb8c0401),
	.w7(32'hbb8d7577),
	.w8(32'hbb96f8d0),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947c309),
	.w1(32'h39f1f0ec),
	.w2(32'h3a98eeaa),
	.w3(32'hb911ed7d),
	.w4(32'h3a0575ec),
	.w5(32'h3a3e1d09),
	.w6(32'h3a1840b4),
	.w7(32'h3a19f190),
	.w8(32'hb9a6c30c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba315e86),
	.w1(32'hb93562f7),
	.w2(32'h3a0ce687),
	.w3(32'h3a4dbf69),
	.w4(32'h3ab2d200),
	.w5(32'h3a04e96a),
	.w6(32'hb9aaf75f),
	.w7(32'hb9dadc0c),
	.w8(32'hb8d819c0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7188c62),
	.w1(32'hb93e4fea),
	.w2(32'hb7a2406d),
	.w3(32'h396fc5be),
	.w4(32'h3a1136c4),
	.w5(32'hb83c41db),
	.w6(32'hb8edd835),
	.w7(32'h39b23b25),
	.w8(32'hb8c2bc49),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3561871a),
	.w1(32'hb9d8cca0),
	.w2(32'hb965ffeb),
	.w3(32'hb9357d7b),
	.w4(32'hb8cd6d30),
	.w5(32'h3a83fb78),
	.w6(32'hb9616c24),
	.w7(32'hb9fb57ae),
	.w8(32'h3a266ebe),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37854705),
	.w1(32'h3afd9b3c),
	.w2(32'h39ac2769),
	.w3(32'h3aa2ab27),
	.w4(32'h3ac1d9a2),
	.w5(32'hb9e6b88c),
	.w6(32'hbaa397ae),
	.w7(32'h390bd238),
	.w8(32'hbaa43166),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa74086),
	.w1(32'hb9269109),
	.w2(32'h385eed67),
	.w3(32'hba7aa3a5),
	.w4(32'hba6094f1),
	.w5(32'hbaa86ffe),
	.w6(32'hbb92be30),
	.w7(32'hbb0c843c),
	.w8(32'hbb2f88f8),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998fab1),
	.w1(32'h3a5627c4),
	.w2(32'hba89a7e1),
	.w3(32'h37fa3f8d),
	.w4(32'hb88e569b),
	.w5(32'hbb22fbc2),
	.w6(32'hbb6c5048),
	.w7(32'hbb8d5cdb),
	.w8(32'hbb68e6e3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d3146),
	.w1(32'hb89d35f5),
	.w2(32'h3a0ef3ea),
	.w3(32'hb707b4b1),
	.w4(32'h3a649c46),
	.w5(32'h3a4de76f),
	.w6(32'h3ab07cba),
	.w7(32'h39e313db),
	.w8(32'h3a1527db),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2f6d3),
	.w1(32'hb9ead007),
	.w2(32'h3a30c63e),
	.w3(32'h3a1ca159),
	.w4(32'h3a589814),
	.w5(32'h3a43f382),
	.w6(32'h3b0eab06),
	.w7(32'h3a9c5974),
	.w8(32'h3a2c055b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c890b9),
	.w1(32'hb8a26c09),
	.w2(32'hb923ef65),
	.w3(32'h398f118e),
	.w4(32'h39a83588),
	.w5(32'hba99ab95),
	.w6(32'h39fa675a),
	.w7(32'h39c513ce),
	.w8(32'hb90325e8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cd594),
	.w1(32'hba221911),
	.w2(32'hb9b77b33),
	.w3(32'hb8887a70),
	.w4(32'hb7ac07c3),
	.w5(32'h3a18b666),
	.w6(32'h38d9e75b),
	.w7(32'hb813ca47),
	.w8(32'h39ff01ae),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83f03f),
	.w1(32'h3a6af168),
	.w2(32'h3a83ceff),
	.w3(32'h3a5ddca7),
	.w4(32'h3a515c53),
	.w5(32'h39c5424d),
	.w6(32'hb9a63b94),
	.w7(32'h3a062d5c),
	.w8(32'h3831e58f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9147020),
	.w1(32'hb93b6c3b),
	.w2(32'hba770877),
	.w3(32'h391148fc),
	.w4(32'hba5e58a5),
	.w5(32'h3acaf6f3),
	.w6(32'h394e1fd2),
	.w7(32'hba2391df),
	.w8(32'hba99f88b),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5188c6),
	.w1(32'h3b156c39),
	.w2(32'h3a9b853a),
	.w3(32'h3b839aeb),
	.w4(32'h3b21a7ae),
	.w5(32'hbaf1a11f),
	.w6(32'h39d57c63),
	.w7(32'h3a45c5b7),
	.w8(32'hbaf91c27),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf29bd),
	.w1(32'hbb48ae91),
	.w2(32'hbb80dcfa),
	.w3(32'hba41ace3),
	.w4(32'hbaf9db25),
	.w5(32'hba7e043c),
	.w6(32'hbb3b99ac),
	.w7(32'hbb762cd5),
	.w8(32'hbb80008d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab913aa),
	.w1(32'h3b53657f),
	.w2(32'h3b874780),
	.w3(32'h3b57c390),
	.w4(32'h3b3dd7fc),
	.w5(32'h3b62e1aa),
	.w6(32'h3ab19fdc),
	.w7(32'h3a383f9b),
	.w8(32'hba87a753),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2422ea),
	.w1(32'hbb5bf94c),
	.w2(32'hbb3fc700),
	.w3(32'h3c115a58),
	.w4(32'h3c029353),
	.w5(32'hbaa291e3),
	.w6(32'hbb773bde),
	.w7(32'hbb78bced),
	.w8(32'hba903c62),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a864869),
	.w1(32'h384aaab5),
	.w2(32'hbb23501c),
	.w3(32'hba22f357),
	.w4(32'hbb1fb810),
	.w5(32'hbb85982c),
	.w6(32'hbbb88eeb),
	.w7(32'hbb9eeacf),
	.w8(32'hbbaba835),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6a78f),
	.w1(32'hbba3c7b5),
	.w2(32'hbba9ac55),
	.w3(32'hbb2e2fca),
	.w4(32'hbaff21af),
	.w5(32'h3b21e604),
	.w6(32'hbbaee687),
	.w7(32'hbb9236a3),
	.w8(32'h3b4bd095),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33d153),
	.w1(32'h3b873156),
	.w2(32'h3b3990e6),
	.w3(32'h3bbd9a03),
	.w4(32'h3c16e44d),
	.w5(32'hbac1d5b3),
	.w6(32'h3ba3bb35),
	.w7(32'h3bc01cf9),
	.w8(32'hbb4e9ac2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb53096e),
	.w1(32'hbb33b53e),
	.w2(32'hbb44b161),
	.w3(32'hbac927e2),
	.w4(32'hbb2956bc),
	.w5(32'h394ae3fa),
	.w6(32'hbba07480),
	.w7(32'hbb8b03db),
	.w8(32'hbb100e99),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00be94),
	.w1(32'h3af44b8c),
	.w2(32'hbb2fd7aa),
	.w3(32'h38e0dcf7),
	.w4(32'h3ab63f7e),
	.w5(32'hbb0b882e),
	.w6(32'h3ab7947e),
	.w7(32'h3adb9ffb),
	.w8(32'hbab3b1e0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5c224),
	.w1(32'h38e929df),
	.w2(32'hb9da541e),
	.w3(32'hbb0c7dcf),
	.w4(32'hbab8d57a),
	.w5(32'h3b0d4878),
	.w6(32'hbaf24832),
	.w7(32'hb91935c8),
	.w8(32'hbb2c4551),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0cb24),
	.w1(32'h3ae8d1c4),
	.w2(32'h3b193bd6),
	.w3(32'h3b69818a),
	.w4(32'h3b4c58c0),
	.w5(32'hba4c5877),
	.w6(32'hba3059ca),
	.w7(32'h3b005ba9),
	.w8(32'hbb31b6d0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa97189),
	.w1(32'h3b4738fd),
	.w2(32'h3ab140ee),
	.w3(32'h3b0c6aab),
	.w4(32'hbaa6763c),
	.w5(32'hbb962059),
	.w6(32'h37d99124),
	.w7(32'hba4c0595),
	.w8(32'h38af66f6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38a06b),
	.w1(32'h3a95b038),
	.w2(32'hba7fe94a),
	.w3(32'hbb250412),
	.w4(32'hb8d8bb5e),
	.w5(32'h3b986910),
	.w6(32'h3b627d85),
	.w7(32'h3b042d81),
	.w8(32'h3bcb1460),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f5210),
	.w1(32'hbb209743),
	.w2(32'hbb6757a5),
	.w3(32'h3a83223c),
	.w4(32'hbaec076c),
	.w5(32'h3a470cda),
	.w6(32'hbb07d90d),
	.w7(32'hbb985235),
	.w8(32'hb9a43dd2),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac32b1e),
	.w1(32'h3b4e63ec),
	.w2(32'h3a4bbf76),
	.w3(32'h394f5123),
	.w4(32'hbb15d22e),
	.w5(32'hbaaf70cc),
	.w6(32'hb9f0352f),
	.w7(32'hbaa99b5c),
	.w8(32'hbafe2343),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39889ce9),
	.w1(32'h3aa8c1e4),
	.w2(32'hba4eb601),
	.w3(32'hbb1dc016),
	.w4(32'hbb1909fa),
	.w5(32'hba3b9d7c),
	.w6(32'hbb19c480),
	.w7(32'hbb67803c),
	.w8(32'hba69d211),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ca381b),
	.w1(32'hbab9e2b4),
	.w2(32'h3b89670f),
	.w3(32'hbae9740d),
	.w4(32'hba05a0dc),
	.w5(32'h3b2334a6),
	.w6(32'hbb3f686a),
	.w7(32'h3a2bc6f6),
	.w8(32'h3b901b24),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946ee81),
	.w1(32'hbaa3352c),
	.w2(32'hbadc5db3),
	.w3(32'h3bbc00fe),
	.w4(32'h3b28a58a),
	.w5(32'h3b2085a8),
	.w6(32'h3ad27891),
	.w7(32'hba3d8499),
	.w8(32'hb9a1311f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9235c),
	.w1(32'h3b68b9b0),
	.w2(32'h3bc87cc9),
	.w3(32'h3bc45608),
	.w4(32'h3b822363),
	.w5(32'hba6b3e2d),
	.w6(32'h3b50282b),
	.w7(32'h3b5ee3ba),
	.w8(32'h3b11482e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae87b2),
	.w1(32'hba736417),
	.w2(32'hbae4beb1),
	.w3(32'hbb156d6d),
	.w4(32'hbaa0a15c),
	.w5(32'hb9216b58),
	.w6(32'hbaf3b89d),
	.w7(32'hb9e5eda6),
	.w8(32'hbb552ba8),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7b51),
	.w1(32'hb9f773fb),
	.w2(32'hbacf829e),
	.w3(32'hb9e171a5),
	.w4(32'hbb0a4a5e),
	.w5(32'h3afc1da7),
	.w6(32'hbba1803c),
	.w7(32'hbb983dcd),
	.w8(32'hbba47dd5),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68b273),
	.w1(32'h39ae2172),
	.w2(32'h39405bc3),
	.w3(32'h3b625431),
	.w4(32'h3b1a85da),
	.w5(32'h3a6116b2),
	.w6(32'hbad234dc),
	.w7(32'hbb2e253e),
	.w8(32'h3b0f065e),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921c568),
	.w1(32'hba6cf258),
	.w2(32'hba6f5511),
	.w3(32'h3a4c85e0),
	.w4(32'h3acab09e),
	.w5(32'h3a0f25e7),
	.w6(32'h3b2a4540),
	.w7(32'h3ab90170),
	.w8(32'h3af08afd),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9823167),
	.w1(32'h3a682f34),
	.w2(32'h39e3ae5a),
	.w3(32'hb92a2fc9),
	.w4(32'hbaac28cc),
	.w5(32'hbb8409bc),
	.w6(32'h3a0d29d0),
	.w7(32'hb99568d3),
	.w8(32'hbb970634),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb88b02),
	.w1(32'hbbd382e5),
	.w2(32'hbba88f1d),
	.w3(32'hbba535dd),
	.w4(32'hbb833981),
	.w5(32'hbb47a973),
	.w6(32'hbb9b50e2),
	.w7(32'hbb97f15c),
	.w8(32'hbb57c3f5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f18aa),
	.w1(32'h390ee9bb),
	.w2(32'h3a26247d),
	.w3(32'hbada5aca),
	.w4(32'hbaef13c3),
	.w5(32'hbb9b1941),
	.w6(32'hbb179ea6),
	.w7(32'hb9bcc220),
	.w8(32'hbb85e8f1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb900164),
	.w1(32'hbb8e2528),
	.w2(32'hbb8f4ff0),
	.w3(32'hbb8d144e),
	.w4(32'hbb71b3d2),
	.w5(32'h3b447842),
	.w6(32'hbb253e82),
	.w7(32'hbaf74f91),
	.w8(32'h3a3571e4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9acf4a),
	.w1(32'h3a3d5a10),
	.w2(32'hbb4d3271),
	.w3(32'h3b0c51b0),
	.w4(32'h3ad52546),
	.w5(32'h39b2b050),
	.w6(32'hbb6acc0b),
	.w7(32'hbb9c54e2),
	.w8(32'hbab4997a),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4f0f02),
	.w1(32'h3b44325b),
	.w2(32'h3b1ffeef),
	.w3(32'h3a865d25),
	.w4(32'hb9c22660),
	.w5(32'h3ad26680),
	.w6(32'hbacf8ff3),
	.w7(32'hbadd9f7b),
	.w8(32'hb9cecd30),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39512a7f),
	.w1(32'hba467c6b),
	.w2(32'h3b15f47b),
	.w3(32'hbb8ac556),
	.w4(32'hb7d8b67b),
	.w5(32'hbb0d5462),
	.w6(32'hbb224fd1),
	.w7(32'hb875f137),
	.w8(32'hbb209b8f),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule